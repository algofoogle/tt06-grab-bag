magic
tech sky130A
magscale 1 2
timestamp 1712719843
<< metal1 >>
rect 29432 44410 29632 44420
rect 29432 44350 29502 44410
rect 29562 44350 29632 44410
rect 17660 43260 17860 43266
rect 17660 41610 17860 43060
rect 17660 41410 19910 41610
rect 19710 8190 19910 41410
rect 19704 7990 19710 8190
rect 19910 7990 19916 8190
rect 29432 7686 29632 44350
rect 29432 7486 30410 7686
rect 29432 7480 29632 7486
rect 11598 7037 11604 7237
rect 11804 7037 30116 7237
rect 2102 5937 2108 6137
rect 2308 5937 28688 6137
rect 30204 6090 30404 7486
rect 29920 5892 30404 6090
rect 19710 4770 19910 4776
rect 29916 4770 30116 5357
rect 19910 4570 30116 4770
rect 19710 4564 19910 4570
rect 29916 2070 30116 4570
rect 31270 2070 31470 2076
rect 29916 1870 31270 2070
rect 31270 1864 31470 1870
<< via1 >>
rect 29502 44350 29562 44410
rect 17660 43060 17860 43260
rect 19710 7990 19910 8190
rect 11604 7037 11804 7237
rect 2108 5937 2308 6137
rect 19710 4570 19910 4770
rect 31270 1870 31470 2070
<< metal2 >>
rect 29502 44590 29562 44592
rect 29495 44534 29504 44590
rect 29560 44534 29569 44590
rect 29502 44410 29562 44534
rect 29502 44344 29562 44350
rect 17660 43700 17860 43709
rect 17660 43260 17860 43500
rect 17654 43060 17660 43260
rect 17860 43060 17866 43260
rect 19710 8190 19910 8196
rect 11604 7237 11804 7243
rect 11147 7037 11156 7237
rect 11356 7037 11604 7237
rect 11604 7031 11804 7037
rect 2108 6137 2308 6143
rect 1611 5937 1620 6137
rect 1820 5937 2108 6137
rect 2108 5931 2308 5937
rect 19710 4770 19910 7990
rect 19704 4570 19710 4770
rect 19910 4570 19916 4770
rect 31264 1870 31270 2070
rect 31470 1870 31476 2070
rect 31270 1660 31470 1870
rect 31270 1451 31470 1460
<< via2 >>
rect 29504 44534 29560 44590
rect 17660 43500 17860 43700
rect 11156 7037 11356 7237
rect 1620 5937 1820 6137
rect 31270 1460 31470 1660
<< metal3 >>
rect 29494 44752 29500 44816
rect 29564 44752 29570 44816
rect 29502 44595 29562 44752
rect 29499 44590 29565 44595
rect 29499 44534 29504 44590
rect 29560 44534 29565 44590
rect 29499 44529 29565 44534
rect 17660 44090 17860 44096
rect 17660 43705 17860 43890
rect 17655 43700 17865 43705
rect 17655 43500 17660 43700
rect 17860 43500 17865 43700
rect 17655 43495 17865 43500
rect 11151 7237 11361 7242
rect 10664 7037 10670 7237
rect 10870 7037 11156 7237
rect 11356 7037 11361 7237
rect 11151 7032 11361 7037
rect 1615 6137 1825 6142
rect 1078 5937 1084 6137
rect 1284 5937 1620 6137
rect 1820 5937 1825 6137
rect 1615 5932 1825 5937
rect 31265 1660 31475 1665
rect 31265 1460 31270 1660
rect 31470 1460 31475 1660
rect 31265 1455 31475 1460
rect 31270 1240 31470 1455
rect 31270 1034 31470 1040
<< via3 >>
rect 29500 44752 29564 44816
rect 17660 43890 17860 44090
rect 10670 7037 10870 7237
rect 1084 5937 1284 6137
rect 31270 1040 31470 1240
<< metal4 >>
rect 798 44438 858 45152
rect 1534 44438 1594 45152
rect 2270 44438 2330 45152
rect 3006 44438 3066 45152
rect 3742 44438 3802 45152
rect 4478 44438 4538 45152
rect 5214 44438 5274 45152
rect 5950 44438 6010 45152
rect 6686 44438 6746 45152
rect 7422 44438 7482 45152
rect 8158 44438 8218 45152
rect 8894 44438 8954 45152
rect 9630 44438 9690 45152
rect 10366 44438 10426 45152
rect 11102 44438 11162 45152
rect 11838 44438 11898 45152
rect 12574 44438 12634 45152
rect 13310 44438 13370 45152
rect 14046 44438 14106 45152
rect 14782 44438 14842 45152
rect 15518 44438 15578 45152
rect 16254 44438 16314 45152
rect 16990 44438 17050 45152
rect 17726 44620 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44817 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29499 44816 29565 44817
rect 29499 44752 29500 44816
rect 29564 44752 29565 44816
rect 29499 44751 29565 44752
rect 200 6137 500 44152
rect 748 43926 17168 44438
rect 17660 44091 17860 44620
rect 17659 44090 17861 44091
rect 9800 7237 10100 43926
rect 17659 43890 17660 44090
rect 17860 43890 17861 44090
rect 17659 43889 17861 43890
rect 10669 7237 10871 7238
rect 9800 7037 10670 7237
rect 10870 7037 10871 7237
rect 1083 6137 1285 6138
rect 200 5937 1084 6137
rect 1284 5937 1285 6137
rect 200 1000 500 5937
rect 1083 5936 1285 5937
rect 9800 1000 10100 7037
rect 10669 7036 10871 7037
rect 31269 1240 31471 1241
rect 31269 1040 31270 1240
rect 31470 1040 31471 1240
rect 31269 1039 31471 1040
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31306 46 31435 1039
rect 31312 0 31432 46
use inverter  inverter_0
timestamp 1712241802
transform 1 0 28896 0 1 4427
box -410 547 1220 2810
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
