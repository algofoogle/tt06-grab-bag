magic
tech sky130A
magscale 1 2
timestamp 1713486661
<< viali >>
rect 1225 17289 1259 17323
rect 2053 17289 2087 17323
rect 4077 17289 4111 17323
rect 4721 17289 4755 17323
rect 5917 17289 5951 17323
rect 7297 17289 7331 17323
rect 8125 17289 8159 17323
rect 8861 17289 8895 17323
rect 5273 17221 5307 17255
rect 6561 17221 6595 17255
rect 7665 17221 7699 17255
rect 12725 17221 12759 17255
rect 13553 17221 13587 17255
rect 13829 17221 13863 17255
rect 2973 17153 3007 17187
rect 8493 17153 8527 17187
rect 11529 17153 11563 17187
rect 11621 17153 11655 17187
rect 12449 17153 12483 17187
rect 16221 17153 16255 17187
rect 1501 17085 1535 17119
rect 1869 17085 1903 17119
rect 2237 17085 2271 17119
rect 3801 17085 3835 17119
rect 4261 17085 4295 17119
rect 4905 17085 4939 17119
rect 6837 17085 6871 17119
rect 7113 17085 7147 17119
rect 7481 17085 7515 17119
rect 7941 17085 7975 17119
rect 8585 17085 8619 17119
rect 9045 17085 9079 17119
rect 9137 17085 9171 17119
rect 9781 17085 9815 17119
rect 9873 17085 9907 17119
rect 10793 17085 10827 17119
rect 11437 17085 11471 17119
rect 13369 17085 13403 17119
rect 13737 17085 13771 17119
rect 14013 17085 14047 17119
rect 14289 17085 14323 17119
rect 14565 17085 14599 17119
rect 16497 17085 16531 17119
rect 2697 17017 2731 17051
rect 3249 17017 3283 17051
rect 5089 17017 5123 17051
rect 6193 17017 6227 17051
rect 6561 17017 6595 17051
rect 6745 17017 6779 17051
rect 12265 17017 12299 17051
rect 14832 17017 14866 17051
rect 1685 16949 1719 16983
rect 2329 16949 2363 16983
rect 2789 16949 2823 16983
rect 9321 16949 9355 16983
rect 9597 16949 9631 16983
rect 10057 16949 10091 16983
rect 10149 16949 10183 16983
rect 11069 16949 11103 16983
rect 11897 16949 11931 16983
rect 12357 16949 12391 16983
rect 14105 16949 14139 16983
rect 15945 16949 15979 16983
rect 2421 16745 2455 16779
rect 5273 16745 5307 16779
rect 6377 16745 6411 16779
rect 6561 16745 6595 16779
rect 7389 16745 7423 16779
rect 10425 16745 10459 16779
rect 1308 16677 1342 16711
rect 6745 16677 6779 16711
rect 7757 16677 7791 16711
rect 2881 16609 2915 16643
rect 3065 16609 3099 16643
rect 3413 16609 3447 16643
rect 4813 16609 4847 16643
rect 5089 16609 5123 16643
rect 5549 16609 5583 16643
rect 6009 16609 6043 16643
rect 9330 16609 9364 16643
rect 9597 16609 9631 16643
rect 9873 16609 9907 16643
rect 10333 16609 10367 16643
rect 11253 16609 11287 16643
rect 11529 16609 11563 16643
rect 11785 16609 11819 16643
rect 13277 16609 13311 16643
rect 13553 16609 13587 16643
rect 13829 16609 13863 16643
rect 14085 16609 14119 16643
rect 15485 16609 15519 16643
rect 15761 16609 15795 16643
rect 16497 16609 16531 16643
rect 17141 16609 17175 16643
rect 1041 16541 1075 16575
rect 3157 16541 3191 16575
rect 6101 16541 6135 16575
rect 7849 16541 7883 16575
rect 7941 16541 7975 16575
rect 10609 16541 10643 16575
rect 16589 16541 16623 16575
rect 16681 16541 16715 16575
rect 7113 16473 7147 16507
rect 9965 16473 9999 16507
rect 11437 16473 11471 16507
rect 12909 16473 12943 16507
rect 13737 16473 13771 16507
rect 16957 16473 16991 16507
rect 3065 16405 3099 16439
rect 4537 16405 4571 16439
rect 4629 16405 4663 16439
rect 5365 16405 5399 16439
rect 6745 16405 6779 16439
rect 8217 16405 8251 16439
rect 9689 16405 9723 16439
rect 13093 16405 13127 16439
rect 15209 16405 15243 16439
rect 15301 16405 15335 16439
rect 15577 16405 15611 16439
rect 16129 16405 16163 16439
rect 7021 16201 7055 16235
rect 7297 16201 7331 16235
rect 10701 16201 10735 16235
rect 13553 16201 13587 16235
rect 3065 16133 3099 16167
rect 7941 16133 7975 16167
rect 11161 16133 11195 16167
rect 12633 16133 12667 16167
rect 14381 16133 14415 16167
rect 4629 16065 4663 16099
rect 6469 16065 6503 16099
rect 9321 16065 9355 16099
rect 11253 16065 11287 16099
rect 11621 16065 11655 16099
rect 12265 16065 12299 16099
rect 14013 16065 14047 16099
rect 14197 16065 14231 16099
rect 15025 16065 15059 16099
rect 15669 16065 15703 16099
rect 1225 15997 1259 16031
rect 2881 15997 2915 16031
rect 4813 15997 4847 16031
rect 5080 15997 5114 16031
rect 6561 15997 6595 16031
rect 7481 15997 7515 16031
rect 7665 15997 7699 16031
rect 7757 15997 7791 16031
rect 7941 15997 7975 16031
rect 8033 15997 8067 16031
rect 8769 15997 8803 16031
rect 8953 15997 8987 16031
rect 9045 15997 9079 16031
rect 10977 15997 11011 16031
rect 12449 15997 12483 16031
rect 12725 15997 12759 16031
rect 13093 15997 13127 16031
rect 13277 15997 13311 16031
rect 13369 15997 13403 16031
rect 13921 15997 13955 16031
rect 1492 15929 1526 15963
rect 4384 15929 4418 15963
rect 6653 15929 6687 15963
rect 9588 15929 9622 15963
rect 11713 15929 11747 15963
rect 11805 15929 11839 15963
rect 14565 15929 14599 15963
rect 15209 15929 15243 15963
rect 15914 15929 15948 15963
rect 2605 15861 2639 15895
rect 3249 15861 3283 15895
rect 6193 15861 6227 15895
rect 8125 15861 8159 15895
rect 8585 15861 8619 15895
rect 10793 15861 10827 15895
rect 12173 15861 12207 15895
rect 12909 15861 12943 15895
rect 15117 15861 15151 15895
rect 15577 15861 15611 15895
rect 17049 15861 17083 15895
rect 1409 15657 1443 15691
rect 2053 15657 2087 15691
rect 2145 15657 2179 15691
rect 3341 15657 3375 15691
rect 6009 15657 6043 15691
rect 8033 15657 8067 15691
rect 9597 15657 9631 15691
rect 13277 15657 13311 15691
rect 15025 15657 15059 15691
rect 15669 15657 15703 15691
rect 2881 15589 2915 15623
rect 4629 15589 4663 15623
rect 7297 15589 7331 15623
rect 11805 15589 11839 15623
rect 1593 15521 1627 15555
rect 1961 15521 1995 15555
rect 2421 15521 2455 15555
rect 3157 15521 3191 15555
rect 3801 15521 3835 15555
rect 4077 15521 4111 15555
rect 4353 15521 4387 15555
rect 5089 15521 5123 15555
rect 5181 15521 5215 15555
rect 5457 15521 5491 15555
rect 5825 15521 5859 15555
rect 6101 15521 6135 15555
rect 6285 15521 6319 15555
rect 7113 15521 7147 15555
rect 7389 15521 7423 15555
rect 7573 15521 7607 15555
rect 7665 15521 7699 15555
rect 7757 15521 7791 15555
rect 9229 15521 9263 15555
rect 9413 15521 9447 15555
rect 9873 15521 9907 15555
rect 10149 15521 10183 15555
rect 11161 15521 11195 15555
rect 11713 15521 11747 15555
rect 11897 15521 11931 15555
rect 12817 15521 12851 15555
rect 12909 15521 12943 15555
rect 13553 15521 13587 15555
rect 13921 15521 13955 15555
rect 14197 15521 14231 15555
rect 14473 15521 14507 15555
rect 14841 15521 14875 15555
rect 15485 15521 15519 15555
rect 15945 15521 15979 15555
rect 16957 15521 16991 15555
rect 17233 15521 17267 15555
rect 1869 15453 1903 15487
rect 4997 15453 5031 15487
rect 5273 15453 5307 15487
rect 6837 15453 6871 15487
rect 9689 15453 9723 15487
rect 11345 15453 11379 15487
rect 11437 15453 11471 15487
rect 12541 15453 12575 15487
rect 13001 15453 13035 15487
rect 14749 15453 14783 15487
rect 1777 15385 1811 15419
rect 2513 15385 2547 15419
rect 3065 15385 3099 15419
rect 3617 15385 3651 15419
rect 10057 15385 10091 15419
rect 13369 15385 13403 15419
rect 14105 15385 14139 15419
rect 14657 15385 14691 15419
rect 17049 15385 17083 15419
rect 2881 15317 2915 15351
rect 3893 15317 3927 15351
rect 4169 15317 4203 15351
rect 4537 15317 4571 15351
rect 4813 15317 4847 15351
rect 5641 15317 5675 15351
rect 6193 15317 6227 15351
rect 6929 15317 6963 15351
rect 9045 15317 9079 15351
rect 10977 15317 11011 15351
rect 12909 15317 12943 15351
rect 13737 15317 13771 15351
rect 14289 15317 14323 15351
rect 15761 15317 15795 15351
rect 16865 15317 16899 15351
rect 2697 15113 2731 15147
rect 2881 15113 2915 15147
rect 7573 15113 7607 15147
rect 7849 15113 7883 15147
rect 8217 15113 8251 15147
rect 8585 15113 8619 15147
rect 8769 15113 8803 15147
rect 13737 15113 13771 15147
rect 14657 15113 14691 15147
rect 2237 15045 2271 15079
rect 3249 15045 3283 15079
rect 4169 15045 4203 15079
rect 14013 15045 14047 15079
rect 3525 14977 3559 15011
rect 4905 14977 4939 15011
rect 5114 14977 5148 15011
rect 5641 14977 5675 15011
rect 6193 14977 6227 15011
rect 15853 14977 15887 15011
rect 857 14909 891 14943
rect 3433 14909 3467 14943
rect 3617 14909 3651 14943
rect 3709 14909 3743 14943
rect 3893 14909 3927 14943
rect 4077 14909 4111 14943
rect 4261 14909 4295 14943
rect 4353 14909 4387 14943
rect 4629 14909 4663 14943
rect 6009 14909 6043 14943
rect 7021 14909 7055 14943
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 8401 14909 8435 14943
rect 8585 14909 8619 14943
rect 11345 14909 11379 14943
rect 12909 14909 12943 14943
rect 13185 14909 13219 14943
rect 13553 14909 13587 14943
rect 13829 14909 13863 14943
rect 14289 14909 14323 14943
rect 15485 14909 15519 14943
rect 1124 14841 1158 14875
rect 3065 14841 3099 14875
rect 5524 14841 5558 14875
rect 7297 14841 7331 14875
rect 12642 14841 12676 14875
rect 16098 14841 16132 14875
rect 2855 14773 2889 14807
rect 4997 14773 5031 14807
rect 5273 14773 5307 14807
rect 5365 14773 5399 14807
rect 5733 14773 5767 14807
rect 6837 14773 6871 14807
rect 7205 14773 7239 14807
rect 7389 14773 7423 14807
rect 11253 14773 11287 14807
rect 11529 14773 11563 14807
rect 13001 14773 13035 14807
rect 14657 14773 14691 14807
rect 14841 14773 14875 14807
rect 15669 14773 15703 14807
rect 17233 14773 17267 14807
rect 1875 14569 1909 14603
rect 2421 14569 2455 14603
rect 4261 14569 4295 14603
rect 7573 14569 7607 14603
rect 9137 14569 9171 14603
rect 12541 14569 12575 14603
rect 13835 14569 13869 14603
rect 1685 14501 1719 14535
rect 1777 14501 1811 14535
rect 1961 14501 1995 14535
rect 4537 14501 4571 14535
rect 4997 14501 5031 14535
rect 5365 14501 5399 14535
rect 6101 14501 6135 14535
rect 6561 14501 6595 14535
rect 7849 14501 7883 14535
rect 8125 14501 8159 14535
rect 8217 14501 8251 14535
rect 14534 14501 14568 14535
rect 1409 14433 1443 14467
rect 2053 14433 2087 14467
rect 2697 14433 2731 14467
rect 2789 14433 2823 14467
rect 3893 14433 3927 14467
rect 4629 14433 4663 14467
rect 6929 14433 6963 14467
rect 7021 14433 7055 14467
rect 7389 14433 7423 14467
rect 8585 14433 8619 14467
rect 8977 14433 9011 14467
rect 9505 14433 9539 14467
rect 10333 14433 10367 14467
rect 10609 14433 10643 14467
rect 10977 14433 11011 14467
rect 11897 14423 11931 14457
rect 12081 14433 12115 14467
rect 12817 14433 12851 14467
rect 13737 14433 13771 14467
rect 13921 14433 13955 14467
rect 14013 14433 14047 14467
rect 14289 14433 14323 14467
rect 15945 14433 15979 14467
rect 1685 14365 1719 14399
rect 2605 14365 2639 14399
rect 2881 14365 2915 14399
rect 3617 14365 3651 14399
rect 6009 14365 6043 14399
rect 10517 14365 10551 14399
rect 6561 14297 6595 14331
rect 9689 14297 9723 14331
rect 10149 14297 10183 14331
rect 12173 14297 12207 14331
rect 13001 14297 13035 14331
rect 15669 14297 15703 14331
rect 15761 14297 15795 14331
rect 1501 14229 1535 14263
rect 5549 14229 5583 14263
rect 5825 14229 5859 14263
rect 7389 14229 7423 14263
rect 10609 14229 10643 14263
rect 11161 14229 11195 14263
rect 11713 14229 11747 14263
rect 12541 14229 12575 14263
rect 12725 14229 12759 14263
rect 3801 14025 3835 14059
rect 4813 14025 4847 14059
rect 6653 14025 6687 14059
rect 7205 14025 7239 14059
rect 7389 14025 7423 14059
rect 11069 14025 11103 14059
rect 11989 14025 12023 14059
rect 13645 14025 13679 14059
rect 13921 14025 13955 14059
rect 2605 13957 2639 13991
rect 8401 13957 8435 13991
rect 10701 13957 10735 13991
rect 15761 13957 15795 13991
rect 16681 13957 16715 13991
rect 2973 13889 3007 13923
rect 4169 13889 4203 13923
rect 6193 13889 6227 13923
rect 11621 13889 11655 13923
rect 12909 13889 12943 13923
rect 13553 13889 13587 13923
rect 13737 13889 13771 13923
rect 16129 13889 16163 13923
rect 16405 13889 16439 13923
rect 2789 13821 2823 13855
rect 3249 13821 3283 13855
rect 3525 13821 3559 13855
rect 3709 13821 3743 13855
rect 3985 13821 4019 13855
rect 4077 13821 4111 13855
rect 4262 13821 4296 13855
rect 4445 13821 4479 13855
rect 4721 13821 4755 13855
rect 4997 13821 5031 13855
rect 5273 13821 5307 13855
rect 5549 13821 5583 13855
rect 5641 13821 5675 13855
rect 6285 13821 6319 13855
rect 6653 13821 6687 13855
rect 6929 13821 6963 13855
rect 7389 13821 7423 13855
rect 7757 13821 7791 13855
rect 7849 13821 7883 13855
rect 8585 13821 8619 13855
rect 8861 13821 8895 13855
rect 9781 13821 9815 13855
rect 11897 13821 11931 13855
rect 12173 13821 12207 13855
rect 12265 13821 12299 13855
rect 12541 13821 12575 13855
rect 12725 13821 12759 13855
rect 13185 13821 13219 13855
rect 13829 13821 13863 13855
rect 14381 13821 14415 13855
rect 14648 13821 14682 13855
rect 16037 13821 16071 13855
rect 16865 13821 16899 13855
rect 17141 13821 17175 13855
rect 3617 13753 3651 13787
rect 9689 13753 9723 13787
rect 10149 13753 10183 13787
rect 11053 13753 11087 13787
rect 11253 13753 11287 13787
rect 11437 13753 11471 13787
rect 14105 13753 14139 13787
rect 14289 13753 14323 13787
rect 3433 13685 3467 13719
rect 4629 13685 4663 13719
rect 6837 13685 6871 13719
rect 7113 13685 7147 13719
rect 9045 13685 9079 13719
rect 9413 13685 9447 13719
rect 10517 13685 10551 13719
rect 10885 13685 10919 13719
rect 11713 13685 11747 13719
rect 12449 13685 12483 13719
rect 13001 13685 13035 13719
rect 16957 13685 16991 13719
rect 3341 13481 3375 13515
rect 3617 13481 3651 13515
rect 3893 13481 3927 13515
rect 5825 13481 5859 13515
rect 7665 13481 7699 13515
rect 9505 13481 9539 13515
rect 9689 13481 9723 13515
rect 10701 13481 10735 13515
rect 12817 13481 12851 13515
rect 15761 13481 15795 13515
rect 16865 13481 16899 13515
rect 2865 13413 2899 13447
rect 3065 13413 3099 13447
rect 4261 13413 4295 13447
rect 6561 13413 6595 13447
rect 6837 13413 6871 13447
rect 7297 13413 7331 13447
rect 8217 13413 8251 13447
rect 9321 13413 9355 13447
rect 13369 13413 13403 13447
rect 13737 13413 13771 13447
rect 14473 13413 14507 13447
rect 1216 13345 1250 13379
rect 2605 13329 2639 13363
rect 3157 13345 3191 13379
rect 3433 13345 3467 13379
rect 4077 13345 4111 13379
rect 4537 13345 4571 13379
rect 5641 13345 5675 13379
rect 6009 13345 6043 13379
rect 6929 13345 6963 13379
rect 8493 13345 8527 13379
rect 8585 13345 8619 13379
rect 8953 13345 8987 13379
rect 9873 13345 9907 13379
rect 10149 13345 10183 13379
rect 10517 13345 10551 13379
rect 11161 13345 11195 13379
rect 11345 13345 11379 13379
rect 13645 13345 13679 13379
rect 14105 13345 14139 13379
rect 15945 13345 15979 13379
rect 16313 13345 16347 13379
rect 16773 13345 16807 13379
rect 17049 13345 17083 13379
rect 17325 13345 17359 13379
rect 949 13277 983 13311
rect 5365 13277 5399 13311
rect 10057 13277 10091 13311
rect 14841 13277 14875 13311
rect 15117 13277 15151 13311
rect 16497 13277 16531 13311
rect 10977 13209 11011 13243
rect 16589 13209 16623 13243
rect 2329 13141 2363 13175
rect 2421 13141 2455 13175
rect 2697 13141 2731 13175
rect 2881 13141 2915 13175
rect 4721 13141 4755 13175
rect 7849 13141 7883 13175
rect 10425 13141 10459 13175
rect 14657 13141 14691 13175
rect 16129 13141 16163 13175
rect 17141 13141 17175 13175
rect 1317 12937 1351 12971
rect 2881 12937 2915 12971
rect 6101 12937 6135 12971
rect 7113 12937 7147 12971
rect 11989 12937 12023 12971
rect 17233 12937 17267 12971
rect 4629 12869 4663 12903
rect 11897 12869 11931 12903
rect 1593 12801 1627 12835
rect 5181 12801 5215 12835
rect 6561 12801 6595 12835
rect 6653 12801 6687 12835
rect 12449 12801 12483 12835
rect 12817 12801 12851 12835
rect 12909 12801 12943 12835
rect 15117 12801 15151 12835
rect 1317 12733 1351 12767
rect 1501 12733 1535 12767
rect 1777 12733 1811 12767
rect 1869 12733 1903 12767
rect 2513 12733 2547 12767
rect 3249 12733 3283 12767
rect 5089 12733 5123 12767
rect 5457 12733 5491 12767
rect 6469 12733 6503 12767
rect 6929 12733 6963 12767
rect 9689 12733 9723 12767
rect 10701 12733 10735 12767
rect 11093 12733 11127 12767
rect 11713 12733 11747 12767
rect 12173 12709 12207 12743
rect 12633 12733 12667 12767
rect 12725 12733 12759 12767
rect 13737 12733 13771 12767
rect 13829 12733 13863 12767
rect 14105 12733 14139 12767
rect 14841 12733 14875 12767
rect 15853 12733 15887 12767
rect 16120 12733 16154 12767
rect 1593 12665 1627 12699
rect 3516 12665 3550 12699
rect 8585 12665 8619 12699
rect 9965 12665 9999 12699
rect 10241 12665 10275 12699
rect 10333 12665 10367 12699
rect 2881 12597 2915 12631
rect 3065 12597 3099 12631
rect 4905 12597 4939 12631
rect 8493 12597 8527 12631
rect 9505 12597 9539 12631
rect 11253 12597 11287 12631
rect 13553 12597 13587 12631
rect 3157 12393 3191 12427
rect 3617 12393 3651 12427
rect 4491 12393 4525 12427
rect 7941 12393 7975 12427
rect 8401 12393 8435 12427
rect 13829 12393 13863 12427
rect 7573 12325 7607 12359
rect 7711 12325 7745 12359
rect 14013 12325 14047 12359
rect 14810 12325 14844 12359
rect 1124 12257 1158 12291
rect 2973 12257 3007 12291
rect 3525 12257 3559 12291
rect 3801 12257 3835 12291
rect 4813 12257 4847 12291
rect 6009 12257 6043 12291
rect 6193 12257 6227 12291
rect 6285 12257 6319 12291
rect 7205 12257 7239 12291
rect 7389 12257 7423 12291
rect 7481 12257 7515 12291
rect 8125 12257 8159 12291
rect 8585 12257 8619 12291
rect 11437 12257 11471 12291
rect 11704 12257 11738 12291
rect 13737 12257 13771 12291
rect 13921 12257 13955 12291
rect 16681 12257 16715 12291
rect 17141 12257 17175 12291
rect 17233 12257 17267 12291
rect 857 12189 891 12223
rect 4721 12189 4755 12223
rect 5089 12189 5123 12223
rect 6561 12189 6595 12223
rect 7849 12189 7883 12223
rect 8309 12189 8343 12223
rect 14473 12189 14507 12223
rect 14565 12189 14599 12223
rect 16773 12189 16807 12223
rect 5825 12121 5859 12155
rect 14289 12121 14323 12155
rect 2237 12053 2271 12087
rect 3433 12053 3467 12087
rect 12817 12053 12851 12087
rect 15945 12053 15979 12087
rect 16313 12053 16347 12087
rect 16957 12053 16991 12087
rect 1409 11849 1443 11883
rect 1777 11849 1811 11883
rect 1961 11849 1995 11883
rect 3985 11849 4019 11883
rect 8033 11849 8067 11883
rect 8585 11849 8619 11883
rect 9045 11849 9079 11883
rect 9413 11849 9447 11883
rect 11897 11849 11931 11883
rect 13001 11849 13035 11883
rect 13921 11849 13955 11883
rect 14105 11849 14139 11883
rect 14381 11849 14415 11883
rect 16681 11849 16715 11883
rect 9137 11781 9171 11815
rect 12173 11781 12207 11815
rect 13553 11781 13587 11815
rect 2237 11713 2271 11747
rect 4629 11713 4663 11747
rect 8953 11713 8987 11747
rect 11989 11713 12023 11747
rect 1409 11645 1443 11679
rect 1593 11645 1627 11679
rect 2421 11645 2455 11679
rect 2513 11645 2547 11679
rect 3893 11645 3927 11679
rect 4169 11645 4203 11679
rect 4353 11645 4387 11679
rect 4537 11645 4571 11679
rect 7389 11645 7423 11679
rect 7573 11645 7607 11679
rect 7665 11645 7699 11679
rect 7757 11645 7791 11679
rect 7849 11645 7883 11679
rect 8769 11645 8803 11679
rect 9045 11645 9079 11679
rect 9321 11645 9355 11679
rect 9413 11645 9447 11679
rect 9873 11645 9907 11679
rect 10057 11645 10091 11679
rect 10149 11645 10183 11679
rect 11253 11645 11287 11679
rect 11621 11645 11655 11679
rect 11713 11645 11747 11679
rect 11897 11645 11931 11679
rect 12265 11645 12299 11679
rect 12725 11645 12759 11679
rect 14657 11645 14691 11679
rect 14841 11645 14875 11679
rect 15301 11645 15335 11679
rect 2145 11577 2179 11611
rect 4261 11577 4295 11611
rect 6377 11577 6411 11611
rect 9597 11577 9631 11611
rect 10517 11577 10551 11611
rect 11989 11577 12023 11611
rect 13185 11577 13219 11611
rect 13921 11577 13955 11611
rect 14565 11577 14599 11611
rect 15568 11577 15602 11611
rect 1945 11509 1979 11543
rect 2237 11509 2271 11543
rect 3709 11509 3743 11543
rect 9689 11509 9723 11543
rect 11437 11509 11471 11543
rect 12541 11509 12575 11543
rect 12817 11509 12851 11543
rect 12985 11509 13019 11543
rect 14197 11509 14231 11543
rect 14360 11509 14394 11543
rect 15025 11509 15059 11543
rect 1685 11305 1719 11339
rect 4261 11305 4295 11339
rect 4629 11305 4663 11339
rect 7757 11305 7791 11339
rect 8033 11305 8067 11339
rect 8677 11305 8711 11339
rect 9229 11305 9263 11339
rect 15669 11305 15703 11339
rect 16129 11305 16163 11339
rect 2872 11237 2906 11271
rect 12449 11237 12483 11271
rect 1869 11169 1903 11203
rect 2053 11169 2087 11203
rect 2145 11169 2179 11203
rect 2605 11169 2639 11203
rect 4353 11169 4387 11203
rect 4445 11169 4479 11203
rect 4997 11169 5031 11203
rect 5181 11169 5215 11203
rect 5273 11169 5307 11203
rect 5825 11169 5859 11203
rect 6745 11169 6779 11203
rect 7021 11169 7055 11203
rect 7389 11169 7423 11203
rect 7481 11169 7515 11203
rect 7849 11169 7883 11203
rect 8033 11169 8067 11203
rect 8861 11169 8895 11203
rect 9137 11169 9171 11203
rect 9597 11169 9631 11203
rect 10609 11169 10643 11203
rect 10793 11169 10827 11203
rect 11621 11169 11655 11203
rect 14197 11169 14231 11203
rect 15577 11169 15611 11203
rect 15945 11169 15979 11203
rect 16313 11169 16347 11203
rect 16497 11169 16531 11203
rect 16589 11169 16623 11203
rect 16773 11169 16807 11203
rect 2421 11101 2455 11135
rect 9045 11101 9079 11135
rect 9505 11101 9539 11135
rect 10425 11101 10459 11135
rect 11437 11101 11471 11135
rect 12265 11101 12299 11135
rect 15669 11101 15703 11135
rect 2237 11033 2271 11067
rect 3985 11033 4019 11067
rect 4077 11033 4111 11067
rect 6837 11033 6871 11067
rect 7205 11033 7239 11067
rect 7297 11033 7331 11067
rect 16957 11033 16991 11067
rect 2329 10965 2363 10999
rect 4721 10965 4755 10999
rect 4997 10965 5031 10999
rect 5457 10965 5491 10999
rect 6009 10965 6043 10999
rect 8861 10965 8895 10999
rect 9597 10965 9631 10999
rect 15347 10965 15381 10999
rect 15853 10965 15887 10999
rect 4537 10761 4571 10795
rect 5089 10761 5123 10795
rect 7021 10761 7055 10795
rect 7849 10761 7883 10795
rect 13553 10761 13587 10795
rect 14749 10761 14783 10795
rect 14933 10761 14967 10795
rect 5457 10693 5491 10727
rect 14381 10693 14415 10727
rect 4077 10625 4111 10659
rect 4905 10625 4939 10659
rect 6009 10625 6043 10659
rect 6745 10625 6779 10659
rect 13001 10625 13035 10659
rect 16405 10625 16439 10659
rect 1501 10557 1535 10591
rect 1685 10557 1719 10591
rect 4353 10557 4387 10591
rect 4721 10557 4755 10591
rect 5641 10557 5675 10591
rect 6101 10557 6135 10591
rect 6285 10557 6319 10591
rect 7205 10557 7239 10591
rect 7573 10557 7607 10591
rect 7665 10557 7699 10591
rect 10241 10557 10275 10591
rect 12817 10557 12851 10591
rect 13093 10557 13127 10591
rect 13277 10557 13311 10591
rect 13737 10557 13771 10591
rect 13921 10557 13955 10591
rect 15393 10557 15427 10591
rect 15669 10557 15703 10591
rect 16497 10557 16531 10591
rect 5181 10489 5215 10523
rect 5825 10489 5859 10523
rect 6377 10489 6411 10523
rect 6469 10489 6503 10523
rect 6607 10489 6641 10523
rect 7297 10489 7331 10523
rect 7389 10489 7423 10523
rect 8677 10489 8711 10523
rect 13185 10489 13219 10523
rect 14749 10489 14783 10523
rect 15025 10489 15059 10523
rect 15209 10489 15243 10523
rect 1593 10421 1627 10455
rect 5733 10421 5767 10455
rect 12633 10421 12667 10455
rect 15485 10421 15519 10455
rect 16865 10421 16899 10455
rect 3801 10217 3835 10251
rect 4169 10217 4203 10251
rect 4353 10217 4387 10251
rect 4905 10217 4939 10251
rect 5457 10217 5491 10251
rect 6025 10217 6059 10251
rect 6929 10217 6963 10251
rect 7941 10217 7975 10251
rect 9321 10217 9355 10251
rect 10241 10217 10275 10251
rect 12357 10217 12391 10251
rect 12725 10217 12759 10251
rect 13645 10217 13679 10251
rect 14381 10217 14415 10251
rect 16681 10217 16715 10251
rect 2596 10149 2630 10183
rect 5825 10149 5859 10183
rect 7113 10149 7147 10183
rect 10609 10149 10643 10183
rect 11222 10149 11256 10183
rect 16865 10149 16899 10183
rect 1124 10081 1158 10115
rect 2329 10081 2363 10115
rect 3985 10081 4019 10115
rect 4077 10081 4111 10115
rect 4537 10081 4571 10115
rect 5089 10081 5123 10115
rect 5273 10081 5307 10115
rect 5365 10081 5399 10115
rect 6469 10081 6503 10115
rect 7297 10081 7331 10115
rect 7389 10081 7423 10115
rect 7573 10081 7607 10115
rect 8217 10081 8251 10115
rect 8355 10081 8389 10115
rect 8953 10081 8987 10115
rect 9229 10081 9263 10115
rect 9505 10081 9539 10115
rect 9689 10081 9723 10115
rect 9781 10081 9815 10115
rect 10057 10081 10091 10115
rect 10333 10081 10367 10115
rect 10517 10081 10551 10115
rect 10701 10081 10735 10115
rect 10977 10081 11011 10115
rect 12633 10081 12667 10115
rect 12909 10081 12943 10115
rect 13461 10081 13495 10115
rect 14197 10081 14231 10115
rect 15393 10081 15427 10115
rect 15669 10081 15703 10115
rect 15853 10081 15887 10115
rect 15945 10081 15979 10115
rect 16313 10081 16347 10115
rect 16773 10081 16807 10115
rect 16957 10081 16991 10115
rect 17049 10081 17083 10115
rect 857 10013 891 10047
rect 4445 10013 4479 10047
rect 4629 10013 4663 10047
rect 5641 10013 5675 10047
rect 6561 10013 6595 10047
rect 7481 10013 7515 10047
rect 8125 10013 8159 10047
rect 8493 10013 8527 10047
rect 8585 10013 8619 10047
rect 9137 10013 9171 10047
rect 14013 10013 14047 10047
rect 16221 10013 16255 10047
rect 3709 9945 3743 9979
rect 6193 9945 6227 9979
rect 15301 9945 15335 9979
rect 2237 9877 2271 9911
rect 4537 9877 4571 9911
rect 6009 9877 6043 9911
rect 6745 9877 6779 9911
rect 8769 9877 8803 9911
rect 8953 9877 8987 9911
rect 10057 9877 10091 9911
rect 12449 9877 12483 9911
rect 15485 9877 15519 9911
rect 17141 9877 17175 9911
rect 4261 9673 4295 9707
rect 11897 9673 11931 9707
rect 12449 9673 12483 9707
rect 13185 9673 13219 9707
rect 2513 9605 2547 9639
rect 3985 9605 4019 9639
rect 10425 9605 10459 9639
rect 16221 9605 16255 9639
rect 2697 9537 2731 9571
rect 6929 9537 6963 9571
rect 16773 9537 16807 9571
rect 857 9469 891 9503
rect 2329 9469 2363 9503
rect 2605 9469 2639 9503
rect 3801 9469 3835 9503
rect 4077 9469 4111 9503
rect 4261 9469 4295 9503
rect 6193 9469 6227 9503
rect 6469 9469 6503 9503
rect 6653 9469 6687 9503
rect 9137 9469 9171 9503
rect 9781 9469 9815 9503
rect 10057 9469 10091 9503
rect 10149 9469 10183 9503
rect 10241 9469 10275 9503
rect 10517 9469 10551 9503
rect 12265 9469 12299 9503
rect 12357 9469 12391 9503
rect 12633 9445 12667 9479
rect 13369 9469 13403 9503
rect 13553 9469 13587 9503
rect 14105 9469 14139 9503
rect 14289 9469 14323 9503
rect 14381 9469 14415 9503
rect 14473 9469 14507 9503
rect 14841 9469 14875 9503
rect 16497 9469 16531 9503
rect 1124 9401 1158 9435
rect 6561 9401 6595 9435
rect 6771 9401 6805 9435
rect 9939 9401 9973 9435
rect 10773 9401 10807 9435
rect 12541 9401 12575 9435
rect 13737 9401 13771 9435
rect 14749 9401 14783 9435
rect 15086 9401 15120 9435
rect 2237 9333 2271 9367
rect 4905 9333 4939 9367
rect 6285 9333 6319 9367
rect 9321 9333 9355 9367
rect 12081 9333 12115 9367
rect 12817 9333 12851 9367
rect 13921 9333 13955 9367
rect 3157 9129 3191 9163
rect 6193 9129 6227 9163
rect 7481 9129 7515 9163
rect 10701 9129 10735 9163
rect 15117 9129 15151 9163
rect 15853 9129 15887 9163
rect 7021 9061 7055 9095
rect 8953 9061 8987 9095
rect 10977 9061 11011 9095
rect 11172 9061 11206 9095
rect 11345 9061 11379 9095
rect 11589 9061 11623 9095
rect 11805 9061 11839 9095
rect 1777 8993 1811 9027
rect 2044 8993 2078 9027
rect 4373 8993 4407 9027
rect 4629 8993 4663 9027
rect 5917 8993 5951 9027
rect 6101 8993 6135 9027
rect 6377 8993 6411 9027
rect 6561 8993 6595 9027
rect 6837 8993 6871 9027
rect 6929 8993 6963 9027
rect 7139 8993 7173 9027
rect 7389 8993 7423 9027
rect 8033 8993 8067 9027
rect 9229 8993 9263 9027
rect 9321 8993 9355 9027
rect 9413 8993 9447 9027
rect 9597 8993 9631 9027
rect 10169 8993 10203 9027
rect 10333 8993 10367 9027
rect 10425 8993 10459 9027
rect 10517 8993 10551 9027
rect 12357 8993 12391 9027
rect 12541 8993 12575 9027
rect 12909 8993 12943 9027
rect 13829 8993 13863 9027
rect 14105 8993 14139 9027
rect 14749 8993 14783 9027
rect 15201 8993 15235 9027
rect 15945 8993 15979 9027
rect 17049 8993 17083 9027
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 7297 8925 7331 8959
rect 8309 8925 8343 8959
rect 13185 8925 13219 8959
rect 16681 8925 16715 8959
rect 16957 8925 16991 8959
rect 3249 8857 3283 8891
rect 12541 8857 12575 8891
rect 14933 8857 14967 8891
rect 6101 8789 6135 8823
rect 6653 8789 6687 8823
rect 11437 8789 11471 8823
rect 11621 8789 11655 8823
rect 17233 8789 17267 8823
rect 857 8585 891 8619
rect 5549 8585 5583 8619
rect 5733 8585 5767 8619
rect 6285 8585 6319 8619
rect 7665 8585 7699 8619
rect 9505 8585 9539 8619
rect 9781 8585 9815 8619
rect 17325 8585 17359 8619
rect 6653 8517 6687 8551
rect 7113 8517 7147 8551
rect 5089 8449 5123 8483
rect 5825 8449 5859 8483
rect 6469 8449 6503 8483
rect 6929 8449 6963 8483
rect 7389 8449 7423 8483
rect 8493 8449 8527 8483
rect 13829 8449 13863 8483
rect 15945 8449 15979 8483
rect 2237 8381 2271 8415
rect 4813 8381 4847 8415
rect 5181 8381 5215 8415
rect 5549 8381 5583 8415
rect 6009 8381 6043 8415
rect 6101 8381 6135 8415
rect 6377 8381 6411 8415
rect 7021 8381 7055 8415
rect 7297 8381 7331 8415
rect 7481 8381 7515 8415
rect 7849 8381 7883 8415
rect 8125 8381 8159 8415
rect 8769 8381 8803 8415
rect 9413 8381 9447 8415
rect 9597 8381 9631 8415
rect 9965 8381 9999 8415
rect 10057 8381 10091 8415
rect 10425 8381 10459 8415
rect 11713 8381 11747 8415
rect 13553 8381 13587 8415
rect 13737 8381 13771 8415
rect 13921 8381 13955 8415
rect 14105 8381 14139 8415
rect 1992 8313 2026 8347
rect 3801 8313 3835 8347
rect 8033 8313 8067 8347
rect 11253 8313 11287 8347
rect 11437 8313 11471 8347
rect 16212 8313 16246 8347
rect 10149 8245 10183 8279
rect 10333 8245 10367 8279
rect 11069 8245 11103 8279
rect 11529 8245 11563 8279
rect 14289 8245 14323 8279
rect 3249 8041 3283 8075
rect 6127 8041 6161 8075
rect 6745 8041 6779 8075
rect 15301 8041 15335 8075
rect 16329 8041 16363 8075
rect 16589 8041 16623 8075
rect 4629 7973 4663 8007
rect 5917 7973 5951 8007
rect 6377 7973 6411 8007
rect 6593 7973 6627 8007
rect 15485 7973 15519 8007
rect 16129 7973 16163 8007
rect 1593 7905 1627 7939
rect 2145 7905 2179 7939
rect 2789 7905 2823 7939
rect 2973 7905 3007 7939
rect 3065 7905 3099 7939
rect 4077 7905 4111 7939
rect 4353 7905 4387 7939
rect 5089 7905 5123 7939
rect 5365 7905 5399 7939
rect 10333 7905 10367 7939
rect 10517 7905 10551 7939
rect 10793 7905 10827 7939
rect 11161 7905 11195 7939
rect 11437 7905 11471 7939
rect 11713 7905 11747 7939
rect 11897 7905 11931 7939
rect 12173 7905 12207 7939
rect 12265 7905 12299 7939
rect 12449 7905 12483 7939
rect 12541 7905 12575 7939
rect 13461 7905 13495 7939
rect 13649 7905 13683 7939
rect 13829 7905 13863 7939
rect 14013 7905 14047 7939
rect 14289 7905 14323 7939
rect 14473 7905 14507 7939
rect 14565 7905 14599 7939
rect 14657 7905 14691 7939
rect 14841 7905 14875 7939
rect 15209 7905 15243 7939
rect 15393 7905 15427 7939
rect 15669 7905 15703 7939
rect 16773 7905 16807 7939
rect 1869 7837 1903 7871
rect 2053 7837 2087 7871
rect 4997 7837 5031 7871
rect 8125 7837 8159 7871
rect 8401 7837 8435 7871
rect 12081 7837 12115 7871
rect 13737 7837 13771 7871
rect 1685 7769 1719 7803
rect 2513 7769 2547 7803
rect 4537 7769 4571 7803
rect 5549 7769 5583 7803
rect 6285 7769 6319 7803
rect 10609 7769 10643 7803
rect 12725 7769 12759 7803
rect 16497 7769 16531 7803
rect 1777 7701 1811 7735
rect 2605 7701 2639 7735
rect 4261 7701 4295 7735
rect 5089 7701 5123 7735
rect 5273 7701 5307 7735
rect 6101 7701 6135 7735
rect 6561 7701 6595 7735
rect 10425 7701 10459 7735
rect 11253 7701 11287 7735
rect 11621 7701 11655 7735
rect 14197 7701 14231 7735
rect 15025 7701 15059 7735
rect 15853 7701 15887 7735
rect 16313 7701 16347 7735
rect 2053 7497 2087 7531
rect 4353 7497 4387 7531
rect 4629 7497 4663 7531
rect 5181 7497 5215 7531
rect 5549 7497 5583 7531
rect 6101 7497 6135 7531
rect 10149 7497 10183 7531
rect 10701 7497 10735 7531
rect 12081 7497 12115 7531
rect 12357 7497 12391 7531
rect 2329 7429 2363 7463
rect 4169 7429 4203 7463
rect 14013 7429 14047 7463
rect 14565 7429 14599 7463
rect 15393 7429 15427 7463
rect 3709 7361 3743 7395
rect 4445 7361 4479 7395
rect 11253 7361 11287 7395
rect 11345 7361 11379 7395
rect 11529 7361 11563 7395
rect 13921 7361 13955 7395
rect 14473 7361 14507 7395
rect 1961 7293 1995 7327
rect 2145 7293 2179 7327
rect 2237 7293 2271 7327
rect 2421 7293 2455 7327
rect 2513 7293 2547 7327
rect 2697 7293 2731 7327
rect 2881 7293 2915 7327
rect 3801 7293 3835 7327
rect 3985 7293 4019 7327
rect 4537 7293 4571 7327
rect 4629 7293 4663 7327
rect 4813 7293 4847 7327
rect 4997 7293 5031 7327
rect 5365 7293 5399 7327
rect 5641 7293 5675 7327
rect 5917 7293 5951 7327
rect 6377 7293 6411 7327
rect 8585 7293 8619 7327
rect 8769 7293 8803 7327
rect 8861 7293 8895 7327
rect 8953 7293 8987 7327
rect 9137 7293 9171 7327
rect 9229 7293 9263 7327
rect 9321 7293 9355 7327
rect 9505 7293 9539 7327
rect 9965 7293 9999 7327
rect 10241 7293 10275 7327
rect 10425 7293 10459 7327
rect 10517 7293 10551 7327
rect 11437 7293 11471 7327
rect 12265 7293 12299 7327
rect 12541 7293 12575 7327
rect 14197 7293 14231 7327
rect 14749 7293 14783 7327
rect 15209 7293 15243 7327
rect 15485 7293 15519 7327
rect 16681 7293 16715 7327
rect 16865 7293 16899 7327
rect 4261 7225 4295 7259
rect 16773 7225 16807 7259
rect 5825 7157 5859 7191
rect 6561 7157 6595 7191
rect 8401 7157 8435 7191
rect 9689 7157 9723 7191
rect 10333 7157 10367 7191
rect 11069 7157 11103 7191
rect 14381 7157 14415 7191
rect 14933 7157 14967 7191
rect 15025 7157 15059 7191
rect 16589 6885 16623 6919
rect 1124 6817 1158 6851
rect 2697 6817 2731 6851
rect 3617 6817 3651 6851
rect 3801 6817 3835 6851
rect 3985 6817 4019 6851
rect 4261 6817 4295 6851
rect 4353 6817 4387 6851
rect 4721 6817 4755 6851
rect 4905 6817 4939 6851
rect 7297 6817 7331 6851
rect 7849 6817 7883 6851
rect 8033 6817 8067 6851
rect 8401 6817 8435 6851
rect 9781 6817 9815 6851
rect 10609 6817 10643 6851
rect 10977 6817 11011 6851
rect 11161 6817 11195 6851
rect 11299 6817 11333 6851
rect 11529 6817 11563 6851
rect 11713 6817 11747 6851
rect 13829 6817 13863 6851
rect 16405 6817 16439 6851
rect 857 6749 891 6783
rect 7021 6749 7055 6783
rect 7113 6749 7147 6783
rect 7205 6749 7239 6783
rect 8125 6749 8159 6783
rect 8217 6749 8251 6783
rect 8585 6749 8619 6783
rect 9413 6749 9447 6783
rect 9689 6749 9723 6783
rect 10241 6749 10275 6783
rect 10425 6749 10459 6783
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 11437 6749 11471 6783
rect 16221 6749 16255 6783
rect 2237 6681 2271 6715
rect 3985 6681 4019 6715
rect 4629 6681 4663 6715
rect 14013 6681 14047 6715
rect 2881 6613 2915 6647
rect 4261 6613 4295 6647
rect 4721 6613 4755 6647
rect 7481 6613 7515 6647
rect 9965 6613 9999 6647
rect 8401 6409 8435 6443
rect 8769 6409 8803 6443
rect 9137 6409 9171 6443
rect 11069 6409 11103 6443
rect 11437 6409 11471 6443
rect 14473 6409 14507 6443
rect 5825 6341 5859 6375
rect 7849 6341 7883 6375
rect 16405 6341 16439 6375
rect 6101 6273 6135 6307
rect 7481 6273 7515 6307
rect 8861 6273 8895 6307
rect 11529 6273 11563 6307
rect 13829 6273 13863 6307
rect 14289 6273 14323 6307
rect 15117 6273 15151 6307
rect 16681 6273 16715 6307
rect 2789 6205 2823 6239
rect 6009 6205 6043 6239
rect 7205 6205 7239 6239
rect 7389 6205 7423 6239
rect 7573 6205 7607 6239
rect 7757 6205 7791 6239
rect 8033 6205 8067 6239
rect 8585 6205 8619 6239
rect 8953 6205 8987 6239
rect 11253 6205 11287 6239
rect 11897 6205 11931 6239
rect 12817 6205 12851 6239
rect 13553 6205 13587 6239
rect 13737 6205 13771 6239
rect 13921 6205 13955 6239
rect 14105 6205 14139 6239
rect 14381 6205 14415 6239
rect 14657 6205 14691 6239
rect 15393 6205 15427 6239
rect 16037 6205 16071 6239
rect 16221 6205 16255 6239
rect 16313 6205 16347 6239
rect 16497 6205 16531 6239
rect 16589 6205 16623 6239
rect 17049 6205 17083 6239
rect 7021 6137 7055 6171
rect 2605 6069 2639 6103
rect 6331 6069 6365 6103
rect 12081 6069 12115 6103
rect 12633 6069 12667 6103
rect 14841 6069 14875 6103
rect 16129 6069 16163 6103
rect 16865 6069 16899 6103
rect 2605 5865 2639 5899
rect 2881 5865 2915 5899
rect 4307 5865 4341 5899
rect 3709 5797 3743 5831
rect 9873 5797 9907 5831
rect 1124 5729 1158 5763
rect 2513 5729 2547 5763
rect 2697 5729 2731 5763
rect 2789 5729 2823 5763
rect 3065 5729 3099 5763
rect 3433 5729 3467 5763
rect 3617 5729 3651 5763
rect 3985 5729 4019 5763
rect 6009 5729 6043 5763
rect 6285 5729 6319 5763
rect 6377 5729 6411 5763
rect 6561 5729 6595 5763
rect 7113 5729 7147 5763
rect 9413 5729 9447 5763
rect 10057 5729 10091 5763
rect 10333 5729 10367 5763
rect 11989 5729 12023 5763
rect 12173 5729 12207 5763
rect 12265 5729 12299 5763
rect 12357 5729 12391 5763
rect 12909 5729 12943 5763
rect 13001 5729 13035 5763
rect 13277 5729 13311 5763
rect 13553 5729 13587 5763
rect 13645 5729 13679 5763
rect 13921 5729 13955 5763
rect 14841 5729 14875 5763
rect 15117 5729 15151 5763
rect 15393 5729 15427 5763
rect 15577 5729 15611 5763
rect 15761 5729 15795 5763
rect 15945 5729 15979 5763
rect 16313 5729 16347 5763
rect 16497 5729 16531 5763
rect 16681 5729 16715 5763
rect 16957 5729 16991 5763
rect 17141 5729 17175 5763
rect 857 5661 891 5695
rect 3709 5661 3743 5695
rect 3893 5661 3927 5695
rect 4077 5661 4111 5695
rect 6193 5661 6227 5695
rect 7389 5661 7423 5695
rect 9137 5661 9171 5695
rect 12725 5661 12759 5695
rect 15669 5661 15703 5695
rect 3065 5593 3099 5627
rect 9597 5593 9631 5627
rect 14657 5593 14691 5627
rect 16221 5593 16255 5627
rect 16773 5593 16807 5627
rect 2237 5525 2271 5559
rect 3249 5525 3283 5559
rect 5825 5525 5859 5559
rect 6929 5525 6963 5559
rect 7297 5525 7331 5559
rect 9229 5525 9263 5559
rect 9689 5525 9723 5559
rect 10149 5525 10183 5559
rect 12633 5525 12667 5559
rect 13185 5525 13219 5559
rect 13369 5525 13403 5559
rect 13829 5525 13863 5559
rect 14933 5525 14967 5559
rect 15209 5525 15243 5559
rect 16957 5525 16991 5559
rect 949 5321 983 5355
rect 2053 5321 2087 5355
rect 2881 5321 2915 5355
rect 3433 5321 3467 5355
rect 5641 5321 5675 5355
rect 7573 5321 7607 5355
rect 13645 5321 13679 5355
rect 2421 5253 2455 5287
rect 4261 5253 4295 5287
rect 8861 5253 8895 5287
rect 9413 5253 9447 5287
rect 11345 5253 11379 5287
rect 3801 5185 3835 5219
rect 5181 5185 5215 5219
rect 5273 5185 5307 5219
rect 6193 5185 6227 5219
rect 6469 5185 6503 5219
rect 10609 5185 10643 5219
rect 11437 5185 11471 5219
rect 12173 5185 12207 5219
rect 14105 5185 14139 5219
rect 857 5117 891 5151
rect 1041 5117 1075 5151
rect 1317 5117 1351 5151
rect 1409 5117 1443 5151
rect 2329 5117 2363 5151
rect 2605 5117 2639 5151
rect 3617 5117 3651 5151
rect 3709 5117 3743 5151
rect 3893 5117 3927 5151
rect 4077 5117 4111 5151
rect 4905 5117 4939 5151
rect 5089 5117 5123 5151
rect 5457 5117 5491 5151
rect 7297 5117 7331 5151
rect 7389 5117 7423 5151
rect 7665 5117 7699 5151
rect 8401 5117 8435 5151
rect 8585 5117 8619 5151
rect 8677 5117 8711 5151
rect 8953 5117 8987 5151
rect 9045 5117 9079 5151
rect 9321 5117 9355 5151
rect 9597 5117 9631 5151
rect 9689 5117 9723 5151
rect 10333 5117 10367 5151
rect 10517 5117 10551 5151
rect 10701 5117 10735 5151
rect 10885 5117 10919 5151
rect 10977 5117 11011 5151
rect 11161 5117 11195 5151
rect 11897 5117 11931 5151
rect 12081 5117 12115 5151
rect 12265 5117 12299 5151
rect 12449 5117 12483 5151
rect 12909 5117 12943 5151
rect 13553 5117 13587 5151
rect 13829 5117 13863 5151
rect 13921 5117 13955 5151
rect 1593 5049 1627 5083
rect 1777 5049 1811 5083
rect 2021 5049 2055 5083
rect 2237 5049 2271 5083
rect 2513 5049 2547 5083
rect 2849 5049 2883 5083
rect 3065 5049 3099 5083
rect 12633 5049 12667 5083
rect 1225 4981 1259 5015
rect 1869 4981 1903 5015
rect 2697 4981 2731 5015
rect 7113 4981 7147 5015
rect 9229 4981 9263 5015
rect 9873 4981 9907 5015
rect 10149 4981 10183 5015
rect 12725 4981 12759 5015
rect 1685 4777 1719 4811
rect 3065 4777 3099 4811
rect 11345 4777 11379 4811
rect 11989 4777 12023 4811
rect 11621 4709 11655 4743
rect 11805 4709 11839 4743
rect 14657 4709 14691 4743
rect 1409 4641 1443 4675
rect 1777 4641 1811 4675
rect 3341 4641 3375 4675
rect 3433 4641 3467 4675
rect 4905 4641 4939 4675
rect 5089 4641 5123 4675
rect 5181 4641 5215 4675
rect 5273 4641 5307 4675
rect 5457 4641 5491 4675
rect 5825 4651 5859 4685
rect 6009 4641 6043 4675
rect 6193 4641 6227 4675
rect 6377 4641 6411 4675
rect 6929 4641 6963 4675
rect 7205 4641 7239 4675
rect 7665 4641 7699 4675
rect 8033 4641 8067 4675
rect 8229 4641 8263 4675
rect 9597 4641 9631 4675
rect 9873 4641 9907 4675
rect 9977 4641 10011 4675
rect 10149 4641 10183 4675
rect 11529 4641 11563 4675
rect 12357 4641 12391 4675
rect 13737 4641 13771 4675
rect 14841 4641 14875 4675
rect 14933 4641 14967 4675
rect 15117 4641 15151 4675
rect 16589 4641 16623 4675
rect 3065 4573 3099 4607
rect 3249 4573 3283 4607
rect 6101 4573 6135 4607
rect 7021 4573 7055 4607
rect 7389 4573 7423 4607
rect 7849 4573 7883 4607
rect 7941 4573 7975 4607
rect 9413 4573 9447 4607
rect 9781 4573 9815 4607
rect 12081 4573 12115 4607
rect 13829 4573 13863 4607
rect 13921 4573 13955 4607
rect 14013 4573 14047 4607
rect 16681 4573 16715 4607
rect 1225 4437 1259 4471
rect 3617 4437 3651 4471
rect 5641 4437 5675 4471
rect 6561 4437 6595 4471
rect 7481 4437 7515 4471
rect 14197 4437 14231 4471
rect 14473 4437 14507 4471
rect 15025 4437 15059 4471
rect 16221 4437 16255 4471
rect 4629 4233 4663 4267
rect 6193 4233 6227 4267
rect 11437 4233 11471 4267
rect 13553 4233 13587 4267
rect 7573 4165 7607 4199
rect 16129 4165 16163 4199
rect 3249 4097 3283 4131
rect 7665 4097 7699 4131
rect 11345 4097 11379 4131
rect 12633 4097 12667 4131
rect 12909 4097 12943 4131
rect 14473 4097 14507 4131
rect 14657 4097 14691 4131
rect 14749 4097 14783 4131
rect 16221 4097 16255 4131
rect 857 4029 891 4063
rect 2513 4029 2547 4063
rect 2697 4029 2731 4063
rect 3516 4029 3550 4063
rect 5641 4029 5675 4063
rect 5733 4029 5767 4063
rect 5825 4029 5859 4063
rect 6009 4029 6043 4063
rect 6101 4029 6135 4063
rect 6377 4029 6411 4063
rect 7389 4029 7423 4063
rect 9597 4029 9631 4063
rect 9781 4029 9815 4063
rect 11069 4029 11103 4063
rect 11621 4029 11655 4063
rect 12357 4029 12391 4063
rect 13001 4029 13035 4063
rect 13093 4029 13127 4063
rect 13185 4029 13219 4063
rect 13829 4029 13863 4063
rect 13921 4029 13955 4063
rect 14013 4029 14047 4063
rect 14197 4029 14231 4063
rect 14565 4029 14599 4063
rect 15301 4029 15335 4063
rect 15393 4029 15427 4063
rect 15669 4029 15703 4063
rect 15853 4029 15887 4063
rect 16037 4029 16071 4063
rect 16313 4029 16347 4063
rect 16773 4029 16807 4063
rect 16957 4029 16991 4063
rect 17325 4029 17359 4063
rect 1124 3961 1158 3995
rect 2881 3961 2915 3995
rect 15761 3961 15795 3995
rect 17233 3961 17267 3995
rect 2237 3893 2271 3927
rect 2329 3893 2363 3927
rect 2973 3893 3007 3927
rect 5365 3893 5399 3927
rect 6561 3893 6595 3927
rect 7205 3893 7239 3927
rect 9781 3893 9815 3927
rect 13369 3893 13403 3927
rect 14289 3893 14323 3927
rect 15117 3893 15151 3927
rect 2237 3689 2271 3723
rect 2789 3689 2823 3723
rect 13921 3689 13955 3723
rect 5273 3621 5307 3655
rect 6101 3621 6135 3655
rect 6285 3621 6319 3655
rect 8953 3621 8987 3655
rect 9505 3621 9539 3655
rect 12081 3621 12115 3655
rect 2053 3553 2087 3587
rect 2329 3553 2363 3587
rect 2421 3553 2455 3587
rect 2605 3553 2639 3587
rect 2881 3553 2915 3587
rect 3801 3553 3835 3587
rect 5457 3553 5491 3587
rect 6377 3553 6411 3587
rect 7849 3553 7883 3587
rect 7941 3553 7975 3587
rect 8033 3553 8067 3587
rect 8217 3553 8251 3587
rect 9137 3553 9171 3587
rect 9781 3553 9815 3587
rect 9873 3553 9907 3587
rect 9965 3553 9999 3587
rect 10149 3553 10183 3587
rect 10333 3553 10367 3587
rect 10517 3553 10551 3587
rect 12173 3553 12207 3587
rect 12441 3553 12475 3587
rect 12633 3553 12667 3587
rect 13093 3553 13127 3587
rect 13277 3553 13311 3587
rect 13369 3553 13403 3587
rect 13461 3553 13495 3587
rect 13829 3553 13863 3587
rect 14013 3553 14047 3587
rect 14473 3553 14507 3587
rect 14749 3553 14783 3587
rect 16497 3553 16531 3587
rect 16773 3553 16807 3587
rect 3525 3485 3559 3519
rect 10425 3485 10459 3519
rect 10609 3485 10643 3519
rect 10793 3485 10827 3519
rect 14197 3485 14231 3519
rect 14289 3485 14323 3519
rect 14381 3485 14415 3519
rect 15025 3485 15059 3519
rect 16405 3485 16439 3519
rect 5641 3417 5675 3451
rect 6561 3417 6595 3451
rect 9321 3417 9355 3451
rect 11713 3417 11747 3451
rect 12357 3417 12391 3451
rect 16129 3417 16163 3451
rect 1869 3349 1903 3383
rect 2421 3349 2455 3383
rect 5917 3349 5951 3383
rect 7573 3349 7607 3383
rect 11621 3349 11655 3383
rect 12541 3349 12575 3383
rect 13737 3349 13771 3383
rect 14657 3349 14691 3383
rect 16865 3349 16899 3383
rect 17233 3349 17267 3383
rect 2145 3145 2179 3179
rect 7205 3145 7239 3179
rect 16865 3145 16899 3179
rect 1777 3009 1811 3043
rect 3985 3009 4019 3043
rect 6661 3009 6695 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 9781 3009 9815 3043
rect 9873 3009 9907 3043
rect 13553 3009 13587 3043
rect 13829 3009 13863 3043
rect 14013 3009 14047 3043
rect 15577 3009 15611 3043
rect 17049 3009 17083 3043
rect 1685 2941 1719 2975
rect 2145 2941 2179 2975
rect 2329 2941 2363 2975
rect 3709 2941 3743 2975
rect 3893 2941 3927 2975
rect 4169 2941 4203 2975
rect 4629 2941 4663 2975
rect 4721 2941 4755 2975
rect 5273 2941 5307 2975
rect 5457 2941 5491 2975
rect 5733 2941 5767 2975
rect 5825 2941 5859 2975
rect 5917 2941 5951 2975
rect 6035 2941 6069 2975
rect 6193 2941 6227 2975
rect 6377 2941 6411 2975
rect 6469 2941 6503 2975
rect 6561 2941 6595 2975
rect 7021 2941 7055 2975
rect 7297 2941 7331 2975
rect 7757 2941 7791 2975
rect 7849 2941 7883 2975
rect 9597 2941 9631 2975
rect 9689 2941 9723 2975
rect 11805 2941 11839 2975
rect 11989 2941 12023 2975
rect 12081 2941 12115 2975
rect 12265 2941 12299 2975
rect 12357 2941 12391 2975
rect 13185 2941 13219 2975
rect 13737 2941 13771 2975
rect 13921 2941 13955 2975
rect 15301 2941 15335 2975
rect 16405 2941 16439 2975
rect 16773 2941 16807 2975
rect 17141 2941 17175 2975
rect 17325 2941 17359 2975
rect 5365 2873 5399 2907
rect 14381 2873 14415 2907
rect 14565 2873 14599 2907
rect 17049 2873 17083 2907
rect 2053 2805 2087 2839
rect 3801 2805 3835 2839
rect 4353 2805 4387 2839
rect 4445 2805 4479 2839
rect 5549 2805 5583 2839
rect 6837 2805 6871 2839
rect 7481 2805 7515 2839
rect 8125 2805 8159 2839
rect 9413 2805 9447 2839
rect 13369 2805 13403 2839
rect 14197 2805 14231 2839
rect 16589 2805 16623 2839
rect 17325 2805 17359 2839
rect 3249 2601 3283 2635
rect 5825 2601 5859 2635
rect 11161 2601 11195 2635
rect 16329 2601 16363 2635
rect 17141 2601 17175 2635
rect 3157 2533 3191 2567
rect 7481 2533 7515 2567
rect 7665 2533 7699 2567
rect 11069 2533 11103 2567
rect 16129 2533 16163 2567
rect 17049 2533 17083 2567
rect 1041 2465 1075 2499
rect 3065 2465 3099 2499
rect 3433 2465 3467 2499
rect 4077 2465 4111 2499
rect 4261 2465 4295 2499
rect 6009 2465 6043 2499
rect 6193 2465 6227 2499
rect 6561 2465 6595 2499
rect 9045 2465 9079 2499
rect 9137 2465 9171 2499
rect 9321 2465 9355 2499
rect 9413 2465 9447 2499
rect 11345 2465 11379 2499
rect 12440 2465 12474 2499
rect 12541 2465 12575 2499
rect 12817 2465 12851 2499
rect 14289 2465 14323 2499
rect 14464 2465 14498 2499
rect 14565 2465 14599 2499
rect 14749 2465 14783 2499
rect 14933 2465 14967 2499
rect 15117 2465 15151 2499
rect 15301 2465 15335 2499
rect 15393 2465 15427 2499
rect 15577 2465 15611 2499
rect 15669 2465 15703 2499
rect 16865 2465 16899 2499
rect 17141 2465 17175 2499
rect 17325 2465 17359 2499
rect 1133 2397 1167 2431
rect 6285 2397 6319 2431
rect 14381 2397 14415 2431
rect 14841 2397 14875 2431
rect 15485 2397 15519 2431
rect 1409 2329 1443 2363
rect 6377 2329 6411 2363
rect 12265 2329 12299 2363
rect 13001 2329 13035 2363
rect 3341 2261 3375 2295
rect 4077 2261 4111 2295
rect 7297 2261 7331 2295
rect 8861 2261 8895 2295
rect 11529 2261 11563 2295
rect 12725 2261 12759 2295
rect 14105 2261 14139 2295
rect 15301 2261 15335 2295
rect 15853 2261 15887 2295
rect 16313 2261 16347 2295
rect 16497 2261 16531 2295
rect 16681 2261 16715 2295
rect 3433 2057 3467 2091
rect 6101 2057 6135 2091
rect 10793 2057 10827 2091
rect 15485 2057 15519 2091
rect 16957 2057 16991 2091
rect 17141 2057 17175 2091
rect 3617 1989 3651 2023
rect 5273 1989 5307 2023
rect 5365 1989 5399 2023
rect 6469 1989 6503 2023
rect 9137 1989 9171 2023
rect 10517 1989 10551 2023
rect 11161 1989 11195 2023
rect 12541 1989 12575 2023
rect 14105 1989 14139 2023
rect 14657 1989 14691 2023
rect 1501 1921 1535 1955
rect 4353 1921 4387 1955
rect 6929 1921 6963 1955
rect 7113 1921 7147 1955
rect 7389 1921 7423 1955
rect 9597 1921 9631 1955
rect 11989 1921 12023 1955
rect 12265 1921 12299 1955
rect 13645 1921 13679 1955
rect 13737 1921 13771 1955
rect 13921 1921 13955 1955
rect 15117 1921 15151 1955
rect 1409 1853 1443 1887
rect 1961 1853 1995 1887
rect 2145 1853 2179 1887
rect 2237 1853 2271 1887
rect 2513 1853 2547 1887
rect 2789 1853 2823 1887
rect 2973 1853 3007 1887
rect 3709 1853 3743 1887
rect 3801 1853 3835 1887
rect 3985 1853 4019 1887
rect 4077 1853 4111 1887
rect 4629 1853 4663 1887
rect 4721 1853 4755 1887
rect 4997 1853 5031 1887
rect 5181 1853 5215 1887
rect 5457 1853 5491 1887
rect 6285 1853 6319 1887
rect 6377 1853 6411 1887
rect 6561 1853 6595 1887
rect 6837 1853 6871 1887
rect 7021 1853 7055 1887
rect 7665 1853 7699 1887
rect 8401 1853 8435 1887
rect 8677 1853 8711 1887
rect 8861 1853 8895 1887
rect 9045 1853 9079 1887
rect 9321 1853 9355 1887
rect 9505 1853 9539 1887
rect 9689 1853 9723 1887
rect 9781 1853 9815 1887
rect 9965 1853 9999 1887
rect 10425 1853 10459 1887
rect 10701 1853 10735 1887
rect 10977 1853 11011 1887
rect 11345 1853 11379 1887
rect 12357 1853 12391 1887
rect 12909 1853 12943 1887
rect 13001 1853 13035 1887
rect 13093 1853 13127 1887
rect 13277 1853 13311 1887
rect 13829 1853 13863 1887
rect 14381 1853 14415 1887
rect 14473 1853 14507 1887
rect 14657 1853 14691 1887
rect 15025 1853 15059 1887
rect 15301 1853 15335 1887
rect 15853 1853 15887 1887
rect 16129 1853 16163 1887
rect 16313 1853 16347 1887
rect 16589 1853 16623 1887
rect 16681 1853 16715 1887
rect 17049 1853 17083 1887
rect 17141 1853 17175 1887
rect 17319 1853 17353 1887
rect 3479 1819 3513 1853
rect 3249 1785 3283 1819
rect 15945 1785 15979 1819
rect 16037 1785 16071 1819
rect 1777 1717 1811 1751
rect 2145 1717 2179 1751
rect 2329 1717 2363 1751
rect 2697 1717 2731 1751
rect 2973 1717 3007 1751
rect 4261 1717 4295 1751
rect 4537 1717 4571 1751
rect 4905 1717 4939 1751
rect 7297 1717 7331 1751
rect 8585 1717 8619 1751
rect 10149 1717 10183 1751
rect 10241 1717 10275 1751
rect 12633 1717 12667 1751
rect 14289 1717 14323 1751
rect 14841 1717 14875 1751
rect 15669 1717 15703 1751
rect 16405 1717 16439 1751
rect 2421 1513 2455 1547
rect 2973 1513 3007 1547
rect 3709 1513 3743 1547
rect 7021 1513 7055 1547
rect 12633 1513 12667 1547
rect 15025 1513 15059 1547
rect 15761 1513 15795 1547
rect 2237 1445 2271 1479
rect 2605 1445 2639 1479
rect 2805 1445 2839 1479
rect 3801 1445 3835 1479
rect 11897 1445 11931 1479
rect 13185 1445 13219 1479
rect 16221 1445 16255 1479
rect 16865 1445 16899 1479
rect 1317 1377 1351 1411
rect 1685 1377 1719 1411
rect 2053 1377 2087 1411
rect 3249 1377 3283 1411
rect 3341 1377 3375 1411
rect 3985 1377 4019 1411
rect 4077 1377 4111 1411
rect 4169 1377 4203 1411
rect 4353 1377 4387 1411
rect 4813 1377 4847 1411
rect 5549 1377 5583 1411
rect 6009 1377 6043 1411
rect 6285 1377 6319 1411
rect 6469 1377 6503 1411
rect 6929 1377 6963 1411
rect 7021 1377 7055 1411
rect 7205 1377 7239 1411
rect 7481 1377 7515 1411
rect 7665 1377 7699 1411
rect 7941 1377 7975 1411
rect 8125 1377 8159 1411
rect 9045 1377 9079 1411
rect 9229 1377 9263 1411
rect 9689 1377 9723 1411
rect 9781 1377 9815 1411
rect 9873 1377 9907 1411
rect 10057 1377 10091 1411
rect 10333 1377 10367 1411
rect 10609 1377 10643 1411
rect 11253 1377 11287 1411
rect 12357 1377 12391 1411
rect 12817 1377 12851 1411
rect 13001 1377 13035 1411
rect 13369 1377 13403 1411
rect 13553 1377 13587 1411
rect 13921 1377 13955 1411
rect 14105 1377 14139 1411
rect 14381 1377 14415 1411
rect 14565 1377 14599 1411
rect 14841 1377 14875 1411
rect 15393 1377 15427 1411
rect 17049 1377 17083 1411
rect 3433 1309 3467 1343
rect 3525 1309 3559 1343
rect 4721 1309 4755 1343
rect 5181 1309 5215 1343
rect 6101 1309 6135 1343
rect 6193 1309 6227 1343
rect 7297 1309 7331 1343
rect 7757 1309 7791 1343
rect 7849 1309 7883 1343
rect 8309 1309 8343 1343
rect 9321 1309 9355 1343
rect 10517 1309 10551 1343
rect 10977 1309 11011 1343
rect 12081 1309 12115 1343
rect 13093 1309 13127 1343
rect 13645 1309 13679 1343
rect 14197 1309 14231 1343
rect 14289 1309 14323 1343
rect 15301 1309 15335 1343
rect 16681 1309 16715 1343
rect 3893 1241 3927 1275
rect 8861 1241 8895 1275
rect 10149 1241 10183 1275
rect 10425 1241 10459 1275
rect 13737 1241 13771 1275
rect 14749 1241 14783 1275
rect 1133 1173 1167 1207
rect 1501 1173 1535 1207
rect 2789 1173 2823 1207
rect 4261 1173 4295 1207
rect 5365 1173 5399 1207
rect 5825 1173 5859 1207
rect 6653 1173 6687 1207
rect 6745 1173 6779 1207
rect 9413 1173 9447 1207
rect 11069 1173 11103 1207
rect 11437 1173 11471 1207
rect 11621 1173 11655 1207
rect 12173 1173 12207 1207
rect 12541 1173 12575 1207
rect 16313 1173 16347 1207
rect 2513 969 2547 1003
rect 9873 969 9907 1003
rect 10517 969 10551 1003
rect 11069 969 11103 1003
rect 11621 969 11655 1003
rect 12725 969 12759 1003
rect 14381 969 14415 1003
rect 14933 969 14967 1003
rect 15301 969 15335 1003
rect 16313 969 16347 1003
rect 17049 969 17083 1003
rect 2697 901 2731 935
rect 13093 901 13127 935
rect 13185 833 13219 867
rect 15761 833 15795 867
rect 16681 833 16715 867
rect 1133 765 1167 799
rect 1593 765 1627 799
rect 2237 765 2271 799
rect 2513 765 2547 799
rect 2881 765 2915 799
rect 3525 765 3559 799
rect 3893 765 3927 799
rect 4629 765 4663 799
rect 5365 765 5399 799
rect 6101 765 6135 799
rect 6837 765 6871 799
rect 7297 765 7331 799
rect 8217 765 8251 799
rect 8493 765 8527 799
rect 9597 765 9631 799
rect 9781 765 9815 799
rect 10057 765 10091 799
rect 10977 765 11011 799
rect 11253 765 11287 799
rect 11805 765 11839 799
rect 11989 765 12023 799
rect 12449 765 12483 799
rect 12909 765 12943 799
rect 13645 765 13679 799
rect 14289 765 14323 799
rect 14565 765 14599 799
rect 14841 765 14875 799
rect 15117 765 15151 799
rect 16865 765 16899 799
rect 2421 697 2455 731
rect 10241 697 10275 731
rect 10425 697 10459 731
rect 14749 697 14783 731
rect 15485 697 15519 731
rect 16221 697 16255 731
rect 949 629 983 663
rect 1317 629 1351 663
rect 3341 629 3375 663
rect 3709 629 3743 663
rect 4445 629 4479 663
rect 5181 629 5215 663
rect 5917 629 5951 663
rect 6653 629 6687 663
rect 7481 629 7515 663
rect 8033 629 8067 663
rect 8585 629 8619 663
rect 9505 629 9539 663
rect 11437 629 11471 663
rect 12173 629 12207 663
rect 13737 629 13771 663
<< metal1 >>
rect 12802 17620 12808 17672
rect 12860 17660 12866 17672
rect 14090 17660 14096 17672
rect 12860 17632 14096 17660
rect 12860 17620 12866 17632
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 11790 17592 11796 17604
rect 7340 17564 11796 17592
rect 7340 17552 7346 17564
rect 11790 17552 11796 17564
rect 11848 17592 11854 17604
rect 14826 17592 14832 17604
rect 11848 17564 14832 17592
rect 11848 17552 11854 17564
rect 14826 17552 14832 17564
rect 14884 17552 14890 17604
rect 2958 17484 2964 17536
rect 3016 17524 3022 17536
rect 7190 17524 7196 17536
rect 3016 17496 7196 17524
rect 3016 17484 3022 17496
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 11422 17484 11428 17536
rect 11480 17524 11486 17536
rect 12986 17524 12992 17536
rect 11480 17496 12992 17524
rect 11480 17484 11486 17496
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 13630 17484 13636 17536
rect 13688 17524 13694 17536
rect 14550 17524 14556 17536
rect 13688 17496 14556 17524
rect 13688 17484 13694 17496
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 552 17434 17664 17456
rect 552 17382 1366 17434
rect 1418 17382 1430 17434
rect 1482 17382 1494 17434
rect 1546 17382 1558 17434
rect 1610 17382 1622 17434
rect 1674 17382 1686 17434
rect 1738 17382 7366 17434
rect 7418 17382 7430 17434
rect 7482 17382 7494 17434
rect 7546 17382 7558 17434
rect 7610 17382 7622 17434
rect 7674 17382 7686 17434
rect 7738 17382 13366 17434
rect 13418 17382 13430 17434
rect 13482 17382 13494 17434
rect 13546 17382 13558 17434
rect 13610 17382 13622 17434
rect 13674 17382 13686 17434
rect 13738 17382 17664 17434
rect 552 17360 17664 17382
rect 1210 17280 1216 17332
rect 1268 17280 1274 17332
rect 2038 17280 2044 17332
rect 2096 17280 2102 17332
rect 2866 17280 2872 17332
rect 2924 17280 2930 17332
rect 3694 17280 3700 17332
rect 3752 17320 3758 17332
rect 4065 17323 4123 17329
rect 4065 17320 4077 17323
rect 3752 17292 4077 17320
rect 3752 17280 3758 17292
rect 4065 17289 4077 17292
rect 4111 17289 4123 17323
rect 4065 17283 4123 17289
rect 4522 17280 4528 17332
rect 4580 17320 4586 17332
rect 4709 17323 4767 17329
rect 4709 17320 4721 17323
rect 4580 17292 4721 17320
rect 4580 17280 4586 17292
rect 4709 17289 4721 17292
rect 4755 17289 4767 17323
rect 4709 17283 4767 17289
rect 5350 17280 5356 17332
rect 5408 17320 5414 17332
rect 5905 17323 5963 17329
rect 5905 17320 5917 17323
rect 5408 17292 5917 17320
rect 5408 17280 5414 17292
rect 5905 17289 5917 17292
rect 5951 17289 5963 17323
rect 5905 17283 5963 17289
rect 6178 17280 6184 17332
rect 6236 17320 6242 17332
rect 6236 17292 6960 17320
rect 6236 17280 6242 17292
rect 2884 17252 2912 17280
rect 5261 17255 5319 17261
rect 5261 17252 5273 17255
rect 2884 17224 5273 17252
rect 5261 17221 5273 17224
rect 5307 17221 5319 17255
rect 5261 17215 5319 17221
rect 6549 17255 6607 17261
rect 6549 17221 6561 17255
rect 6595 17252 6607 17255
rect 6730 17252 6736 17264
rect 6595 17224 6736 17252
rect 6595 17221 6607 17224
rect 6549 17215 6607 17221
rect 6730 17212 6736 17224
rect 6788 17212 6794 17264
rect 6932 17252 6960 17292
rect 7006 17280 7012 17332
rect 7064 17320 7070 17332
rect 7285 17323 7343 17329
rect 7285 17320 7297 17323
rect 7064 17292 7297 17320
rect 7064 17280 7070 17292
rect 7285 17289 7297 17292
rect 7331 17289 7343 17323
rect 7285 17283 7343 17289
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 8113 17323 8171 17329
rect 8113 17320 8125 17323
rect 7892 17292 8125 17320
rect 7892 17280 7898 17292
rect 8113 17289 8125 17292
rect 8159 17289 8171 17323
rect 8113 17283 8171 17289
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 8849 17323 8907 17329
rect 8849 17320 8861 17323
rect 8720 17292 8861 17320
rect 8720 17280 8726 17292
rect 8849 17289 8861 17292
rect 8895 17289 8907 17323
rect 8849 17283 8907 17289
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 11204 17292 13676 17320
rect 11204 17280 11210 17292
rect 7653 17255 7711 17261
rect 7653 17252 7665 17255
rect 6932 17224 7665 17252
rect 7653 17221 7665 17224
rect 7699 17221 7711 17255
rect 12713 17255 12771 17261
rect 12713 17252 12725 17255
rect 7653 17215 7711 17221
rect 11532 17224 12725 17252
rect 1504 17156 2912 17184
rect 1504 17125 1532 17156
rect 1489 17119 1547 17125
rect 1489 17085 1501 17119
rect 1535 17085 1547 17119
rect 1489 17079 1547 17085
rect 1857 17119 1915 17125
rect 1857 17085 1869 17119
rect 1903 17085 1915 17119
rect 1857 17079 1915 17085
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17116 2283 17119
rect 2774 17116 2780 17128
rect 2271 17088 2780 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 1872 17048 1900 17079
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 2884 17116 2912 17156
rect 2958 17144 2964 17196
rect 3016 17144 3022 17196
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 7282 17184 7288 17196
rect 3712 17156 7288 17184
rect 3068 17116 3096 17144
rect 2884 17088 3096 17116
rect 2685 17051 2743 17057
rect 1872 17020 2360 17048
rect 1670 16940 1676 16992
rect 1728 16940 1734 16992
rect 2332 16989 2360 17020
rect 2685 17017 2697 17051
rect 2731 17048 2743 17051
rect 3237 17051 3295 17057
rect 3237 17048 3249 17051
rect 2731 17020 3249 17048
rect 2731 17017 2743 17020
rect 2685 17011 2743 17017
rect 3237 17017 3249 17020
rect 3283 17017 3295 17051
rect 3237 17011 3295 17017
rect 2317 16983 2375 16989
rect 2317 16949 2329 16983
rect 2363 16949 2375 16983
rect 2317 16943 2375 16949
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 3712 16980 3740 17156
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 11532 17193 11560 17224
rect 12713 17221 12725 17224
rect 12759 17221 12771 17255
rect 12713 17215 12771 17221
rect 12986 17212 12992 17264
rect 13044 17252 13050 17264
rect 13541 17255 13599 17261
rect 13541 17252 13553 17255
rect 13044 17224 13553 17252
rect 13044 17212 13050 17224
rect 13541 17221 13553 17224
rect 13587 17221 13599 17255
rect 13541 17215 13599 17221
rect 8481 17187 8539 17193
rect 8481 17184 8493 17187
rect 7392 17156 8493 17184
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17085 3847 17119
rect 3789 17079 3847 17085
rect 3804 17048 3832 17079
rect 4246 17076 4252 17128
rect 4304 17076 4310 17128
rect 4890 17076 4896 17128
rect 4948 17076 4954 17128
rect 6822 17076 6828 17128
rect 6880 17076 6886 17128
rect 7098 17076 7104 17128
rect 7156 17076 7162 17128
rect 5077 17051 5135 17057
rect 5077 17048 5089 17051
rect 3804 17020 5089 17048
rect 3804 16992 3832 17020
rect 5077 17017 5089 17020
rect 5123 17017 5135 17051
rect 5077 17011 5135 17017
rect 6181 17051 6239 17057
rect 6181 17017 6193 17051
rect 6227 17048 6239 17051
rect 6454 17048 6460 17060
rect 6227 17020 6460 17048
rect 6227 17017 6239 17020
rect 6181 17011 6239 17017
rect 6454 17008 6460 17020
rect 6512 17008 6518 17060
rect 6546 17008 6552 17060
rect 6604 17008 6610 17060
rect 6733 17051 6791 17057
rect 6733 17017 6745 17051
rect 6779 17048 6791 17051
rect 7392 17048 7420 17156
rect 8481 17153 8493 17156
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 11664 17156 12449 17184
rect 11664 17144 11670 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17085 7527 17119
rect 7469 17079 7527 17085
rect 6779 17020 7420 17048
rect 6779 17017 6791 17020
rect 6733 17011 6791 17017
rect 2823 16952 3740 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 3786 16940 3792 16992
rect 3844 16940 3850 16992
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 5442 16980 5448 16992
rect 4304 16952 5448 16980
rect 4304 16940 4310 16952
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 6362 16940 6368 16992
rect 6420 16980 6426 16992
rect 7484 16980 7512 17079
rect 7926 17076 7932 17128
rect 7984 17076 7990 17128
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17085 8631 17119
rect 8573 17079 8631 17085
rect 8588 16992 8616 17079
rect 9030 17076 9036 17128
rect 9088 17076 9094 17128
rect 9125 17119 9183 17125
rect 9125 17085 9137 17119
rect 9171 17085 9183 17119
rect 9125 17079 9183 17085
rect 9140 17048 9168 17079
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 9548 17088 9781 17116
rect 9548 17076 9554 17088
rect 9769 17085 9781 17088
rect 9815 17085 9827 17119
rect 9769 17079 9827 17085
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17116 9919 17119
rect 10318 17116 10324 17128
rect 9907 17088 10324 17116
rect 9907 17085 9919 17088
rect 9861 17079 9919 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 10778 17076 10784 17128
rect 10836 17076 10842 17128
rect 11422 17076 11428 17128
rect 11480 17076 11486 17128
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 13357 17119 13415 17125
rect 12032 17088 13216 17116
rect 12032 17076 12038 17088
rect 12253 17051 12311 17057
rect 9140 17020 11928 17048
rect 6420 16952 7512 16980
rect 6420 16940 6426 16952
rect 8570 16940 8576 16992
rect 8628 16940 8634 16992
rect 9306 16940 9312 16992
rect 9364 16940 9370 16992
rect 9398 16940 9404 16992
rect 9456 16980 9462 16992
rect 9585 16983 9643 16989
rect 9585 16980 9597 16983
rect 9456 16952 9597 16980
rect 9456 16940 9462 16952
rect 9585 16949 9597 16952
rect 9631 16949 9643 16983
rect 9585 16943 9643 16949
rect 10042 16940 10048 16992
rect 10100 16940 10106 16992
rect 10134 16940 10140 16992
rect 10192 16940 10198 16992
rect 11054 16940 11060 16992
rect 11112 16940 11118 16992
rect 11900 16989 11928 17020
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 12710 17048 12716 17060
rect 12299 17020 12716 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12710 17008 12716 17020
rect 12768 17048 12774 17060
rect 13188 17048 13216 17088
rect 13357 17085 13369 17119
rect 13403 17116 13415 17119
rect 13446 17116 13452 17128
rect 13403 17088 13452 17116
rect 13403 17085 13415 17088
rect 13357 17079 13415 17085
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 13648 17116 13676 17292
rect 15286 17280 15292 17332
rect 15344 17320 15350 17332
rect 16206 17320 16212 17332
rect 15344 17292 16212 17320
rect 15344 17280 15350 17292
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 13814 17212 13820 17264
rect 13872 17212 13878 17264
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 16172 17156 16221 17184
rect 16172 17144 16178 17156
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13648 17088 13737 17116
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 14016 17048 14044 17079
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 14148 17088 14289 17116
rect 14148 17076 14154 17088
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 14553 17119 14611 17125
rect 14553 17116 14565 17119
rect 14424 17088 14565 17116
rect 14424 17076 14430 17088
rect 14553 17085 14565 17088
rect 14599 17085 14611 17119
rect 14553 17079 14611 17085
rect 15378 17076 15384 17128
rect 15436 17116 15442 17128
rect 16485 17119 16543 17125
rect 16485 17116 16497 17119
rect 15436 17088 16497 17116
rect 15436 17076 15442 17088
rect 16485 17085 16497 17088
rect 16531 17085 16543 17119
rect 16485 17079 16543 17085
rect 12768 17020 13124 17048
rect 13188 17020 14044 17048
rect 14820 17051 14878 17057
rect 12768 17008 12774 17020
rect 11885 16983 11943 16989
rect 11885 16949 11897 16983
rect 11931 16949 11943 16983
rect 11885 16943 11943 16949
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 12345 16983 12403 16989
rect 12345 16980 12357 16983
rect 12124 16952 12357 16980
rect 12124 16940 12130 16952
rect 12345 16949 12357 16952
rect 12391 16949 12403 16983
rect 13096 16980 13124 17020
rect 14820 17017 14832 17051
rect 14866 17048 14878 17051
rect 15102 17048 15108 17060
rect 14866 17020 15108 17048
rect 14866 17017 14878 17020
rect 14820 17011 14878 17017
rect 15102 17008 15108 17020
rect 15160 17008 15166 17060
rect 14093 16983 14151 16989
rect 14093 16980 14105 16983
rect 13096 16952 14105 16980
rect 12345 16943 12403 16949
rect 14093 16949 14105 16952
rect 14139 16949 14151 16983
rect 14093 16943 14151 16949
rect 15838 16940 15844 16992
rect 15896 16980 15902 16992
rect 15933 16983 15991 16989
rect 15933 16980 15945 16983
rect 15896 16952 15945 16980
rect 15896 16940 15902 16952
rect 15933 16949 15945 16952
rect 15979 16949 15991 16983
rect 15933 16943 15991 16949
rect 552 16890 17664 16912
rect 552 16838 4366 16890
rect 4418 16838 4430 16890
rect 4482 16838 4494 16890
rect 4546 16838 4558 16890
rect 4610 16838 4622 16890
rect 4674 16838 4686 16890
rect 4738 16838 10366 16890
rect 10418 16838 10430 16890
rect 10482 16838 10494 16890
rect 10546 16838 10558 16890
rect 10610 16838 10622 16890
rect 10674 16838 10686 16890
rect 10738 16838 16366 16890
rect 16418 16838 16430 16890
rect 16482 16838 16494 16890
rect 16546 16838 16558 16890
rect 16610 16838 16622 16890
rect 16674 16838 16686 16890
rect 16738 16838 17664 16890
rect 552 16816 17664 16838
rect 1670 16736 1676 16788
rect 1728 16736 1734 16788
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 3786 16776 3792 16788
rect 2455 16748 3792 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 3786 16736 3792 16748
rect 3844 16736 3850 16788
rect 5261 16779 5319 16785
rect 5261 16745 5273 16779
rect 5307 16776 5319 16779
rect 5534 16776 5540 16788
rect 5307 16748 5540 16776
rect 5307 16745 5319 16748
rect 5261 16739 5319 16745
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 6362 16736 6368 16788
rect 6420 16736 6426 16788
rect 6546 16736 6552 16788
rect 6604 16736 6610 16788
rect 7377 16779 7435 16785
rect 7377 16776 7389 16779
rect 6656 16748 7389 16776
rect 1296 16711 1354 16717
rect 1296 16677 1308 16711
rect 1342 16708 1354 16711
rect 1688 16708 1716 16736
rect 6656 16708 6684 16748
rect 7377 16745 7389 16748
rect 7423 16745 7435 16779
rect 7377 16739 7435 16745
rect 9306 16736 9312 16788
rect 9364 16736 9370 16788
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 10413 16779 10471 16785
rect 10413 16776 10425 16779
rect 10192 16748 10425 16776
rect 10192 16736 10198 16748
rect 10413 16745 10425 16748
rect 10459 16745 10471 16779
rect 10413 16739 10471 16745
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 13722 16776 13728 16788
rect 12860 16748 13728 16776
rect 12860 16736 12866 16748
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 14516 16748 15792 16776
rect 14516 16736 14522 16748
rect 1342 16680 1716 16708
rect 4816 16680 6684 16708
rect 6733 16711 6791 16717
rect 1342 16677 1354 16680
rect 1296 16671 1354 16677
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 2869 16643 2927 16649
rect 2869 16640 2881 16643
rect 2832 16612 2881 16640
rect 2832 16600 2838 16612
rect 2869 16609 2881 16612
rect 2915 16640 2927 16643
rect 2958 16640 2964 16652
rect 2915 16612 2964 16640
rect 2915 16609 2927 16612
rect 2869 16603 2927 16609
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3050 16600 3056 16652
rect 3108 16600 3114 16652
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 4816 16649 4844 16680
rect 6733 16677 6745 16711
rect 6779 16677 6791 16711
rect 6733 16671 6791 16677
rect 7745 16711 7803 16717
rect 7745 16677 7757 16711
rect 7791 16708 7803 16711
rect 9214 16708 9220 16720
rect 7791 16680 9220 16708
rect 7791 16677 7803 16680
rect 7745 16671 7803 16677
rect 3401 16643 3459 16649
rect 3401 16640 3413 16643
rect 3292 16612 3413 16640
rect 3292 16600 3298 16612
rect 3401 16609 3413 16612
rect 3447 16609 3459 16643
rect 3401 16603 3459 16609
rect 4801 16643 4859 16649
rect 4801 16609 4813 16643
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 5077 16643 5135 16649
rect 5077 16609 5089 16643
rect 5123 16609 5135 16643
rect 5077 16603 5135 16609
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16640 5595 16643
rect 5902 16640 5908 16652
rect 5583 16612 5908 16640
rect 5583 16609 5595 16612
rect 5537 16603 5595 16609
rect 842 16532 848 16584
rect 900 16572 906 16584
rect 1029 16575 1087 16581
rect 1029 16572 1041 16575
rect 900 16544 1041 16572
rect 900 16532 906 16544
rect 1029 16541 1041 16544
rect 1075 16541 1087 16575
rect 3145 16575 3203 16581
rect 3145 16572 3157 16575
rect 1029 16535 1087 16541
rect 2792 16544 3157 16572
rect 2792 16448 2820 16544
rect 3145 16541 3157 16544
rect 3191 16541 3203 16575
rect 3145 16535 3203 16541
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 5092 16572 5120 16603
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 5994 16600 6000 16652
rect 6052 16600 6058 16652
rect 6270 16600 6276 16652
rect 6328 16640 6334 16652
rect 6748 16640 6776 16671
rect 9214 16668 9220 16680
rect 9272 16668 9278 16720
rect 9324 16649 9352 16736
rect 14366 16708 14372 16720
rect 9600 16680 14372 16708
rect 9600 16652 9628 16680
rect 9318 16643 9376 16649
rect 6328 16612 6776 16640
rect 6932 16612 8248 16640
rect 6328 16600 6334 16612
rect 4304 16544 5120 16572
rect 6089 16575 6147 16581
rect 4304 16532 4310 16544
rect 6089 16541 6101 16575
rect 6135 16572 6147 16575
rect 6178 16572 6184 16584
rect 6135 16544 6184 16572
rect 6135 16541 6147 16544
rect 6089 16535 6147 16541
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 6362 16504 6368 16516
rect 4172 16476 6368 16504
rect 2774 16396 2780 16448
rect 2832 16396 2838 16448
rect 3053 16439 3111 16445
rect 3053 16405 3065 16439
rect 3099 16436 3111 16439
rect 4172 16436 4200 16476
rect 6362 16464 6368 16476
rect 6420 16464 6426 16516
rect 3099 16408 4200 16436
rect 3099 16405 3111 16408
rect 3053 16399 3111 16405
rect 4246 16396 4252 16448
rect 4304 16436 4310 16448
rect 4525 16439 4583 16445
rect 4525 16436 4537 16439
rect 4304 16408 4537 16436
rect 4304 16396 4310 16408
rect 4525 16405 4537 16408
rect 4571 16405 4583 16439
rect 4525 16399 4583 16405
rect 4614 16396 4620 16448
rect 4672 16396 4678 16448
rect 5350 16396 5356 16448
rect 5408 16396 5414 16448
rect 6733 16439 6791 16445
rect 6733 16405 6745 16439
rect 6779 16436 6791 16439
rect 6932 16436 6960 16612
rect 7006 16532 7012 16584
rect 7064 16572 7070 16584
rect 7837 16575 7895 16581
rect 7837 16572 7849 16575
rect 7064 16544 7849 16572
rect 7064 16532 7070 16544
rect 7837 16541 7849 16544
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 7101 16507 7159 16513
rect 7101 16473 7113 16507
rect 7147 16504 7159 16507
rect 7374 16504 7380 16516
rect 7147 16476 7380 16504
rect 7147 16473 7159 16476
rect 7101 16467 7159 16473
rect 7374 16464 7380 16476
rect 7432 16464 7438 16516
rect 6779 16408 6960 16436
rect 6779 16405 6791 16408
rect 6733 16399 6791 16405
rect 7006 16396 7012 16448
rect 7064 16436 7070 16448
rect 7944 16436 7972 16535
rect 8220 16445 8248 16612
rect 9318 16609 9330 16643
rect 9364 16609 9376 16643
rect 9318 16603 9376 16609
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 9861 16643 9919 16649
rect 9861 16609 9873 16643
rect 9907 16640 9919 16643
rect 9907 16612 9996 16640
rect 9907 16609 9919 16612
rect 9861 16603 9919 16609
rect 9968 16513 9996 16612
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 10321 16643 10379 16649
rect 10321 16640 10333 16643
rect 10100 16612 10333 16640
rect 10100 16600 10106 16612
rect 10321 16609 10333 16612
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11532 16649 11560 16680
rect 11241 16643 11299 16649
rect 11241 16640 11253 16643
rect 11112 16612 11253 16640
rect 11112 16600 11118 16612
rect 11241 16609 11253 16612
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16609 11575 16643
rect 11773 16643 11831 16649
rect 11773 16640 11785 16643
rect 11517 16603 11575 16609
rect 11624 16612 11785 16640
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 11624 16572 11652 16612
rect 11773 16609 11785 16612
rect 11819 16609 11831 16643
rect 11773 16603 11831 16609
rect 13170 16600 13176 16652
rect 13228 16640 13234 16652
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 13228 16612 13277 16640
rect 13228 16600 13234 16612
rect 13265 16609 13277 16612
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 13354 16600 13360 16652
rect 13412 16640 13418 16652
rect 13832 16649 13860 16680
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13412 16612 13553 16640
rect 13412 16600 13418 16612
rect 13541 16609 13553 16612
rect 13587 16609 13599 16643
rect 13541 16603 13599 16609
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16609 13875 16643
rect 14073 16643 14131 16649
rect 14073 16640 14085 16643
rect 13817 16603 13875 16609
rect 13924 16612 14085 16640
rect 13446 16572 13452 16584
rect 10597 16535 10655 16541
rect 11440 16544 11652 16572
rect 12912 16544 13452 16572
rect 9953 16507 10011 16513
rect 9953 16473 9965 16507
rect 9999 16473 10011 16507
rect 9953 16467 10011 16473
rect 7064 16408 7972 16436
rect 8205 16439 8263 16445
rect 7064 16396 7070 16408
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 8570 16436 8576 16448
rect 8251 16408 8576 16436
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 8570 16396 8576 16408
rect 8628 16436 8634 16448
rect 9214 16436 9220 16448
rect 8628 16408 9220 16436
rect 8628 16396 8634 16408
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 9674 16396 9680 16448
rect 9732 16396 9738 16448
rect 10612 16436 10640 16535
rect 11440 16513 11468 16544
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16473 11483 16507
rect 11425 16467 11483 16473
rect 11514 16464 11520 16516
rect 11572 16464 11578 16516
rect 12912 16513 12940 16544
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 13924 16572 13952 16612
rect 14073 16609 14085 16612
rect 14119 16609 14131 16643
rect 14073 16603 14131 16609
rect 14550 16600 14556 16652
rect 14608 16640 14614 16652
rect 15764 16649 15792 16748
rect 16206 16736 16212 16788
rect 16264 16736 16270 16788
rect 16224 16708 16252 16736
rect 16224 16680 17172 16708
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 14608 16612 15485 16640
rect 14608 16600 14614 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 17144 16649 17172 16680
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 16080 16612 16497 16640
rect 16080 16600 16086 16612
rect 16485 16609 16497 16612
rect 16531 16640 16543 16643
rect 17129 16643 17187 16649
rect 16531 16612 16988 16640
rect 16531 16609 16543 16612
rect 16485 16603 16543 16609
rect 13832 16544 13952 16572
rect 12897 16507 12955 16513
rect 12897 16473 12909 16507
rect 12943 16473 12955 16507
rect 12897 16467 12955 16473
rect 13725 16507 13783 16513
rect 13725 16473 13737 16507
rect 13771 16504 13783 16507
rect 13832 16504 13860 16544
rect 14826 16532 14832 16584
rect 14884 16532 14890 16584
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 16577 16575 16635 16581
rect 16577 16572 16589 16575
rect 15896 16544 16589 16572
rect 15896 16532 15902 16544
rect 16577 16541 16589 16544
rect 16623 16541 16635 16575
rect 16577 16535 16635 16541
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 13771 16476 13860 16504
rect 13771 16473 13783 16476
rect 13725 16467 13783 16473
rect 11532 16436 11560 16464
rect 10612 16408 11560 16436
rect 12526 16396 12532 16448
rect 12584 16436 12590 16448
rect 12912 16436 12940 16467
rect 12584 16408 12940 16436
rect 12584 16396 12590 16408
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 14182 16436 14188 16448
rect 13136 16408 14188 16436
rect 13136 16396 13142 16408
rect 14182 16396 14188 16408
rect 14240 16396 14246 16448
rect 14844 16436 14872 16532
rect 15010 16464 15016 16516
rect 15068 16504 15074 16516
rect 16684 16504 16712 16535
rect 16960 16513 16988 16612
rect 17129 16609 17141 16643
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 15068 16476 16712 16504
rect 16945 16507 17003 16513
rect 15068 16464 15074 16476
rect 16945 16473 16957 16507
rect 16991 16473 17003 16507
rect 16945 16467 17003 16473
rect 15197 16439 15255 16445
rect 15197 16436 15209 16439
rect 14844 16408 15209 16436
rect 15197 16405 15209 16408
rect 15243 16405 15255 16439
rect 15197 16399 15255 16405
rect 15286 16396 15292 16448
rect 15344 16396 15350 16448
rect 15562 16396 15568 16448
rect 15620 16396 15626 16448
rect 16114 16396 16120 16448
rect 16172 16396 16178 16448
rect 552 16346 17664 16368
rect 552 16294 1366 16346
rect 1418 16294 1430 16346
rect 1482 16294 1494 16346
rect 1546 16294 1558 16346
rect 1610 16294 1622 16346
rect 1674 16294 1686 16346
rect 1738 16294 7366 16346
rect 7418 16294 7430 16346
rect 7482 16294 7494 16346
rect 7546 16294 7558 16346
rect 7610 16294 7622 16346
rect 7674 16294 7686 16346
rect 7738 16294 13366 16346
rect 13418 16294 13430 16346
rect 13482 16294 13494 16346
rect 13546 16294 13558 16346
rect 13610 16294 13622 16346
rect 13674 16294 13686 16346
rect 13738 16294 17664 16346
rect 552 16272 17664 16294
rect 6730 16192 6736 16244
rect 6788 16192 6794 16244
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 7009 16235 7067 16241
rect 7009 16232 7021 16235
rect 6880 16204 7021 16232
rect 6880 16192 6886 16204
rect 7009 16201 7021 16204
rect 7055 16201 7067 16235
rect 7009 16195 7067 16201
rect 7190 16192 7196 16244
rect 7248 16192 7254 16244
rect 7282 16192 7288 16244
rect 7340 16192 7346 16244
rect 9582 16232 9588 16244
rect 9324 16204 9588 16232
rect 3053 16167 3111 16173
rect 3053 16133 3065 16167
rect 3099 16164 3111 16167
rect 3234 16164 3240 16176
rect 3099 16136 3240 16164
rect 3099 16133 3111 16136
rect 3053 16127 3111 16133
rect 3234 16124 3240 16136
rect 3292 16124 3298 16176
rect 2774 16096 2780 16108
rect 2599 16068 2780 16096
rect 842 15988 848 16040
rect 900 16028 906 16040
rect 1213 16031 1271 16037
rect 1213 16028 1225 16031
rect 900 16000 1225 16028
rect 900 15988 906 16000
rect 1213 15997 1225 16000
rect 1259 16028 1271 16031
rect 2599 16028 2627 16068
rect 2774 16056 2780 16068
rect 2832 16096 2838 16108
rect 4617 16099 4675 16105
rect 2832 16068 3188 16096
rect 2832 16056 2838 16068
rect 1259 16000 2627 16028
rect 2869 16031 2927 16037
rect 1259 15997 1271 16000
rect 1213 15991 1271 15997
rect 2869 15997 2881 16031
rect 2915 16028 2927 16031
rect 3050 16028 3056 16040
rect 2915 16000 3056 16028
rect 2915 15997 2927 16000
rect 2869 15991 2927 15997
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 3160 16028 3188 16068
rect 4617 16065 4629 16099
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 4632 16028 4660 16059
rect 6454 16056 6460 16108
rect 6512 16056 6518 16108
rect 6748 16096 6776 16192
rect 7208 16164 7236 16192
rect 7929 16167 7987 16173
rect 7929 16164 7941 16167
rect 7208 16136 7941 16164
rect 7929 16133 7941 16136
rect 7975 16133 7987 16167
rect 7929 16127 7987 16133
rect 9324 16105 9352 16204
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 10689 16235 10747 16241
rect 10689 16201 10701 16235
rect 10735 16232 10747 16235
rect 10778 16232 10784 16244
rect 10735 16204 10784 16232
rect 10735 16201 10747 16204
rect 10689 16195 10747 16201
rect 10778 16192 10784 16204
rect 10836 16232 10842 16244
rect 11514 16232 11520 16244
rect 10836 16204 11520 16232
rect 10836 16192 10842 16204
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 12342 16232 12348 16244
rect 12268 16204 12348 16232
rect 11146 16124 11152 16176
rect 11204 16164 11210 16176
rect 12268 16164 12296 16204
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 13541 16235 13599 16241
rect 13541 16232 13553 16235
rect 13320 16204 13553 16232
rect 13320 16192 13326 16204
rect 13541 16201 13553 16204
rect 13587 16201 13599 16235
rect 13541 16195 13599 16201
rect 11204 16136 12296 16164
rect 11204 16124 11210 16136
rect 12618 16124 12624 16176
rect 12676 16164 12682 16176
rect 13078 16164 13084 16176
rect 12676 16136 13084 16164
rect 12676 16124 12682 16136
rect 13078 16124 13084 16136
rect 13136 16124 13142 16176
rect 14369 16167 14427 16173
rect 14369 16164 14381 16167
rect 14016 16136 14381 16164
rect 9309 16099 9367 16105
rect 6748 16068 8064 16096
rect 4801 16031 4859 16037
rect 4801 16028 4813 16031
rect 3160 16000 4813 16028
rect 4801 15997 4813 16000
rect 4847 15997 4859 16031
rect 4801 15991 4859 15997
rect 5068 16031 5126 16037
rect 5068 15997 5080 16031
rect 5114 16028 5126 16031
rect 5350 16028 5356 16040
rect 5114 16000 5356 16028
rect 5114 15997 5126 16000
rect 5068 15991 5126 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 6549 16031 6607 16037
rect 6549 16028 6561 16031
rect 5552 16000 6561 16028
rect 5552 15972 5580 16000
rect 6549 15997 6561 16000
rect 6595 15997 6607 16031
rect 6549 15991 6607 15997
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 15997 7527 16031
rect 7469 15991 7527 15997
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 16028 7803 16031
rect 7834 16028 7840 16040
rect 7791 16000 7840 16028
rect 7791 15997 7803 16000
rect 7745 15991 7803 15997
rect 1486 15969 1492 15972
rect 1480 15923 1492 15969
rect 1486 15920 1492 15923
rect 1544 15920 1550 15972
rect 4372 15963 4430 15969
rect 2608 15932 4292 15960
rect 2608 15904 2636 15932
rect 2590 15852 2596 15904
rect 2648 15852 2654 15904
rect 3234 15852 3240 15904
rect 3292 15852 3298 15904
rect 4264 15892 4292 15932
rect 4372 15929 4384 15963
rect 4418 15960 4430 15963
rect 4614 15960 4620 15972
rect 4418 15932 4620 15960
rect 4418 15929 4430 15932
rect 4372 15923 4430 15929
rect 4614 15920 4620 15932
rect 4672 15920 4678 15972
rect 5534 15920 5540 15972
rect 5592 15920 5598 15972
rect 5626 15920 5632 15972
rect 5684 15960 5690 15972
rect 6641 15963 6699 15969
rect 6641 15960 6653 15963
rect 5684 15932 6653 15960
rect 5684 15920 5690 15932
rect 6641 15929 6653 15932
rect 6687 15929 6699 15963
rect 6641 15923 6699 15929
rect 7484 15904 7512 15991
rect 7668 15960 7696 15991
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 7926 15988 7932 16040
rect 7984 15988 7990 16040
rect 8036 16037 8064 16068
rect 9309 16065 9321 16099
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16096 11299 16099
rect 11422 16096 11428 16108
rect 11287 16068 11428 16096
rect 11287 16065 11299 16068
rect 11241 16059 11299 16065
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 11606 16056 11612 16108
rect 11664 16056 11670 16108
rect 12250 16056 12256 16108
rect 12308 16056 12314 16108
rect 12452 16068 13216 16096
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8202 15988 8208 16040
rect 8260 15988 8266 16040
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 8941 16031 8999 16037
rect 8941 15997 8953 16031
rect 8987 15997 8999 16031
rect 8941 15991 8999 15997
rect 9033 16031 9091 16037
rect 9033 15997 9045 16031
rect 9079 16028 9091 16031
rect 9398 16028 9404 16040
rect 9079 16000 9404 16028
rect 9079 15997 9091 16000
rect 9033 15991 9091 15997
rect 8220 15960 8248 15988
rect 7668 15932 8248 15960
rect 8772 15960 8800 15991
rect 8846 15960 8852 15972
rect 8772 15932 8852 15960
rect 8846 15920 8852 15932
rect 8904 15920 8910 15972
rect 8956 15960 8984 15991
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 12452 16037 12480 16068
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 11020 16000 12449 16028
rect 11020 15988 11026 16000
rect 12437 15997 12449 16000
rect 12483 16028 12495 16031
rect 12483 16000 12537 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12710 15988 12716 16040
rect 12768 15988 12774 16040
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 15997 13139 16031
rect 13081 15991 13139 15997
rect 9306 15960 9312 15972
rect 8956 15932 9312 15960
rect 9306 15920 9312 15932
rect 9364 15920 9370 15972
rect 9576 15963 9634 15969
rect 9576 15929 9588 15963
rect 9622 15960 9634 15963
rect 9674 15960 9680 15972
rect 9622 15932 9680 15960
rect 9622 15929 9634 15932
rect 9576 15923 9634 15929
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 11698 15920 11704 15972
rect 11756 15920 11762 15972
rect 11793 15963 11851 15969
rect 11793 15929 11805 15963
rect 11839 15960 11851 15963
rect 12802 15960 12808 15972
rect 11839 15932 12808 15960
rect 11839 15929 11851 15932
rect 11793 15923 11851 15929
rect 12802 15920 12808 15932
rect 12860 15920 12866 15972
rect 13096 15904 13124 15991
rect 13188 15960 13216 16068
rect 13814 16056 13820 16108
rect 13872 16096 13878 16108
rect 14016 16105 14044 16136
rect 14369 16133 14381 16136
rect 14415 16133 14427 16167
rect 14369 16127 14427 16133
rect 14458 16124 14464 16176
rect 14516 16164 14522 16176
rect 14516 16136 15700 16164
rect 14516 16124 14522 16136
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13872 16068 14013 16096
rect 13872 16056 13878 16068
rect 14001 16065 14013 16068
rect 14047 16065 14059 16099
rect 14001 16059 14059 16065
rect 14185 16099 14243 16105
rect 14185 16065 14197 16099
rect 14231 16096 14243 16099
rect 15010 16096 15016 16108
rect 14231 16068 15016 16096
rect 14231 16065 14243 16068
rect 14185 16059 14243 16065
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 15672 16105 15700 16136
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 13262 15988 13268 16040
rect 13320 15988 13326 16040
rect 13357 16031 13415 16037
rect 13357 15997 13369 16031
rect 13403 16028 13415 16031
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 13403 16000 13921 16028
rect 13403 15997 13415 16000
rect 13357 15991 13415 15997
rect 13909 15997 13921 16000
rect 13955 16028 13967 16031
rect 15286 16028 15292 16040
rect 13955 16000 15292 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 15562 15988 15568 16040
rect 15620 15988 15626 16040
rect 14553 15963 14611 15969
rect 13188 15932 14320 15960
rect 14292 15904 14320 15932
rect 14553 15929 14565 15963
rect 14599 15960 14611 15963
rect 14826 15960 14832 15972
rect 14599 15932 14832 15960
rect 14599 15929 14611 15932
rect 14553 15923 14611 15929
rect 14826 15920 14832 15932
rect 14884 15920 14890 15972
rect 15194 15920 15200 15972
rect 15252 15960 15258 15972
rect 15580 15960 15608 15988
rect 15252 15932 15608 15960
rect 15252 15920 15258 15932
rect 15746 15920 15752 15972
rect 15804 15960 15810 15972
rect 15902 15963 15960 15969
rect 15902 15960 15914 15963
rect 15804 15932 15914 15960
rect 15804 15920 15810 15932
rect 15902 15929 15914 15932
rect 15948 15929 15960 15963
rect 15902 15923 15960 15929
rect 5718 15892 5724 15904
rect 4264 15864 5724 15892
rect 5718 15852 5724 15864
rect 5776 15852 5782 15904
rect 6178 15852 6184 15904
rect 6236 15852 6242 15904
rect 7466 15852 7472 15904
rect 7524 15852 7530 15904
rect 8113 15895 8171 15901
rect 8113 15861 8125 15895
rect 8159 15892 8171 15895
rect 8478 15892 8484 15904
rect 8159 15864 8484 15892
rect 8159 15861 8171 15864
rect 8113 15855 8171 15861
rect 8478 15852 8484 15864
rect 8536 15852 8542 15904
rect 8573 15895 8631 15901
rect 8573 15861 8585 15895
rect 8619 15892 8631 15895
rect 8938 15892 8944 15904
rect 8619 15864 8944 15892
rect 8619 15861 8631 15864
rect 8573 15855 8631 15861
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 10778 15852 10784 15904
rect 10836 15852 10842 15904
rect 12158 15852 12164 15904
rect 12216 15852 12222 15904
rect 12894 15852 12900 15904
rect 12952 15852 12958 15904
rect 13078 15852 13084 15904
rect 13136 15892 13142 15904
rect 13906 15892 13912 15904
rect 13136 15864 13912 15892
rect 13136 15852 13142 15864
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 14274 15852 14280 15904
rect 14332 15852 14338 15904
rect 15105 15895 15163 15901
rect 15105 15861 15117 15895
rect 15151 15892 15163 15895
rect 15470 15892 15476 15904
rect 15151 15864 15476 15892
rect 15151 15861 15163 15864
rect 15105 15855 15163 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 15562 15852 15568 15904
rect 15620 15852 15626 15904
rect 17034 15852 17040 15904
rect 17092 15852 17098 15904
rect 552 15802 17664 15824
rect 552 15750 4366 15802
rect 4418 15750 4430 15802
rect 4482 15750 4494 15802
rect 4546 15750 4558 15802
rect 4610 15750 4622 15802
rect 4674 15750 4686 15802
rect 4738 15750 10366 15802
rect 10418 15750 10430 15802
rect 10482 15750 10494 15802
rect 10546 15750 10558 15802
rect 10610 15750 10622 15802
rect 10674 15750 10686 15802
rect 10738 15750 16366 15802
rect 16418 15750 16430 15802
rect 16482 15750 16494 15802
rect 16546 15750 16558 15802
rect 16610 15750 16622 15802
rect 16674 15750 16686 15802
rect 16738 15750 17664 15802
rect 552 15728 17664 15750
rect 1397 15691 1455 15697
rect 1397 15657 1409 15691
rect 1443 15688 1455 15691
rect 1486 15688 1492 15700
rect 1443 15660 1492 15688
rect 1443 15657 1455 15660
rect 1397 15651 1455 15657
rect 1486 15648 1492 15660
rect 1544 15648 1550 15700
rect 2038 15648 2044 15700
rect 2096 15648 2102 15700
rect 2133 15691 2191 15697
rect 2133 15657 2145 15691
rect 2179 15657 2191 15691
rect 2133 15651 2191 15657
rect 2148 15620 2176 15651
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 2648 15660 3188 15688
rect 2648 15648 2654 15660
rect 2774 15620 2780 15632
rect 1596 15592 2176 15620
rect 2424 15592 2780 15620
rect 1596 15561 1624 15592
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15521 1639 15555
rect 1949 15555 2007 15561
rect 1949 15552 1961 15555
rect 1581 15515 1639 15521
rect 1780 15524 1961 15552
rect 1780 15425 1808 15524
rect 1949 15521 1961 15524
rect 1995 15521 2007 15555
rect 1949 15515 2007 15521
rect 2038 15512 2044 15564
rect 2096 15512 2102 15564
rect 2424 15561 2452 15592
rect 2774 15580 2780 15592
rect 2832 15620 2838 15632
rect 2869 15623 2927 15629
rect 2869 15620 2881 15623
rect 2832 15592 2881 15620
rect 2832 15580 2838 15592
rect 2869 15589 2881 15592
rect 2915 15589 2927 15623
rect 2869 15583 2927 15589
rect 3050 15580 3056 15632
rect 3108 15580 3114 15632
rect 2409 15555 2467 15561
rect 2409 15521 2421 15555
rect 2455 15521 2467 15555
rect 2409 15515 2467 15521
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15484 1915 15487
rect 2056 15484 2084 15512
rect 1903 15456 2084 15484
rect 1903 15453 1915 15456
rect 1857 15447 1915 15453
rect 1765 15419 1823 15425
rect 1765 15385 1777 15419
rect 1811 15416 1823 15419
rect 2501 15419 2559 15425
rect 2501 15416 2513 15419
rect 1811 15388 2513 15416
rect 1811 15385 1823 15388
rect 1765 15379 1823 15385
rect 2501 15385 2513 15388
rect 2547 15416 2559 15419
rect 2682 15416 2688 15428
rect 2547 15388 2688 15416
rect 2547 15385 2559 15388
rect 2501 15379 2559 15385
rect 2682 15376 2688 15388
rect 2740 15376 2746 15428
rect 3068 15425 3096 15580
rect 3160 15561 3188 15660
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 3292 15660 3341 15688
rect 3292 15648 3298 15660
rect 3329 15657 3341 15660
rect 3375 15688 3387 15691
rect 3970 15688 3976 15700
rect 3375 15660 3976 15688
rect 3375 15657 3387 15660
rect 3329 15651 3387 15657
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4890 15648 4896 15700
rect 4948 15688 4954 15700
rect 4948 15660 5396 15688
rect 4948 15648 4954 15660
rect 3804 15592 4200 15620
rect 3804 15561 3832 15592
rect 4172 15564 4200 15592
rect 4614 15580 4620 15632
rect 4672 15620 4678 15632
rect 4982 15620 4988 15632
rect 4672 15592 4988 15620
rect 4672 15580 4678 15592
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 5258 15620 5264 15632
rect 5093 15592 5264 15620
rect 3145 15555 3203 15561
rect 3145 15521 3157 15555
rect 3191 15521 3203 15555
rect 3145 15515 3203 15521
rect 3789 15555 3847 15561
rect 3789 15521 3801 15555
rect 3835 15521 3847 15555
rect 3789 15515 3847 15521
rect 4062 15512 4068 15564
rect 4120 15512 4126 15564
rect 4154 15512 4160 15564
rect 4212 15512 4218 15564
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 5093 15561 5121 15592
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 5368 15620 5396 15660
rect 5810 15648 5816 15700
rect 5868 15688 5874 15700
rect 5997 15691 6055 15697
rect 5997 15688 6009 15691
rect 5868 15660 6009 15688
rect 5868 15648 5874 15660
rect 5997 15657 6009 15660
rect 6043 15688 6055 15691
rect 6270 15688 6276 15700
rect 6043 15660 6276 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 6362 15648 6368 15700
rect 6420 15688 6426 15700
rect 6420 15660 7880 15688
rect 6420 15648 6426 15660
rect 5368 15592 6132 15620
rect 4341 15555 4399 15561
rect 4341 15552 4353 15555
rect 4304 15524 4353 15552
rect 4304 15512 4310 15524
rect 4341 15521 4353 15524
rect 4387 15521 4399 15555
rect 4341 15515 4399 15521
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15521 5135 15555
rect 5077 15515 5135 15521
rect 5169 15555 5227 15561
rect 5169 15521 5181 15555
rect 5215 15521 5227 15555
rect 5169 15515 5227 15521
rect 3878 15444 3884 15496
rect 3936 15484 3942 15496
rect 4985 15487 5043 15493
rect 4985 15484 4997 15487
rect 3936 15456 4997 15484
rect 3936 15444 3942 15456
rect 4985 15453 4997 15456
rect 5031 15453 5043 15487
rect 5184 15484 5212 15515
rect 5350 15512 5356 15564
rect 5408 15552 5414 15564
rect 5445 15555 5503 15561
rect 5445 15552 5457 15555
rect 5408 15524 5457 15552
rect 5408 15512 5414 15524
rect 5445 15521 5457 15524
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 5718 15512 5724 15564
rect 5776 15552 5782 15564
rect 6104 15561 6132 15592
rect 6454 15580 6460 15632
rect 6512 15620 6518 15632
rect 7285 15623 7343 15629
rect 6512 15592 7236 15620
rect 6512 15580 6518 15592
rect 5813 15555 5871 15561
rect 5813 15552 5825 15555
rect 5776 15524 5825 15552
rect 5776 15512 5782 15524
rect 5813 15521 5825 15524
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 6089 15555 6147 15561
rect 6089 15521 6101 15555
rect 6135 15521 6147 15555
rect 6089 15515 6147 15521
rect 4985 15447 5043 15453
rect 5117 15456 5212 15484
rect 5261 15487 5319 15493
rect 3053 15419 3111 15425
rect 3053 15385 3065 15419
rect 3099 15385 3111 15419
rect 3053 15379 3111 15385
rect 3605 15419 3663 15425
rect 3605 15385 3617 15419
rect 3651 15416 3663 15419
rect 3786 15416 3792 15428
rect 3651 15388 3792 15416
rect 3651 15385 3663 15388
rect 3605 15379 3663 15385
rect 3786 15376 3792 15388
rect 3844 15376 3850 15428
rect 5117 15416 5145 15456
rect 5261 15453 5273 15487
rect 5307 15453 5319 15487
rect 5828 15484 5856 15515
rect 6270 15512 6276 15564
rect 6328 15512 6334 15564
rect 7101 15555 7159 15561
rect 7101 15521 7113 15555
rect 7147 15521 7159 15555
rect 7208 15552 7236 15592
rect 7285 15589 7297 15623
rect 7331 15620 7343 15623
rect 7466 15620 7472 15632
rect 7331 15592 7472 15620
rect 7331 15589 7343 15592
rect 7285 15583 7343 15589
rect 7466 15580 7472 15592
rect 7524 15620 7530 15632
rect 7852 15620 7880 15660
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 7984 15660 8033 15688
rect 7984 15648 7990 15660
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 9306 15648 9312 15700
rect 9364 15648 9370 15700
rect 9585 15691 9643 15697
rect 9585 15657 9597 15691
rect 9631 15688 9643 15691
rect 9631 15660 9904 15688
rect 9631 15657 9643 15660
rect 9585 15651 9643 15657
rect 9324 15620 9352 15648
rect 9876 15620 9904 15660
rect 10962 15648 10968 15700
rect 11020 15648 11026 15700
rect 13078 15688 13084 15700
rect 11164 15660 13084 15688
rect 10980 15620 11008 15648
rect 7524 15592 7604 15620
rect 7852 15592 9260 15620
rect 9324 15592 9674 15620
rect 7524 15580 7530 15592
rect 7576 15561 7604 15592
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 7208 15524 7389 15552
rect 7101 15515 7159 15521
rect 7377 15521 7389 15524
rect 7423 15521 7435 15555
rect 7377 15515 7435 15521
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15521 7619 15555
rect 7561 15515 7619 15521
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15552 7803 15555
rect 8754 15552 8760 15564
rect 7791 15524 8760 15552
rect 7791 15521 7803 15524
rect 7745 15515 7803 15521
rect 6638 15484 6644 15496
rect 5828 15456 6644 15484
rect 5261 15447 5319 15453
rect 5276 15416 5304 15447
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15453 6883 15487
rect 7116 15484 7144 15515
rect 7190 15484 7196 15496
rect 7116 15456 7196 15484
rect 6825 15447 6883 15453
rect 5000 15388 5145 15416
rect 5184 15388 5304 15416
rect 6840 15416 6868 15447
rect 7190 15444 7196 15456
rect 7248 15444 7254 15496
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 7668 15484 7696 15515
rect 7340 15456 7696 15484
rect 7340 15444 7346 15456
rect 7760 15416 7788 15515
rect 8754 15512 8760 15524
rect 8812 15512 8818 15564
rect 9232 15561 9260 15592
rect 9217 15555 9275 15561
rect 9217 15521 9229 15555
rect 9263 15552 9275 15555
rect 9401 15555 9459 15561
rect 9401 15552 9413 15555
rect 9263 15524 9413 15552
rect 9263 15521 9275 15524
rect 9217 15515 9275 15521
rect 9401 15521 9413 15524
rect 9447 15521 9459 15555
rect 9646 15552 9674 15592
rect 9876 15592 11008 15620
rect 9876 15561 9904 15592
rect 9861 15555 9919 15561
rect 9646 15524 9812 15552
rect 9401 15515 9459 15521
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9677 15487 9735 15493
rect 9677 15484 9689 15487
rect 9180 15456 9689 15484
rect 9180 15444 9186 15456
rect 9677 15453 9689 15456
rect 9723 15453 9735 15487
rect 9784 15484 9812 15524
rect 9861 15521 9873 15555
rect 9907 15521 9919 15555
rect 9861 15515 9919 15521
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 10100 15524 10149 15552
rect 10100 15512 10106 15524
rect 10137 15521 10149 15524
rect 10183 15521 10195 15555
rect 10137 15515 10195 15521
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 11164 15561 11192 15660
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 13170 15648 13176 15700
rect 13228 15688 13234 15700
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 13228 15660 13277 15688
rect 13228 15648 13234 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 15010 15648 15016 15700
rect 15068 15648 15074 15700
rect 15562 15648 15568 15700
rect 15620 15648 15626 15700
rect 15657 15691 15715 15697
rect 15657 15657 15669 15691
rect 15703 15688 15715 15691
rect 15746 15688 15752 15700
rect 15703 15660 15752 15688
rect 15703 15657 15715 15660
rect 15657 15651 15715 15657
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 16114 15648 16120 15700
rect 16172 15648 16178 15700
rect 17034 15648 17040 15700
rect 17092 15648 17098 15700
rect 11793 15623 11851 15629
rect 11793 15589 11805 15623
rect 11839 15620 11851 15623
rect 11974 15620 11980 15632
rect 11839 15592 11980 15620
rect 11839 15589 11851 15592
rect 11793 15583 11851 15589
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 12158 15580 12164 15632
rect 12216 15620 12222 15632
rect 12216 15592 13584 15620
rect 12216 15580 12222 15592
rect 11149 15555 11207 15561
rect 11149 15552 11161 15555
rect 10284 15524 11161 15552
rect 10284 15512 10290 15524
rect 11149 15521 11161 15524
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 11514 15512 11520 15564
rect 11572 15552 11578 15564
rect 11701 15555 11759 15561
rect 11701 15552 11713 15555
rect 11572 15524 11713 15552
rect 11572 15512 11578 15524
rect 11701 15521 11713 15524
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15552 11943 15555
rect 12342 15552 12348 15564
rect 11931 15524 12348 15552
rect 11931 15521 11943 15524
rect 11885 15515 11943 15521
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 12710 15552 12716 15564
rect 12452 15524 12716 15552
rect 11330 15484 11336 15496
rect 9784 15456 11336 15484
rect 9677 15447 9735 15453
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15484 11483 15487
rect 12452 15484 12480 15524
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 12805 15555 12863 15561
rect 12805 15521 12817 15555
rect 12851 15521 12863 15555
rect 12805 15515 12863 15521
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 13078 15552 13084 15564
rect 12943 15524 13084 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 11471 15456 12480 15484
rect 12529 15487 12587 15493
rect 11471 15453 11483 15456
rect 11425 15447 11483 15453
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 6840 15388 7788 15416
rect 5000 15360 5028 15388
rect 5184 15360 5212 15388
rect 9950 15376 9956 15428
rect 10008 15376 10014 15428
rect 10045 15419 10103 15425
rect 10045 15385 10057 15419
rect 10091 15416 10103 15419
rect 11146 15416 11152 15428
rect 10091 15388 11152 15416
rect 10091 15385 10103 15388
rect 10045 15379 10103 15385
rect 11146 15376 11152 15388
rect 11204 15376 11210 15428
rect 11606 15376 11612 15428
rect 11664 15416 11670 15428
rect 12544 15416 12572 15447
rect 12820 15428 12848 15515
rect 13078 15512 13084 15524
rect 13136 15512 13142 15564
rect 13556 15561 13584 15592
rect 14200 15592 15240 15620
rect 13541 15555 13599 15561
rect 13541 15521 13553 15555
rect 13587 15521 13599 15555
rect 13541 15515 13599 15521
rect 13906 15512 13912 15564
rect 13964 15512 13970 15564
rect 14200 15561 14228 15592
rect 15212 15564 15240 15592
rect 14185 15555 14243 15561
rect 14185 15521 14197 15555
rect 14231 15521 14243 15555
rect 14185 15515 14243 15521
rect 14274 15512 14280 15564
rect 14332 15552 14338 15564
rect 14461 15555 14519 15561
rect 14461 15552 14473 15555
rect 14332 15524 14473 15552
rect 14332 15512 14338 15524
rect 14461 15521 14473 15524
rect 14507 15521 14519 15555
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 14461 15515 14519 15521
rect 14568 15524 14841 15552
rect 14568 15496 14596 15524
rect 14829 15521 14841 15524
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 15194 15512 15200 15564
rect 15252 15512 15258 15564
rect 15473 15555 15531 15561
rect 15473 15521 15485 15555
rect 15519 15552 15531 15555
rect 15580 15552 15608 15648
rect 15519 15524 15608 15552
rect 15933 15555 15991 15561
rect 15519 15521 15531 15524
rect 15473 15515 15531 15521
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 16132 15552 16160 15648
rect 15979 15524 16160 15552
rect 16945 15555 17003 15561
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 16945 15521 16957 15555
rect 16991 15552 17003 15555
rect 17052 15552 17080 15648
rect 17221 15555 17279 15561
rect 17221 15552 17233 15555
rect 16991 15524 17233 15552
rect 16991 15521 17003 15524
rect 16945 15515 17003 15521
rect 17221 15521 17233 15524
rect 17267 15521 17279 15555
rect 17221 15515 17279 15521
rect 12986 15444 12992 15496
rect 13044 15444 13050 15496
rect 14550 15444 14556 15496
rect 14608 15444 14614 15496
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 16022 15484 16028 15496
rect 14783 15456 16028 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 11664 15388 12572 15416
rect 11664 15376 11670 15388
rect 12802 15376 12808 15428
rect 12860 15376 12866 15428
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 13357 15419 13415 15425
rect 13357 15416 13369 15419
rect 13320 15388 13369 15416
rect 13320 15376 13326 15388
rect 13357 15385 13369 15388
rect 13403 15385 13415 15419
rect 13357 15379 13415 15385
rect 13446 15376 13452 15428
rect 13504 15416 13510 15428
rect 13906 15416 13912 15428
rect 13504 15388 13912 15416
rect 13504 15376 13510 15388
rect 13906 15376 13912 15388
rect 13964 15416 13970 15428
rect 14093 15419 14151 15425
rect 14093 15416 14105 15419
rect 13964 15388 14105 15416
rect 13964 15376 13970 15388
rect 14093 15385 14105 15388
rect 14139 15385 14151 15419
rect 14093 15379 14151 15385
rect 14182 15376 14188 15428
rect 14240 15416 14246 15428
rect 14645 15419 14703 15425
rect 14645 15416 14657 15419
rect 14240 15388 14657 15416
rect 14240 15376 14246 15388
rect 14645 15385 14657 15388
rect 14691 15385 14703 15419
rect 14645 15379 14703 15385
rect 15470 15376 15476 15428
rect 15528 15416 15534 15428
rect 17037 15419 17095 15425
rect 17037 15416 17049 15419
rect 15528 15388 17049 15416
rect 15528 15376 15534 15388
rect 2866 15308 2872 15360
rect 2924 15308 2930 15360
rect 3510 15308 3516 15360
rect 3568 15348 3574 15360
rect 3881 15351 3939 15357
rect 3881 15348 3893 15351
rect 3568 15320 3893 15348
rect 3568 15308 3574 15320
rect 3881 15317 3893 15320
rect 3927 15317 3939 15351
rect 3881 15311 3939 15317
rect 4154 15308 4160 15360
rect 4212 15308 4218 15360
rect 4246 15308 4252 15360
rect 4304 15348 4310 15360
rect 4525 15351 4583 15357
rect 4525 15348 4537 15351
rect 4304 15320 4537 15348
rect 4304 15308 4310 15320
rect 4525 15317 4537 15320
rect 4571 15317 4583 15351
rect 4525 15311 4583 15317
rect 4798 15308 4804 15360
rect 4856 15308 4862 15360
rect 4982 15308 4988 15360
rect 5040 15308 5046 15360
rect 5166 15308 5172 15360
rect 5224 15308 5230 15360
rect 5626 15308 5632 15360
rect 5684 15308 5690 15360
rect 6181 15351 6239 15357
rect 6181 15317 6193 15351
rect 6227 15348 6239 15351
rect 6917 15351 6975 15357
rect 6917 15348 6929 15351
rect 6227 15320 6929 15348
rect 6227 15317 6239 15320
rect 6181 15311 6239 15317
rect 6917 15317 6929 15320
rect 6963 15317 6975 15351
rect 6917 15311 6975 15317
rect 7926 15308 7932 15360
rect 7984 15348 7990 15360
rect 8570 15348 8576 15360
rect 7984 15320 8576 15348
rect 7984 15308 7990 15320
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 8846 15308 8852 15360
rect 8904 15348 8910 15360
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 8904 15320 9045 15348
rect 8904 15308 8910 15320
rect 9033 15317 9045 15320
rect 9079 15348 9091 15351
rect 9968 15348 9996 15376
rect 15948 15360 15976 15388
rect 17037 15385 17049 15388
rect 17083 15385 17095 15419
rect 17037 15379 17095 15385
rect 9079 15320 9996 15348
rect 9079 15317 9091 15320
rect 9033 15311 9091 15317
rect 10134 15308 10140 15360
rect 10192 15348 10198 15360
rect 10965 15351 11023 15357
rect 10965 15348 10977 15351
rect 10192 15320 10977 15348
rect 10192 15308 10198 15320
rect 10965 15317 10977 15320
rect 11011 15317 11023 15351
rect 10965 15311 11023 15317
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 12768 15320 12909 15348
rect 12768 15308 12774 15320
rect 12897 15317 12909 15320
rect 12943 15317 12955 15351
rect 12897 15311 12955 15317
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13044 15320 13737 15348
rect 13044 15308 13050 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 15102 15308 15108 15360
rect 15160 15348 15166 15360
rect 15749 15351 15807 15357
rect 15749 15348 15761 15351
rect 15160 15320 15761 15348
rect 15160 15308 15166 15320
rect 15749 15317 15761 15320
rect 15795 15317 15807 15351
rect 15749 15311 15807 15317
rect 15930 15308 15936 15360
rect 15988 15308 15994 15360
rect 16850 15308 16856 15360
rect 16908 15308 16914 15360
rect 552 15258 17664 15280
rect 552 15206 1366 15258
rect 1418 15206 1430 15258
rect 1482 15206 1494 15258
rect 1546 15206 1558 15258
rect 1610 15206 1622 15258
rect 1674 15206 1686 15258
rect 1738 15206 7366 15258
rect 7418 15206 7430 15258
rect 7482 15206 7494 15258
rect 7546 15206 7558 15258
rect 7610 15206 7622 15258
rect 7674 15206 7686 15258
rect 7738 15206 13366 15258
rect 13418 15206 13430 15258
rect 13482 15206 13494 15258
rect 13546 15206 13558 15258
rect 13610 15206 13622 15258
rect 13674 15206 13686 15258
rect 13738 15206 17664 15258
rect 552 15184 17664 15206
rect 2682 15104 2688 15156
rect 2740 15104 2746 15156
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 2958 15144 2964 15156
rect 2915 15116 2964 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 2958 15104 2964 15116
rect 3016 15144 3022 15156
rect 3510 15144 3516 15156
rect 3016 15116 3516 15144
rect 3016 15104 3022 15116
rect 3510 15104 3516 15116
rect 3568 15104 3574 15156
rect 5166 15144 5172 15156
rect 4080 15116 5172 15144
rect 2225 15079 2283 15085
rect 2225 15045 2237 15079
rect 2271 15076 2283 15079
rect 2271 15048 3004 15076
rect 2271 15045 2283 15048
rect 2225 15039 2283 15045
rect 842 14900 848 14952
rect 900 14900 906 14952
rect 1112 14875 1170 14881
rect 1112 14841 1124 14875
rect 1158 14872 1170 14875
rect 1394 14872 1400 14884
rect 1158 14844 1400 14872
rect 1158 14841 1170 14844
rect 1112 14835 1170 14841
rect 1394 14832 1400 14844
rect 1452 14832 1458 14884
rect 2038 14764 2044 14816
rect 2096 14804 2102 14816
rect 2843 14807 2901 14813
rect 2843 14804 2855 14807
rect 2096 14776 2855 14804
rect 2096 14764 2102 14776
rect 2843 14773 2855 14776
rect 2889 14773 2901 14807
rect 2976 14804 3004 15048
rect 3142 15036 3148 15088
rect 3200 15076 3206 15088
rect 3237 15079 3295 15085
rect 3237 15076 3249 15079
rect 3200 15048 3249 15076
rect 3200 15036 3206 15048
rect 3237 15045 3249 15048
rect 3283 15045 3295 15079
rect 3237 15039 3295 15045
rect 3510 14968 3516 15020
rect 3568 14968 3574 15020
rect 4080 15008 4108 15116
rect 5166 15104 5172 15116
rect 5224 15104 5230 15156
rect 5994 15104 6000 15156
rect 6052 15144 6058 15156
rect 6546 15144 6552 15156
rect 6052 15116 6552 15144
rect 6052 15104 6058 15116
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 7561 15147 7619 15153
rect 7561 15113 7573 15147
rect 7607 15144 7619 15147
rect 7650 15144 7656 15156
rect 7607 15116 7656 15144
rect 7607 15113 7619 15116
rect 7561 15107 7619 15113
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 7837 15147 7895 15153
rect 7837 15113 7849 15147
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8251 15116 8340 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 4157 15079 4215 15085
rect 4157 15045 4169 15079
rect 4203 15076 4215 15079
rect 4246 15076 4252 15088
rect 4203 15048 4252 15076
rect 4203 15045 4215 15048
rect 4157 15039 4215 15045
rect 4246 15036 4252 15048
rect 4304 15036 4310 15088
rect 4816 15048 6316 15076
rect 4816 15008 4844 15048
rect 3620 14980 4108 15008
rect 3418 14900 3424 14952
rect 3476 14900 3482 14952
rect 3620 14949 3648 14980
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 3697 14943 3755 14949
rect 3697 14909 3709 14943
rect 3743 14940 3755 14943
rect 3881 14943 3939 14949
rect 3881 14940 3893 14943
rect 3743 14912 3893 14940
rect 3743 14909 3755 14912
rect 3697 14903 3755 14909
rect 3881 14909 3893 14912
rect 3927 14909 3939 14943
rect 3881 14903 3939 14909
rect 3970 14900 3976 14952
rect 4028 14900 4034 14952
rect 4080 14949 4108 14980
rect 4264 14980 4844 15008
rect 4065 14943 4123 14949
rect 4065 14909 4077 14943
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 4264 14949 4292 14980
rect 4890 14968 4896 15020
rect 4948 14968 4954 15020
rect 5102 15011 5160 15017
rect 5102 14977 5114 15011
rect 5148 15008 5160 15011
rect 5534 15008 5540 15020
rect 5148 14980 5540 15008
rect 5148 14977 5160 14980
rect 5102 14971 5160 14977
rect 5534 14968 5540 14980
rect 5592 15008 5598 15020
rect 5629 15011 5687 15017
rect 5629 15008 5641 15011
rect 5592 14980 5641 15008
rect 5592 14968 5598 14980
rect 5629 14977 5641 14980
rect 5675 15008 5687 15011
rect 6086 15008 6092 15020
rect 5675 14980 6092 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 6086 14968 6092 14980
rect 6144 14968 6150 15020
rect 6178 14968 6184 15020
rect 6236 14968 6242 15020
rect 6288 15008 6316 15048
rect 6638 15036 6644 15088
rect 6696 15076 6702 15088
rect 7852 15076 7880 15107
rect 8018 15076 8024 15088
rect 6696 15048 7696 15076
rect 7852 15048 8024 15076
rect 6696 15036 6702 15048
rect 7374 15008 7380 15020
rect 6288 14980 7380 15008
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 4212 14912 4261 14940
rect 4212 14900 4218 14912
rect 4249 14909 4261 14912
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14940 4675 14943
rect 5258 14940 5264 14952
rect 4663 14912 5264 14940
rect 4663 14909 4675 14912
rect 4617 14903 4675 14909
rect 3053 14875 3111 14881
rect 3053 14841 3065 14875
rect 3099 14872 3111 14875
rect 3786 14872 3792 14884
rect 3099 14844 3792 14872
rect 3099 14841 3111 14844
rect 3053 14835 3111 14841
rect 3786 14832 3792 14844
rect 3844 14832 3850 14884
rect 3988 14872 4016 14900
rect 4356 14872 4384 14903
rect 5258 14900 5264 14912
rect 5316 14940 5322 14952
rect 5810 14940 5816 14952
rect 5316 14912 5816 14940
rect 5316 14900 5322 14912
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 5997 14943 6055 14949
rect 5997 14909 6009 14943
rect 6043 14940 6055 14943
rect 6270 14940 6276 14952
rect 6043 14912 6276 14940
rect 6043 14909 6055 14912
rect 5997 14903 6055 14909
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 6546 14900 6552 14952
rect 6604 14940 6610 14952
rect 6730 14940 6736 14952
rect 6604 14912 6736 14940
rect 6604 14900 6610 14912
rect 6730 14900 6736 14912
rect 6788 14940 6794 14952
rect 6914 14940 6920 14952
rect 6788 14912 6920 14940
rect 6788 14900 6794 14912
rect 6914 14900 6920 14912
rect 6972 14940 6978 14952
rect 7668 14949 7696 15048
rect 8018 15036 8024 15048
rect 8076 15036 8082 15088
rect 7009 14943 7067 14949
rect 7009 14940 7021 14943
rect 6972 14912 7021 14940
rect 6972 14900 6978 14912
rect 7009 14909 7021 14912
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 7742 14900 7748 14952
rect 7800 14942 7806 14952
rect 8312 14950 8340 15116
rect 8570 15104 8576 15156
rect 8628 15104 8634 15156
rect 8754 15104 8760 15156
rect 8812 15104 8818 15156
rect 13446 15144 13452 15156
rect 9646 15116 13452 15144
rect 8386 15036 8392 15088
rect 8444 15036 8450 15088
rect 8588 15076 8616 15104
rect 9646 15076 9674 15116
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 13725 15147 13783 15153
rect 13725 15113 13737 15147
rect 13771 15144 13783 15147
rect 13906 15144 13912 15156
rect 13771 15116 13912 15144
rect 13771 15113 13783 15116
rect 13725 15107 13783 15113
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 14645 15147 14703 15153
rect 14645 15113 14657 15147
rect 14691 15144 14703 15147
rect 15010 15144 15016 15156
rect 14691 15116 15016 15144
rect 14691 15113 14703 15116
rect 14645 15107 14703 15113
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 15378 15104 15384 15156
rect 15436 15104 15442 15156
rect 8588 15048 9674 15076
rect 11790 15036 11796 15088
rect 11848 15036 11854 15088
rect 12894 15036 12900 15088
rect 12952 15076 12958 15088
rect 14001 15079 14059 15085
rect 14001 15076 14013 15079
rect 12952 15048 14013 15076
rect 12952 15036 12958 15048
rect 14001 15045 14013 15048
rect 14047 15076 14059 15079
rect 14550 15076 14556 15088
rect 14047 15048 14556 15076
rect 14047 15045 14059 15048
rect 14001 15039 14059 15045
rect 8404 15008 8432 15036
rect 10042 15008 10048 15020
rect 8404 14980 10048 15008
rect 10042 14968 10048 14980
rect 10100 14968 10106 15020
rect 8312 14949 8432 14950
rect 7929 14943 7987 14949
rect 7800 14940 7880 14942
rect 7929 14940 7941 14943
rect 7800 14914 7941 14940
rect 7800 14900 7806 14914
rect 7852 14912 7941 14914
rect 7929 14909 7941 14912
rect 7975 14909 7987 14943
rect 8312 14943 8447 14949
rect 8312 14922 8401 14943
rect 7929 14903 7987 14909
rect 8389 14909 8401 14922
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 8570 14900 8576 14952
rect 8628 14900 8634 14952
rect 8846 14900 8852 14952
rect 8904 14940 8910 14952
rect 9582 14940 9588 14952
rect 8904 14912 9588 14940
rect 8904 14900 8910 14912
rect 9582 14900 9588 14912
rect 9640 14940 9646 14952
rect 11333 14943 11391 14949
rect 9640 14912 11284 14940
rect 9640 14900 9646 14912
rect 3988 14844 4384 14872
rect 5512 14875 5570 14881
rect 5512 14841 5524 14875
rect 5558 14872 5570 14875
rect 6362 14872 6368 14884
rect 5558 14844 6368 14872
rect 5558 14841 5570 14844
rect 5512 14835 5570 14841
rect 6362 14832 6368 14844
rect 6420 14832 6426 14884
rect 7285 14875 7343 14881
rect 7285 14841 7297 14875
rect 7331 14872 7343 14875
rect 8202 14872 8208 14884
rect 7331 14844 8208 14872
rect 7331 14841 7343 14844
rect 7285 14835 7343 14841
rect 8202 14832 8208 14844
rect 8260 14872 8266 14884
rect 8260 14844 9904 14872
rect 8260 14832 8266 14844
rect 9876 14816 9904 14844
rect 3694 14804 3700 14816
rect 2976 14776 3700 14804
rect 2843 14767 2901 14773
rect 3694 14764 3700 14776
rect 3752 14804 3758 14816
rect 4614 14804 4620 14816
rect 3752 14776 4620 14804
rect 3752 14764 3758 14776
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 4982 14764 4988 14816
rect 5040 14764 5046 14816
rect 5258 14764 5264 14816
rect 5316 14764 5322 14816
rect 5350 14764 5356 14816
rect 5408 14764 5414 14816
rect 5721 14807 5779 14813
rect 5721 14773 5733 14807
rect 5767 14804 5779 14807
rect 5994 14804 6000 14816
rect 5767 14776 6000 14804
rect 5767 14773 5779 14776
rect 5721 14767 5779 14773
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6546 14764 6552 14816
rect 6604 14804 6610 14816
rect 6825 14807 6883 14813
rect 6825 14804 6837 14807
rect 6604 14776 6837 14804
rect 6604 14764 6610 14776
rect 6825 14773 6837 14776
rect 6871 14773 6883 14807
rect 6825 14767 6883 14773
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 7156 14776 7205 14804
rect 7156 14764 7162 14776
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7193 14767 7251 14773
rect 7374 14764 7380 14816
rect 7432 14764 7438 14816
rect 9858 14764 9864 14816
rect 9916 14764 9922 14816
rect 11256 14813 11284 14912
rect 11333 14909 11345 14943
rect 11379 14940 11391 14943
rect 11808 14940 11836 15036
rect 14200 15020 14228 15048
rect 14550 15036 14556 15048
rect 14608 15036 14614 15088
rect 14734 15036 14740 15088
rect 14792 15076 14798 15088
rect 15396 15076 15424 15104
rect 14792 15048 15424 15076
rect 14792 15036 14798 15048
rect 13262 14968 13268 15020
rect 13320 14968 13326 15020
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 15841 15011 15899 15017
rect 15841 15008 15853 15011
rect 14424 14980 15853 15008
rect 14424 14968 14430 14980
rect 15841 14977 15853 14980
rect 15887 14977 15899 15011
rect 15841 14971 15899 14977
rect 11379 14912 11836 14940
rect 11379 14909 11391 14912
rect 11333 14903 11391 14909
rect 11882 14900 11888 14952
rect 11940 14940 11946 14952
rect 12250 14940 12256 14952
rect 11940 14912 12256 14940
rect 11940 14900 11946 14912
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 12406 14912 12756 14940
rect 12406 14884 12434 14912
rect 12342 14872 12348 14884
rect 11532 14844 12348 14872
rect 11241 14807 11299 14813
rect 11241 14773 11253 14807
rect 11287 14804 11299 14807
rect 11422 14804 11428 14816
rect 11287 14776 11428 14804
rect 11287 14773 11299 14776
rect 11241 14767 11299 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 11532 14813 11560 14844
rect 12342 14832 12348 14844
rect 12400 14844 12434 14884
rect 12618 14872 12624 14884
rect 12676 14881 12682 14884
rect 12588 14844 12624 14872
rect 12400 14832 12406 14844
rect 12618 14832 12624 14844
rect 12676 14835 12688 14881
rect 12728 14872 12756 14912
rect 12894 14900 12900 14952
rect 12952 14900 12958 14952
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14909 13231 14943
rect 13280 14940 13308 14968
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13280 14912 13553 14940
rect 13173 14903 13231 14909
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 13188 14872 13216 14903
rect 12728 14844 13216 14872
rect 12676 14832 12682 14835
rect 13446 14832 13452 14884
rect 13504 14832 13510 14884
rect 13832 14872 13860 14903
rect 13998 14900 14004 14952
rect 14056 14940 14062 14952
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 14056 14912 14289 14940
rect 14056 14900 14062 14912
rect 14277 14909 14289 14912
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 14550 14900 14556 14952
rect 14608 14900 14614 14952
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 14844 14912 15485 14940
rect 13906 14872 13912 14884
rect 13832 14844 13912 14872
rect 13906 14832 13912 14844
rect 13964 14872 13970 14884
rect 14568 14872 14596 14900
rect 13964 14844 14596 14872
rect 13964 14832 13970 14844
rect 11517 14807 11575 14813
rect 11517 14773 11529 14807
rect 11563 14773 11575 14807
rect 11517 14767 11575 14773
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 12989 14807 13047 14813
rect 12989 14804 13001 14807
rect 11756 14776 13001 14804
rect 11756 14764 11762 14776
rect 12989 14773 13001 14776
rect 13035 14804 13047 14807
rect 13078 14804 13084 14816
rect 13035 14776 13084 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13464 14804 13492 14832
rect 14090 14804 14096 14816
rect 13464 14776 14096 14804
rect 14090 14764 14096 14776
rect 14148 14804 14154 14816
rect 14844 14813 14872 14912
rect 15473 14909 15485 14912
rect 15519 14909 15531 14943
rect 15473 14903 15531 14909
rect 16086 14875 16144 14881
rect 16086 14872 16098 14875
rect 15672 14844 16098 14872
rect 15672 14813 15700 14844
rect 16086 14841 16098 14844
rect 16132 14841 16144 14875
rect 16086 14835 16144 14841
rect 14645 14807 14703 14813
rect 14645 14804 14657 14807
rect 14148 14776 14657 14804
rect 14148 14764 14154 14776
rect 14645 14773 14657 14776
rect 14691 14773 14703 14807
rect 14645 14767 14703 14773
rect 14829 14807 14887 14813
rect 14829 14773 14841 14807
rect 14875 14773 14887 14807
rect 14829 14767 14887 14773
rect 15657 14807 15715 14813
rect 15657 14773 15669 14807
rect 15703 14773 15715 14807
rect 15657 14767 15715 14773
rect 17034 14764 17040 14816
rect 17092 14804 17098 14816
rect 17221 14807 17279 14813
rect 17221 14804 17233 14807
rect 17092 14776 17233 14804
rect 17092 14764 17098 14776
rect 17221 14773 17233 14776
rect 17267 14773 17279 14807
rect 17221 14767 17279 14773
rect 552 14714 17664 14736
rect 552 14662 4366 14714
rect 4418 14662 4430 14714
rect 4482 14662 4494 14714
rect 4546 14662 4558 14714
rect 4610 14662 4622 14714
rect 4674 14662 4686 14714
rect 4738 14662 10366 14714
rect 10418 14662 10430 14714
rect 10482 14662 10494 14714
rect 10546 14662 10558 14714
rect 10610 14662 10622 14714
rect 10674 14662 10686 14714
rect 10738 14662 16366 14714
rect 16418 14662 16430 14714
rect 16482 14662 16494 14714
rect 16546 14662 16558 14714
rect 16610 14662 16622 14714
rect 16674 14662 16686 14714
rect 16738 14662 17664 14714
rect 552 14640 17664 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 1863 14603 1921 14609
rect 1863 14600 1875 14603
rect 1452 14572 1875 14600
rect 1452 14560 1458 14572
rect 1863 14569 1875 14572
rect 1909 14569 1921 14603
rect 1863 14563 1921 14569
rect 2409 14603 2467 14609
rect 2409 14569 2421 14603
rect 2455 14600 2467 14603
rect 2866 14600 2872 14612
rect 2455 14572 2872 14600
rect 2455 14569 2467 14572
rect 2409 14563 2467 14569
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 3568 14572 4261 14600
rect 3568 14560 3574 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 5074 14600 5080 14612
rect 4249 14563 4307 14569
rect 4387 14572 5080 14600
rect 1673 14535 1731 14541
rect 1673 14501 1685 14535
rect 1719 14532 1731 14535
rect 1765 14535 1823 14541
rect 1765 14532 1777 14535
rect 1719 14504 1777 14532
rect 1719 14501 1731 14504
rect 1673 14495 1731 14501
rect 1765 14501 1777 14504
rect 1811 14501 1823 14535
rect 1765 14495 1823 14501
rect 1949 14535 2007 14541
rect 1949 14501 1961 14535
rect 1995 14532 2007 14535
rect 1995 14504 3096 14532
rect 1995 14501 2007 14504
rect 1949 14495 2007 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 1964 14464 1992 14495
rect 1443 14436 1992 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2038 14424 2044 14476
rect 2096 14424 2102 14476
rect 2498 14424 2504 14476
rect 2556 14464 2562 14476
rect 2682 14464 2688 14476
rect 2556 14436 2688 14464
rect 2556 14424 2562 14436
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 2792 14473 2820 14504
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14433 2835 14467
rect 2958 14464 2964 14476
rect 2777 14427 2835 14433
rect 2884 14436 2964 14464
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1762 14396 1768 14408
rect 1719 14368 1768 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 2056 14396 2084 14424
rect 1872 14368 2084 14396
rect 1872 14272 1900 14368
rect 2590 14356 2596 14408
rect 2648 14356 2654 14408
rect 2884 14405 2912 14436
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14365 2927 14399
rect 3068 14396 3096 14504
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 3881 14467 3939 14473
rect 3881 14464 3893 14467
rect 3844 14436 3893 14464
rect 3844 14424 3850 14436
rect 3881 14433 3893 14436
rect 3927 14464 3939 14467
rect 4387 14464 4415 14572
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5316 14572 6960 14600
rect 5316 14560 5322 14572
rect 4522 14492 4528 14544
rect 4580 14492 4586 14544
rect 4985 14535 5043 14541
rect 4985 14501 4997 14535
rect 5031 14532 5043 14535
rect 5092 14532 5120 14560
rect 5031 14504 5120 14532
rect 5353 14535 5411 14541
rect 5031 14501 5043 14504
rect 4985 14495 5043 14501
rect 5353 14501 5365 14535
rect 5399 14532 5411 14535
rect 5534 14532 5540 14544
rect 5399 14504 5540 14532
rect 5399 14501 5411 14504
rect 5353 14495 5411 14501
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 6089 14535 6147 14541
rect 6089 14532 6101 14535
rect 5684 14504 6101 14532
rect 5684 14492 5690 14504
rect 6089 14501 6101 14504
rect 6135 14532 6147 14535
rect 6270 14532 6276 14544
rect 6135 14504 6276 14532
rect 6135 14501 6147 14504
rect 6089 14495 6147 14501
rect 6270 14492 6276 14504
rect 6328 14492 6334 14544
rect 6549 14535 6607 14541
rect 6549 14501 6561 14535
rect 6595 14501 6607 14535
rect 6549 14495 6607 14501
rect 3927 14436 4415 14464
rect 3927 14433 3939 14436
rect 3881 14427 3939 14433
rect 4614 14424 4620 14476
rect 4672 14424 4678 14476
rect 5074 14424 5080 14476
rect 5132 14464 5138 14476
rect 5132 14436 5488 14464
rect 5132 14424 5138 14436
rect 3605 14399 3663 14405
rect 3605 14396 3617 14399
rect 2869 14359 2927 14365
rect 2976 14368 3617 14396
rect 2976 14272 3004 14368
rect 3605 14365 3617 14368
rect 3651 14365 3663 14399
rect 3605 14359 3663 14365
rect 4890 14356 4896 14408
rect 4948 14356 4954 14408
rect 5460 14328 5488 14436
rect 5810 14424 5816 14476
rect 5868 14464 5874 14476
rect 6564 14464 6592 14495
rect 6932 14473 6960 14572
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 7432 14572 7573 14600
rect 7432 14560 7438 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 7561 14563 7619 14569
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 8570 14600 8576 14612
rect 7708 14572 8576 14600
rect 7708 14560 7714 14572
rect 7837 14535 7895 14541
rect 7837 14532 7849 14535
rect 7392 14504 7849 14532
rect 7392 14473 7420 14504
rect 7837 14501 7849 14504
rect 7883 14532 7895 14535
rect 7926 14532 7932 14544
rect 7883 14504 7932 14532
rect 7883 14501 7895 14504
rect 7837 14495 7895 14501
rect 7926 14492 7932 14504
rect 7984 14492 7990 14544
rect 8128 14541 8156 14572
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 8812 14572 9137 14600
rect 8812 14560 8818 14572
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 9125 14563 9183 14569
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 12158 14600 12164 14612
rect 9272 14572 12164 14600
rect 9272 14560 9278 14572
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 12529 14603 12587 14609
rect 12529 14600 12541 14603
rect 12400 14572 12541 14600
rect 12400 14560 12406 14572
rect 12529 14569 12541 14572
rect 12575 14569 12587 14603
rect 12529 14563 12587 14569
rect 13823 14603 13881 14609
rect 13823 14569 13835 14603
rect 13869 14600 13881 14603
rect 13869 14572 14136 14600
rect 13869 14569 13881 14572
rect 13823 14563 13881 14569
rect 8113 14535 8171 14541
rect 8113 14501 8125 14535
rect 8159 14501 8171 14535
rect 8113 14495 8171 14501
rect 8205 14535 8263 14541
rect 8205 14501 8217 14535
rect 8251 14532 8263 14535
rect 8251 14504 9260 14532
rect 8251 14501 8263 14504
rect 8205 14495 8263 14501
rect 5868 14436 6592 14464
rect 6917 14467 6975 14473
rect 5868 14424 5874 14436
rect 6917 14433 6929 14467
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14433 7067 14467
rect 7009 14427 7067 14433
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14433 7435 14467
rect 8294 14464 8300 14476
rect 7377 14427 7435 14433
rect 7484 14436 8300 14464
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14396 6055 14399
rect 6362 14396 6368 14408
rect 6043 14368 6368 14396
rect 6043 14365 6055 14368
rect 5997 14359 6055 14365
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 7024 14396 7052 14427
rect 6880 14368 7052 14396
rect 6880 14356 6886 14368
rect 6549 14331 6607 14337
rect 6549 14328 6561 14331
rect 5460 14300 6561 14328
rect 6549 14297 6561 14300
rect 6595 14328 6607 14331
rect 7484 14328 7512 14436
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8444 14436 8585 14464
rect 8444 14424 8450 14436
rect 8573 14433 8585 14436
rect 8619 14433 8631 14467
rect 8573 14427 8631 14433
rect 8965 14467 9023 14473
rect 8965 14433 8977 14467
rect 9011 14464 9023 14467
rect 9122 14464 9128 14476
rect 9011 14436 9128 14464
rect 9011 14433 9023 14436
rect 8965 14427 9023 14433
rect 9122 14424 9128 14436
rect 9180 14424 9186 14476
rect 8852 14408 8904 14414
rect 8662 14356 8668 14408
rect 8720 14407 8726 14408
rect 8720 14379 8852 14407
rect 8720 14356 8726 14379
rect 8852 14350 8904 14356
rect 6595 14300 7512 14328
rect 9232 14328 9260 14504
rect 10336 14504 11008 14532
rect 9490 14424 9496 14476
rect 9548 14424 9554 14476
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 10336 14473 10364 14504
rect 10321 14467 10379 14473
rect 10321 14464 10333 14467
rect 10008 14436 10333 14464
rect 10008 14424 10014 14436
rect 10321 14433 10333 14436
rect 10367 14433 10379 14467
rect 10321 14427 10379 14433
rect 10594 14424 10600 14476
rect 10652 14424 10658 14476
rect 10980 14473 11008 14504
rect 11882 14492 11888 14544
rect 11940 14492 11946 14544
rect 14108 14532 14136 14572
rect 14522 14535 14580 14541
rect 14522 14532 14534 14535
rect 14108 14504 14534 14532
rect 14522 14501 14534 14504
rect 14568 14501 14580 14535
rect 14522 14495 14580 14501
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 11330 14464 11336 14476
rect 11011 14436 11336 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 11900 14463 11928 14492
rect 12069 14467 12127 14473
rect 11885 14457 11943 14463
rect 11885 14423 11897 14457
rect 11931 14423 11943 14457
rect 12069 14433 12081 14467
rect 12115 14464 12127 14467
rect 12342 14464 12348 14476
rect 12115 14436 12348 14464
rect 12115 14433 12127 14436
rect 12069 14427 12127 14433
rect 12342 14424 12348 14436
rect 12400 14424 12406 14476
rect 12805 14467 12863 14473
rect 12805 14433 12817 14467
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 13725 14467 13783 14473
rect 13725 14433 13737 14467
rect 13771 14464 13783 14467
rect 13814 14464 13820 14476
rect 13771 14436 13820 14464
rect 13771 14433 13783 14436
rect 13725 14427 13783 14433
rect 11885 14417 11943 14423
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14396 10563 14399
rect 10870 14396 10876 14408
rect 10551 14368 10876 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 11606 14396 11612 14408
rect 10980 14368 11612 14396
rect 9677 14331 9735 14337
rect 9677 14328 9689 14331
rect 9232 14300 9689 14328
rect 6595 14297 6607 14300
rect 6549 14291 6607 14297
rect 9677 14297 9689 14300
rect 9723 14328 9735 14331
rect 9766 14328 9772 14340
rect 9723 14300 9772 14328
rect 9723 14297 9735 14300
rect 9677 14291 9735 14297
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 9858 14288 9864 14340
rect 9916 14328 9922 14340
rect 10137 14331 10195 14337
rect 10137 14328 10149 14331
rect 9916 14300 10149 14328
rect 9916 14288 9922 14300
rect 10137 14297 10149 14300
rect 10183 14297 10195 14331
rect 10980 14328 11008 14368
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 12084 14368 12480 14396
rect 12084 14328 12112 14368
rect 10137 14291 10195 14297
rect 10520 14300 11008 14328
rect 11072 14300 12112 14328
rect 12161 14331 12219 14337
rect 1489 14263 1547 14269
rect 1489 14229 1501 14263
rect 1535 14260 1547 14263
rect 1854 14260 1860 14272
rect 1535 14232 1860 14260
rect 1535 14229 1547 14232
rect 1489 14223 1547 14229
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 2958 14220 2964 14272
rect 3016 14220 3022 14272
rect 5534 14220 5540 14272
rect 5592 14220 5598 14272
rect 5810 14220 5816 14272
rect 5868 14220 5874 14272
rect 7377 14263 7435 14269
rect 7377 14229 7389 14263
rect 7423 14260 7435 14263
rect 7834 14260 7840 14272
rect 7423 14232 7840 14260
rect 7423 14229 7435 14232
rect 7377 14223 7435 14229
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 9784 14260 9812 14288
rect 10520 14260 10548 14300
rect 11072 14272 11100 14300
rect 12161 14297 12173 14331
rect 12207 14297 12219 14331
rect 12452 14328 12480 14368
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 12820 14396 12848 14427
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 13906 14424 13912 14476
rect 13964 14424 13970 14476
rect 13998 14424 14004 14476
rect 14056 14424 14062 14476
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14464 14335 14467
rect 14366 14464 14372 14476
rect 14323 14436 14372 14464
rect 14323 14433 14335 14436
rect 14277 14427 14335 14433
rect 12584 14368 12848 14396
rect 12584 14356 12590 14368
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 14292 14396 14320 14427
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 15930 14464 15936 14476
rect 15672 14436 15936 14464
rect 12952 14368 14320 14396
rect 12952 14356 12958 14368
rect 12989 14331 13047 14337
rect 12989 14328 13001 14331
rect 12452 14300 13001 14328
rect 12161 14291 12219 14297
rect 12989 14297 13001 14300
rect 13035 14328 13047 14331
rect 13998 14328 14004 14340
rect 13035 14300 14004 14328
rect 13035 14297 13047 14300
rect 12989 14291 13047 14297
rect 9784 14232 10548 14260
rect 10594 14220 10600 14272
rect 10652 14220 10658 14272
rect 11054 14220 11060 14272
rect 11112 14220 11118 14272
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 11514 14260 11520 14272
rect 11204 14232 11520 14260
rect 11204 14220 11210 14232
rect 11514 14220 11520 14232
rect 11572 14220 11578 14272
rect 11698 14220 11704 14272
rect 11756 14220 11762 14272
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 12176 14260 12204 14291
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 15672 14337 15700 14436
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 15657 14331 15715 14337
rect 15657 14297 15669 14331
rect 15703 14297 15715 14331
rect 15657 14291 15715 14297
rect 15746 14288 15752 14340
rect 15804 14328 15810 14340
rect 16022 14328 16028 14340
rect 15804 14300 16028 14328
rect 15804 14288 15810 14300
rect 16022 14288 16028 14300
rect 16080 14288 16086 14340
rect 11848 14232 12204 14260
rect 11848 14220 11854 14232
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 12529 14263 12587 14269
rect 12529 14260 12541 14263
rect 12492 14232 12541 14260
rect 12492 14220 12498 14232
rect 12529 14229 12541 14232
rect 12575 14229 12587 14263
rect 12529 14223 12587 14229
rect 12710 14220 12716 14272
rect 12768 14220 12774 14272
rect 552 14170 17664 14192
rect 552 14118 1366 14170
rect 1418 14118 1430 14170
rect 1482 14118 1494 14170
rect 1546 14118 1558 14170
rect 1610 14118 1622 14170
rect 1674 14118 1686 14170
rect 1738 14118 7366 14170
rect 7418 14118 7430 14170
rect 7482 14118 7494 14170
rect 7546 14118 7558 14170
rect 7610 14118 7622 14170
rect 7674 14118 7686 14170
rect 7738 14118 13366 14170
rect 13418 14118 13430 14170
rect 13482 14118 13494 14170
rect 13546 14118 13558 14170
rect 13610 14118 13622 14170
rect 13674 14118 13686 14170
rect 13738 14118 17664 14170
rect 552 14096 17664 14118
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 3789 14059 3847 14065
rect 3789 14056 3801 14059
rect 3476 14028 3801 14056
rect 3476 14016 3482 14028
rect 3789 14025 3801 14028
rect 3835 14025 3847 14059
rect 3789 14019 3847 14025
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 4982 14056 4988 14068
rect 4847 14028 4988 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 5350 14016 5356 14068
rect 5408 14016 5414 14068
rect 5810 14056 5816 14068
rect 5552 14028 5816 14056
rect 1854 13948 1860 14000
rect 1912 13988 1918 14000
rect 2593 13991 2651 13997
rect 2593 13988 2605 13991
rect 1912 13960 2605 13988
rect 1912 13948 1918 13960
rect 2593 13957 2605 13960
rect 2639 13957 2651 13991
rect 2593 13951 2651 13957
rect 3620 13960 4660 13988
rect 3620 13932 3648 13960
rect 2498 13880 2504 13932
rect 2556 13920 2562 13932
rect 2961 13923 3019 13929
rect 2961 13920 2973 13923
rect 2556 13892 2973 13920
rect 2556 13880 2562 13892
rect 2961 13889 2973 13892
rect 3007 13889 3019 13923
rect 2961 13883 3019 13889
rect 3602 13880 3608 13932
rect 3660 13880 3666 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 4338 13920 4344 13932
rect 4203 13892 4344 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 2590 13812 2596 13864
rect 2648 13852 2654 13864
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 2648 13824 2789 13852
rect 2648 13812 2654 13824
rect 2777 13821 2789 13824
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 3283 13824 3525 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 3513 13821 3525 13824
rect 3559 13852 3571 13855
rect 3620 13852 3648 13880
rect 3559 13824 3648 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3694 13812 3700 13864
rect 3752 13812 3758 13864
rect 3878 13852 3884 13864
rect 3804 13824 3884 13852
rect 3605 13787 3663 13793
rect 3605 13753 3617 13787
rect 3651 13784 3663 13787
rect 3804 13784 3832 13824
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 3970 13812 3976 13864
rect 4028 13812 4034 13864
rect 4062 13812 4068 13864
rect 4120 13812 4126 13864
rect 4246 13812 4252 13864
rect 4304 13852 4310 13864
rect 4433 13855 4491 13861
rect 4304 13824 4349 13852
rect 4304 13812 4310 13824
rect 4433 13821 4445 13855
rect 4479 13821 4491 13855
rect 4433 13815 4491 13821
rect 3651 13756 3832 13784
rect 3651 13753 3663 13756
rect 3605 13747 3663 13753
rect 3421 13719 3479 13725
rect 3421 13685 3433 13719
rect 3467 13716 3479 13719
rect 4080 13716 4108 13812
rect 4448 13784 4476 13815
rect 4264 13756 4476 13784
rect 4632 13784 4660 13960
rect 5368 13920 5396 14016
rect 5000 13892 5396 13920
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4798 13852 4804 13864
rect 4755 13824 4804 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5000 13861 5028 13892
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13821 5043 13855
rect 4985 13815 5043 13821
rect 5258 13812 5264 13864
rect 5316 13812 5322 13864
rect 5552 13861 5580 14028
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 6638 14016 6644 14068
rect 6696 14016 6702 14068
rect 6822 14016 6828 14068
rect 6880 14016 6886 14068
rect 7190 14016 7196 14068
rect 7248 14016 7254 14068
rect 7377 14059 7435 14065
rect 7377 14025 7389 14059
rect 7423 14025 7435 14059
rect 7377 14019 7435 14025
rect 6454 13988 6460 14000
rect 5920 13960 6460 13988
rect 5920 13920 5948 13960
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 6840 13988 6868 14016
rect 7392 13988 7420 14019
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 9214 14056 9220 14068
rect 8076 14028 9220 14056
rect 8076 14016 8082 14028
rect 8389 13991 8447 13997
rect 8389 13988 8401 13991
rect 6840 13960 7420 13988
rect 8220 13960 8401 13988
rect 8220 13932 8248 13960
rect 8389 13957 8401 13960
rect 8435 13957 8447 13991
rect 8389 13951 8447 13957
rect 5736 13892 5948 13920
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13821 5595 13855
rect 5537 13815 5595 13821
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13852 5687 13855
rect 5736 13852 5764 13892
rect 6086 13880 6092 13932
rect 6144 13920 6150 13932
rect 6181 13923 6239 13929
rect 6181 13920 6193 13923
rect 6144 13892 6193 13920
rect 6144 13880 6150 13892
rect 6181 13889 6193 13892
rect 6227 13889 6239 13923
rect 6181 13883 6239 13889
rect 6288 13892 6960 13920
rect 6288 13864 6316 13892
rect 6270 13852 6276 13864
rect 5675 13824 5764 13852
rect 6231 13824 6276 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 6932 13861 6960 13892
rect 7282 13880 7288 13932
rect 7340 13880 7346 13932
rect 8202 13920 8208 13932
rect 7392 13892 8208 13920
rect 6641 13855 6699 13861
rect 6641 13821 6653 13855
rect 6687 13821 6699 13855
rect 6641 13815 6699 13821
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 7300 13852 7328 13880
rect 7392 13864 7420 13892
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 8754 13920 8760 13932
rect 8352 13892 8760 13920
rect 8352 13880 8358 13892
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 6917 13815 6975 13821
rect 7024 13824 7328 13852
rect 4632 13756 6132 13784
rect 4264 13728 4292 13756
rect 3467 13688 4108 13716
rect 3467 13685 3479 13688
rect 3421 13679 3479 13685
rect 4246 13676 4252 13728
rect 4304 13676 4310 13728
rect 4617 13719 4675 13725
rect 4617 13685 4629 13719
rect 4663 13716 4675 13719
rect 5994 13716 6000 13728
rect 4663 13688 6000 13716
rect 4663 13685 4675 13688
rect 4617 13679 4675 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 6104 13716 6132 13756
rect 6362 13744 6368 13796
rect 6420 13784 6426 13796
rect 6656 13784 6684 13815
rect 6420 13756 6684 13784
rect 6420 13744 6426 13756
rect 6380 13716 6408 13744
rect 6104 13688 6408 13716
rect 6825 13719 6883 13725
rect 6825 13685 6837 13719
rect 6871 13716 6883 13719
rect 7024 13716 7052 13824
rect 7374 13812 7380 13864
rect 7432 13812 7438 13864
rect 7742 13812 7748 13864
rect 7800 13812 7806 13864
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 7926 13852 7932 13864
rect 7883 13824 7932 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 6871 13688 7052 13716
rect 7101 13719 7159 13725
rect 6871 13685 6883 13688
rect 6825 13679 6883 13685
rect 7101 13685 7113 13719
rect 7147 13716 7159 13719
rect 7852 13716 7880 13815
rect 7926 13812 7932 13824
rect 7984 13812 7990 13864
rect 8864 13861 8892 14028
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 10652 14028 11069 14056
rect 10652 14016 10658 14028
rect 11057 14025 11069 14028
rect 11103 14056 11115 14059
rect 11790 14056 11796 14068
rect 11103 14028 11796 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 11790 14016 11796 14028
rect 11848 14056 11854 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11848 14028 11989 14056
rect 11848 14016 11854 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 13633 14059 13691 14065
rect 11977 14019 12035 14025
rect 12084 14028 13584 14056
rect 10689 13991 10747 13997
rect 10689 13957 10701 13991
rect 10735 13988 10747 13991
rect 10962 13988 10968 14000
rect 10735 13960 10968 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 11238 13948 11244 14000
rect 11296 13988 11302 14000
rect 12084 13988 12112 14028
rect 11296 13960 12112 13988
rect 11296 13948 11302 13960
rect 12158 13948 12164 14000
rect 12216 13948 12222 14000
rect 12250 13948 12256 14000
rect 12308 13948 12314 14000
rect 11609 13923 11667 13929
rect 9508 13864 9536 13906
rect 10704 13892 10916 13920
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8404 13824 8585 13852
rect 8404 13784 8432 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 9490 13812 9496 13864
rect 9548 13812 9554 13864
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 9640 13824 9781 13852
rect 9640 13812 9646 13824
rect 9769 13821 9781 13824
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 9122 13784 9128 13796
rect 8404 13756 9128 13784
rect 8404 13728 8432 13756
rect 9122 13744 9128 13756
rect 9180 13744 9186 13796
rect 9674 13744 9680 13796
rect 9732 13744 9738 13796
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10137 13787 10195 13793
rect 10137 13784 10149 13787
rect 10100 13756 10149 13784
rect 10100 13744 10106 13756
rect 10137 13753 10149 13756
rect 10183 13753 10195 13787
rect 10704 13784 10732 13892
rect 10888 13852 10916 13892
rect 11609 13889 11621 13923
rect 11655 13920 11667 13923
rect 12066 13920 12072 13932
rect 11655 13892 12072 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 10888 13824 11836 13852
rect 11054 13793 11060 13796
rect 10137 13747 10195 13753
rect 10520 13756 10732 13784
rect 11041 13787 11060 13793
rect 7147 13688 7880 13716
rect 7147 13685 7159 13688
rect 7101 13679 7159 13685
rect 8386 13676 8392 13728
rect 8444 13676 8450 13728
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 9033 13719 9091 13725
rect 9033 13716 9045 13719
rect 8812 13688 9045 13716
rect 8812 13676 8818 13688
rect 9033 13685 9045 13688
rect 9079 13716 9091 13719
rect 9401 13719 9459 13725
rect 9401 13716 9413 13719
rect 9079 13688 9413 13716
rect 9079 13685 9091 13688
rect 9033 13679 9091 13685
rect 9401 13685 9413 13688
rect 9447 13685 9459 13719
rect 9692 13716 9720 13744
rect 9858 13716 9864 13728
rect 9692 13688 9864 13716
rect 9401 13679 9459 13685
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 10520 13725 10548 13756
rect 11041 13753 11053 13787
rect 11041 13747 11060 13753
rect 11054 13744 11060 13747
rect 11112 13744 11118 13796
rect 11241 13787 11299 13793
rect 11241 13753 11253 13787
rect 11287 13784 11299 13787
rect 11330 13784 11336 13796
rect 11287 13756 11336 13784
rect 11287 13753 11299 13756
rect 11241 13747 11299 13753
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 11425 13787 11483 13793
rect 11425 13753 11437 13787
rect 11471 13784 11483 13787
rect 11606 13784 11612 13796
rect 11471 13756 11612 13784
rect 11471 13753 11483 13756
rect 11425 13747 11483 13753
rect 11606 13744 11612 13756
rect 11664 13744 11670 13796
rect 11808 13784 11836 13824
rect 11882 13812 11888 13864
rect 11940 13812 11946 13864
rect 12176 13861 12204 13948
rect 12268 13861 12296 13948
rect 13556 13929 13584 14028
rect 13633 14025 13645 14059
rect 13679 14056 13691 14059
rect 13722 14056 13728 14068
rect 13679 14028 13728 14056
rect 13679 14025 13691 14028
rect 13633 14019 13691 14025
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14056 13967 14059
rect 14090 14056 14096 14068
rect 13955 14028 14096 14056
rect 13955 14025 13967 14028
rect 13909 14019 13967 14025
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 13998 13988 14004 14000
rect 13740 13960 14004 13988
rect 13740 13929 13768 13960
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 15749 13991 15807 13997
rect 15749 13957 15761 13991
rect 15795 13988 15807 13991
rect 15795 13960 15884 13988
rect 15795 13957 15807 13960
rect 15749 13951 15807 13957
rect 12897 13923 12955 13929
rect 12897 13920 12909 13923
rect 12636 13892 12909 13920
rect 12636 13864 12664 13892
rect 12897 13889 12909 13892
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 13964 13892 14504 13920
rect 13964 13880 13970 13892
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13821 12311 13855
rect 12253 13815 12311 13821
rect 12526 13812 12532 13864
rect 12584 13812 12590 13864
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 13173 13855 13231 13861
rect 13173 13852 13185 13855
rect 12759 13824 13185 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 13173 13821 13185 13824
rect 13219 13852 13231 13855
rect 13817 13855 13875 13861
rect 13219 13824 13768 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13740 13784 13768 13824
rect 13817 13821 13829 13855
rect 13863 13852 13875 13855
rect 13924 13852 13952 13880
rect 13863 13824 13952 13852
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 14366 13812 14372 13864
rect 14424 13812 14430 13864
rect 11808 13756 13032 13784
rect 13740 13756 13952 13784
rect 10505 13719 10563 13725
rect 10505 13716 10517 13719
rect 10284 13688 10517 13716
rect 10284 13676 10290 13688
rect 10505 13685 10517 13688
rect 10551 13685 10563 13719
rect 10505 13679 10563 13685
rect 10594 13676 10600 13728
rect 10652 13716 10658 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10652 13688 10885 13716
rect 10652 13676 10658 13688
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 11348 13716 11376 13744
rect 11701 13719 11759 13725
rect 11701 13716 11713 13719
rect 11348 13688 11713 13716
rect 10873 13679 10931 13685
rect 11701 13685 11713 13688
rect 11747 13685 11759 13719
rect 11701 13679 11759 13685
rect 12434 13676 12440 13728
rect 12492 13676 12498 13728
rect 13004 13725 13032 13756
rect 12989 13719 13047 13725
rect 12989 13685 13001 13719
rect 13035 13716 13047 13719
rect 13814 13716 13820 13728
rect 13035 13688 13820 13716
rect 13035 13685 13047 13688
rect 12989 13679 13047 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 13924 13716 13952 13756
rect 14090 13744 14096 13796
rect 14148 13744 14154 13796
rect 14277 13787 14335 13793
rect 14277 13753 14289 13787
rect 14323 13753 14335 13787
rect 14476 13784 14504 13892
rect 14636 13855 14694 13861
rect 14636 13821 14648 13855
rect 14682 13852 14694 13855
rect 15746 13852 15752 13864
rect 14682 13824 15752 13852
rect 14682 13821 14694 13824
rect 14636 13815 14694 13821
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 15856 13852 15884 13960
rect 15930 13948 15936 14000
rect 15988 13948 15994 14000
rect 16669 13991 16727 13997
rect 16669 13988 16681 13991
rect 16224 13960 16681 13988
rect 15948 13920 15976 13948
rect 16224 13932 16252 13960
rect 16669 13957 16681 13960
rect 16715 13988 16727 13991
rect 17126 13988 17132 14000
rect 16715 13960 17132 13988
rect 16715 13957 16727 13960
rect 16669 13951 16727 13957
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15948 13892 16129 13920
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16206 13880 16212 13932
rect 16264 13880 16270 13932
rect 16390 13880 16396 13932
rect 16448 13880 16454 13932
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 15856 13824 16037 13852
rect 16025 13821 16037 13824
rect 16071 13852 16083 13855
rect 16758 13852 16764 13864
rect 16071 13824 16764 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 16758 13812 16764 13824
rect 16816 13812 16822 13864
rect 16850 13812 16856 13864
rect 16908 13812 16914 13864
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 17052 13824 17141 13852
rect 17052 13796 17080 13824
rect 17129 13821 17141 13824
rect 17175 13821 17187 13855
rect 17129 13815 17187 13821
rect 14734 13784 14740 13796
rect 14476 13756 14740 13784
rect 14277 13747 14335 13753
rect 14292 13716 14320 13747
rect 14734 13744 14740 13756
rect 14792 13744 14798 13796
rect 17034 13744 17040 13796
rect 17092 13744 17098 13796
rect 16945 13719 17003 13725
rect 16945 13716 16957 13719
rect 13924 13688 16957 13716
rect 16945 13685 16957 13688
rect 16991 13716 17003 13719
rect 17402 13716 17408 13728
rect 16991 13688 17408 13716
rect 16991 13685 17003 13688
rect 16945 13679 17003 13685
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 552 13626 17664 13648
rect 552 13574 4366 13626
rect 4418 13574 4430 13626
rect 4482 13574 4494 13626
rect 4546 13574 4558 13626
rect 4610 13574 4622 13626
rect 4674 13574 4686 13626
rect 4738 13574 10366 13626
rect 10418 13574 10430 13626
rect 10482 13574 10494 13626
rect 10546 13574 10558 13626
rect 10610 13574 10622 13626
rect 10674 13574 10686 13626
rect 10738 13574 16366 13626
rect 16418 13574 16430 13626
rect 16482 13574 16494 13626
rect 16546 13574 16558 13626
rect 16610 13574 16622 13626
rect 16674 13574 16686 13626
rect 16738 13574 17664 13626
rect 552 13552 17664 13574
rect 2130 13472 2136 13524
rect 2188 13512 2194 13524
rect 3329 13515 3387 13521
rect 2188 13484 3096 13512
rect 2188 13472 2194 13484
rect 2590 13404 2596 13456
rect 2648 13404 2654 13456
rect 3068 13453 3096 13484
rect 3329 13481 3341 13515
rect 3375 13512 3387 13515
rect 3510 13512 3516 13524
rect 3375 13484 3516 13512
rect 3375 13481 3387 13484
rect 3329 13475 3387 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 3602 13472 3608 13524
rect 3660 13472 3666 13524
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 3970 13512 3976 13524
rect 3927 13484 3976 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 4338 13472 4344 13524
rect 4396 13472 4402 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5644 13484 5825 13512
rect 2853 13447 2911 13453
rect 2853 13413 2865 13447
rect 2899 13444 2911 13447
rect 3053 13447 3111 13453
rect 2899 13413 2912 13444
rect 2853 13407 2912 13413
rect 3053 13413 3065 13447
rect 3099 13413 3111 13447
rect 4249 13447 4307 13453
rect 4249 13444 4261 13447
rect 3053 13407 3111 13413
rect 3712 13416 4261 13444
rect 1210 13385 1216 13388
rect 1204 13339 1216 13385
rect 1210 13336 1216 13339
rect 1268 13336 1274 13388
rect 2608 13369 2636 13404
rect 2593 13363 2651 13369
rect 2593 13329 2605 13363
rect 2639 13329 2651 13363
rect 2593 13323 2651 13329
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 937 13311 995 13317
rect 937 13308 949 13311
rect 900 13280 949 13308
rect 900 13268 906 13280
rect 937 13277 949 13280
rect 983 13277 995 13311
rect 937 13271 995 13277
rect 2884 13240 2912 13407
rect 3068 13376 3096 13407
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 3068 13348 3157 13376
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13345 3479 13379
rect 3421 13339 3479 13345
rect 3436 13240 3464 13339
rect 2332 13212 3464 13240
rect 2332 13184 2360 13212
rect 2314 13132 2320 13184
rect 2372 13132 2378 13184
rect 2406 13132 2412 13184
rect 2464 13132 2470 13184
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 2685 13175 2743 13181
rect 2685 13172 2697 13175
rect 2556 13144 2697 13172
rect 2556 13132 2562 13144
rect 2685 13141 2697 13144
rect 2731 13141 2743 13175
rect 2685 13135 2743 13141
rect 2869 13175 2927 13181
rect 2869 13141 2881 13175
rect 2915 13172 2927 13175
rect 3234 13172 3240 13184
rect 2915 13144 3240 13172
rect 2915 13141 2927 13144
rect 2869 13135 2927 13141
rect 3234 13132 3240 13144
rect 3292 13172 3298 13184
rect 3712 13172 3740 13416
rect 4249 13413 4261 13416
rect 4295 13444 4307 13447
rect 4356 13444 4384 13472
rect 4295 13416 4384 13444
rect 4295 13413 4307 13416
rect 4249 13407 4307 13413
rect 5644 13388 5672 13484
rect 5813 13481 5825 13484
rect 5859 13512 5871 13515
rect 5859 13484 6684 13512
rect 5859 13481 5871 13484
rect 5813 13475 5871 13481
rect 6362 13404 6368 13456
rect 6420 13444 6426 13456
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 6420 13416 6561 13444
rect 6420 13404 6426 13416
rect 6549 13413 6561 13416
rect 6595 13413 6607 13447
rect 6656 13444 6684 13484
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7650 13512 7656 13524
rect 6972 13484 7656 13512
rect 6972 13472 6978 13484
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 9180 13484 9505 13512
rect 9180 13472 9186 13484
rect 9493 13481 9505 13484
rect 9539 13481 9551 13515
rect 9493 13475 9551 13481
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 10042 13512 10048 13524
rect 9723 13484 10048 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10689 13515 10747 13521
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 10870 13512 10876 13524
rect 10735 13484 10876 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 12124 13484 12756 13512
rect 12124 13472 12130 13484
rect 6822 13444 6828 13456
rect 6656 13416 6828 13444
rect 6549 13407 6607 13413
rect 6822 13404 6828 13416
rect 6880 13404 6886 13456
rect 7285 13447 7343 13453
rect 7285 13413 7297 13447
rect 7331 13444 7343 13447
rect 7374 13444 7380 13456
rect 7331 13416 7380 13444
rect 7331 13413 7343 13416
rect 7285 13407 7343 13413
rect 7374 13404 7380 13416
rect 7432 13404 7438 13456
rect 7926 13404 7932 13456
rect 7984 13444 7990 13456
rect 8205 13447 8263 13453
rect 7984 13416 8156 13444
rect 7984 13404 7990 13416
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 4080 13308 4108 13339
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4396 13348 4537 13376
rect 4396 13336 4402 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 4614 13336 4620 13388
rect 4672 13336 4678 13388
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 4948 13348 5488 13376
rect 4948 13336 4954 13348
rect 4632 13308 4660 13336
rect 4080 13280 4660 13308
rect 5350 13268 5356 13320
rect 5408 13268 5414 13320
rect 5460 13308 5488 13348
rect 5626 13336 5632 13388
rect 5684 13336 5690 13388
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6086 13376 6092 13388
rect 6043 13348 6092 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6914 13376 6920 13388
rect 6196 13348 6920 13376
rect 6196 13308 6224 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 8128 13376 8156 13416
rect 8205 13413 8217 13447
rect 8251 13444 8263 13447
rect 8386 13444 8392 13456
rect 8251 13416 8392 13444
rect 8251 13413 8263 13416
rect 8205 13407 8263 13413
rect 8386 13404 8392 13416
rect 8444 13404 8450 13456
rect 9309 13447 9367 13453
rect 9309 13413 9321 13447
rect 9355 13444 9367 13447
rect 9355 13416 9444 13444
rect 9355 13413 9367 13416
rect 9309 13407 9367 13413
rect 9416 13388 9444 13416
rect 9582 13404 9588 13456
rect 9640 13444 9646 13456
rect 10226 13444 10232 13456
rect 9640 13416 10088 13444
rect 9640 13404 9646 13416
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8128 13348 8493 13376
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 8570 13336 8576 13388
rect 8628 13336 8634 13388
rect 8662 13336 8668 13388
rect 8720 13376 8726 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8720 13348 8953 13376
rect 8720 13336 8726 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13345 9919 13379
rect 9861 13339 9919 13345
rect 7834 13308 7840 13320
rect 5460 13280 6224 13308
rect 7590 13280 7840 13308
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 9766 13308 9772 13320
rect 9246 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 4982 13200 4988 13252
rect 5040 13240 5046 13252
rect 5718 13240 5724 13252
rect 5040 13212 5724 13240
rect 5040 13200 5046 13212
rect 5718 13200 5724 13212
rect 5776 13200 5782 13252
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 9876 13240 9904 13339
rect 10060 13317 10088 13416
rect 10152 13416 10232 13444
rect 10152 13385 10180 13416
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 12618 13444 12624 13456
rect 10520 13416 12624 13444
rect 10520 13385 10548 13416
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 12728 13444 12756 13484
rect 12802 13472 12808 13524
rect 12860 13472 12866 13524
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 13078 13512 13084 13524
rect 12952 13484 13084 13512
rect 12952 13472 12958 13484
rect 13078 13472 13084 13484
rect 13136 13472 13142 13524
rect 13280 13484 13768 13512
rect 13280 13444 13308 13484
rect 12728 13416 13308 13444
rect 13354 13404 13360 13456
rect 13412 13404 13418 13456
rect 13740 13453 13768 13484
rect 15746 13472 15752 13524
rect 15804 13472 15810 13524
rect 16853 13515 16911 13521
rect 16853 13481 16865 13515
rect 16899 13481 16911 13515
rect 16853 13475 16911 13481
rect 13725 13447 13783 13453
rect 13725 13413 13737 13447
rect 13771 13413 13783 13447
rect 13725 13407 13783 13413
rect 13998 13404 14004 13456
rect 14056 13444 14062 13456
rect 14461 13447 14519 13453
rect 14461 13444 14473 13447
rect 14056 13416 14473 13444
rect 14056 13404 14062 13416
rect 14461 13413 14473 13416
rect 14507 13444 14519 13447
rect 16868 13444 16896 13475
rect 17126 13472 17132 13524
rect 17184 13472 17190 13524
rect 14507 13416 16896 13444
rect 14507 13413 14519 13416
rect 14461 13407 14519 13413
rect 15580 13388 15608 13416
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10505 13379 10563 13385
rect 10505 13345 10517 13379
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 10594 13336 10600 13388
rect 10652 13376 10658 13388
rect 11149 13379 11207 13385
rect 11149 13376 11161 13379
rect 10652 13348 11161 13376
rect 10652 13336 10658 13348
rect 11149 13345 11161 13348
rect 11195 13345 11207 13379
rect 11149 13339 11207 13345
rect 11330 13336 11336 13388
rect 11388 13336 11394 13388
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 12158 13376 12164 13388
rect 11572 13348 12164 13376
rect 11572 13336 11578 13348
rect 12158 13336 12164 13348
rect 12216 13376 12222 13388
rect 13096 13376 13308 13382
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 12216 13354 13645 13376
rect 12216 13348 13124 13354
rect 13280 13348 13645 13354
rect 12216 13336 12222 13348
rect 13633 13345 13645 13348
rect 13679 13345 13691 13379
rect 13633 13339 13691 13345
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 13872 13348 14105 13376
rect 13872 13336 13878 13348
rect 14093 13345 14105 13348
rect 14139 13376 14151 13379
rect 14918 13376 14924 13388
rect 14139 13348 14924 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 15562 13336 15568 13388
rect 15620 13336 15626 13388
rect 15930 13336 15936 13388
rect 15988 13336 15994 13388
rect 16022 13336 16028 13388
rect 16080 13376 16086 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 16080 13348 16313 13376
rect 16080 13336 16086 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 16390 13336 16396 13388
rect 16448 13376 16454 13388
rect 16448 13348 16620 13376
rect 16448 13336 16454 13348
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 10336 13280 11100 13308
rect 10336 13252 10364 13280
rect 10226 13240 10232 13252
rect 9732 13212 10232 13240
rect 9732 13200 9738 13212
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 10318 13200 10324 13252
rect 10376 13200 10382 13252
rect 10965 13243 11023 13249
rect 10965 13240 10977 13243
rect 10704 13212 10977 13240
rect 10704 13184 10732 13212
rect 10965 13209 10977 13212
rect 11011 13209 11023 13243
rect 10965 13203 11023 13209
rect 3292 13144 3740 13172
rect 4709 13175 4767 13181
rect 3292 13132 3298 13144
rect 4709 13141 4721 13175
rect 4755 13172 4767 13175
rect 5166 13172 5172 13184
rect 4755 13144 5172 13172
rect 4755 13141 4767 13144
rect 4709 13135 4767 13141
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 7837 13175 7895 13181
rect 7837 13141 7849 13175
rect 7883 13172 7895 13175
rect 7926 13172 7932 13184
rect 7883 13144 7932 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 9858 13132 9864 13184
rect 9916 13172 9922 13184
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9916 13144 10425 13172
rect 9916 13132 9922 13144
rect 10413 13141 10425 13144
rect 10459 13172 10471 13175
rect 10594 13172 10600 13184
rect 10459 13144 10600 13172
rect 10459 13141 10471 13144
rect 10413 13135 10471 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 10686 13132 10692 13184
rect 10744 13132 10750 13184
rect 11072 13172 11100 13280
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11480 13280 13202 13308
rect 11480 13268 11486 13280
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 14829 13311 14887 13317
rect 14829 13308 14841 13311
rect 14608 13280 14841 13308
rect 14608 13268 14614 13280
rect 14829 13277 14841 13280
rect 14875 13277 14887 13311
rect 14829 13271 14887 13277
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13277 16543 13311
rect 16592 13308 16620 13348
rect 16758 13336 16764 13388
rect 16816 13336 16822 13388
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13376 17095 13379
rect 17144 13376 17172 13472
rect 17083 13348 17172 13376
rect 17313 13379 17371 13385
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 17313 13345 17325 13379
rect 17359 13345 17371 13379
rect 17313 13339 17371 13345
rect 17328 13308 17356 13339
rect 16592 13280 17356 13308
rect 16485 13271 16543 13277
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 15120 13240 15148 13271
rect 14792 13212 15148 13240
rect 14792 13200 14798 13212
rect 15286 13200 15292 13252
rect 15344 13240 15350 13252
rect 16500 13240 16528 13271
rect 16577 13243 16635 13249
rect 16577 13240 16589 13243
rect 15344 13212 16589 13240
rect 15344 13200 15350 13212
rect 16577 13209 16589 13212
rect 16623 13209 16635 13243
rect 16577 13203 16635 13209
rect 13170 13172 13176 13184
rect 11072 13144 13176 13172
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 14645 13175 14703 13181
rect 14645 13141 14657 13175
rect 14691 13172 14703 13175
rect 15378 13172 15384 13184
rect 14691 13144 15384 13172
rect 14691 13141 14703 13144
rect 14645 13135 14703 13141
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15746 13132 15752 13184
rect 15804 13172 15810 13184
rect 16117 13175 16175 13181
rect 16117 13172 16129 13175
rect 15804 13144 16129 13172
rect 15804 13132 15810 13144
rect 16117 13141 16129 13144
rect 16163 13141 16175 13175
rect 16117 13135 16175 13141
rect 17126 13132 17132 13184
rect 17184 13132 17190 13184
rect 552 13082 17664 13104
rect 552 13030 1366 13082
rect 1418 13030 1430 13082
rect 1482 13030 1494 13082
rect 1546 13030 1558 13082
rect 1610 13030 1622 13082
rect 1674 13030 1686 13082
rect 1738 13030 7366 13082
rect 7418 13030 7430 13082
rect 7482 13030 7494 13082
rect 7546 13030 7558 13082
rect 7610 13030 7622 13082
rect 7674 13030 7686 13082
rect 7738 13030 13366 13082
rect 13418 13030 13430 13082
rect 13482 13030 13494 13082
rect 13546 13030 13558 13082
rect 13610 13030 13622 13082
rect 13674 13030 13686 13082
rect 13738 13030 17664 13082
rect 552 13008 17664 13030
rect 1210 12928 1216 12980
rect 1268 12968 1274 12980
rect 1305 12971 1363 12977
rect 1305 12968 1317 12971
rect 1268 12940 1317 12968
rect 1268 12928 1274 12940
rect 1305 12937 1317 12940
rect 1351 12937 1363 12971
rect 1305 12931 1363 12937
rect 1762 12928 1768 12980
rect 1820 12928 1826 12980
rect 2866 12928 2872 12980
rect 2924 12928 2930 12980
rect 5350 12968 5356 12980
rect 3252 12940 5356 12968
rect 1670 12900 1676 12912
rect 1504 12872 1676 12900
rect 1504 12773 1532 12872
rect 1670 12860 1676 12872
rect 1728 12860 1734 12912
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 1780 12832 1808 12928
rect 3252 12832 3280 12940
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5902 12928 5908 12980
rect 5960 12968 5966 12980
rect 6089 12971 6147 12977
rect 6089 12968 6101 12971
rect 5960 12940 6101 12968
rect 5960 12928 5966 12940
rect 6089 12937 6101 12940
rect 6135 12937 6147 12971
rect 6089 12931 6147 12937
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7101 12971 7159 12977
rect 7101 12968 7113 12971
rect 7064 12940 7113 12968
rect 7064 12928 7070 12940
rect 7101 12937 7113 12940
rect 7147 12937 7159 12971
rect 7101 12931 7159 12937
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 9490 12968 9496 12980
rect 8444 12940 9496 12968
rect 8444 12928 8450 12940
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 9674 12928 9680 12980
rect 9732 12928 9738 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11440 12940 11989 12968
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 9692 12900 9720 12928
rect 4672 12872 6802 12900
rect 4672 12860 4678 12872
rect 1627 12804 1808 12832
rect 1872 12804 3280 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 1305 12767 1363 12773
rect 1305 12733 1317 12767
rect 1351 12733 1363 12767
rect 1305 12727 1363 12733
rect 1489 12767 1547 12773
rect 1489 12733 1501 12767
rect 1535 12733 1547 12767
rect 1489 12727 1547 12733
rect 1320 12696 1348 12727
rect 1581 12699 1639 12705
rect 1581 12696 1593 12699
rect 1320 12668 1593 12696
rect 1581 12665 1593 12668
rect 1627 12665 1639 12699
rect 1688 12696 1716 12804
rect 1762 12724 1768 12776
rect 1820 12724 1826 12776
rect 1872 12773 1900 12804
rect 5166 12792 5172 12844
rect 5224 12792 5230 12844
rect 6546 12792 6552 12844
rect 6604 12792 6610 12844
rect 6638 12792 6644 12844
rect 6696 12792 6702 12844
rect 6774 12832 6802 12872
rect 9646 12872 9720 12900
rect 9646 12832 9674 12872
rect 6774 12804 9674 12832
rect 9772 12844 9824 12850
rect 11440 12844 11468 12940
rect 11977 12937 11989 12940
rect 12023 12968 12035 12971
rect 12023 12940 12940 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 11790 12860 11796 12912
rect 11848 12860 11854 12912
rect 11885 12903 11943 12909
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 11931 12872 12664 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 11422 12792 11428 12844
rect 11480 12792 11486 12844
rect 9772 12786 9824 12792
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12733 1915 12767
rect 1857 12727 1915 12733
rect 1946 12724 1952 12776
rect 2004 12764 2010 12776
rect 2406 12764 2412 12776
rect 2004 12736 2412 12764
rect 2004 12724 2010 12736
rect 2406 12724 2412 12736
rect 2464 12764 2470 12776
rect 2501 12767 2559 12773
rect 2501 12764 2513 12767
rect 2464 12736 2513 12764
rect 2464 12724 2470 12736
rect 2501 12733 2513 12736
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 3283 12736 3648 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 3620 12708 3648 12736
rect 5074 12724 5080 12776
rect 5132 12724 5138 12776
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12733 5503 12767
rect 5445 12727 5503 12733
rect 2590 12696 2596 12708
rect 1688 12668 2596 12696
rect 1581 12659 1639 12665
rect 2590 12656 2596 12668
rect 2648 12696 2654 12708
rect 3510 12705 3516 12708
rect 2648 12668 3464 12696
rect 2648 12656 2654 12668
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2832 12600 2881 12628
rect 2832 12588 2838 12600
rect 2869 12597 2881 12600
rect 2915 12628 2927 12631
rect 2958 12628 2964 12640
rect 2915 12600 2964 12628
rect 2915 12597 2927 12600
rect 2869 12591 2927 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 3050 12588 3056 12640
rect 3108 12588 3114 12640
rect 3436 12628 3464 12668
rect 3504 12659 3516 12705
rect 3510 12656 3516 12659
rect 3568 12656 3574 12708
rect 3602 12656 3608 12708
rect 3660 12656 3666 12708
rect 4154 12656 4160 12708
rect 4212 12656 4218 12708
rect 4172 12628 4200 12656
rect 3436 12600 4200 12628
rect 4890 12588 4896 12640
rect 4948 12588 4954 12640
rect 5460 12628 5488 12727
rect 6270 12724 6276 12776
rect 6328 12764 6334 12776
rect 6457 12767 6515 12773
rect 6457 12764 6469 12767
rect 6328 12736 6469 12764
rect 6328 12724 6334 12736
rect 6457 12733 6469 12736
rect 6503 12733 6515 12767
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6457 12727 6515 12733
rect 6656 12736 6929 12764
rect 6178 12656 6184 12708
rect 6236 12696 6242 12708
rect 6656 12696 6684 12736
rect 6917 12733 6929 12736
rect 6963 12764 6975 12767
rect 7098 12764 7104 12776
rect 6963 12736 7104 12764
rect 6963 12733 6975 12736
rect 6917 12727 6975 12733
rect 7098 12724 7104 12736
rect 7156 12764 7162 12776
rect 8386 12764 8392 12776
rect 7156 12736 8392 12764
rect 7156 12724 7162 12736
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 9582 12724 9588 12776
rect 9640 12764 9646 12776
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 9640 12736 9689 12764
rect 9640 12724 9646 12736
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 10686 12764 10692 12776
rect 9677 12727 9735 12733
rect 9876 12736 10692 12764
rect 6236 12668 6684 12696
rect 6236 12656 6242 12668
rect 6730 12656 6736 12708
rect 6788 12656 6794 12708
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 8294 12696 8300 12708
rect 6880 12668 8300 12696
rect 6880 12656 6886 12668
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 8573 12699 8631 12705
rect 8573 12696 8585 12699
rect 8404 12668 8585 12696
rect 6748 12628 6776 12656
rect 7006 12628 7012 12640
rect 5460 12600 7012 12628
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 8404 12628 8432 12668
rect 8573 12665 8585 12668
rect 8619 12696 8631 12699
rect 9398 12696 9404 12708
rect 8619 12668 9404 12696
rect 8619 12665 8631 12668
rect 8573 12659 8631 12665
rect 9398 12656 9404 12668
rect 9456 12696 9462 12708
rect 9876 12696 9904 12736
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 11081 12767 11139 12773
rect 11081 12733 11093 12767
rect 11127 12764 11139 12767
rect 11701 12767 11759 12773
rect 11701 12764 11713 12767
rect 11127 12736 11713 12764
rect 11127 12733 11139 12736
rect 11081 12727 11139 12733
rect 11701 12733 11713 12736
rect 11747 12764 11759 12767
rect 11808 12764 11836 12860
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 12158 12792 12164 12844
rect 12216 12792 12222 12844
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12832 12495 12835
rect 12526 12832 12532 12844
rect 12483 12804 12532 12832
rect 12483 12801 12495 12804
rect 12437 12795 12495 12801
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 11747 12736 11836 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 9456 12668 9904 12696
rect 9456 12656 9462 12668
rect 9950 12656 9956 12708
rect 10008 12656 10014 12708
rect 10229 12699 10287 12705
rect 10229 12665 10241 12699
rect 10275 12665 10287 12699
rect 10229 12659 10287 12665
rect 7892 12600 8432 12628
rect 8481 12631 8539 12637
rect 7892 12588 7898 12600
rect 8481 12597 8493 12631
rect 8527 12628 8539 12631
rect 8662 12628 8668 12640
rect 8527 12600 8668 12628
rect 8527 12597 8539 12600
rect 8481 12591 8539 12597
rect 8662 12588 8668 12600
rect 8720 12628 8726 12640
rect 9122 12628 9128 12640
rect 8720 12600 9128 12628
rect 8720 12588 8726 12600
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 10244 12628 10272 12659
rect 10318 12656 10324 12708
rect 10376 12656 10382 12708
rect 10870 12656 10876 12708
rect 10928 12696 10934 12708
rect 11992 12696 12020 12792
rect 12176 12749 12204 12792
rect 12636 12776 12664 12872
rect 12802 12792 12808 12844
rect 12860 12792 12866 12844
rect 12912 12841 12940 12940
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 14550 12968 14556 12980
rect 13320 12940 14556 12968
rect 13320 12928 13326 12940
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 16850 12928 16856 12980
rect 16908 12968 16914 12980
rect 17218 12968 17224 12980
rect 16908 12940 17224 12968
rect 16908 12928 16914 12940
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 12897 12795 12955 12801
rect 13004 12804 15117 12832
rect 12161 12743 12219 12749
rect 12161 12709 12173 12743
rect 12207 12709 12219 12743
rect 12618 12724 12624 12776
rect 12676 12724 12682 12776
rect 12713 12767 12771 12773
rect 12713 12733 12725 12767
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 12161 12703 12219 12709
rect 12728 12696 12756 12727
rect 13004 12696 13032 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 13722 12724 13728 12776
rect 13780 12724 13786 12776
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12764 13875 12767
rect 13998 12764 14004 12776
rect 13863 12736 14004 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12764 14151 12767
rect 14274 12764 14280 12776
rect 14139 12736 14280 12764
rect 14139 12733 14151 12736
rect 14093 12727 14151 12733
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 14918 12764 14924 12776
rect 14875 12736 14924 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15841 12767 15899 12773
rect 15841 12764 15853 12767
rect 15252 12736 15853 12764
rect 15252 12724 15258 12736
rect 15841 12733 15853 12736
rect 15887 12733 15899 12767
rect 15841 12727 15899 12733
rect 16108 12767 16166 12773
rect 16108 12733 16120 12767
rect 16154 12764 16166 12767
rect 17126 12764 17132 12776
rect 16154 12736 17132 12764
rect 16154 12733 16166 12736
rect 16108 12727 16166 12733
rect 17126 12724 17132 12736
rect 17184 12724 17190 12776
rect 10928 12668 12020 12696
rect 12636 12668 13032 12696
rect 10928 12656 10934 12668
rect 12636 12640 12664 12668
rect 13078 12656 13084 12708
rect 13136 12696 13142 12708
rect 14182 12696 14188 12708
rect 13136 12668 14188 12696
rect 13136 12656 13142 12668
rect 14182 12656 14188 12668
rect 14240 12696 14246 12708
rect 15286 12696 15292 12708
rect 14240 12668 15292 12696
rect 14240 12656 14246 12668
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 15470 12656 15476 12708
rect 15528 12696 15534 12708
rect 16390 12696 16396 12708
rect 15528 12668 16396 12696
rect 15528 12656 15534 12668
rect 16390 12656 16396 12668
rect 16448 12656 16454 12708
rect 9548 12600 10272 12628
rect 11241 12631 11299 12637
rect 9548 12588 9554 12600
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 11790 12628 11796 12640
rect 11287 12600 11796 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 12618 12588 12624 12640
rect 12676 12588 12682 12640
rect 12802 12588 12808 12640
rect 12860 12628 12866 12640
rect 13541 12631 13599 12637
rect 13541 12628 13553 12631
rect 12860 12600 13553 12628
rect 12860 12588 12866 12600
rect 13541 12597 13553 12600
rect 13587 12628 13599 12631
rect 13630 12628 13636 12640
rect 13587 12600 13636 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 15930 12628 15936 12640
rect 14884 12600 15936 12628
rect 14884 12588 14890 12600
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 552 12538 17664 12560
rect 552 12486 4366 12538
rect 4418 12486 4430 12538
rect 4482 12486 4494 12538
rect 4546 12486 4558 12538
rect 4610 12486 4622 12538
rect 4674 12486 4686 12538
rect 4738 12486 10366 12538
rect 10418 12486 10430 12538
rect 10482 12486 10494 12538
rect 10546 12486 10558 12538
rect 10610 12486 10622 12538
rect 10674 12486 10686 12538
rect 10738 12486 16366 12538
rect 16418 12486 16430 12538
rect 16482 12486 16494 12538
rect 16546 12486 16558 12538
rect 16610 12486 16622 12538
rect 16674 12486 16686 12538
rect 16738 12486 17664 12538
rect 552 12464 17664 12486
rect 2958 12384 2964 12436
rect 3016 12384 3022 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 3510 12424 3516 12436
rect 3191 12396 3516 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 3605 12427 3663 12433
rect 3605 12393 3617 12427
rect 3651 12393 3663 12427
rect 3605 12387 3663 12393
rect 2976 12356 3004 12384
rect 3620 12356 3648 12387
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4479 12427 4537 12433
rect 4479 12424 4491 12427
rect 4212 12396 4491 12424
rect 4212 12384 4218 12396
rect 4479 12393 4491 12396
rect 4525 12424 4537 12427
rect 6822 12424 6828 12436
rect 4525 12396 6828 12424
rect 4525 12393 4537 12396
rect 4479 12387 4537 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7926 12384 7932 12436
rect 7984 12384 7990 12436
rect 8386 12384 8392 12436
rect 8444 12384 8450 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 13262 12424 13268 12436
rect 12584 12396 13268 12424
rect 12584 12384 12590 12396
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 13817 12427 13875 12433
rect 13817 12393 13829 12427
rect 13863 12424 13875 12427
rect 13863 12396 14688 12424
rect 13863 12393 13875 12396
rect 13817 12387 13875 12393
rect 2976 12328 4844 12356
rect 1118 12297 1124 12300
rect 1112 12251 1124 12297
rect 1118 12248 1124 12251
rect 1176 12248 1182 12300
rect 2958 12248 2964 12300
rect 3016 12248 3022 12300
rect 4816 12297 4844 12328
rect 5718 12316 5724 12368
rect 5776 12316 5782 12368
rect 6012 12328 6316 12356
rect 3513 12291 3571 12297
rect 3513 12257 3525 12291
rect 3559 12257 3571 12291
rect 3513 12251 3571 12257
rect 3789 12291 3847 12297
rect 3789 12257 3801 12291
rect 3835 12288 3847 12291
rect 4801 12291 4859 12297
rect 3835 12260 4752 12288
rect 3835 12257 3847 12260
rect 3789 12251 3847 12257
rect 842 12180 848 12232
rect 900 12180 906 12232
rect 2222 12180 2228 12232
rect 2280 12180 2286 12232
rect 3528 12220 3556 12251
rect 4246 12220 4252 12232
rect 3528 12192 4252 12220
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 4724 12229 4752 12260
rect 4801 12257 4813 12291
rect 4847 12257 4859 12291
rect 5736 12288 5764 12316
rect 6012 12297 6040 12328
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 5736 12260 6009 12288
rect 4801 12251 4859 12257
rect 5997 12257 6009 12260
rect 6043 12257 6055 12291
rect 5997 12251 6055 12257
rect 6178 12248 6184 12300
rect 6236 12248 6242 12300
rect 6288 12297 6316 12328
rect 6454 12316 6460 12368
rect 6512 12356 6518 12368
rect 7561 12359 7619 12365
rect 7561 12356 7573 12359
rect 6512 12328 7573 12356
rect 6512 12316 6518 12328
rect 7561 12325 7573 12328
rect 7607 12325 7619 12359
rect 7561 12319 7619 12325
rect 7699 12359 7757 12365
rect 7699 12325 7711 12359
rect 7745 12356 7757 12359
rect 7745 12328 8248 12356
rect 7745 12325 7757 12328
rect 7699 12319 7757 12325
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 6788 12260 7205 12288
rect 6788 12248 6794 12260
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 7340 12260 7389 12288
rect 7340 12248 7346 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12257 7527 12291
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 7469 12251 7527 12257
rect 7944 12260 8125 12288
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12220 5135 12223
rect 6549 12223 6607 12229
rect 5123 12192 6500 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 2240 12152 2268 12180
rect 4724 12152 4752 12183
rect 4982 12152 4988 12164
rect 2240 12124 3547 12152
rect 4724 12124 4988 12152
rect 2130 12044 2136 12096
rect 2188 12084 2194 12096
rect 2225 12087 2283 12093
rect 2225 12084 2237 12087
rect 2188 12056 2237 12084
rect 2188 12044 2194 12056
rect 2225 12053 2237 12056
rect 2271 12053 2283 12087
rect 2225 12047 2283 12053
rect 3418 12044 3424 12096
rect 3476 12044 3482 12096
rect 3519 12084 3547 12124
rect 4982 12112 4988 12124
rect 5040 12152 5046 12164
rect 5813 12155 5871 12161
rect 5813 12152 5825 12155
rect 5040 12124 5825 12152
rect 5040 12112 5046 12124
rect 5813 12121 5825 12124
rect 5859 12121 5871 12155
rect 6472 12152 6500 12192
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 6638 12220 6644 12232
rect 6595 12192 6644 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7098 12152 7104 12164
rect 6472 12124 7104 12152
rect 5813 12115 5871 12121
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 7484 12152 7512 12251
rect 7834 12180 7840 12232
rect 7892 12180 7898 12232
rect 7944 12152 7972 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8220 12288 8248 12328
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 11238 12356 11244 12368
rect 8352 12328 11244 12356
rect 8352 12316 8358 12328
rect 11238 12316 11244 12328
rect 11296 12316 11302 12368
rect 11440 12328 13584 12356
rect 8573 12291 8631 12297
rect 8220 12260 8340 12288
rect 8113 12251 8171 12257
rect 8312 12232 8340 12260
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 9306 12288 9312 12300
rect 8619 12260 9312 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 8294 12180 8300 12232
rect 8352 12180 8358 12232
rect 8588 12220 8616 12251
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11440 12297 11468 12328
rect 11698 12297 11704 12300
rect 11425 12291 11483 12297
rect 11425 12288 11437 12291
rect 11020 12260 11437 12288
rect 11020 12248 11026 12260
rect 11425 12257 11437 12260
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 11692 12251 11704 12297
rect 11698 12248 11704 12251
rect 11756 12248 11762 12300
rect 8404 12192 8616 12220
rect 7484 12124 7972 12152
rect 7944 12096 7972 12124
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 8404 12152 8432 12192
rect 8168 12124 8432 12152
rect 8168 12112 8174 12124
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 8938 12152 8944 12164
rect 8628 12124 8944 12152
rect 8628 12112 8634 12124
rect 8938 12112 8944 12124
rect 8996 12112 9002 12164
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 9456 12124 11468 12152
rect 9456 12112 9462 12124
rect 4890 12084 4896 12096
rect 3519 12056 4896 12084
rect 4890 12044 4896 12056
rect 4948 12084 4954 12096
rect 6546 12084 6552 12096
rect 4948 12056 6552 12084
rect 4948 12044 4954 12056
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 7742 12084 7748 12096
rect 7248 12056 7748 12084
rect 7248 12044 7254 12056
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 7926 12044 7932 12096
rect 7984 12044 7990 12096
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 11330 12084 11336 12096
rect 8536 12056 11336 12084
rect 8536 12044 8542 12056
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 11440 12084 11468 12124
rect 12526 12084 12532 12096
rect 11440 12056 12532 12084
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 12802 12044 12808 12096
rect 12860 12044 12866 12096
rect 13556 12084 13584 12328
rect 13630 12316 13636 12368
rect 13688 12356 13694 12368
rect 14001 12359 14059 12365
rect 14001 12356 14013 12359
rect 13688 12328 14013 12356
rect 13688 12316 13694 12328
rect 14001 12325 14013 12328
rect 14047 12356 14059 12359
rect 14550 12356 14556 12368
rect 14047 12328 14556 12356
rect 14047 12325 14059 12328
rect 14001 12319 14059 12325
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 14660 12356 14688 12396
rect 15470 12384 15476 12436
rect 15528 12384 15534 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17218 12424 17224 12436
rect 17000 12396 17224 12424
rect 17000 12384 17006 12396
rect 17218 12384 17224 12396
rect 17276 12384 17282 12436
rect 14798 12359 14856 12365
rect 14798 12356 14810 12359
rect 14660 12328 14810 12356
rect 14798 12325 14810 12328
rect 14844 12325 14856 12359
rect 14798 12319 14856 12325
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 13814 12288 13820 12300
rect 13771 12260 13820 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 13906 12248 13912 12300
rect 13964 12248 13970 12300
rect 15488 12288 15516 12384
rect 16684 12328 17264 12356
rect 16684 12297 16712 12328
rect 17236 12297 17264 12328
rect 16669 12291 16727 12297
rect 16669 12288 16681 12291
rect 14476 12260 15516 12288
rect 15948 12260 16681 12288
rect 14476 12229 14504 12260
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14274 12112 14280 12164
rect 14332 12112 14338 12164
rect 14568 12084 14596 12183
rect 14918 12084 14924 12096
rect 13556 12056 14924 12084
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15194 12044 15200 12096
rect 15252 12084 15258 12096
rect 15948 12093 15976 12260
rect 16669 12257 16681 12260
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17221 12291 17279 12297
rect 17221 12257 17233 12291
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 16761 12223 16819 12229
rect 16761 12189 16773 12223
rect 16807 12220 16819 12223
rect 17034 12220 17040 12232
rect 16807 12192 17040 12220
rect 16807 12189 16819 12192
rect 16761 12183 16819 12189
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 17144 12220 17172 12251
rect 17402 12220 17408 12232
rect 17144 12192 17408 12220
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 15933 12087 15991 12093
rect 15933 12084 15945 12087
rect 15252 12056 15945 12084
rect 15252 12044 15258 12056
rect 15933 12053 15945 12056
rect 15979 12053 15991 12087
rect 15933 12047 15991 12053
rect 16206 12044 16212 12096
rect 16264 12084 16270 12096
rect 16301 12087 16359 12093
rect 16301 12084 16313 12087
rect 16264 12056 16313 12084
rect 16264 12044 16270 12056
rect 16301 12053 16313 12056
rect 16347 12053 16359 12087
rect 16301 12047 16359 12053
rect 16942 12044 16948 12096
rect 17000 12044 17006 12096
rect 552 11994 17664 12016
rect 552 11942 1366 11994
rect 1418 11942 1430 11994
rect 1482 11942 1494 11994
rect 1546 11942 1558 11994
rect 1610 11942 1622 11994
rect 1674 11942 1686 11994
rect 1738 11942 7366 11994
rect 7418 11942 7430 11994
rect 7482 11942 7494 11994
rect 7546 11942 7558 11994
rect 7610 11942 7622 11994
rect 7674 11942 7686 11994
rect 7738 11942 13366 11994
rect 13418 11942 13430 11994
rect 13482 11942 13494 11994
rect 13546 11942 13558 11994
rect 13610 11942 13622 11994
rect 13674 11942 13686 11994
rect 13738 11942 17664 11994
rect 552 11920 17664 11942
rect 1118 11840 1124 11892
rect 1176 11880 1182 11892
rect 1397 11883 1455 11889
rect 1397 11880 1409 11883
rect 1176 11852 1409 11880
rect 1176 11840 1182 11852
rect 1397 11849 1409 11852
rect 1443 11849 1455 11883
rect 1397 11843 1455 11849
rect 1762 11840 1768 11892
rect 1820 11840 1826 11892
rect 1949 11883 2007 11889
rect 1949 11849 1961 11883
rect 1995 11880 2007 11883
rect 2682 11880 2688 11892
rect 1995 11852 2688 11880
rect 1995 11849 2007 11852
rect 1949 11843 2007 11849
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3200 11852 3985 11880
rect 3200 11840 3206 11852
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 3973 11843 4031 11849
rect 7282 11840 7288 11892
rect 7340 11840 7346 11892
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 7892 11852 8033 11880
rect 7892 11840 7898 11852
rect 8021 11849 8033 11852
rect 8067 11849 8079 11883
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 8021 11843 8079 11849
rect 8128 11852 8585 11880
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 1780 11676 1808 11840
rect 2590 11812 2596 11824
rect 2240 11784 2596 11812
rect 2240 11753 2268 11784
rect 2590 11772 2596 11784
rect 2648 11772 2654 11824
rect 3326 11772 3332 11824
rect 3384 11812 3390 11824
rect 3384 11784 5948 11812
rect 3384 11772 3390 11784
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 1627 11648 1808 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 1412 11608 1440 11639
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2096 11648 2176 11676
rect 2096 11636 2102 11648
rect 2148 11617 2176 11648
rect 2406 11636 2412 11688
rect 2464 11636 2470 11688
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11645 2559 11679
rect 3528 11676 3556 11784
rect 5920 11756 5948 11784
rect 6178 11772 6184 11824
rect 6236 11812 6242 11824
rect 7300 11812 7328 11840
rect 8128 11812 8156 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 8573 11843 8631 11849
rect 9033 11883 9091 11889
rect 9033 11849 9045 11883
rect 9079 11880 9091 11883
rect 9398 11880 9404 11892
rect 9079 11852 9404 11880
rect 9079 11849 9091 11852
rect 9033 11843 9091 11849
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 11885 11883 11943 11889
rect 11885 11880 11897 11883
rect 11756 11852 11897 11880
rect 11756 11840 11762 11852
rect 11885 11849 11897 11852
rect 11931 11849 11943 11883
rect 11885 11843 11943 11849
rect 12989 11883 13047 11889
rect 12989 11849 13001 11883
rect 13035 11880 13047 11883
rect 13078 11880 13084 11892
rect 13035 11852 13084 11880
rect 13035 11849 13047 11852
rect 12989 11843 13047 11849
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 13909 11883 13967 11889
rect 13909 11880 13921 11883
rect 13832 11852 13921 11880
rect 6236 11784 7236 11812
rect 7300 11784 8156 11812
rect 9125 11815 9183 11821
rect 6236 11772 6242 11784
rect 3602 11704 3608 11756
rect 3660 11744 3666 11756
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 3660 11716 4629 11744
rect 3660 11704 3666 11716
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6638 11744 6644 11756
rect 6420 11716 6644 11744
rect 6420 11704 6426 11716
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 7208 11744 7236 11784
rect 9125 11781 9137 11815
rect 9171 11812 9183 11815
rect 9306 11812 9312 11824
rect 9171 11784 9312 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 9306 11772 9312 11784
rect 9364 11772 9370 11824
rect 12161 11815 12219 11821
rect 11716 11784 12112 11812
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 7208 11716 7604 11744
rect 3881 11679 3939 11685
rect 3881 11676 3893 11679
rect 3528 11648 3893 11676
rect 2501 11639 2559 11645
rect 3881 11645 3893 11648
rect 3927 11645 3939 11679
rect 3881 11639 3939 11645
rect 2133 11611 2191 11617
rect 1412 11580 2084 11608
rect 1946 11549 1952 11552
rect 1933 11543 1952 11549
rect 1933 11509 1945 11543
rect 1933 11503 1952 11509
rect 1946 11500 1952 11503
rect 2004 11500 2010 11552
rect 2056 11540 2084 11580
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 2516 11608 2544 11639
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 4028 11648 4169 11676
rect 4028 11636 4034 11648
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4338 11636 4344 11688
rect 4396 11636 4402 11688
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11676 4583 11679
rect 4798 11676 4804 11688
rect 4571 11648 4804 11676
rect 4571 11645 4583 11648
rect 4525 11639 4583 11645
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 6454 11676 6460 11688
rect 5460 11648 6460 11676
rect 2179 11580 2544 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 3418 11568 3424 11620
rect 3476 11608 3482 11620
rect 4249 11611 4307 11617
rect 4249 11608 4261 11611
rect 3476 11580 4261 11608
rect 3476 11568 3482 11580
rect 4249 11577 4261 11580
rect 4295 11608 4307 11611
rect 5460 11608 5488 11648
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 7576 11685 7604 11716
rect 8220 11716 8953 11744
rect 7377 11679 7435 11685
rect 7377 11676 7389 11679
rect 7064 11648 7389 11676
rect 7064 11636 7070 11648
rect 7377 11645 7389 11648
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 7650 11636 7656 11688
rect 7708 11636 7714 11688
rect 7742 11636 7748 11688
rect 7800 11636 7806 11688
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11676 7895 11679
rect 8018 11676 8024 11688
rect 7883 11648 8024 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 4295 11580 5488 11608
rect 4295 11577 4307 11580
rect 4249 11571 4307 11577
rect 6178 11568 6184 11620
rect 6236 11608 6242 11620
rect 6365 11611 6423 11617
rect 6365 11608 6377 11611
rect 6236 11580 6377 11608
rect 6236 11568 6242 11580
rect 6365 11577 6377 11580
rect 6411 11577 6423 11611
rect 6365 11571 6423 11577
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 2056 11512 2237 11540
rect 2225 11509 2237 11512
rect 2271 11509 2283 11543
rect 2225 11503 2283 11509
rect 3697 11543 3755 11549
rect 3697 11509 3709 11543
rect 3743 11540 3755 11543
rect 4154 11540 4160 11552
rect 3743 11512 4160 11540
rect 3743 11509 3755 11512
rect 3697 11503 3755 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4982 11500 4988 11552
rect 5040 11540 5046 11552
rect 5350 11540 5356 11552
rect 5040 11512 5356 11540
rect 5040 11500 5046 11512
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 7374 11500 7380 11552
rect 7432 11540 7438 11552
rect 8220 11540 8248 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9324 11716 10088 11744
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11672 8815 11679
rect 8803 11645 8892 11672
rect 8757 11644 8892 11645
rect 8757 11639 8815 11644
rect 8864 11608 8892 11644
rect 9030 11636 9036 11688
rect 9088 11636 9094 11688
rect 9324 11685 9352 11716
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 9232 11648 9321 11676
rect 9122 11608 9128 11620
rect 8864 11580 9128 11608
rect 9122 11568 9128 11580
rect 9180 11608 9186 11620
rect 9232 11608 9260 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9398 11636 9404 11688
rect 9456 11636 9462 11688
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 9861 11679 9919 11685
rect 9548 11648 9812 11676
rect 9548 11636 9554 11648
rect 9180 11580 9260 11608
rect 9180 11568 9186 11580
rect 9582 11568 9588 11620
rect 9640 11568 9646 11620
rect 9784 11608 9812 11648
rect 9861 11645 9873 11679
rect 9907 11676 9919 11679
rect 9950 11676 9956 11688
rect 9907 11648 9956 11676
rect 9907 11645 9919 11648
rect 9861 11639 9919 11645
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 10060 11685 10088 11716
rect 10226 11704 10232 11756
rect 10284 11744 10290 11756
rect 11716 11744 11744 11784
rect 10284 11716 10640 11744
rect 10284 11704 10290 11716
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10183 11648 10548 11676
rect 10612 11662 10640 11716
rect 11624 11716 11744 11744
rect 11977 11747 12035 11753
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10520 11617 10548 11648
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 11624 11685 11652 11716
rect 11977 11713 11989 11747
rect 12023 11713 12035 11747
rect 12084 11744 12112 11784
rect 12161 11781 12173 11815
rect 12207 11812 12219 11815
rect 13170 11812 13176 11824
rect 12207 11784 13176 11812
rect 12207 11781 12219 11784
rect 12161 11775 12219 11781
rect 13170 11772 13176 11784
rect 13228 11812 13234 11824
rect 13541 11815 13599 11821
rect 13541 11812 13553 11815
rect 13228 11784 13553 11812
rect 13228 11772 13234 11784
rect 13541 11781 13553 11784
rect 13587 11781 13599 11815
rect 13541 11775 13599 11781
rect 13832 11756 13860 11852
rect 13909 11849 13921 11852
rect 13955 11849 13967 11883
rect 13909 11843 13967 11849
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14369 11883 14427 11889
rect 14139 11852 14320 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14292 11812 14320 11852
rect 14369 11849 14381 11883
rect 14415 11880 14427 11883
rect 15562 11880 15568 11892
rect 14415 11852 15568 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 15562 11840 15568 11852
rect 15620 11880 15626 11892
rect 16669 11883 16727 11889
rect 16669 11880 16681 11883
rect 15620 11852 16681 11880
rect 15620 11840 15626 11852
rect 16669 11849 16681 11852
rect 16715 11849 16727 11883
rect 16669 11843 16727 11849
rect 14826 11812 14832 11824
rect 14292 11784 14832 11812
rect 14826 11772 14832 11784
rect 14884 11772 14890 11824
rect 12802 11744 12808 11756
rect 12084 11716 12434 11744
rect 11977 11707 12035 11713
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 11296 11648 11621 11676
rect 11296 11636 11302 11648
rect 11609 11645 11621 11648
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 11698 11636 11704 11688
rect 11756 11636 11762 11688
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11645 11943 11679
rect 11992 11676 12020 11707
rect 12253 11679 12311 11685
rect 11992 11648 12112 11676
rect 11885 11639 11943 11645
rect 10505 11611 10563 11617
rect 9784 11580 10180 11608
rect 10152 11552 10180 11580
rect 10505 11577 10517 11611
rect 10551 11608 10563 11611
rect 11900 11608 11928 11639
rect 12084 11620 12112 11648
rect 12253 11645 12265 11679
rect 12299 11645 12311 11679
rect 12406 11676 12434 11716
rect 12544 11716 12808 11744
rect 12544 11676 12572 11716
rect 12802 11704 12808 11716
rect 12860 11744 12866 11756
rect 12860 11716 13216 11744
rect 12860 11704 12866 11716
rect 12406 11648 12572 11676
rect 12713 11679 12771 11685
rect 12253 11639 12311 11645
rect 12713 11645 12725 11679
rect 12759 11676 12771 11679
rect 13078 11676 13084 11688
rect 12759 11648 13084 11676
rect 12759 11645 12771 11648
rect 12713 11639 12771 11645
rect 11977 11611 12035 11617
rect 11977 11608 11989 11611
rect 10551 11580 11100 11608
rect 11900 11580 11989 11608
rect 10551 11577 10563 11580
rect 10505 11571 10563 11577
rect 11072 11552 11100 11580
rect 11977 11577 11989 11580
rect 12023 11577 12035 11611
rect 11977 11571 12035 11577
rect 12066 11568 12072 11620
rect 12124 11568 12130 11620
rect 7432 11512 8248 11540
rect 7432 11500 7438 11512
rect 9674 11500 9680 11552
rect 9732 11500 9738 11552
rect 10134 11500 10140 11552
rect 10192 11500 10198 11552
rect 11054 11500 11060 11552
rect 11112 11500 11118 11552
rect 11425 11543 11483 11549
rect 11425 11509 11437 11543
rect 11471 11540 11483 11543
rect 11514 11540 11520 11552
rect 11471 11512 11520 11540
rect 11471 11509 11483 11512
rect 11425 11503 11483 11509
rect 11514 11500 11520 11512
rect 11572 11540 11578 11552
rect 12268 11540 12296 11639
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 13188 11617 13216 11716
rect 13814 11704 13820 11756
rect 13872 11704 13878 11756
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 13838 11648 14657 11676
rect 13173 11611 13231 11617
rect 12452 11580 12848 11608
rect 11572 11512 12296 11540
rect 11572 11500 11578 11512
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 12452 11540 12480 11580
rect 12400 11512 12480 11540
rect 12529 11543 12587 11549
rect 12400 11500 12406 11512
rect 12529 11509 12541 11543
rect 12575 11540 12587 11543
rect 12710 11540 12716 11552
rect 12575 11512 12716 11540
rect 12575 11509 12587 11512
rect 12529 11503 12587 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 12820 11549 12848 11580
rect 13173 11577 13185 11611
rect 13219 11577 13231 11611
rect 13173 11571 13231 11577
rect 12805 11543 12863 11549
rect 12805 11509 12817 11543
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 12973 11543 13031 11549
rect 12973 11509 12985 11543
rect 13019 11540 13031 11543
rect 13722 11540 13728 11552
rect 13019 11512 13728 11540
rect 13019 11509 13031 11512
rect 12973 11503 13031 11509
rect 13722 11500 13728 11512
rect 13780 11540 13786 11552
rect 13838 11540 13866 11648
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 14734 11636 14740 11688
rect 14792 11676 14798 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 14792 11648 14841 11676
rect 14792 11636 14798 11648
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 14918 11636 14924 11688
rect 14976 11676 14982 11688
rect 15289 11679 15347 11685
rect 15289 11676 15301 11679
rect 14976 11648 15301 11676
rect 14976 11636 14982 11648
rect 15289 11645 15301 11648
rect 15335 11645 15347 11679
rect 15289 11639 15347 11645
rect 13909 11611 13967 11617
rect 13909 11577 13921 11611
rect 13955 11608 13967 11611
rect 14553 11611 14611 11617
rect 13955 11580 14504 11608
rect 13955 11577 13967 11580
rect 13909 11571 13967 11577
rect 14366 11549 14372 11552
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 13780 11512 14197 11540
rect 13780 11500 13786 11512
rect 14185 11509 14197 11512
rect 14231 11509 14243 11543
rect 14185 11503 14243 11509
rect 14348 11543 14372 11549
rect 14348 11509 14360 11543
rect 14348 11503 14372 11509
rect 14366 11500 14372 11503
rect 14424 11500 14430 11552
rect 14476 11540 14504 11580
rect 14553 11577 14565 11611
rect 14599 11608 14611 11611
rect 15102 11608 15108 11620
rect 14599 11580 15108 11608
rect 14599 11577 14611 11580
rect 14553 11571 14611 11577
rect 15102 11568 15108 11580
rect 15160 11568 15166 11620
rect 15556 11611 15614 11617
rect 15556 11577 15568 11611
rect 15602 11608 15614 11611
rect 16114 11608 16120 11620
rect 15602 11580 16120 11608
rect 15602 11577 15614 11580
rect 15556 11571 15614 11577
rect 16114 11568 16120 11580
rect 16172 11568 16178 11620
rect 15013 11543 15071 11549
rect 15013 11540 15025 11543
rect 14476 11512 15025 11540
rect 15013 11509 15025 11512
rect 15059 11509 15071 11543
rect 15013 11503 15071 11509
rect 552 11450 17664 11472
rect 552 11398 4366 11450
rect 4418 11398 4430 11450
rect 4482 11398 4494 11450
rect 4546 11398 4558 11450
rect 4610 11398 4622 11450
rect 4674 11398 4686 11450
rect 4738 11398 10366 11450
rect 10418 11398 10430 11450
rect 10482 11398 10494 11450
rect 10546 11398 10558 11450
rect 10610 11398 10622 11450
rect 10674 11398 10686 11450
rect 10738 11398 16366 11450
rect 16418 11398 16430 11450
rect 16482 11398 16494 11450
rect 16546 11398 16558 11450
rect 16610 11398 16622 11450
rect 16674 11398 16686 11450
rect 16738 11398 17664 11450
rect 552 11376 17664 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1762 11336 1768 11348
rect 1719 11308 1768 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1762 11296 1768 11308
rect 1820 11336 1826 11348
rect 2406 11336 2412 11348
rect 1820 11308 2412 11336
rect 1820 11296 1826 11308
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 4338 11336 4344 11348
rect 4295 11308 4344 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 4338 11296 4344 11308
rect 4396 11336 4402 11348
rect 4617 11339 4675 11345
rect 4396 11308 4568 11336
rect 4396 11296 4402 11308
rect 842 11228 848 11280
rect 900 11268 906 11280
rect 2860 11271 2918 11277
rect 900 11240 2636 11268
rect 900 11228 906 11240
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11200 1915 11203
rect 1946 11200 1952 11212
rect 1903 11172 1952 11200
rect 1903 11169 1915 11172
rect 1857 11163 1915 11169
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 2608 11209 2636 11240
rect 2860 11237 2872 11271
rect 2906 11268 2918 11271
rect 4062 11268 4068 11280
rect 2906 11240 4068 11268
rect 2906 11237 2918 11240
rect 2860 11231 2918 11237
rect 4062 11228 4068 11240
rect 4120 11228 4126 11280
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 4540 11268 4568 11308
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 4798 11336 4804 11348
rect 4663 11308 4804 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7745 11339 7803 11345
rect 6972 11308 7420 11336
rect 6972 11296 6978 11308
rect 7392 11268 7420 11308
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 7926 11336 7932 11348
rect 7791 11308 7932 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 8018 11296 8024 11348
rect 8076 11296 8082 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 8570 11336 8576 11348
rect 8444 11308 8576 11336
rect 8444 11296 8450 11308
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8665 11339 8723 11345
rect 8665 11305 8677 11339
rect 8711 11336 8723 11339
rect 9030 11336 9036 11348
rect 8711 11308 9036 11336
rect 8711 11305 8723 11308
rect 8665 11299 8723 11305
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 9217 11339 9275 11345
rect 9217 11305 9229 11339
rect 9263 11336 9275 11339
rect 9582 11336 9588 11348
rect 9263 11308 9588 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 10226 11296 10232 11348
rect 10284 11296 10290 11348
rect 11238 11296 11244 11348
rect 11296 11296 11302 11348
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 12342 11336 12348 11348
rect 11756 11308 12348 11336
rect 11756 11296 11762 11308
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 13078 11336 13084 11348
rect 12952 11308 13084 11336
rect 12952 11296 12958 11308
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 15657 11339 15715 11345
rect 15657 11336 15669 11339
rect 13964 11308 15669 11336
rect 13964 11296 13970 11308
rect 15657 11305 15669 11308
rect 15703 11305 15715 11339
rect 15657 11299 15715 11305
rect 16114 11296 16120 11348
rect 16172 11296 16178 11348
rect 16206 11296 16212 11348
rect 16264 11296 16270 11348
rect 16942 11296 16948 11348
rect 17000 11296 17006 11348
rect 8036 11268 8064 11296
rect 4212 11240 4476 11268
rect 4540 11240 5120 11268
rect 4212 11228 4218 11240
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11200 2099 11203
rect 2133 11203 2191 11209
rect 2133 11200 2145 11203
rect 2087 11172 2145 11200
rect 2087 11169 2099 11172
rect 2041 11163 2099 11169
rect 2133 11169 2145 11172
rect 2179 11200 2191 11203
rect 2593 11203 2651 11209
rect 2179 11172 2544 11200
rect 2179 11169 2191 11172
rect 2133 11163 2191 11169
rect 1964 11064 1992 11160
rect 2314 11092 2320 11144
rect 2372 11132 2378 11144
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2372 11104 2421 11132
rect 2372 11092 2378 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2225 11067 2283 11073
rect 2225 11064 2237 11067
rect 1964 11036 2237 11064
rect 2225 11033 2237 11036
rect 2271 11033 2283 11067
rect 2225 11027 2283 11033
rect 2314 10956 2320 11008
rect 2372 10956 2378 11008
rect 2516 10996 2544 11172
rect 2593 11169 2605 11203
rect 2639 11200 2651 11203
rect 3602 11200 3608 11212
rect 2639 11172 3608 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 3602 11160 3608 11172
rect 3660 11160 3666 11212
rect 4448 11209 4476 11240
rect 5092 11212 5120 11240
rect 5184 11240 6592 11268
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11169 4399 11203
rect 4341 11163 4399 11169
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4798 11200 4804 11212
rect 4479 11172 4804 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4356 11132 4384 11163
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 4982 11160 4988 11212
rect 5040 11160 5046 11212
rect 5074 11160 5080 11212
rect 5132 11160 5138 11212
rect 5184 11209 5212 11240
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11169 5319 11203
rect 5810 11200 5816 11212
rect 5261 11163 5319 11169
rect 5552 11172 5816 11200
rect 5276 11132 5304 11163
rect 4212 11104 4384 11132
rect 5184 11104 5304 11132
rect 4212 11092 4218 11104
rect 5184 11076 5212 11104
rect 3973 11067 4031 11073
rect 3973 11033 3985 11067
rect 4019 11064 4031 11067
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 4019 11036 4077 11064
rect 4019 11033 4031 11036
rect 3973 11027 4031 11033
rect 4065 11033 4077 11036
rect 4111 11064 4123 11067
rect 5166 11064 5172 11076
rect 4111 11036 5172 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 5552 11008 5580 11172
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 6362 11132 6368 11144
rect 5776 11104 6368 11132
rect 5776 11092 5782 11104
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 6564 11132 6592 11240
rect 6656 11240 7328 11268
rect 7392 11240 7788 11268
rect 8036 11240 9628 11268
rect 6656 11212 6684 11240
rect 6638 11160 6644 11212
rect 6696 11160 6702 11212
rect 6730 11160 6736 11212
rect 6788 11160 6794 11212
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 7009 11203 7067 11209
rect 7009 11200 7021 11203
rect 6880 11172 7021 11200
rect 6880 11160 6886 11172
rect 7009 11169 7021 11172
rect 7055 11169 7067 11203
rect 7300 11200 7328 11240
rect 7374 11200 7380 11212
rect 7300 11172 7380 11200
rect 7009 11163 7067 11169
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11169 7527 11203
rect 7760 11198 7788 11240
rect 7837 11203 7895 11209
rect 7837 11198 7849 11203
rect 7760 11170 7849 11198
rect 7469 11163 7527 11169
rect 7837 11169 7849 11170
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 7484 11132 7512 11163
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 8849 11203 8907 11209
rect 8849 11200 8861 11203
rect 8076 11172 8861 11200
rect 8076 11160 8082 11172
rect 8849 11169 8861 11172
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11200 9183 11203
rect 9214 11200 9220 11212
rect 9171 11172 9220 11200
rect 9171 11169 9183 11172
rect 9125 11163 9183 11169
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 9600 11209 9628 11240
rect 9585 11203 9643 11209
rect 9585 11169 9597 11203
rect 9631 11169 9643 11203
rect 10244 11200 10272 11296
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 10244 11172 10609 11200
rect 9585 11163 9643 11169
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11200 10839 11203
rect 11256 11200 11284 11296
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 12437 11271 12495 11277
rect 12437 11268 12449 11271
rect 11388 11240 12449 11268
rect 11388 11228 11394 11240
rect 12437 11237 12449 11240
rect 12483 11237 12495 11271
rect 14734 11268 14740 11280
rect 12437 11231 12495 11237
rect 14108 11240 14740 11268
rect 14108 11212 14136 11240
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 16224 11268 16252 11296
rect 16224 11240 16528 11268
rect 10827 11172 11284 11200
rect 10827 11169 10839 11172
rect 10781 11163 10839 11169
rect 11606 11160 11612 11212
rect 11664 11160 11670 11212
rect 12710 11160 12716 11212
rect 12768 11200 12774 11212
rect 14090 11200 14096 11212
rect 12768 11172 14096 11200
rect 12768 11160 12774 11172
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 14185 11203 14243 11209
rect 14185 11169 14197 11203
rect 14231 11200 14243 11203
rect 14918 11200 14924 11212
rect 14231 11172 14924 11200
rect 14231 11169 14243 11172
rect 14185 11163 14243 11169
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 15160 11172 15577 11200
rect 15160 11160 15166 11172
rect 15565 11169 15577 11172
rect 15611 11169 15623 11203
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 15565 11163 15623 11169
rect 15764 11172 15945 11200
rect 8110 11132 8116 11144
rect 6564 11104 7328 11132
rect 7484 11104 8116 11132
rect 7300 11073 7328 11104
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 6825 11067 6883 11073
rect 6825 11033 6837 11067
rect 6871 11064 6883 11067
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 6871 11036 7205 11064
rect 6871 11033 6883 11036
rect 6825 11027 6883 11033
rect 7193 11033 7205 11036
rect 7239 11033 7251 11067
rect 7193 11027 7251 11033
rect 7285 11067 7343 11073
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 8570 11064 8576 11076
rect 7331 11036 8576 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 3326 10996 3332 11008
rect 2516 10968 3332 10996
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 4709 10999 4767 11005
rect 4709 10996 4721 10999
rect 3752 10968 4721 10996
rect 3752 10956 3758 10968
rect 4709 10965 4721 10968
rect 4755 10965 4767 10999
rect 4709 10959 4767 10965
rect 4985 10999 5043 11005
rect 4985 10965 4997 10999
rect 5031 10996 5043 10999
rect 5350 10996 5356 11008
rect 5031 10968 5356 10996
rect 5031 10965 5043 10968
rect 4985 10959 5043 10965
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 5445 10999 5503 11005
rect 5445 10965 5457 10999
rect 5491 10996 5503 10999
rect 5534 10996 5540 11008
rect 5491 10968 5540 10996
rect 5491 10965 5503 10968
rect 5445 10959 5503 10965
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 5997 10999 6055 11005
rect 5997 10965 6009 10999
rect 6043 10996 6055 10999
rect 6454 10996 6460 11008
rect 6043 10968 6460 10996
rect 6043 10965 6055 10968
rect 5997 10959 6055 10965
rect 6454 10956 6460 10968
rect 6512 10996 6518 11008
rect 6730 10996 6736 11008
rect 6512 10968 6736 10996
rect 6512 10956 6518 10968
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 7208 10996 7236 11027
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 9048 11064 9076 11095
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 9493 11135 9551 11141
rect 9493 11132 9505 11135
rect 9364 11104 9505 11132
rect 9364 11092 9370 11104
rect 9493 11101 9505 11104
rect 9539 11101 9551 11135
rect 9493 11095 9551 11101
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 10008 11104 10425 11132
rect 10008 11092 10014 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 11112 11104 11437 11132
rect 11112 11092 11118 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 12250 11092 12256 11144
rect 12308 11092 12314 11144
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 15010 11132 15016 11144
rect 14608 11104 15016 11132
rect 14608 11092 14614 11104
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 13630 11064 13636 11076
rect 9048 11036 13636 11064
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 14274 11024 14280 11076
rect 14332 11064 14338 11076
rect 15672 11064 15700 11095
rect 14332 11036 15700 11064
rect 14332 11024 14338 11036
rect 8849 10999 8907 11005
rect 8849 10996 8861 10999
rect 7208 10968 8861 10996
rect 8849 10965 8861 10968
rect 8895 10965 8907 10999
rect 8849 10959 8907 10965
rect 9582 10956 9588 11008
rect 9640 10956 9646 11008
rect 10134 10956 10140 11008
rect 10192 10996 10198 11008
rect 11146 10996 11152 11008
rect 10192 10968 11152 10996
rect 10192 10956 10198 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 14292 10996 14320 11024
rect 12124 10968 14320 10996
rect 12124 10956 12130 10968
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 15335 10999 15393 11005
rect 15335 10996 15347 10999
rect 14608 10968 15347 10996
rect 14608 10956 14614 10968
rect 15335 10965 15347 10968
rect 15381 10996 15393 10999
rect 15764 10996 15792 11172
rect 15933 11169 15945 11172
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 16298 11160 16304 11212
rect 16356 11160 16362 11212
rect 16500 11209 16528 11240
rect 16485 11203 16543 11209
rect 16485 11169 16497 11203
rect 16531 11169 16543 11203
rect 16485 11163 16543 11169
rect 16574 11160 16580 11212
rect 16632 11160 16638 11212
rect 16761 11203 16819 11209
rect 16761 11169 16773 11203
rect 16807 11200 16819 11203
rect 16960 11200 16988 11296
rect 16807 11172 16988 11200
rect 16807 11169 16819 11172
rect 16761 11163 16819 11169
rect 16945 11067 17003 11073
rect 16945 11033 16957 11067
rect 16991 11064 17003 11067
rect 17494 11064 17500 11076
rect 16991 11036 17500 11064
rect 16991 11033 17003 11036
rect 16945 11027 17003 11033
rect 17494 11024 17500 11036
rect 17552 11024 17558 11076
rect 15381 10968 15792 10996
rect 15381 10965 15393 10968
rect 15335 10959 15393 10965
rect 15838 10956 15844 11008
rect 15896 10956 15902 11008
rect 552 10906 17664 10928
rect 552 10854 1366 10906
rect 1418 10854 1430 10906
rect 1482 10854 1494 10906
rect 1546 10854 1558 10906
rect 1610 10854 1622 10906
rect 1674 10854 1686 10906
rect 1738 10854 7366 10906
rect 7418 10854 7430 10906
rect 7482 10854 7494 10906
rect 7546 10854 7558 10906
rect 7610 10854 7622 10906
rect 7674 10854 7686 10906
rect 7738 10854 13366 10906
rect 13418 10854 13430 10906
rect 13482 10854 13494 10906
rect 13546 10854 13558 10906
rect 13610 10854 13622 10906
rect 13674 10854 13686 10906
rect 13738 10854 17664 10906
rect 552 10832 17664 10854
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4304 10764 4537 10792
rect 4304 10752 4310 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5810 10792 5816 10804
rect 5123 10764 5816 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 6914 10752 6920 10804
rect 6972 10752 6978 10804
rect 7006 10752 7012 10804
rect 7064 10752 7070 10804
rect 7837 10795 7895 10801
rect 7837 10761 7849 10795
rect 7883 10761 7895 10795
rect 7837 10755 7895 10761
rect 4338 10684 4344 10736
rect 4396 10684 4402 10736
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10724 5503 10727
rect 6454 10724 6460 10736
rect 5491 10696 6460 10724
rect 5491 10693 5503 10696
rect 5445 10687 5503 10693
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 6932 10724 6960 10752
rect 7852 10724 7880 10755
rect 8018 10752 8024 10804
rect 8076 10792 8082 10804
rect 9398 10792 9404 10804
rect 8076 10764 9404 10792
rect 8076 10752 8082 10764
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 9582 10752 9588 10804
rect 9640 10792 9646 10804
rect 12802 10792 12808 10804
rect 9640 10764 12808 10792
rect 9640 10752 9646 10764
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13541 10795 13599 10801
rect 13541 10792 13553 10795
rect 13228 10764 13553 10792
rect 13228 10752 13234 10764
rect 13541 10761 13553 10764
rect 13587 10761 13599 10795
rect 13541 10755 13599 10761
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 13964 10764 14749 10792
rect 13964 10752 13970 10764
rect 14737 10761 14749 10764
rect 14783 10792 14795 10795
rect 14826 10792 14832 10804
rect 14783 10764 14832 10792
rect 14783 10761 14795 10764
rect 14737 10755 14795 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 16298 10792 16304 10804
rect 14967 10764 16304 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 6604 10684 6618 10724
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4356 10656 4384 10684
rect 4120 10628 4384 10656
rect 4893 10659 4951 10665
rect 4120 10616 4126 10628
rect 4893 10625 4905 10659
rect 4939 10656 4951 10659
rect 5258 10656 5264 10668
rect 4939 10628 5264 10656
rect 4939 10625 4951 10628
rect 4893 10619 4951 10625
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5997 10659 6055 10665
rect 5368 10628 5764 10656
rect 1489 10591 1547 10597
rect 1489 10557 1501 10591
rect 1535 10557 1547 10591
rect 1489 10551 1547 10557
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 1762 10588 1768 10600
rect 1719 10560 1768 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 1504 10520 1532 10551
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 2314 10548 2320 10600
rect 2372 10548 2378 10600
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4264 10560 4353 10588
rect 2332 10520 2360 10548
rect 1504 10492 2360 10520
rect 4264 10464 4292 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 4672 10560 4721 10588
rect 4672 10548 4678 10560
rect 4709 10557 4721 10560
rect 4755 10557 4767 10591
rect 4709 10551 4767 10557
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5368 10588 5396 10628
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5132 10560 5396 10588
rect 5552 10560 5641 10588
rect 5132 10548 5138 10560
rect 5169 10523 5227 10529
rect 5169 10489 5181 10523
rect 5215 10520 5227 10523
rect 5258 10520 5264 10532
rect 5215 10492 5264 10520
rect 5215 10489 5227 10492
rect 5169 10483 5227 10489
rect 5258 10480 5264 10492
rect 5316 10520 5322 10532
rect 5552 10520 5580 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5736 10588 5764 10628
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 6362 10656 6368 10668
rect 6043 10628 6368 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6089 10591 6147 10597
rect 6089 10588 6101 10591
rect 5736 10560 6101 10588
rect 5629 10551 5687 10557
rect 6089 10557 6101 10560
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 6273 10591 6331 10597
rect 6273 10557 6285 10591
rect 6319 10557 6331 10591
rect 6273 10551 6331 10557
rect 5813 10523 5871 10529
rect 5813 10520 5825 10523
rect 5316 10492 5580 10520
rect 5644 10492 5825 10520
rect 5316 10480 5322 10492
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 4246 10412 4252 10464
rect 4304 10412 4310 10464
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5644 10452 5672 10492
rect 5813 10489 5825 10492
rect 5859 10489 5871 10523
rect 5813 10483 5871 10489
rect 6288 10464 6316 10551
rect 6362 10480 6368 10532
rect 6420 10480 6426 10532
rect 6454 10480 6460 10532
rect 6512 10480 6518 10532
rect 6590 10529 6618 10684
rect 6932 10696 7880 10724
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 6932 10656 6960 10696
rect 7098 10656 7104 10668
rect 6779 10628 6960 10656
rect 7024 10628 7104 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 6822 10548 6828 10600
rect 6880 10548 6886 10600
rect 7024 10582 7052 10628
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7484 10600 7512 10696
rect 7926 10684 7932 10736
rect 7984 10724 7990 10736
rect 8570 10724 8576 10736
rect 7984 10696 8576 10724
rect 7984 10684 7990 10696
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 11238 10724 11244 10736
rect 9088 10696 11244 10724
rect 9088 10684 9094 10696
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 14369 10727 14427 10733
rect 11388 10696 14320 10724
rect 11388 10684 11394 10696
rect 8110 10656 8116 10668
rect 7668 10628 8116 10656
rect 7193 10591 7251 10597
rect 7193 10582 7205 10591
rect 7024 10557 7205 10582
rect 7239 10557 7251 10591
rect 7024 10554 7251 10557
rect 7193 10551 7251 10554
rect 7466 10548 7472 10600
rect 7524 10548 7530 10600
rect 7668 10597 7696 10628
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 9646 10628 11008 10656
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10557 7711 10591
rect 9646 10588 9674 10628
rect 7653 10551 7711 10557
rect 8266 10560 9674 10588
rect 10229 10591 10287 10597
rect 6590 10523 6653 10529
rect 6590 10492 6607 10523
rect 6595 10489 6607 10492
rect 6641 10520 6653 10523
rect 6730 10520 6736 10532
rect 6641 10492 6736 10520
rect 6641 10489 6653 10492
rect 6595 10483 6653 10489
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 6840 10520 6868 10548
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 6840 10492 7297 10520
rect 7285 10489 7297 10492
rect 7331 10489 7343 10523
rect 7285 10483 7343 10489
rect 7374 10480 7380 10532
rect 7432 10480 7438 10532
rect 5408 10424 5672 10452
rect 5408 10412 5414 10424
rect 5718 10412 5724 10464
rect 5776 10412 5782 10464
rect 6270 10412 6276 10464
rect 6328 10412 6334 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7576 10452 7604 10551
rect 7156 10424 7604 10452
rect 7156 10412 7162 10424
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 8266 10452 8294 10560
rect 10229 10557 10241 10591
rect 10275 10588 10287 10591
rect 10870 10588 10876 10600
rect 10275 10560 10876 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 10980 10588 11008 10628
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 12989 10659 13047 10665
rect 12768 10628 12940 10656
rect 12768 10616 12774 10628
rect 11698 10588 11704 10600
rect 10980 10560 11704 10588
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10557 12863 10591
rect 12912 10588 12940 10628
rect 12989 10625 13001 10659
rect 13035 10656 13047 10659
rect 13998 10656 14004 10668
rect 13035 10628 14004 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 14292 10656 14320 10696
rect 14369 10693 14381 10727
rect 14415 10724 14427 10727
rect 15194 10724 15200 10736
rect 14415 10696 15200 10724
rect 14415 10693 14427 10696
rect 14369 10687 14427 10693
rect 15194 10684 15200 10696
rect 15252 10724 15258 10736
rect 15838 10724 15844 10736
rect 15252 10696 15844 10724
rect 15252 10684 15258 10696
rect 15838 10684 15844 10696
rect 15896 10684 15902 10736
rect 15286 10656 15292 10668
rect 14292 10628 15292 10656
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 15562 10616 15568 10668
rect 15620 10616 15626 10668
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 16393 10659 16451 10665
rect 16393 10656 16405 10659
rect 16264 10628 16405 10656
rect 16264 10616 16270 10628
rect 16393 10625 16405 10628
rect 16439 10625 16451 10659
rect 16393 10619 16451 10625
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 12912 10560 13093 10588
rect 12805 10551 12863 10557
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10588 13323 10591
rect 13354 10588 13360 10600
rect 13311 10560 13360 10588
rect 13311 10557 13323 10560
rect 13265 10551 13323 10557
rect 8665 10523 8723 10529
rect 8665 10520 8677 10523
rect 8496 10492 8677 10520
rect 8496 10464 8524 10492
rect 8665 10489 8677 10492
rect 8711 10489 8723 10523
rect 8665 10483 8723 10489
rect 9030 10480 9036 10532
rect 9088 10520 9094 10532
rect 12820 10520 12848 10551
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 13814 10588 13820 10600
rect 13771 10560 13820 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 14090 10588 14096 10600
rect 13955 10560 14096 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 15381 10591 15439 10597
rect 15381 10588 15393 10591
rect 14752 10560 15393 10588
rect 13173 10523 13231 10529
rect 13173 10520 13185 10523
rect 9088 10492 12434 10520
rect 12820 10492 13185 10520
rect 9088 10480 9094 10492
rect 7708 10424 8294 10452
rect 7708 10412 7714 10424
rect 8478 10412 8484 10464
rect 8536 10412 8542 10464
rect 8570 10412 8576 10464
rect 8628 10452 8634 10464
rect 10226 10452 10232 10464
rect 8628 10424 10232 10452
rect 8628 10412 8634 10424
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 12406 10452 12434 10492
rect 13173 10489 13185 10492
rect 13219 10520 13231 10523
rect 14366 10520 14372 10532
rect 13219 10492 14372 10520
rect 13219 10489 13231 10492
rect 13173 10483 13231 10489
rect 14366 10480 14372 10492
rect 14424 10480 14430 10532
rect 14752 10529 14780 10560
rect 15381 10557 15393 10560
rect 15427 10557 15439 10591
rect 15580 10588 15608 10616
rect 15657 10591 15715 10597
rect 15657 10588 15669 10591
rect 15580 10560 15669 10588
rect 15381 10551 15439 10557
rect 15657 10557 15669 10560
rect 15703 10588 15715 10591
rect 15838 10588 15844 10600
rect 15703 10560 15844 10588
rect 15703 10557 15715 10560
rect 15657 10551 15715 10557
rect 15838 10548 15844 10560
rect 15896 10548 15902 10600
rect 16485 10591 16543 10597
rect 16485 10588 16497 10591
rect 16224 10560 16497 10588
rect 14737 10523 14795 10529
rect 14737 10489 14749 10523
rect 14783 10489 14795 10523
rect 14737 10483 14795 10489
rect 15013 10523 15071 10529
rect 15013 10489 15025 10523
rect 15059 10489 15071 10523
rect 15013 10483 15071 10489
rect 12621 10455 12679 10461
rect 12621 10452 12633 10455
rect 12406 10424 12633 10452
rect 12621 10421 12633 10424
rect 12667 10421 12679 10455
rect 12621 10415 12679 10421
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 15028 10452 15056 10483
rect 15102 10480 15108 10532
rect 15160 10520 15166 10532
rect 15197 10523 15255 10529
rect 15197 10520 15209 10523
rect 15160 10492 15209 10520
rect 15160 10480 15166 10492
rect 15197 10489 15209 10492
rect 15243 10489 15255 10523
rect 15197 10483 15255 10489
rect 13596 10424 15056 10452
rect 15212 10452 15240 10483
rect 16224 10464 16252 10560
rect 16485 10557 16497 10560
rect 16531 10557 16543 10591
rect 16485 10551 16543 10557
rect 15473 10455 15531 10461
rect 15473 10452 15485 10455
rect 15212 10424 15485 10452
rect 13596 10412 13602 10424
rect 15473 10421 15485 10424
rect 15519 10421 15531 10455
rect 15473 10415 15531 10421
rect 16206 10412 16212 10464
rect 16264 10412 16270 10464
rect 16853 10455 16911 10461
rect 16853 10421 16865 10455
rect 16899 10452 16911 10455
rect 16942 10452 16948 10464
rect 16899 10424 16948 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 552 10362 17664 10384
rect 552 10310 4366 10362
rect 4418 10310 4430 10362
rect 4482 10310 4494 10362
rect 4546 10310 4558 10362
rect 4610 10310 4622 10362
rect 4674 10310 4686 10362
rect 4738 10310 10366 10362
rect 10418 10310 10430 10362
rect 10482 10310 10494 10362
rect 10546 10310 10558 10362
rect 10610 10310 10622 10362
rect 10674 10310 10686 10362
rect 10738 10310 16366 10362
rect 16418 10310 16430 10362
rect 16482 10310 16494 10362
rect 16546 10310 16558 10362
rect 16610 10310 16622 10362
rect 16674 10310 16686 10362
rect 16738 10310 17664 10362
rect 552 10288 17664 10310
rect 3789 10251 3847 10257
rect 3789 10217 3801 10251
rect 3835 10248 3847 10251
rect 3970 10248 3976 10260
rect 3835 10220 3976 10248
rect 3835 10217 3847 10220
rect 3789 10211 3847 10217
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4154 10208 4160 10260
rect 4212 10208 4218 10260
rect 4341 10251 4399 10257
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 4706 10248 4712 10260
rect 4387 10220 4712 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 4893 10251 4951 10257
rect 4893 10217 4905 10251
rect 4939 10248 4951 10251
rect 4982 10248 4988 10260
rect 4939 10220 4988 10248
rect 4939 10217 4951 10220
rect 4893 10211 4951 10217
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5074 10208 5080 10260
rect 5132 10208 5138 10260
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5408 10220 5457 10248
rect 5408 10208 5414 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 6013 10251 6071 10257
rect 6013 10248 6025 10251
rect 5960 10220 6025 10248
rect 5960 10208 5966 10220
rect 6013 10217 6025 10220
rect 6059 10217 6071 10251
rect 6013 10211 6071 10217
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6420 10220 6929 10248
rect 6420 10208 6426 10220
rect 6917 10217 6929 10220
rect 6963 10217 6975 10251
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 6917 10211 6975 10217
rect 7024 10220 7941 10248
rect 2584 10183 2642 10189
rect 860 10152 2360 10180
rect 860 10056 888 10152
rect 1112 10115 1170 10121
rect 1112 10081 1124 10115
rect 1158 10112 1170 10115
rect 1578 10112 1584 10124
rect 1158 10084 1584 10112
rect 1158 10081 1170 10084
rect 1112 10075 1170 10081
rect 1578 10072 1584 10084
rect 1636 10072 1642 10124
rect 2332 10121 2360 10152
rect 2584 10149 2596 10183
rect 2630 10180 2642 10183
rect 5092 10180 5120 10208
rect 5813 10183 5871 10189
rect 5813 10180 5825 10183
rect 2630 10152 5120 10180
rect 5184 10152 5825 10180
rect 2630 10149 2642 10152
rect 2584 10143 2642 10149
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10081 2375 10115
rect 2317 10075 2375 10081
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3936 10084 3985 10112
rect 3936 10072 3942 10084
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 4062 10072 4068 10124
rect 4120 10072 4126 10124
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10112 4583 10115
rect 4798 10112 4804 10124
rect 4571 10084 4804 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 5074 10072 5080 10124
rect 5132 10072 5138 10124
rect 842 10004 848 10056
rect 900 10004 906 10056
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4396 10016 4445 10044
rect 4396 10004 4402 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10044 4675 10047
rect 5184 10044 5212 10152
rect 5813 10149 5825 10152
rect 5859 10149 5871 10183
rect 7024 10180 7052 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 9122 10208 9128 10260
rect 9180 10248 9186 10260
rect 9309 10251 9367 10257
rect 9309 10248 9321 10251
rect 9180 10220 9321 10248
rect 9180 10208 9186 10220
rect 9309 10217 9321 10220
rect 9355 10248 9367 10251
rect 10229 10251 10287 10257
rect 10229 10248 10241 10251
rect 9355 10220 10241 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 10229 10217 10241 10220
rect 10275 10217 10287 10251
rect 10229 10211 10287 10217
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 11330 10248 11336 10260
rect 10468 10220 11336 10248
rect 10468 10208 10474 10220
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 12400 10208 12434 10248
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12713 10251 12771 10257
rect 12713 10248 12725 10251
rect 12584 10220 12725 10248
rect 12584 10208 12590 10220
rect 12713 10217 12725 10220
rect 12759 10217 12771 10251
rect 12713 10211 12771 10217
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13633 10251 13691 10257
rect 13633 10248 13645 10251
rect 12860 10220 13645 10248
rect 12860 10208 12866 10220
rect 13633 10217 13645 10220
rect 13679 10248 13691 10251
rect 13814 10248 13820 10260
rect 13679 10220 13820 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14369 10251 14427 10257
rect 14369 10217 14381 10251
rect 14415 10248 14427 10251
rect 15194 10248 15200 10260
rect 14415 10220 15200 10248
rect 14415 10217 14427 10220
rect 14369 10211 14427 10217
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 16669 10251 16727 10257
rect 15344 10220 16436 10248
rect 15344 10208 15350 10220
rect 5813 10143 5871 10149
rect 5920 10152 7052 10180
rect 7101 10183 7159 10189
rect 5258 10072 5264 10124
rect 5316 10072 5322 10124
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5718 10112 5724 10124
rect 5399 10084 5724 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5718 10072 5724 10084
rect 5776 10112 5782 10124
rect 5920 10112 5948 10152
rect 7101 10149 7113 10183
rect 7147 10180 7159 10183
rect 7466 10180 7472 10192
rect 7147 10152 7472 10180
rect 7147 10149 7159 10152
rect 7101 10143 7159 10149
rect 7466 10140 7472 10152
rect 7524 10180 7530 10192
rect 10597 10183 10655 10189
rect 10597 10180 10609 10183
rect 7524 10152 7604 10180
rect 7524 10140 7530 10152
rect 5776 10084 5948 10112
rect 6457 10115 6515 10121
rect 5776 10072 5782 10084
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 6822 10112 6828 10124
rect 6503 10084 6828 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7576 10121 7604 10152
rect 8220 10152 9628 10180
rect 8220 10121 8248 10152
rect 8956 10121 8984 10152
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 7248 10084 7297 10112
rect 7248 10072 7254 10084
rect 7285 10081 7297 10084
rect 7331 10112 7343 10115
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 7331 10084 7389 10112
rect 7331 10081 7343 10084
rect 7285 10075 7343 10081
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 7561 10115 7619 10121
rect 7561 10081 7573 10115
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10081 8263 10115
rect 8205 10075 8263 10081
rect 8343 10115 8401 10121
rect 8343 10081 8355 10115
rect 8389 10112 8401 10115
rect 8941 10115 8999 10121
rect 8389 10084 8892 10112
rect 8389 10081 8401 10084
rect 8343 10075 8401 10081
rect 4663 10016 5212 10044
rect 5629 10047 5687 10053
rect 4663 10013 4675 10016
rect 4617 10007 4675 10013
rect 5629 10013 5641 10047
rect 5675 10044 5687 10047
rect 6086 10044 6092 10056
rect 5675 10016 6092 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 3697 9979 3755 9985
rect 3697 9945 3709 9979
rect 3743 9976 3755 9979
rect 4246 9976 4252 9988
rect 3743 9948 4252 9976
rect 3743 9945 3755 9948
rect 3697 9939 3755 9945
rect 4246 9936 4252 9948
rect 4304 9976 4310 9988
rect 4632 9976 4660 10007
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6328 10016 6561 10044
rect 6328 10004 6334 10016
rect 6549 10013 6561 10016
rect 6595 10044 6607 10047
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 6595 10016 7481 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 4304 9948 4660 9976
rect 4304 9936 4310 9948
rect 5166 9936 5172 9988
rect 5224 9976 5230 9988
rect 6181 9979 6239 9985
rect 5224 9948 6040 9976
rect 5224 9936 5230 9948
rect 2225 9911 2283 9917
rect 2225 9877 2237 9911
rect 2271 9908 2283 9911
rect 2682 9908 2688 9920
rect 2271 9880 2688 9908
rect 2271 9877 2283 9880
rect 2225 9871 2283 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4525 9911 4583 9917
rect 4525 9908 4537 9911
rect 4212 9880 4537 9908
rect 4212 9868 4218 9880
rect 4525 9877 4537 9880
rect 4571 9908 4583 9911
rect 4798 9908 4804 9920
rect 4571 9880 4804 9908
rect 4571 9877 4583 9880
rect 4525 9871 4583 9877
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 6012 9917 6040 9948
rect 6181 9945 6193 9979
rect 6227 9976 6239 9979
rect 8496 9976 8524 10007
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 6227 9948 8524 9976
rect 8864 9976 8892 10084
rect 8941 10081 8953 10115
rect 8987 10081 8999 10115
rect 8941 10075 8999 10081
rect 9214 10072 9220 10124
rect 9272 10072 9278 10124
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10112 9551 10115
rect 9600 10112 9628 10152
rect 10336 10152 10609 10180
rect 10336 10124 10364 10152
rect 10597 10149 10609 10152
rect 10643 10149 10655 10183
rect 10597 10143 10655 10149
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 11210 10183 11268 10189
rect 11210 10180 11222 10183
rect 10836 10152 11222 10180
rect 10836 10140 10842 10152
rect 11210 10149 11222 10152
rect 11256 10149 11268 10183
rect 11210 10143 11268 10149
rect 11606 10140 11612 10192
rect 11664 10180 11670 10192
rect 12406 10180 12434 10208
rect 16408 10180 16436 10220
rect 16669 10217 16681 10251
rect 16715 10248 16727 10251
rect 17586 10248 17592 10260
rect 16715 10220 17592 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 16853 10183 16911 10189
rect 16853 10180 16865 10183
rect 11664 10152 12112 10180
rect 12406 10152 16344 10180
rect 16408 10152 16865 10180
rect 11664 10140 11670 10152
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9539 10084 9689 10112
rect 9539 10081 9551 10084
rect 9493 10075 9551 10081
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 10008 10084 10057 10112
rect 10008 10072 10014 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10318 10072 10324 10124
rect 10376 10072 10382 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10468 10084 10517 10112
rect 10468 10072 10474 10084
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10686 10072 10692 10124
rect 10744 10072 10750 10124
rect 10962 10072 10968 10124
rect 11020 10072 11026 10124
rect 12084 10112 12112 10152
rect 12912 10121 12940 10152
rect 12621 10115 12679 10121
rect 12621 10112 12633 10115
rect 11072 10084 12020 10112
rect 12084 10084 12633 10112
rect 9122 10004 9128 10056
rect 9180 10004 9186 10056
rect 9232 10044 9260 10072
rect 11072 10044 11100 10084
rect 9232 10016 11100 10044
rect 11992 10044 12020 10084
rect 12621 10081 12633 10084
rect 12667 10081 12679 10115
rect 12621 10075 12679 10081
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 13464 10044 13492 10075
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 13596 10084 14197 10112
rect 13596 10072 13602 10084
rect 14185 10081 14197 10084
rect 14231 10081 14243 10115
rect 14185 10075 14243 10081
rect 14458 10072 14464 10124
rect 14516 10112 14522 10124
rect 15286 10112 15292 10124
rect 14516 10084 15292 10112
rect 14516 10072 14522 10084
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15396 10121 15424 10152
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10081 15439 10115
rect 15381 10075 15439 10081
rect 15657 10115 15715 10121
rect 15657 10081 15669 10115
rect 15703 10112 15715 10115
rect 15746 10112 15752 10124
rect 15703 10084 15752 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 16316 10121 16344 10152
rect 16853 10149 16865 10152
rect 16899 10149 16911 10183
rect 16853 10143 16911 10149
rect 15841 10115 15899 10121
rect 15841 10081 15853 10115
rect 15887 10081 15899 10115
rect 15841 10075 15899 10081
rect 15933 10115 15991 10121
rect 15933 10081 15945 10115
rect 15979 10112 15991 10115
rect 16301 10115 16359 10121
rect 15979 10084 16068 10112
rect 15979 10081 15991 10084
rect 15933 10075 15991 10081
rect 13906 10044 13912 10056
rect 11992 10016 13912 10044
rect 13906 10004 13912 10016
rect 13964 10004 13970 10056
rect 14001 10047 14059 10053
rect 14001 10013 14013 10047
rect 14047 10044 14059 10047
rect 14734 10044 14740 10056
rect 14047 10016 14740 10044
rect 14047 10013 14059 10016
rect 14001 10007 14059 10013
rect 14734 10004 14740 10016
rect 14792 10044 14798 10056
rect 15102 10044 15108 10056
rect 14792 10016 15108 10044
rect 14792 10004 14798 10016
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15856 10044 15884 10075
rect 16040 10056 16068 10084
rect 16301 10081 16313 10115
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 16758 10072 16764 10124
rect 16816 10072 16822 10124
rect 16945 10115 17003 10121
rect 16945 10081 16957 10115
rect 16991 10081 17003 10115
rect 16945 10075 17003 10081
rect 15304 10016 15884 10044
rect 12342 9976 12348 9988
rect 8864 9948 11008 9976
rect 6227 9945 6239 9948
rect 6181 9939 6239 9945
rect 5997 9911 6055 9917
rect 5997 9877 6009 9911
rect 6043 9877 6055 9911
rect 5997 9871 6055 9877
rect 6733 9911 6791 9917
rect 6733 9877 6745 9911
rect 6779 9908 6791 9911
rect 7098 9908 7104 9920
rect 6779 9880 7104 9908
rect 6779 9877 6791 9880
rect 6733 9871 6791 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 7984 9880 8769 9908
rect 7984 9868 7990 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8864 9908 8892 9948
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8864 9880 8953 9908
rect 8757 9871 8815 9877
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 8941 9871 8999 9877
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9950 9908 9956 9920
rect 9732 9880 9956 9908
rect 9732 9868 9738 9880
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 10042 9868 10048 9920
rect 10100 9868 10106 9920
rect 10410 9868 10416 9920
rect 10468 9908 10474 9920
rect 10778 9908 10784 9920
rect 10468 9880 10784 9908
rect 10468 9868 10474 9880
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 10980 9908 11008 9948
rect 11900 9948 12348 9976
rect 11900 9908 11928 9948
rect 12342 9936 12348 9948
rect 12400 9976 12406 9988
rect 15304 9985 15332 10016
rect 16022 10004 16028 10056
rect 16080 10044 16086 10056
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 16080 10016 16221 10044
rect 16080 10004 16086 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16960 10044 16988 10075
rect 17034 10072 17040 10124
rect 17092 10072 17098 10124
rect 16960 10016 17172 10044
rect 16209 10007 16267 10013
rect 15289 9979 15347 9985
rect 15289 9976 15301 9979
rect 12400 9948 15301 9976
rect 12400 9936 12406 9948
rect 15289 9945 15301 9948
rect 15335 9945 15347 9979
rect 15289 9939 15347 9945
rect 17144 9920 17172 10016
rect 10980 9880 11928 9908
rect 12434 9868 12440 9920
rect 12492 9868 12498 9920
rect 15470 9868 15476 9920
rect 15528 9868 15534 9920
rect 17126 9868 17132 9920
rect 17184 9868 17190 9920
rect 552 9818 17664 9840
rect 552 9766 1366 9818
rect 1418 9766 1430 9818
rect 1482 9766 1494 9818
rect 1546 9766 1558 9818
rect 1610 9766 1622 9818
rect 1674 9766 1686 9818
rect 1738 9766 7366 9818
rect 7418 9766 7430 9818
rect 7482 9766 7494 9818
rect 7546 9766 7558 9818
rect 7610 9766 7622 9818
rect 7674 9766 7686 9818
rect 7738 9766 13366 9818
rect 13418 9766 13430 9818
rect 13482 9766 13494 9818
rect 13546 9766 13558 9818
rect 13610 9766 13622 9818
rect 13674 9766 13686 9818
rect 13738 9766 17664 9818
rect 552 9744 17664 9766
rect 4154 9664 4160 9716
rect 4212 9664 4218 9716
rect 4249 9707 4307 9713
rect 4249 9673 4261 9707
rect 4295 9704 4307 9707
rect 5258 9704 5264 9716
rect 4295 9676 5264 9704
rect 4295 9673 4307 9676
rect 4249 9667 4307 9673
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 9766 9704 9772 9716
rect 5868 9676 9772 9704
rect 5868 9664 5874 9676
rect 9766 9664 9772 9676
rect 9824 9704 9830 9716
rect 11606 9704 11612 9716
rect 9824 9676 11612 9704
rect 9824 9664 9830 9676
rect 11606 9664 11612 9676
rect 11664 9704 11670 9716
rect 11885 9707 11943 9713
rect 11885 9704 11897 9707
rect 11664 9676 11897 9704
rect 11664 9664 11670 9676
rect 11885 9673 11897 9676
rect 11931 9673 11943 9707
rect 11885 9667 11943 9673
rect 12342 9664 12348 9716
rect 12400 9704 12406 9716
rect 12437 9707 12495 9713
rect 12437 9704 12449 9707
rect 12400 9676 12449 9704
rect 12400 9664 12406 9676
rect 12437 9673 12449 9676
rect 12483 9673 12495 9707
rect 12437 9667 12495 9673
rect 13173 9707 13231 9713
rect 13173 9673 13185 9707
rect 13219 9673 13231 9707
rect 13173 9667 13231 9673
rect 2501 9639 2559 9645
rect 2501 9636 2513 9639
rect 1964 9608 2513 9636
rect 1964 9580 1992 9608
rect 2501 9605 2513 9608
rect 2547 9636 2559 9639
rect 3878 9636 3884 9648
rect 2547 9608 3884 9636
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 3973 9639 4031 9645
rect 3973 9605 3985 9639
rect 4019 9636 4031 9639
rect 4172 9636 4200 9664
rect 4019 9608 4200 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 5718 9596 5724 9648
rect 5776 9636 5782 9648
rect 6638 9636 6644 9648
rect 5776 9608 6644 9636
rect 5776 9596 5782 9608
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 6822 9596 6828 9648
rect 6880 9636 6886 9648
rect 7190 9636 7196 9648
rect 6880 9608 7196 9636
rect 6880 9596 6886 9608
rect 7190 9596 7196 9608
rect 7248 9596 7254 9648
rect 9122 9596 9128 9648
rect 9180 9636 9186 9648
rect 10226 9636 10232 9648
rect 9180 9608 10232 9636
rect 9180 9596 9186 9608
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 10410 9596 10416 9648
rect 10468 9596 10474 9648
rect 13188 9636 13216 9667
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 13964 9676 17448 9704
rect 13964 9664 13970 9676
rect 13102 9608 13216 9636
rect 1946 9528 1952 9580
rect 2004 9528 2010 9580
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2280 9540 2697 9568
rect 2280 9528 2286 9540
rect 2685 9537 2697 9540
rect 2731 9568 2743 9571
rect 3510 9568 3516 9580
rect 2731 9540 3516 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 5166 9568 5172 9580
rect 3804 9540 5172 9568
rect 3804 9512 3832 9540
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 6380 9540 6929 9568
rect 6380 9512 6408 9540
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9950 9568 9956 9580
rect 9364 9540 9956 9568
rect 9364 9528 9370 9540
rect 9950 9528 9956 9540
rect 10008 9568 10014 9580
rect 13102 9568 13130 9608
rect 14274 9596 14280 9648
rect 14332 9596 14338 9648
rect 16209 9639 16267 9645
rect 16209 9605 16221 9639
rect 16255 9636 16267 9639
rect 17034 9636 17040 9648
rect 16255 9608 17040 9636
rect 16255 9605 16267 9608
rect 16209 9599 16267 9605
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 10008 9540 10088 9568
rect 10008 9528 10014 9540
rect 842 9460 848 9512
rect 900 9460 906 9512
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2593 9503 2651 9509
rect 2593 9500 2605 9503
rect 2363 9472 2605 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2593 9469 2605 9472
rect 2639 9469 2651 9503
rect 2593 9463 2651 9469
rect 1112 9435 1170 9441
rect 1112 9401 1124 9435
rect 1158 9432 1170 9435
rect 1854 9432 1860 9444
rect 1158 9404 1860 9432
rect 1158 9401 1170 9404
rect 1112 9395 1170 9401
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 2608 9364 2636 9463
rect 3786 9460 3792 9512
rect 3844 9460 3850 9512
rect 4062 9460 4068 9512
rect 4120 9460 4126 9512
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4212 9472 4261 9500
rect 4212 9460 4218 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 5258 9500 5264 9512
rect 4580 9472 5264 9500
rect 4580 9460 4586 9472
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4614 9432 4620 9444
rect 3936 9404 4620 9432
rect 3936 9392 3942 9404
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 4724 9364 4752 9472
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 6178 9460 6184 9512
rect 6236 9460 6242 9512
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 6454 9460 6460 9512
rect 6512 9460 6518 9512
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 9030 9500 9036 9512
rect 6696 9472 9036 9500
rect 6696 9460 6702 9472
rect 9030 9460 9036 9472
rect 9088 9500 9094 9512
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 9088 9472 9137 9500
rect 9088 9460 9094 9472
rect 9125 9469 9137 9472
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9766 9460 9772 9512
rect 9824 9460 9830 9512
rect 10060 9509 10088 9540
rect 12360 9540 13130 9568
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 10134 9460 10140 9512
rect 10192 9460 10198 9512
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9500 10287 9503
rect 10318 9500 10324 9512
rect 10275 9472 10324 9500
rect 10275 9469 10287 9472
rect 10229 9463 10287 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9500 10563 9503
rect 11054 9500 11060 9512
rect 10551 9472 11060 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 12250 9500 12256 9512
rect 11756 9472 12256 9500
rect 11756 9460 11762 9472
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 12360 9509 12388 9540
rect 13262 9528 13268 9580
rect 13320 9568 13326 9580
rect 14292 9568 14320 9596
rect 17420 9580 17448 9676
rect 16761 9571 16819 9577
rect 16761 9568 16773 9571
rect 13320 9540 13584 9568
rect 13320 9528 13326 9540
rect 12345 9503 12403 9509
rect 12345 9469 12357 9503
rect 12391 9469 12403 9503
rect 12345 9463 12403 9469
rect 12621 9479 12679 9485
rect 6549 9435 6607 9441
rect 6549 9432 6561 9435
rect 6196 9404 6561 9432
rect 6196 9376 6224 9404
rect 6549 9401 6561 9404
rect 6595 9401 6607 9435
rect 6549 9395 6607 9401
rect 6730 9392 6736 9444
rect 6788 9441 6794 9444
rect 6788 9435 6817 9441
rect 6805 9401 6817 9435
rect 9927 9435 9985 9441
rect 9927 9432 9939 9435
rect 6788 9395 6817 9401
rect 6932 9404 9939 9432
rect 6788 9392 6794 9395
rect 6932 9376 6960 9404
rect 9927 9401 9939 9404
rect 9973 9432 9985 9435
rect 10761 9435 10819 9441
rect 9973 9404 10272 9432
rect 9973 9401 9985 9404
rect 9927 9395 9985 9401
rect 10244 9376 10272 9404
rect 10761 9401 10773 9435
rect 10807 9401 10819 9435
rect 10761 9395 10819 9401
rect 2271 9336 4752 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 4890 9324 4896 9376
rect 4948 9324 4954 9376
rect 6178 9324 6184 9376
rect 6236 9324 6242 9376
rect 6270 9324 6276 9376
rect 6328 9324 6334 9376
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 6914 9364 6920 9376
rect 6696 9336 6920 9364
rect 6696 9324 6702 9336
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 9306 9364 9312 9376
rect 7340 9336 9312 9364
rect 7340 9324 7346 9336
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 10226 9324 10232 9376
rect 10284 9324 10290 9376
rect 10787 9364 10815 9395
rect 12360 9376 12388 9463
rect 12621 9445 12633 9479
rect 12667 9445 12679 9479
rect 12802 9460 12808 9512
rect 12860 9500 12866 9512
rect 13556 9509 13584 9540
rect 14108 9540 14320 9568
rect 16224 9540 16773 9568
rect 14108 9509 14136 9540
rect 16224 9512 16252 9540
rect 16761 9537 16773 9540
rect 16807 9537 16819 9571
rect 16761 9531 16819 9537
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 13357 9503 13415 9509
rect 13357 9500 13369 9503
rect 12860 9472 13369 9500
rect 12860 9460 12866 9472
rect 13357 9469 13369 9472
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 14274 9460 14280 9512
rect 14332 9460 14338 9512
rect 14366 9460 14372 9512
rect 14424 9460 14430 9512
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 14918 9500 14924 9512
rect 14875 9472 14924 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 16206 9460 16212 9512
rect 16264 9460 16270 9512
rect 16485 9503 16543 9509
rect 16485 9469 16497 9503
rect 16531 9469 16543 9503
rect 16485 9463 16543 9469
rect 12621 9444 12679 9445
rect 12529 9435 12587 9441
rect 12529 9401 12541 9435
rect 12575 9401 12587 9435
rect 12529 9395 12587 9401
rect 11054 9364 11060 9376
rect 10787 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11204 9336 12081 9364
rect 11204 9324 11210 9336
rect 12069 9333 12081 9336
rect 12115 9333 12127 9367
rect 12069 9327 12127 9333
rect 12342 9324 12348 9376
rect 12400 9324 12406 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12544 9364 12572 9395
rect 12618 9392 12624 9444
rect 12676 9392 12682 9444
rect 13725 9435 13783 9441
rect 13725 9432 13737 9435
rect 12820 9404 13737 9432
rect 12820 9376 12848 9404
rect 13725 9401 13737 9404
rect 13771 9401 13783 9435
rect 13725 9395 13783 9401
rect 14737 9435 14795 9441
rect 14737 9401 14749 9435
rect 14783 9432 14795 9435
rect 15074 9435 15132 9441
rect 15074 9432 15086 9435
rect 14783 9404 15086 9432
rect 14783 9401 14795 9404
rect 14737 9395 14795 9401
rect 15074 9401 15086 9404
rect 15120 9401 15132 9435
rect 16500 9432 16528 9463
rect 16500 9404 16896 9432
rect 15074 9395 15132 9401
rect 16868 9376 16896 9404
rect 12492 9336 12572 9364
rect 12492 9324 12498 9336
rect 12802 9324 12808 9376
rect 12860 9324 12866 9376
rect 13909 9367 13967 9373
rect 13909 9333 13921 9367
rect 13955 9364 13967 9367
rect 13998 9364 14004 9376
rect 13955 9336 14004 9364
rect 13955 9333 13967 9336
rect 13909 9327 13967 9333
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 14550 9364 14556 9376
rect 14424 9336 14556 9364
rect 14424 9324 14430 9336
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 552 9274 17664 9296
rect 552 9222 4366 9274
rect 4418 9222 4430 9274
rect 4482 9222 4494 9274
rect 4546 9222 4558 9274
rect 4610 9222 4622 9274
rect 4674 9222 4686 9274
rect 4738 9222 10366 9274
rect 10418 9222 10430 9274
rect 10482 9222 10494 9274
rect 10546 9222 10558 9274
rect 10610 9222 10622 9274
rect 10674 9222 10686 9274
rect 10738 9222 16366 9274
rect 16418 9222 16430 9274
rect 16482 9222 16494 9274
rect 16546 9222 16558 9274
rect 16610 9222 16622 9274
rect 16674 9222 16686 9274
rect 16738 9222 17664 9274
rect 552 9200 17664 9222
rect 3145 9163 3203 9169
rect 3145 9129 3157 9163
rect 3191 9160 3203 9163
rect 4154 9160 4160 9172
rect 3191 9132 4160 9160
rect 3191 9129 3203 9132
rect 3145 9123 3203 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4890 9120 4896 9172
rect 4948 9120 4954 9172
rect 6178 9120 6184 9172
rect 6236 9120 6242 9172
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 6512 9132 7481 9160
rect 6512 9120 6518 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 9950 9120 9956 9172
rect 10008 9120 10014 9172
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10689 9163 10747 9169
rect 10192 9132 10640 9160
rect 10192 9120 10198 9132
rect 1780 9064 4660 9092
rect 842 8984 848 9036
rect 900 9024 906 9036
rect 1780 9033 1808 9064
rect 1765 9027 1823 9033
rect 1765 9024 1777 9027
rect 900 8996 1777 9024
rect 900 8984 906 8996
rect 1765 8993 1777 8996
rect 1811 8993 1823 9027
rect 1765 8987 1823 8993
rect 2032 9027 2090 9033
rect 2032 8993 2044 9027
rect 2078 9024 2090 9027
rect 2590 9024 2596 9036
rect 2078 8996 2596 9024
rect 2078 8993 2090 8996
rect 2032 8987 2090 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 3786 9024 3792 9036
rect 3620 8996 3792 9024
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8888 3295 8891
rect 3620 8888 3648 8996
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 4632 9033 4660 9064
rect 4361 9027 4419 9033
rect 4361 8993 4373 9027
rect 4407 9024 4419 9027
rect 4617 9027 4675 9033
rect 4407 8996 4568 9024
rect 4407 8993 4419 8996
rect 4361 8987 4419 8993
rect 4540 8956 4568 8996
rect 4617 8993 4629 9027
rect 4663 9024 4675 9027
rect 4908 9024 4936 9120
rect 7009 9095 7067 9101
rect 6104 9064 6868 9092
rect 4663 8996 4936 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 6104 9033 6132 9064
rect 6840 9036 6868 9064
rect 7009 9061 7021 9095
rect 7055 9092 7067 9095
rect 7282 9092 7288 9104
rect 7055 9064 7288 9092
rect 7055 9061 7067 9064
rect 7009 9055 7067 9061
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 8938 9052 8944 9104
rect 8996 9052 9002 9104
rect 9122 9052 9128 9104
rect 9180 9092 9186 9104
rect 9968 9092 9996 9120
rect 10612 9092 10640 9132
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 11054 9160 11060 9172
rect 10735 9132 11060 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 13872 9132 14228 9160
rect 13872 9120 13878 9132
rect 10965 9095 11023 9101
rect 10965 9092 10977 9095
rect 9180 9064 9628 9092
rect 9968 9064 10272 9092
rect 10612 9064 10977 9092
rect 9180 9052 9186 9064
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5592 8996 5917 9024
rect 5592 8984 5598 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 8993 6147 9027
rect 6089 8987 6147 8993
rect 4709 8959 4767 8965
rect 4540 8928 4660 8956
rect 3283 8860 3648 8888
rect 4632 8888 4660 8928
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 4798 8956 4804 8968
rect 4755 8928 4804 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5166 8956 5172 8968
rect 5031 8928 5172 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 5920 8956 5948 8987
rect 6362 8984 6368 9036
rect 6420 8984 6426 9036
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 9024 6607 9027
rect 6730 9024 6736 9036
rect 6595 8996 6736 9024
rect 6595 8993 6607 8996
rect 6549 8987 6607 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6822 8984 6828 9036
rect 6880 8984 6886 9036
rect 6914 8984 6920 9036
rect 6972 8984 6978 9036
rect 7127 9027 7185 9033
rect 7127 9024 7139 9027
rect 7024 8996 7139 9024
rect 5920 8928 6408 8956
rect 6270 8888 6276 8900
rect 4632 8860 6276 8888
rect 3283 8857 3295 8860
rect 3237 8851 3295 8857
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 6380 8888 6408 8928
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 7024 8956 7052 8996
rect 7127 8993 7139 8996
rect 7173 8993 7185 9027
rect 7127 8987 7185 8993
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 6696 8928 7052 8956
rect 6696 8916 6702 8928
rect 7282 8916 7288 8968
rect 7340 8916 7346 8968
rect 6380 8860 6776 8888
rect 6086 8780 6092 8832
rect 6144 8780 6150 8832
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 6512 8792 6653 8820
rect 6512 8780 6518 8792
rect 6641 8789 6653 8792
rect 6687 8789 6699 8823
rect 6748 8820 6776 8860
rect 7098 8848 7104 8900
rect 7156 8888 7162 8900
rect 7392 8888 7420 8987
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 7892 8996 8033 9024
rect 7892 8984 7898 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 9232 8956 9260 8987
rect 9306 8984 9312 9036
rect 9364 8984 9370 9036
rect 9600 9033 9628 9064
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 9585 9027 9643 9033
rect 9585 8993 9597 9027
rect 9631 9024 9643 9027
rect 9631 8996 9996 9024
rect 9631 8993 9643 8996
rect 9585 8987 9643 8993
rect 9416 8956 9444 8987
rect 9766 8956 9772 8968
rect 8343 8928 8524 8956
rect 9232 8928 9352 8956
rect 9416 8928 9772 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8496 8900 8524 8928
rect 7156 8860 7420 8888
rect 7156 8848 7162 8860
rect 8478 8848 8484 8900
rect 8536 8848 8542 8900
rect 9324 8888 9352 8928
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 9968 8956 9996 8996
rect 10042 8984 10048 9036
rect 10100 9022 10106 9036
rect 10157 9027 10215 9033
rect 10157 9024 10169 9027
rect 10152 9022 10169 9024
rect 10100 8994 10169 9022
rect 10100 8984 10106 8994
rect 10157 8993 10169 8994
rect 10203 8993 10215 9027
rect 10244 9024 10272 9064
rect 10965 9061 10977 9064
rect 11011 9061 11023 9095
rect 11160 9095 11218 9101
rect 11160 9092 11172 9095
rect 10965 9055 11023 9061
rect 11096 9064 11172 9092
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 10244 8996 10333 9024
rect 10157 8987 10215 8993
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 10410 8984 10416 9036
rect 10468 8984 10474 9036
rect 10502 8984 10508 9036
rect 10560 8984 10566 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 11096 9024 11124 9064
rect 11160 9061 11172 9064
rect 11206 9061 11218 9095
rect 11160 9055 11218 9061
rect 11330 9052 11336 9104
rect 11388 9092 11394 9104
rect 11577 9095 11635 9101
rect 11577 9092 11589 9095
rect 11388 9064 11589 9092
rect 11388 9052 11394 9064
rect 11577 9061 11589 9064
rect 11623 9061 11635 9095
rect 11577 9055 11635 9061
rect 11698 9052 11704 9104
rect 11756 9092 11762 9104
rect 11793 9095 11851 9101
rect 11793 9092 11805 9095
rect 11756 9064 11805 9092
rect 11756 9052 11762 9064
rect 11793 9061 11805 9064
rect 11839 9061 11851 9095
rect 12434 9092 12440 9104
rect 11793 9055 11851 9061
rect 12360 9064 12440 9092
rect 12066 9024 12072 9036
rect 10836 8996 11124 9024
rect 11225 9008 12072 9024
rect 11164 8996 12072 9008
rect 10836 8984 10842 8996
rect 11164 8980 11253 8996
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 12360 9033 12388 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 8993 12403 9027
rect 12345 8987 12403 8993
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 9024 12587 9027
rect 12710 9024 12716 9036
rect 12575 8996 12716 9024
rect 12575 8993 12587 8996
rect 12529 8987 12587 8993
rect 11164 8956 11192 8980
rect 12544 8956 12572 8987
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 12802 9008 12808 9060
rect 12860 9024 12866 9060
rect 13170 9052 13176 9104
rect 13228 9092 13234 9104
rect 13906 9092 13912 9104
rect 13228 9064 13912 9092
rect 13228 9052 13234 9064
rect 13906 9052 13912 9064
rect 13964 9092 13970 9104
rect 13964 9064 14136 9092
rect 13964 9052 13970 9064
rect 12897 9027 12955 9033
rect 12897 9024 12909 9027
rect 12860 9008 12909 9024
rect 12820 8996 12909 9008
rect 12897 8993 12909 8996
rect 12943 9024 12955 9027
rect 13814 9024 13820 9036
rect 12943 8996 13820 9024
rect 12943 8993 12955 8996
rect 12897 8987 12955 8993
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 14108 9033 14136 9064
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 8993 14151 9027
rect 14200 9024 14228 9132
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 15105 9163 15163 9169
rect 15105 9160 15117 9163
rect 14332 9132 15117 9160
rect 14332 9120 14338 9132
rect 15105 9129 15117 9132
rect 15151 9129 15163 9163
rect 15105 9123 15163 9129
rect 15841 9163 15899 9169
rect 15841 9129 15853 9163
rect 15887 9160 15899 9163
rect 16758 9160 16764 9172
rect 15887 9132 16764 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 16758 9120 16764 9132
rect 16816 9120 16822 9172
rect 17034 9120 17040 9172
rect 17092 9120 17098 9172
rect 14550 9024 14556 9036
rect 14200 8996 14556 9024
rect 14093 8987 14151 8993
rect 14550 8984 14556 8996
rect 14608 9024 14614 9036
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 14608 8996 14749 9024
rect 14608 8984 14614 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 15189 9027 15247 9033
rect 15189 9024 15201 9027
rect 14737 8987 14795 8993
rect 15120 8996 15201 9024
rect 9968 8928 11192 8956
rect 11348 8928 12572 8956
rect 11348 8888 11376 8928
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 12860 8928 13185 8956
rect 12860 8916 12866 8928
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 9324 8860 11376 8888
rect 9324 8820 9352 8860
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 12529 8891 12587 8897
rect 12529 8888 12541 8891
rect 12308 8860 12541 8888
rect 12308 8848 12314 8860
rect 12529 8857 12541 8860
rect 12575 8888 12587 8891
rect 12575 8860 14412 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 6748 8792 9352 8820
rect 6641 8783 6699 8789
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 9732 8792 11437 8820
rect 9732 8780 9738 8792
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11425 8783 11483 8789
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 12618 8820 12624 8832
rect 11655 8792 12624 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 14384 8820 14412 8860
rect 14458 8848 14464 8900
rect 14516 8888 14522 8900
rect 14921 8891 14979 8897
rect 14921 8888 14933 8891
rect 14516 8860 14933 8888
rect 14516 8848 14522 8860
rect 14921 8857 14933 8860
rect 14967 8857 14979 8891
rect 14921 8851 14979 8857
rect 15120 8820 15148 8996
rect 15189 8993 15201 8996
rect 15235 8993 15247 9027
rect 15189 8987 15247 8993
rect 15746 8984 15752 9036
rect 15804 8984 15810 9036
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16850 9024 16856 9036
rect 15979 8996 16856 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 17052 9033 17080 9120
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 8993 17095 9027
rect 17037 8987 17095 8993
rect 15764 8956 15792 8984
rect 16022 8956 16028 8968
rect 15764 8928 16028 8956
rect 16022 8916 16028 8928
rect 16080 8956 16086 8968
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 16080 8928 16681 8956
rect 16080 8916 16086 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 16945 8959 17003 8965
rect 16945 8925 16957 8959
rect 16991 8956 17003 8959
rect 17126 8956 17132 8968
rect 16991 8928 17132 8956
rect 16991 8925 17003 8928
rect 16945 8919 17003 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 15194 8820 15200 8832
rect 14384 8792 15200 8820
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 17126 8780 17132 8832
rect 17184 8820 17190 8832
rect 17221 8823 17279 8829
rect 17221 8820 17233 8823
rect 17184 8792 17233 8820
rect 17184 8780 17190 8792
rect 17221 8789 17233 8792
rect 17267 8820 17279 8823
rect 17402 8820 17408 8832
rect 17267 8792 17408 8820
rect 17267 8789 17279 8792
rect 17221 8783 17279 8789
rect 17402 8780 17408 8792
rect 17460 8780 17466 8832
rect 552 8730 17664 8752
rect 552 8678 1366 8730
rect 1418 8678 1430 8730
rect 1482 8678 1494 8730
rect 1546 8678 1558 8730
rect 1610 8678 1622 8730
rect 1674 8678 1686 8730
rect 1738 8678 7366 8730
rect 7418 8678 7430 8730
rect 7482 8678 7494 8730
rect 7546 8678 7558 8730
rect 7610 8678 7622 8730
rect 7674 8678 7686 8730
rect 7738 8678 13366 8730
rect 13418 8678 13430 8730
rect 13482 8678 13494 8730
rect 13546 8678 13558 8730
rect 13610 8678 13622 8730
rect 13674 8678 13686 8730
rect 13738 8678 17664 8730
rect 552 8656 17664 8678
rect 845 8619 903 8625
rect 845 8585 857 8619
rect 891 8616 903 8619
rect 3142 8616 3148 8628
rect 891 8588 3148 8616
rect 891 8585 903 8588
rect 845 8579 903 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 5534 8576 5540 8628
rect 5592 8576 5598 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 6086 8576 6092 8628
rect 6144 8616 6150 8628
rect 6273 8619 6331 8625
rect 6273 8616 6285 8619
rect 6144 8588 6285 8616
rect 6144 8576 6150 8588
rect 6273 8585 6285 8588
rect 6319 8585 6331 8619
rect 6273 8579 6331 8585
rect 6822 8576 6828 8628
rect 6880 8576 6886 8628
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7653 8619 7711 8625
rect 7653 8616 7665 8619
rect 6972 8588 7665 8616
rect 6972 8576 6978 8588
rect 7653 8585 7665 8588
rect 7699 8585 7711 8619
rect 7653 8579 7711 8585
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9364 8588 9505 8616
rect 9364 8576 9370 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 9766 8576 9772 8628
rect 9824 8576 9830 8628
rect 12342 8576 12348 8628
rect 12400 8616 12406 8628
rect 13170 8616 13176 8628
rect 12400 8588 13176 8616
rect 12400 8576 12406 8588
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 16908 8588 17325 8616
rect 16908 8576 16914 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 2746 8520 5856 8548
rect 842 8440 848 8492
rect 900 8440 906 8492
rect 860 8412 888 8440
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 860 8384 2237 8412
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 1980 8347 2038 8353
rect 1980 8313 1992 8347
rect 2026 8344 2038 8347
rect 2746 8344 2774 8520
rect 3970 8440 3976 8492
rect 4028 8480 4034 8492
rect 5828 8489 5856 8520
rect 5902 8508 5908 8560
rect 5960 8548 5966 8560
rect 6641 8551 6699 8557
rect 5960 8520 6592 8548
rect 5960 8508 5966 8520
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 4028 8452 5089 8480
rect 4028 8440 4034 8452
rect 5077 8449 5089 8452
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 6457 8483 6515 8489
rect 6457 8480 6469 8483
rect 5813 8443 5871 8449
rect 6012 8452 6469 8480
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 4801 8415 4859 8421
rect 3936 8384 4186 8412
rect 3936 8372 3942 8384
rect 4801 8381 4813 8415
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 5626 8412 5632 8424
rect 5583 8384 5632 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 2026 8316 2774 8344
rect 2026 8313 2038 8316
rect 1980 8307 2038 8313
rect 3786 8304 3792 8356
rect 3844 8304 3850 8356
rect 4816 8344 4844 8375
rect 5184 8344 5212 8375
rect 5626 8372 5632 8384
rect 5684 8412 5690 8424
rect 5902 8412 5908 8424
rect 5684 8384 5908 8412
rect 5684 8372 5690 8384
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 6012 8421 6040 8452
rect 6457 8449 6469 8452
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 5997 8415 6055 8421
rect 5997 8381 6009 8415
rect 6043 8381 6055 8415
rect 5997 8375 6055 8381
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8412 6423 8415
rect 6564 8412 6592 8520
rect 6641 8517 6653 8551
rect 6687 8517 6699 8551
rect 6840 8548 6868 8576
rect 7101 8551 7159 8557
rect 7101 8548 7113 8551
rect 6840 8520 7113 8548
rect 6641 8511 6699 8517
rect 7101 8517 7113 8520
rect 7147 8548 7159 8551
rect 7147 8520 7328 8548
rect 7147 8517 7159 8520
rect 7101 8511 7159 8517
rect 6411 8384 6592 8412
rect 6411 8381 6423 8384
rect 6365 8375 6423 8381
rect 4816 8316 5212 8344
rect 6104 8344 6132 8375
rect 6546 8344 6552 8356
rect 6104 8316 6552 8344
rect 5184 8288 5212 8316
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 6656 8344 6684 8511
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6788 8452 6929 8480
rect 6788 8440 6794 8452
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7006 8372 7012 8424
rect 7064 8372 7070 8424
rect 7300 8421 7328 8520
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 7852 8480 7880 8576
rect 10778 8508 10784 8560
rect 10836 8548 10842 8560
rect 11422 8548 11428 8560
rect 10836 8520 11428 8548
rect 10836 8508 10842 8520
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 7852 8452 8493 8480
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 7466 8372 7472 8424
rect 7524 8372 7530 8424
rect 7834 8414 7840 8424
rect 7760 8412 7840 8414
rect 7668 8386 7840 8412
rect 7668 8384 7788 8386
rect 6656 8316 7328 8344
rect 5166 8236 5172 8288
rect 5224 8236 5230 8288
rect 7300 8276 7328 8316
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 7668 8344 7696 8384
rect 7834 8372 7840 8386
rect 7892 8372 7898 8424
rect 7432 8316 7696 8344
rect 7432 8304 7438 8316
rect 7944 8276 7972 8452
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 9674 8480 9680 8492
rect 8481 8443 8539 8449
rect 8680 8452 9680 8480
rect 8110 8372 8116 8424
rect 8168 8412 8174 8424
rect 8680 8412 8708 8452
rect 8168 8384 8708 8412
rect 8757 8415 8815 8421
rect 8168 8372 8174 8384
rect 8757 8381 8769 8415
rect 8803 8412 8815 8415
rect 9122 8412 9128 8424
rect 8803 8384 9128 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9600 8421 9628 8452
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 10318 8480 10324 8492
rect 10060 8452 10324 8480
rect 10060 8424 10088 8452
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 12250 8480 12256 8492
rect 10428 8452 12256 8480
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 9416 8344 9444 8375
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 10042 8372 10048 8424
rect 10100 8372 10106 8424
rect 10428 8421 10456 8452
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 14976 8452 15945 8480
rect 14976 8440 14982 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8381 10471 8415
rect 10413 8375 10471 8381
rect 11698 8372 11704 8424
rect 11756 8412 11762 8424
rect 13541 8415 13599 8421
rect 11756 8384 11928 8412
rect 11756 8372 11762 8384
rect 9968 8344 9996 8372
rect 11900 8356 11928 8384
rect 13541 8381 13553 8415
rect 13587 8381 13599 8415
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 13541 8375 13599 8381
rect 13648 8384 13737 8412
rect 10226 8344 10232 8356
rect 8076 8316 9996 8344
rect 10152 8316 10232 8344
rect 8076 8304 8082 8316
rect 10152 8285 10180 8316
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 11241 8347 11299 8353
rect 11241 8313 11253 8347
rect 11287 8313 11299 8347
rect 11241 8307 11299 8313
rect 10137 8279 10195 8285
rect 10137 8276 10149 8279
rect 7300 8248 7972 8276
rect 10115 8248 10149 8276
rect 10137 8245 10149 8248
rect 10183 8245 10195 8279
rect 10137 8239 10195 8245
rect 10321 8279 10379 8285
rect 10321 8245 10333 8279
rect 10367 8276 10379 8279
rect 10962 8276 10968 8288
rect 10367 8248 10968 8276
rect 10367 8245 10379 8248
rect 10321 8239 10379 8245
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 11054 8236 11060 8288
rect 11112 8236 11118 8288
rect 11256 8276 11284 8307
rect 11422 8304 11428 8356
rect 11480 8304 11486 8356
rect 11882 8304 11888 8356
rect 11940 8304 11946 8356
rect 13556 8288 13584 8375
rect 13648 8288 13676 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 13725 8375 13783 8381
rect 13832 8384 13921 8412
rect 13832 8288 13860 8384
rect 13909 8381 13921 8384
rect 13955 8381 13967 8415
rect 13909 8375 13967 8381
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8412 14151 8415
rect 14182 8412 14188 8424
rect 14139 8384 14188 8412
rect 14139 8381 14151 8384
rect 14093 8375 14151 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 16200 8347 16258 8353
rect 14200 8316 14412 8344
rect 14200 8288 14228 8316
rect 14384 8288 14412 8316
rect 16200 8313 16212 8347
rect 16246 8344 16258 8347
rect 16758 8344 16764 8356
rect 16246 8316 16764 8344
rect 16246 8313 16258 8316
rect 16200 8307 16258 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 11517 8279 11575 8285
rect 11517 8276 11529 8279
rect 11256 8248 11529 8276
rect 11517 8245 11529 8248
rect 11563 8276 11575 8279
rect 12158 8276 12164 8288
rect 11563 8248 12164 8276
rect 11563 8245 11575 8248
rect 11517 8239 11575 8245
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 13538 8236 13544 8288
rect 13596 8236 13602 8288
rect 13630 8236 13636 8288
rect 13688 8236 13694 8288
rect 13814 8236 13820 8288
rect 13872 8236 13878 8288
rect 14182 8236 14188 8288
rect 14240 8236 14246 8288
rect 14274 8236 14280 8288
rect 14332 8236 14338 8288
rect 14366 8236 14372 8288
rect 14424 8236 14430 8288
rect 552 8186 17664 8208
rect 552 8134 4366 8186
rect 4418 8134 4430 8186
rect 4482 8134 4494 8186
rect 4546 8134 4558 8186
rect 4610 8134 4622 8186
rect 4674 8134 4686 8186
rect 4738 8134 10366 8186
rect 10418 8134 10430 8186
rect 10482 8134 10494 8186
rect 10546 8134 10558 8186
rect 10610 8134 10622 8186
rect 10674 8134 10686 8186
rect 10738 8134 16366 8186
rect 16418 8134 16430 8186
rect 16482 8134 16494 8186
rect 16546 8134 16558 8186
rect 16610 8134 16622 8186
rect 16674 8134 16686 8186
rect 16738 8134 17664 8186
rect 552 8112 17664 8134
rect 2222 8032 2228 8084
rect 2280 8032 2286 8084
rect 2682 8032 2688 8084
rect 2740 8032 2746 8084
rect 3234 8032 3240 8084
rect 3292 8032 3298 8084
rect 4246 8032 4252 8084
rect 4304 8032 4310 8084
rect 6115 8075 6173 8081
rect 6115 8041 6127 8075
rect 6161 8072 6173 8075
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6161 8044 6745 8072
rect 6161 8041 6173 8044
rect 6115 8035 6173 8041
rect 6733 8041 6745 8044
rect 6779 8072 6791 8075
rect 7006 8072 7012 8084
rect 6779 8044 7012 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 10192 8044 12296 8072
rect 10192 8032 10198 8044
rect 2240 8004 2268 8032
rect 2148 7976 2268 8004
rect 2700 8004 2728 8032
rect 2700 7976 3096 8004
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7936 1639 7939
rect 1946 7936 1952 7948
rect 1627 7908 1952 7936
rect 1627 7905 1639 7908
rect 1581 7899 1639 7905
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 2148 7945 2176 7976
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7905 2191 7939
rect 2133 7899 2191 7905
rect 2222 7896 2228 7948
rect 2280 7896 2286 7948
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 2590 7936 2596 7948
rect 2372 7908 2596 7936
rect 2372 7896 2378 7908
rect 2590 7896 2596 7908
rect 2648 7936 2654 7948
rect 3068 7945 3096 7976
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 2648 7908 2789 7936
rect 2648 7896 2654 7908
rect 2777 7905 2789 7908
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 2961 7939 3019 7945
rect 2961 7905 2973 7939
rect 3007 7905 3019 7939
rect 2961 7899 3019 7905
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 1854 7828 1860 7880
rect 1912 7828 1918 7880
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7837 2099 7871
rect 2240 7868 2268 7896
rect 2976 7868 3004 7899
rect 3142 7896 3148 7948
rect 3200 7936 3206 7948
rect 4062 7936 4068 7948
rect 3200 7908 4068 7936
rect 3200 7896 3206 7908
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4264 7936 4292 8032
rect 4617 8007 4675 8013
rect 4617 7973 4629 8007
rect 4663 8004 4675 8007
rect 5166 8004 5172 8016
rect 4663 7976 5172 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 5902 7964 5908 8016
rect 5960 7964 5966 8016
rect 6365 8007 6423 8013
rect 6365 8004 6377 8007
rect 6104 7976 6377 8004
rect 4338 7936 4344 7948
rect 4264 7908 4344 7936
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4948 7908 5089 7936
rect 4948 7896 4954 7908
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 5077 7899 5135 7905
rect 5258 7896 5264 7948
rect 5316 7936 5322 7948
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 5316 7908 5365 7936
rect 5316 7896 5322 7908
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 5534 7896 5540 7948
rect 5592 7896 5598 7948
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 2240 7840 3004 7868
rect 4540 7840 4997 7868
rect 2041 7831 2099 7837
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7800 1731 7803
rect 1946 7800 1952 7812
rect 1719 7772 1952 7800
rect 1719 7769 1731 7772
rect 1673 7763 1731 7769
rect 1946 7760 1952 7772
rect 2004 7800 2010 7812
rect 2056 7800 2084 7831
rect 2004 7772 2084 7800
rect 2501 7803 2559 7809
rect 2004 7760 2010 7772
rect 2501 7769 2513 7803
rect 2547 7800 2559 7803
rect 3510 7800 3516 7812
rect 2547 7772 3516 7800
rect 2547 7769 2559 7772
rect 2501 7763 2559 7769
rect 3510 7760 3516 7772
rect 3568 7760 3574 7812
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 4540 7809 4568 7840
rect 4985 7837 4997 7840
rect 5031 7868 5043 7871
rect 5552 7868 5580 7896
rect 6104 7880 6132 7976
rect 6365 7973 6377 7976
rect 6411 7973 6423 8007
rect 6365 7967 6423 7973
rect 6581 8007 6639 8013
rect 6581 7973 6593 8007
rect 6627 8004 6639 8007
rect 8110 8004 8116 8016
rect 6627 7976 8116 8004
rect 6627 7973 6639 7976
rect 6581 7967 6639 7973
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 9214 8004 9220 8016
rect 8352 7976 9220 8004
rect 8352 7964 8358 7976
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 12268 8004 12296 8044
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 13872 8044 14688 8072
rect 13872 8032 13878 8044
rect 10796 7976 12204 8004
rect 8018 7896 8024 7948
rect 8076 7936 8082 7948
rect 10796 7945 10824 7976
rect 12176 7948 12204 7976
rect 12268 7976 14504 8004
rect 10321 7939 10379 7945
rect 8076 7908 8156 7936
rect 8076 7896 8082 7908
rect 5031 7840 5580 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 6086 7828 6092 7880
rect 6144 7828 6150 7880
rect 8128 7877 8156 7908
rect 10321 7905 10333 7939
rect 10367 7905 10379 7939
rect 10321 7899 10379 7905
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 10551 7908 10793 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7936 11207 7939
rect 11238 7936 11244 7948
rect 11195 7908 11244 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 10336 7868 10364 7899
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 11425 7939 11483 7945
rect 11425 7905 11437 7939
rect 11471 7936 11483 7939
rect 11701 7939 11759 7945
rect 11701 7936 11713 7939
rect 11471 7908 11713 7936
rect 11471 7905 11483 7908
rect 11425 7899 11483 7905
rect 11701 7905 11713 7908
rect 11747 7905 11759 7939
rect 11701 7899 11759 7905
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 8435 7840 8524 7868
rect 10336 7840 10824 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 4525 7803 4583 7809
rect 4525 7800 4537 7803
rect 4028 7772 4537 7800
rect 4028 7760 4034 7772
rect 4525 7769 4537 7772
rect 4571 7769 4583 7803
rect 5537 7803 5595 7809
rect 5537 7800 5549 7803
rect 4525 7763 4583 7769
rect 5092 7772 5549 7800
rect 1762 7692 1768 7744
rect 1820 7692 1826 7744
rect 2590 7692 2596 7744
rect 2648 7692 2654 7744
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7732 4307 7735
rect 4982 7732 4988 7744
rect 4295 7704 4988 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 5092 7741 5120 7772
rect 5537 7769 5549 7772
rect 5583 7800 5595 7803
rect 6104 7800 6132 7828
rect 5583 7772 6132 7800
rect 6273 7803 6331 7809
rect 5583 7769 5595 7772
rect 5537 7763 5595 7769
rect 6273 7769 6285 7803
rect 6319 7800 6331 7803
rect 7098 7800 7104 7812
rect 6319 7772 7104 7800
rect 6319 7769 6331 7772
rect 6273 7763 6331 7769
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 8496 7744 8524 7840
rect 10796 7812 10824 7840
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 11900 7868 11928 7899
rect 12158 7896 12164 7948
rect 12216 7896 12222 7948
rect 12268 7945 12296 7976
rect 13648 7948 13676 7976
rect 12253 7939 12311 7945
rect 12253 7905 12265 7939
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7905 12495 7939
rect 12437 7899 12495 7905
rect 11572 7840 11928 7868
rect 12069 7871 12127 7877
rect 11572 7828 11578 7840
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 12452 7868 12480 7899
rect 12526 7896 12532 7948
rect 12584 7896 12590 7948
rect 13170 7896 13176 7948
rect 13228 7896 13234 7948
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 13538 7936 13544 7948
rect 13495 7908 13544 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 13630 7896 13636 7948
rect 13688 7945 13694 7948
rect 13688 7899 13695 7945
rect 13688 7896 13694 7899
rect 13814 7896 13820 7948
rect 13872 7896 13878 7948
rect 14001 7939 14059 7945
rect 14001 7905 14013 7939
rect 14047 7936 14059 7939
rect 14182 7936 14188 7948
rect 14047 7908 14188 7936
rect 14047 7905 14059 7908
rect 14001 7899 14059 7905
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 14476 7945 14504 7976
rect 14277 7939 14335 7945
rect 14277 7905 14289 7939
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14461 7939 14519 7945
rect 14461 7905 14473 7939
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 13188 7868 13216 7896
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 12452 7840 12756 7868
rect 13188 7840 13737 7868
rect 12069 7831 12127 7837
rect 10597 7803 10655 7809
rect 10597 7800 10609 7803
rect 10060 7772 10609 7800
rect 10060 7744 10088 7772
rect 10597 7769 10609 7772
rect 10643 7769 10655 7803
rect 10597 7763 10655 7769
rect 10778 7760 10784 7812
rect 10836 7760 10842 7812
rect 11698 7800 11704 7812
rect 11256 7772 11704 7800
rect 5077 7735 5135 7741
rect 5077 7701 5089 7735
rect 5123 7701 5135 7735
rect 5077 7695 5135 7701
rect 5258 7692 5264 7744
rect 5316 7692 5322 7744
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 6089 7735 6147 7741
rect 6089 7732 6101 7735
rect 5500 7704 6101 7732
rect 5500 7692 5506 7704
rect 6089 7701 6101 7704
rect 6135 7701 6147 7735
rect 6089 7695 6147 7701
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 8478 7732 8484 7744
rect 6604 7704 8484 7732
rect 6604 7692 6610 7704
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 10042 7692 10048 7744
rect 10100 7692 10106 7744
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 10686 7692 10692 7744
rect 10744 7732 10750 7744
rect 11256 7741 11284 7772
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 11241 7735 11299 7741
rect 11241 7732 11253 7735
rect 10744 7704 11253 7732
rect 10744 7692 10750 7704
rect 11241 7701 11253 7704
rect 11287 7701 11299 7735
rect 11241 7695 11299 7701
rect 11606 7692 11612 7744
rect 11664 7692 11670 7744
rect 12084 7732 12112 7831
rect 12728 7809 12756 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 12713 7803 12771 7809
rect 12713 7769 12725 7803
rect 12759 7800 12771 7803
rect 13538 7800 13544 7812
rect 12759 7772 13544 7800
rect 12759 7769 12771 7772
rect 12713 7763 12771 7769
rect 13538 7760 13544 7772
rect 13596 7800 13602 7812
rect 14292 7800 14320 7899
rect 14550 7896 14556 7948
rect 14608 7896 14614 7948
rect 14660 7945 14688 8044
rect 15194 8032 15200 8084
rect 15252 8032 15258 8084
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 16317 8075 16375 8081
rect 16317 8072 16329 8075
rect 15335 8044 16329 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 16317 8041 16329 8044
rect 16363 8041 16375 8075
rect 16317 8035 16375 8041
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 16758 8072 16764 8084
rect 16623 8044 16764 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 15212 8004 15240 8032
rect 15473 8007 15531 8013
rect 15473 8004 15485 8007
rect 15212 7976 15485 8004
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 14734 7896 14740 7948
rect 14792 7936 14798 7948
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 14792 7908 14841 7936
rect 14792 7896 14798 7908
rect 14829 7905 14841 7908
rect 14875 7936 14887 7939
rect 14918 7936 14924 7948
rect 14875 7908 14924 7936
rect 14875 7905 14887 7908
rect 14829 7899 14887 7905
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 15194 7896 15200 7948
rect 15252 7896 15258 7948
rect 15396 7945 15424 7976
rect 15473 7973 15485 7976
rect 15519 7973 15531 8007
rect 15473 7967 15531 7973
rect 15746 7964 15752 8016
rect 15804 8004 15810 8016
rect 16117 8007 16175 8013
rect 16117 8004 16129 8007
rect 15804 7976 16129 8004
rect 15804 7964 15810 7976
rect 16117 7973 16129 7976
rect 16163 7973 16175 8007
rect 16117 7967 16175 7973
rect 15381 7939 15439 7945
rect 15381 7905 15393 7939
rect 15427 7905 15439 7939
rect 15381 7899 15439 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7905 15715 7939
rect 16761 7939 16819 7945
rect 16761 7936 16773 7939
rect 15657 7899 15715 7905
rect 16500 7908 16773 7936
rect 13596 7772 14320 7800
rect 13596 7760 13602 7772
rect 14642 7760 14648 7812
rect 14700 7800 14706 7812
rect 15672 7800 15700 7899
rect 16500 7809 16528 7908
rect 16761 7905 16773 7908
rect 16807 7905 16819 7939
rect 16761 7899 16819 7905
rect 14700 7772 15700 7800
rect 16485 7803 16543 7809
rect 14700 7760 14706 7772
rect 16485 7769 16497 7803
rect 16531 7769 16543 7803
rect 16485 7763 16543 7769
rect 12342 7732 12348 7744
rect 12084 7704 12348 7732
rect 12342 7692 12348 7704
rect 12400 7732 12406 7744
rect 13814 7732 13820 7744
rect 12400 7704 13820 7732
rect 12400 7692 12406 7704
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14185 7735 14243 7741
rect 14185 7701 14197 7735
rect 14231 7732 14243 7735
rect 14918 7732 14924 7744
rect 14231 7704 14924 7732
rect 14231 7701 14243 7704
rect 14185 7695 14243 7701
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15010 7692 15016 7744
rect 15068 7692 15074 7744
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 15887 7704 16313 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 16301 7701 16313 7704
rect 16347 7701 16359 7735
rect 16301 7695 16359 7701
rect 552 7642 17664 7664
rect 552 7590 1366 7642
rect 1418 7590 1430 7642
rect 1482 7590 1494 7642
rect 1546 7590 1558 7642
rect 1610 7590 1622 7642
rect 1674 7590 1686 7642
rect 1738 7590 7366 7642
rect 7418 7590 7430 7642
rect 7482 7590 7494 7642
rect 7546 7590 7558 7642
rect 7610 7590 7622 7642
rect 7674 7590 7686 7642
rect 7738 7590 13366 7642
rect 13418 7590 13430 7642
rect 13482 7590 13494 7642
rect 13546 7590 13558 7642
rect 13610 7590 13622 7642
rect 13674 7590 13686 7642
rect 13738 7590 17664 7642
rect 552 7568 17664 7590
rect 1854 7488 1860 7540
rect 1912 7488 1918 7540
rect 1946 7488 1952 7540
rect 2004 7528 2010 7540
rect 2041 7531 2099 7537
rect 2041 7528 2053 7531
rect 2004 7500 2053 7528
rect 2004 7488 2010 7500
rect 2041 7497 2053 7500
rect 2087 7497 2099 7531
rect 2041 7491 2099 7497
rect 2590 7488 2596 7540
rect 2648 7488 2654 7540
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 4304 7500 4353 7528
rect 4304 7488 4310 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4341 7491 4399 7497
rect 4540 7500 4629 7528
rect 1872 7460 1900 7488
rect 2317 7463 2375 7469
rect 2317 7460 2329 7463
rect 1872 7432 2329 7460
rect 1872 7324 1900 7432
rect 2317 7429 2329 7432
rect 2363 7429 2375 7463
rect 2317 7423 2375 7429
rect 2608 7392 2636 7488
rect 4154 7420 4160 7472
rect 4212 7420 4218 7472
rect 2148 7364 2636 7392
rect 3697 7395 3755 7401
rect 2148 7333 2176 7364
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 3743 7364 4445 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 4433 7361 4445 7364
rect 4479 7392 4491 7395
rect 4540 7392 4568 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 4617 7491 4675 7497
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5169 7531 5227 7537
rect 5169 7528 5181 7531
rect 5040 7500 5181 7528
rect 5040 7488 5046 7500
rect 5169 7497 5181 7500
rect 5215 7528 5227 7531
rect 5442 7528 5448 7540
rect 5215 7500 5448 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 5537 7531 5595 7537
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 5810 7528 5816 7540
rect 5583 7500 5816 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6089 7531 6147 7537
rect 6089 7528 6101 7531
rect 5960 7500 6101 7528
rect 5960 7488 5966 7500
rect 6089 7497 6101 7500
rect 6135 7497 6147 7531
rect 6089 7491 6147 7497
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 9490 7528 9496 7540
rect 6512 7500 9496 7528
rect 6512 7488 6518 7500
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 9732 7500 10088 7528
rect 9732 7488 9738 7500
rect 5258 7420 5264 7472
rect 5316 7460 5322 7472
rect 7926 7460 7932 7472
rect 5316 7432 7932 7460
rect 5316 7420 5322 7432
rect 7926 7420 7932 7432
rect 7984 7420 7990 7472
rect 9766 7460 9772 7472
rect 8680 7432 9772 7460
rect 4479 7364 4568 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5224 7364 5948 7392
rect 5224 7352 5230 7364
rect 1949 7327 2007 7333
rect 1949 7324 1961 7327
rect 1872 7296 1961 7324
rect 1949 7293 1961 7296
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7293 2191 7327
rect 2133 7287 2191 7293
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2314 7324 2320 7336
rect 2271 7296 2320 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7293 2467 7327
rect 2409 7287 2467 7293
rect 1762 7148 1768 7200
rect 1820 7188 1826 7200
rect 2038 7188 2044 7200
rect 1820 7160 2044 7188
rect 1820 7148 1826 7160
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 2222 7148 2228 7200
rect 2280 7188 2286 7200
rect 2424 7188 2452 7287
rect 2498 7284 2504 7336
rect 2556 7284 2562 7336
rect 2682 7284 2688 7336
rect 2740 7284 2746 7336
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 3789 7327 3847 7333
rect 3789 7324 3801 7327
rect 2915 7296 3801 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 3789 7293 3801 7296
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 3234 7216 3240 7268
rect 3292 7216 3298 7268
rect 3804 7256 3832 7287
rect 3970 7284 3976 7336
rect 4028 7284 4034 7336
rect 4525 7327 4583 7333
rect 4525 7324 4537 7327
rect 4080 7296 4537 7324
rect 3878 7256 3884 7268
rect 3804 7228 3884 7256
rect 3878 7216 3884 7228
rect 3936 7256 3942 7268
rect 4080 7256 4108 7296
rect 4525 7293 4537 7296
rect 4571 7293 4583 7327
rect 4525 7287 4583 7293
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 3936 7228 4108 7256
rect 4249 7259 4307 7265
rect 3936 7216 3942 7228
rect 4249 7225 4261 7259
rect 4295 7256 4307 7259
rect 4338 7256 4344 7268
rect 4295 7228 4344 7256
rect 4295 7225 4307 7228
rect 4249 7219 4307 7225
rect 4338 7216 4344 7228
rect 4396 7216 4402 7268
rect 2280 7160 2452 7188
rect 3252 7188 3280 7216
rect 4632 7188 4660 7287
rect 4816 7256 4844 7287
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4948 7296 4997 7324
rect 4948 7284 4954 7296
rect 4985 7293 4997 7296
rect 5031 7324 5043 7327
rect 5353 7327 5411 7333
rect 5353 7324 5365 7327
rect 5031 7296 5365 7324
rect 5031 7293 5043 7296
rect 4985 7287 5043 7293
rect 5353 7293 5365 7296
rect 5399 7293 5411 7327
rect 5353 7287 5411 7293
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5920 7333 5948 7364
rect 5994 7352 6000 7404
rect 6052 7352 6058 7404
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5592 7296 5641 7324
rect 5592 7284 5598 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7293 5963 7327
rect 6012 7324 6040 7352
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 6012 7296 6377 7324
rect 5905 7287 5963 7293
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 6564 7256 6592 7352
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8168 7296 8585 7324
rect 8168 7284 8174 7296
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8680 7324 8708 7432
rect 9766 7420 9772 7432
rect 9824 7420 9830 7472
rect 10060 7460 10088 7500
rect 10134 7488 10140 7540
rect 10192 7488 10198 7540
rect 10410 7488 10416 7540
rect 10468 7488 10474 7540
rect 10686 7488 10692 7540
rect 10744 7488 10750 7540
rect 11606 7488 11612 7540
rect 11664 7488 11670 7540
rect 11698 7488 11704 7540
rect 11756 7488 11762 7540
rect 12069 7531 12127 7537
rect 12069 7497 12081 7531
rect 12115 7528 12127 7531
rect 12158 7528 12164 7540
rect 12115 7500 12164 7528
rect 12115 7497 12127 7500
rect 12069 7491 12127 7497
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12342 7488 12348 7540
rect 12400 7488 12406 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 12894 7528 12900 7540
rect 12492 7500 12900 7528
rect 12492 7488 12498 7500
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 14734 7528 14740 7540
rect 13872 7500 14740 7528
rect 13872 7488 13878 7500
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 10318 7460 10324 7472
rect 10060 7432 10324 7460
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 10428 7460 10456 7488
rect 10428 7432 11376 7460
rect 9048 7364 9674 7392
rect 9048 7340 9076 7364
rect 8956 7333 9076 7340
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 8680 7296 8769 7324
rect 8573 7287 8631 7293
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 8849 7327 8907 7333
rect 8849 7293 8861 7327
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 8941 7327 9076 7333
rect 8941 7293 8953 7327
rect 8987 7312 9076 7327
rect 8987 7293 8999 7312
rect 8941 7287 8999 7293
rect 4816 7228 4936 7256
rect 4908 7200 4936 7228
rect 5828 7228 6592 7256
rect 6840 7256 6868 7284
rect 8772 7256 8800 7287
rect 6840 7228 8800 7256
rect 3252 7160 4660 7188
rect 2280 7148 2286 7160
rect 4890 7148 4896 7200
rect 4948 7148 4954 7200
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 5828 7197 5856 7228
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 5224 7160 5825 7188
rect 5224 7148 5230 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5813 7151 5871 7157
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6420 7160 6561 7188
rect 6420 7148 6426 7160
rect 6549 7157 6561 7160
rect 6595 7188 6607 7191
rect 7098 7188 7104 7200
rect 6595 7160 7104 7188
rect 6595 7157 6607 7160
rect 6549 7151 6607 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 8389 7191 8447 7197
rect 8389 7157 8401 7191
rect 8435 7188 8447 7191
rect 8570 7188 8576 7200
rect 8435 7160 8576 7188
rect 8435 7157 8447 7160
rect 8389 7151 8447 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 8864 7188 8892 7287
rect 8956 7256 8984 7287
rect 9122 7284 9128 7336
rect 9180 7284 9186 7336
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9324 7256 9352 7287
rect 9490 7284 9496 7336
rect 9548 7284 9554 7336
rect 9646 7324 9674 7364
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11348 7401 11376 7432
rect 11241 7395 11299 7401
rect 11241 7392 11253 7395
rect 11112 7364 11253 7392
rect 11112 7352 11118 7364
rect 11241 7361 11253 7364
rect 11287 7361 11299 7395
rect 11241 7355 11299 7361
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7361 11391 7395
rect 11333 7355 11391 7361
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7392 11575 7395
rect 11624 7392 11652 7488
rect 11716 7460 11744 7488
rect 14001 7463 14059 7469
rect 14001 7460 14013 7463
rect 11716 7432 14013 7460
rect 14001 7429 14013 7432
rect 14047 7460 14059 7463
rect 14553 7463 14611 7469
rect 14553 7460 14565 7463
rect 14047 7432 14565 7460
rect 14047 7429 14059 7432
rect 14001 7423 14059 7429
rect 14553 7429 14565 7432
rect 14599 7460 14611 7463
rect 15381 7463 15439 7469
rect 15381 7460 15393 7463
rect 14599 7432 15393 7460
rect 14599 7429 14611 7432
rect 14553 7423 14611 7429
rect 15381 7429 15393 7432
rect 15427 7429 15439 7463
rect 15381 7423 15439 7429
rect 15562 7420 15568 7472
rect 15620 7460 15626 7472
rect 15746 7460 15752 7472
rect 15620 7432 15752 7460
rect 15620 7420 15626 7432
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 11563 7364 11652 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 12032 7364 13921 7392
rect 12032 7352 12038 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14366 7352 14372 7404
rect 14424 7392 14430 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 14424 7364 14473 7392
rect 14424 7352 14430 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 14918 7352 14924 7404
rect 14976 7352 14982 7404
rect 15010 7352 15016 7404
rect 15068 7352 15074 7404
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9646 7296 9965 7324
rect 9953 7293 9965 7296
rect 9999 7324 10011 7327
rect 10229 7327 10287 7333
rect 10229 7324 10241 7327
rect 9999 7296 10241 7324
rect 9999 7293 10011 7296
rect 9953 7287 10011 7293
rect 10229 7293 10241 7296
rect 10275 7293 10287 7327
rect 10229 7287 10287 7293
rect 10413 7327 10471 7333
rect 10413 7293 10425 7327
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10428 7256 10456 7287
rect 10502 7284 10508 7336
rect 10560 7284 10566 7336
rect 11425 7327 11483 7333
rect 10980 7272 11192 7300
rect 11425 7293 11437 7327
rect 11471 7324 11483 7327
rect 11606 7324 11612 7336
rect 11471 7296 11612 7324
rect 11471 7293 11483 7296
rect 11425 7287 11483 7293
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7293 12311 7327
rect 12253 7287 12311 7293
rect 10980 7256 11008 7272
rect 8956 7228 9168 7256
rect 9324 7228 10180 7256
rect 10428 7228 11008 7256
rect 11164 7256 11192 7272
rect 12268 7256 12296 7287
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 12400 7296 12541 7324
rect 12400 7284 12406 7296
rect 12529 7293 12541 7296
rect 12575 7324 12587 7327
rect 12894 7324 12900 7336
rect 12575 7296 12900 7324
rect 12575 7293 12587 7296
rect 12529 7287 12587 7293
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 14185 7327 14243 7333
rect 14185 7293 14197 7327
rect 14231 7324 14243 7327
rect 14274 7324 14280 7336
rect 14231 7296 14280 7324
rect 14231 7293 14243 7296
rect 14185 7287 14243 7293
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7324 14795 7327
rect 14936 7324 14964 7352
rect 14783 7296 14964 7324
rect 15028 7324 15056 7352
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 15028 7296 15209 7324
rect 14783 7293 14795 7296
rect 14737 7287 14795 7293
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 15378 7284 15384 7336
rect 15436 7324 15442 7336
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 15436 7296 15485 7324
rect 15436 7284 15442 7296
rect 15473 7293 15485 7296
rect 15519 7324 15531 7327
rect 15562 7324 15568 7336
rect 15519 7296 15568 7324
rect 15519 7293 15531 7296
rect 15473 7287 15531 7293
rect 15562 7284 15568 7296
rect 15620 7284 15626 7336
rect 15654 7284 15660 7336
rect 15712 7324 15718 7336
rect 16206 7324 16212 7336
rect 15712 7296 16212 7324
rect 15712 7284 15718 7296
rect 16206 7284 16212 7296
rect 16264 7324 16270 7336
rect 16669 7327 16727 7333
rect 16669 7324 16681 7327
rect 16264 7296 16681 7324
rect 16264 7284 16270 7296
rect 16669 7293 16681 7296
rect 16715 7293 16727 7327
rect 16669 7287 16727 7293
rect 16853 7327 16911 7333
rect 16853 7293 16865 7327
rect 16899 7324 16911 7327
rect 17218 7324 17224 7336
rect 16899 7296 17224 7324
rect 16899 7293 16911 7296
rect 16853 7287 16911 7293
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 16761 7259 16819 7265
rect 16761 7256 16773 7259
rect 11164 7228 16773 7256
rect 9140 7200 9168 7228
rect 10152 7200 10180 7228
rect 16761 7225 16773 7228
rect 16807 7225 16819 7259
rect 16761 7219 16819 7225
rect 9030 7188 9036 7200
rect 8864 7160 9036 7188
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9122 7148 9128 7200
rect 9180 7148 9186 7200
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 9364 7160 9689 7188
rect 9364 7148 9370 7160
rect 9677 7157 9689 7160
rect 9723 7157 9735 7191
rect 9677 7151 9735 7157
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10321 7191 10379 7197
rect 10321 7188 10333 7191
rect 10192 7160 10333 7188
rect 10192 7148 10198 7160
rect 10321 7157 10333 7160
rect 10367 7157 10379 7191
rect 10321 7151 10379 7157
rect 11054 7148 11060 7200
rect 11112 7148 11118 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 14369 7191 14427 7197
rect 14369 7188 14381 7191
rect 13228 7160 14381 7188
rect 13228 7148 13234 7160
rect 14369 7157 14381 7160
rect 14415 7157 14427 7191
rect 14369 7151 14427 7157
rect 14918 7148 14924 7200
rect 14976 7148 14982 7200
rect 15010 7148 15016 7200
rect 15068 7148 15074 7200
rect 552 7098 17664 7120
rect 552 7046 4366 7098
rect 4418 7046 4430 7098
rect 4482 7046 4494 7098
rect 4546 7046 4558 7098
rect 4610 7046 4622 7098
rect 4674 7046 4686 7098
rect 4738 7046 10366 7098
rect 10418 7046 10430 7098
rect 10482 7046 10494 7098
rect 10546 7046 10558 7098
rect 10610 7046 10622 7098
rect 10674 7046 10686 7098
rect 10738 7046 16366 7098
rect 16418 7046 16430 7098
rect 16482 7046 16494 7098
rect 16546 7046 16558 7098
rect 16610 7046 16622 7098
rect 16674 7046 16686 7098
rect 16738 7046 17664 7098
rect 552 7024 17664 7046
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 4338 6984 4344 6996
rect 3936 6956 4344 6984
rect 3936 6944 3942 6956
rect 4338 6944 4344 6956
rect 4396 6944 4402 6996
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 9030 6984 9036 6996
rect 6052 6956 9036 6984
rect 6052 6944 6058 6956
rect 3510 6876 3516 6928
rect 3568 6916 3574 6928
rect 3568 6888 4108 6916
rect 3568 6876 3574 6888
rect 1112 6851 1170 6857
rect 1112 6817 1124 6851
rect 1158 6848 1170 6851
rect 1854 6848 1860 6860
rect 1158 6820 1860 6848
rect 1158 6817 1170 6820
rect 1112 6811 1170 6817
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 2498 6848 2504 6860
rect 2240 6820 2504 6848
rect 842 6740 848 6792
rect 900 6740 906 6792
rect 2240 6721 2268 6820
rect 2498 6808 2504 6820
rect 2556 6848 2562 6860
rect 3620 6857 3648 6888
rect 2685 6851 2743 6857
rect 2685 6848 2697 6851
rect 2556 6820 2697 6848
rect 2556 6808 2562 6820
rect 2685 6817 2697 6820
rect 2731 6817 2743 6851
rect 2685 6811 2743 6817
rect 3605 6851 3663 6857
rect 3605 6817 3617 6851
rect 3651 6817 3663 6851
rect 3605 6811 3663 6817
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 3878 6848 3884 6860
rect 3835 6820 3884 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 3973 6851 4031 6857
rect 3973 6817 3985 6851
rect 4019 6817 4031 6851
rect 4080 6848 4108 6888
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4212 6888 4752 6916
rect 4212 6876 4218 6888
rect 4249 6851 4307 6857
rect 4249 6848 4261 6851
rect 4080 6820 4261 6848
rect 3973 6811 4031 6817
rect 4249 6817 4261 6820
rect 4295 6817 4307 6851
rect 4249 6811 4307 6817
rect 3988 6780 4016 6811
rect 4338 6808 4344 6860
rect 4396 6808 4402 6860
rect 4724 6857 4752 6888
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 7006 6916 7012 6928
rect 5316 6888 7012 6916
rect 5316 6876 5322 6888
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 8110 6916 8116 6928
rect 7248 6888 8116 6916
rect 7248 6876 7254 6888
rect 8110 6876 8116 6888
rect 8168 6916 8174 6928
rect 8168 6888 8248 6916
rect 8168 6876 8174 6888
rect 4709 6851 4767 6857
rect 4709 6817 4721 6851
rect 4755 6817 4767 6851
rect 4709 6811 4767 6817
rect 4893 6851 4951 6857
rect 4893 6817 4905 6851
rect 4939 6817 4951 6851
rect 4893 6811 4951 6817
rect 4908 6780 4936 6811
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 7837 6851 7895 6857
rect 7340 6820 7788 6848
rect 7340 6808 7346 6820
rect 7760 6792 7788 6820
rect 7837 6817 7849 6851
rect 7883 6817 7895 6851
rect 7837 6811 7895 6817
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6817 8079 6851
rect 8220 6848 8248 6888
rect 8404 6857 8432 6956
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 10962 6944 10968 6996
rect 11020 6984 11026 6996
rect 15194 6984 15200 6996
rect 11020 6956 15200 6984
rect 11020 6944 11026 6956
rect 15194 6944 15200 6956
rect 15252 6984 15258 6996
rect 15378 6984 15384 6996
rect 15252 6956 15384 6984
rect 15252 6944 15258 6956
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 8570 6876 8576 6928
rect 8628 6916 8634 6928
rect 9490 6916 9496 6928
rect 8628 6888 9496 6916
rect 8628 6876 8634 6888
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 11882 6916 11888 6928
rect 10060 6888 10640 6916
rect 10060 6860 10088 6888
rect 8021 6811 8079 6817
rect 8128 6820 8248 6848
rect 8389 6851 8447 6857
rect 3988 6752 4292 6780
rect 2225 6715 2283 6721
rect 2225 6681 2237 6715
rect 2271 6681 2283 6715
rect 2225 6675 2283 6681
rect 3973 6715 4031 6721
rect 3973 6681 3985 6715
rect 4019 6712 4031 6715
rect 4062 6712 4068 6724
rect 4019 6684 4068 6712
rect 4019 6681 4031 6684
rect 3973 6675 4031 6681
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 4264 6712 4292 6752
rect 4540 6752 4936 6780
rect 4540 6712 4568 6752
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 7098 6740 7104 6792
rect 7156 6740 7162 6792
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6780 7251 6783
rect 7466 6780 7472 6792
rect 7239 6752 7472 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7742 6740 7748 6792
rect 7800 6740 7806 6792
rect 7852 6780 7880 6811
rect 7926 6780 7932 6792
rect 7852 6752 7932 6780
rect 4264 6684 4568 6712
rect 4617 6715 4675 6721
rect 4264 6656 4292 6684
rect 4617 6681 4629 6715
rect 4663 6712 4675 6715
rect 4798 6712 4804 6724
rect 4663 6684 4804 6712
rect 4663 6681 4675 6684
rect 4617 6675 4675 6681
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 7852 6712 7880 6752
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 6564 6684 7880 6712
rect 6564 6656 6592 6684
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3602 6644 3608 6656
rect 2915 6616 3608 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 4246 6604 4252 6656
rect 4304 6604 4310 6656
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4396 6616 4721 6644
rect 4396 6604 4402 6616
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 6546 6604 6552 6656
rect 6604 6604 6610 6656
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 7926 6644 7932 6656
rect 7515 6616 7932 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8036 6644 8064 6811
rect 8128 6789 8156 6820
rect 8389 6817 8401 6851
rect 8435 6817 8447 6851
rect 8389 6811 8447 6817
rect 9122 6808 9128 6860
rect 9180 6848 9186 6860
rect 9769 6851 9827 6857
rect 9769 6848 9781 6851
rect 9180 6820 9781 6848
rect 9180 6808 9186 6820
rect 9769 6817 9781 6820
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 10042 6808 10048 6860
rect 10100 6808 10106 6860
rect 10134 6808 10140 6860
rect 10192 6808 10198 6860
rect 10612 6857 10640 6888
rect 11164 6888 11888 6916
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 11164 6857 11192 6888
rect 11882 6876 11888 6888
rect 11940 6876 11946 6928
rect 13262 6876 13268 6928
rect 13320 6876 13326 6928
rect 14090 6876 14096 6928
rect 14148 6916 14154 6928
rect 14366 6916 14372 6928
rect 14148 6888 14372 6916
rect 14148 6876 14154 6888
rect 14366 6876 14372 6888
rect 14424 6876 14430 6928
rect 14642 6876 14648 6928
rect 14700 6876 14706 6928
rect 16206 6876 16212 6928
rect 16264 6916 16270 6928
rect 16482 6916 16488 6928
rect 16264 6888 16488 6916
rect 16264 6876 16270 6888
rect 16482 6876 16488 6888
rect 16540 6916 16546 6928
rect 16577 6919 16635 6925
rect 16577 6916 16589 6919
rect 16540 6888 16589 6916
rect 16540 6876 16546 6888
rect 16577 6885 16589 6888
rect 16623 6885 16635 6919
rect 16577 6879 16635 6885
rect 11330 6857 11336 6860
rect 11149 6851 11207 6857
rect 11149 6817 11161 6851
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 11287 6851 11336 6857
rect 11287 6817 11299 6851
rect 11333 6817 11336 6851
rect 11287 6811 11336 6817
rect 11330 6808 11336 6811
rect 11388 6808 11394 6860
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 11701 6851 11759 6857
rect 11701 6817 11713 6851
rect 11747 6817 11759 6851
rect 13280 6848 13308 6876
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13280 6820 13829 6848
rect 11701 6811 11759 6817
rect 13817 6817 13829 6820
rect 13863 6817 13875 6851
rect 13817 6811 13875 6817
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8220 6712 8248 6743
rect 8570 6740 8576 6792
rect 8628 6740 8634 6792
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9272 6752 9413 6780
rect 9272 6740 9278 6752
rect 9401 6749 9413 6752
rect 9447 6780 9459 6783
rect 9490 6780 9496 6792
rect 9447 6752 9496 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 10152 6780 10180 6808
rect 9723 6752 10180 6780
rect 10229 6783 10287 6789
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 10229 6749 10241 6783
rect 10275 6780 10287 6783
rect 10318 6780 10324 6792
rect 10275 6752 10324 6780
rect 10275 6749 10287 6752
rect 10229 6743 10287 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 11054 6780 11060 6792
rect 10735 6752 11060 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11422 6740 11428 6792
rect 11480 6740 11486 6792
rect 9766 6712 9772 6724
rect 8220 6684 9772 6712
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 8478 6644 8484 6656
rect 8036 6616 8484 6644
rect 8478 6604 8484 6616
rect 8536 6644 8542 6656
rect 9953 6647 10011 6653
rect 9953 6644 9965 6647
rect 8536 6616 9965 6644
rect 8536 6604 8542 6616
rect 9953 6613 9965 6616
rect 9999 6644 10011 6647
rect 11532 6644 11560 6811
rect 11716 6724 11744 6811
rect 14660 6780 14688 6876
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16114 6848 16120 6860
rect 15988 6820 16120 6848
rect 15988 6808 15994 6820
rect 16114 6808 16120 6820
rect 16172 6848 16178 6860
rect 16393 6851 16451 6857
rect 16393 6848 16405 6851
rect 16172 6820 16405 6848
rect 16172 6808 16178 6820
rect 16393 6817 16405 6820
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 14016 6752 14688 6780
rect 11698 6672 11704 6724
rect 11756 6672 11762 6724
rect 14016 6721 14044 6752
rect 14918 6740 14924 6792
rect 14976 6780 14982 6792
rect 16209 6783 16267 6789
rect 16209 6780 16221 6783
rect 14976 6752 16221 6780
rect 14976 6740 14982 6752
rect 16209 6749 16221 6752
rect 16255 6749 16267 6783
rect 16209 6743 16267 6749
rect 14001 6715 14059 6721
rect 14001 6681 14013 6715
rect 14047 6681 14059 6715
rect 14001 6675 14059 6681
rect 14366 6672 14372 6724
rect 14424 6712 14430 6724
rect 14826 6712 14832 6724
rect 14424 6684 14832 6712
rect 14424 6672 14430 6684
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 12158 6644 12164 6656
rect 9999 6616 12164 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 12526 6604 12532 6656
rect 12584 6644 12590 6656
rect 13078 6644 13084 6656
rect 12584 6616 13084 6644
rect 12584 6604 12590 6616
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 552 6554 17664 6576
rect 552 6502 1366 6554
rect 1418 6502 1430 6554
rect 1482 6502 1494 6554
rect 1546 6502 1558 6554
rect 1610 6502 1622 6554
rect 1674 6502 1686 6554
rect 1738 6502 7366 6554
rect 7418 6502 7430 6554
rect 7482 6502 7494 6554
rect 7546 6502 7558 6554
rect 7610 6502 7622 6554
rect 7674 6502 7686 6554
rect 7738 6502 13366 6554
rect 13418 6502 13430 6554
rect 13482 6502 13494 6554
rect 13546 6502 13558 6554
rect 13610 6502 13622 6554
rect 13674 6502 13686 6554
rect 13738 6502 17664 6554
rect 552 6480 17664 6502
rect 3694 6400 3700 6452
rect 3752 6440 3758 6452
rect 6454 6440 6460 6452
rect 3752 6412 6460 6440
rect 3752 6400 3758 6412
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 7064 6412 8401 6440
rect 7064 6400 7070 6412
rect 8389 6409 8401 6412
rect 8435 6409 8447 6443
rect 8389 6403 8447 6409
rect 8570 6400 8576 6452
rect 8628 6400 8634 6452
rect 8757 6443 8815 6449
rect 8757 6409 8769 6443
rect 8803 6409 8815 6443
rect 8757 6403 8815 6409
rect 5810 6332 5816 6384
rect 5868 6372 5874 6384
rect 5868 6344 6132 6372
rect 5868 6332 5874 6344
rect 6104 6313 6132 6344
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 6328 6344 7849 6372
rect 6328 6332 6334 6344
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 7837 6335 7895 6341
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6273 6147 6307
rect 6822 6304 6828 6316
rect 6089 6267 6147 6273
rect 6288 6276 6828 6304
rect 2590 6236 2596 6248
rect 2240 6208 2596 6236
rect 2240 6180 2268 6208
rect 2590 6196 2596 6208
rect 2648 6236 2654 6248
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 2648 6208 2789 6236
rect 2648 6196 2654 6208
rect 2777 6205 2789 6208
rect 2823 6205 2835 6239
rect 2777 6199 2835 6205
rect 5997 6239 6055 6245
rect 5997 6205 6009 6239
rect 6043 6236 6055 6239
rect 6288 6236 6316 6276
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7156 6276 7481 6304
rect 7156 6264 7162 6276
rect 7469 6273 7481 6276
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 7668 6276 8156 6304
rect 7190 6236 7196 6248
rect 6043 6208 6316 6236
rect 6380 6208 7196 6236
rect 6043 6205 6055 6208
rect 5997 6199 6055 6205
rect 2222 6128 2228 6180
rect 2280 6128 2286 6180
rect 6380 6168 6408 6208
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7374 6196 7380 6248
rect 7432 6196 7438 6248
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6236 7619 6239
rect 7668 6236 7696 6276
rect 8128 6248 8156 6276
rect 7607 6208 7696 6236
rect 7607 6205 7619 6208
rect 7561 6199 7619 6205
rect 2424 6140 6408 6168
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 2424 6100 2452 6140
rect 7006 6128 7012 6180
rect 7064 6128 7070 6180
rect 7668 6168 7696 6208
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 7116 6140 7696 6168
rect 2096 6072 2452 6100
rect 2096 6060 2102 6072
rect 2498 6060 2504 6112
rect 2556 6100 2562 6112
rect 2593 6103 2651 6109
rect 2593 6100 2605 6103
rect 2556 6072 2605 6100
rect 2556 6060 2562 6072
rect 2593 6069 2605 6072
rect 2639 6069 2651 6103
rect 2593 6063 2651 6069
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 6178 6100 6184 6112
rect 5776 6072 6184 6100
rect 5776 6060 5782 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6319 6103 6377 6109
rect 6319 6069 6331 6103
rect 6365 6100 6377 6103
rect 7116 6100 7144 6140
rect 6365 6072 7144 6100
rect 6365 6069 6377 6072
rect 6319 6063 6377 6069
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 7760 6100 7788 6199
rect 8036 6168 8064 6199
rect 8110 6196 8116 6248
rect 8168 6196 8174 6248
rect 8588 6245 8616 6400
rect 8772 6372 8800 6403
rect 9122 6400 9128 6452
rect 9180 6400 9186 6452
rect 9398 6400 9404 6452
rect 9456 6400 9462 6452
rect 9766 6400 9772 6452
rect 9824 6400 9830 6452
rect 11054 6400 11060 6452
rect 11112 6400 11118 6452
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 11425 6443 11483 6449
rect 11425 6440 11437 6443
rect 11296 6412 11437 6440
rect 11296 6400 11302 6412
rect 11425 6409 11437 6412
rect 11471 6409 11483 6443
rect 12250 6440 12256 6452
rect 11425 6403 11483 6409
rect 11560 6412 12256 6440
rect 8938 6372 8944 6384
rect 8772 6344 8944 6372
rect 8938 6332 8944 6344
rect 8996 6372 9002 6384
rect 9416 6372 9444 6400
rect 8996 6344 9444 6372
rect 9784 6372 9812 6400
rect 11330 6372 11336 6384
rect 9784 6344 11336 6372
rect 8996 6332 9002 6344
rect 11330 6332 11336 6344
rect 11388 6372 11394 6384
rect 11560 6372 11588 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 14461 6443 14519 6449
rect 13004 6412 13860 6440
rect 13004 6372 13032 6412
rect 11388 6344 11588 6372
rect 11624 6344 13032 6372
rect 13832 6372 13860 6412
rect 14461 6409 14473 6443
rect 14507 6440 14519 6443
rect 15562 6440 15568 6452
rect 14507 6412 15568 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 15838 6400 15844 6452
rect 15896 6440 15902 6452
rect 16206 6440 16212 6452
rect 15896 6412 16212 6440
rect 15896 6400 15902 6412
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 16393 6375 16451 6381
rect 16393 6372 16405 6375
rect 13832 6344 16405 6372
rect 11388 6332 11394 6344
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 11422 6304 11428 6316
rect 8895 6276 11428 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 8864 6236 8892 6267
rect 11422 6264 11428 6276
rect 11480 6304 11486 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11480 6276 11529 6304
rect 11480 6264 11486 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 8720 6208 8892 6236
rect 8941 6239 8999 6245
rect 8720 6196 8726 6208
rect 8941 6205 8953 6239
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 8956 6168 8984 6199
rect 9950 6196 9956 6248
rect 10008 6236 10014 6248
rect 10318 6236 10324 6248
rect 10008 6208 10324 6236
rect 10008 6196 10014 6208
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 10962 6196 10968 6248
rect 11020 6236 11026 6248
rect 11241 6239 11299 6245
rect 11241 6236 11253 6239
rect 11020 6208 11253 6236
rect 11020 6196 11026 6208
rect 11241 6205 11253 6208
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 11624 6168 11652 6344
rect 16393 6341 16405 6344
rect 16439 6341 16451 6375
rect 16393 6335 16451 6341
rect 12084 6276 13584 6304
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 11885 6239 11943 6245
rect 11885 6236 11897 6239
rect 11848 6208 11897 6236
rect 11848 6196 11854 6208
rect 11885 6205 11897 6208
rect 11931 6205 11943 6239
rect 11885 6199 11943 6205
rect 8036 6140 11652 6168
rect 7248 6072 7788 6100
rect 7248 6060 7254 6072
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 11698 6100 11704 6112
rect 8076 6072 11704 6100
rect 8076 6060 8082 6072
rect 11698 6060 11704 6072
rect 11756 6100 11762 6112
rect 12084 6109 12112 6276
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 12802 6236 12808 6248
rect 12308 6208 12808 6236
rect 12308 6196 12314 6208
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 13556 6245 13584 6276
rect 13814 6264 13820 6316
rect 13872 6264 13878 6316
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 14323 6276 14688 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 13725 6239 13783 6245
rect 13725 6205 13737 6239
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6236 13967 6239
rect 14093 6239 14151 6245
rect 13955 6208 14044 6236
rect 13955 6205 13967 6208
rect 13909 6199 13967 6205
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 13740 6168 13768 6199
rect 12216 6140 13768 6168
rect 12216 6128 12222 6140
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11756 6072 12081 6100
rect 11756 6060 11762 6072
rect 12069 6069 12081 6072
rect 12115 6069 12127 6103
rect 12069 6063 12127 6069
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 12621 6103 12679 6109
rect 12621 6100 12633 6103
rect 12308 6072 12633 6100
rect 12308 6060 12314 6072
rect 12621 6069 12633 6072
rect 12667 6100 12679 6103
rect 14016 6100 14044 6208
rect 14093 6205 14105 6239
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 14108 6168 14136 6199
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 14240 6208 14381 6236
rect 14240 6196 14246 6208
rect 14369 6205 14381 6208
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 14550 6196 14556 6248
rect 14608 6196 14614 6248
rect 14660 6245 14688 6276
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 15105 6307 15163 6313
rect 15105 6304 15117 6307
rect 14884 6276 15117 6304
rect 14884 6264 14890 6276
rect 15105 6273 15117 6276
rect 15151 6273 15163 6307
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 15105 6267 15163 6273
rect 15304 6276 16681 6304
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 14568 6168 14596 6196
rect 14108 6140 14596 6168
rect 15194 6128 15200 6180
rect 15252 6168 15258 6180
rect 15304 6168 15332 6276
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6205 15439 6239
rect 15381 6199 15439 6205
rect 15252 6140 15332 6168
rect 15396 6168 15424 6199
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15620 6208 16037 6236
rect 15620 6196 15626 6208
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16114 6196 16120 6248
rect 16172 6236 16178 6248
rect 16500 6245 16528 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 16209 6239 16267 6245
rect 16209 6236 16221 6239
rect 16172 6208 16221 6236
rect 16172 6196 16178 6208
rect 16209 6205 16221 6208
rect 16255 6236 16267 6239
rect 16301 6239 16359 6245
rect 16301 6236 16313 6239
rect 16255 6208 16313 6236
rect 16255 6205 16267 6208
rect 16209 6199 16267 6205
rect 16301 6205 16313 6208
rect 16347 6205 16359 6239
rect 16301 6199 16359 6205
rect 16485 6239 16543 6245
rect 16485 6205 16497 6239
rect 16531 6205 16543 6239
rect 16485 6199 16543 6205
rect 16574 6196 16580 6248
rect 16632 6196 16638 6248
rect 17037 6239 17095 6245
rect 17037 6205 17049 6239
rect 17083 6236 17095 6239
rect 17218 6236 17224 6248
rect 17083 6208 17224 6236
rect 17083 6205 17095 6208
rect 17037 6199 17095 6205
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 15396 6140 15608 6168
rect 15252 6128 15258 6140
rect 15580 6112 15608 6140
rect 12667 6072 14044 6100
rect 12667 6069 12679 6072
rect 12621 6063 12679 6069
rect 14826 6060 14832 6112
rect 14884 6060 14890 6112
rect 15562 6060 15568 6112
rect 15620 6060 15626 6112
rect 16114 6060 16120 6112
rect 16172 6060 16178 6112
rect 16850 6060 16856 6112
rect 16908 6060 16914 6112
rect 552 6010 17664 6032
rect 552 5958 4366 6010
rect 4418 5958 4430 6010
rect 4482 5958 4494 6010
rect 4546 5958 4558 6010
rect 4610 5958 4622 6010
rect 4674 5958 4686 6010
rect 4738 5958 10366 6010
rect 10418 5958 10430 6010
rect 10482 5958 10494 6010
rect 10546 5958 10558 6010
rect 10610 5958 10622 6010
rect 10674 5958 10686 6010
rect 10738 5958 16366 6010
rect 16418 5958 16430 6010
rect 16482 5958 16494 6010
rect 16546 5958 16558 6010
rect 16610 5958 16622 6010
rect 16674 5958 16686 6010
rect 16738 5958 17664 6010
rect 552 5936 17664 5958
rect 1854 5856 1860 5908
rect 1912 5896 1918 5908
rect 2593 5899 2651 5905
rect 2593 5896 2605 5899
rect 1912 5868 2605 5896
rect 1912 5856 1918 5868
rect 2593 5865 2605 5868
rect 2639 5865 2651 5899
rect 2593 5859 2651 5865
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 3326 5896 3332 5908
rect 2915 5868 3332 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4295 5899 4353 5905
rect 4295 5896 4307 5899
rect 4028 5868 4307 5896
rect 4028 5856 4034 5868
rect 4295 5865 4307 5868
rect 4341 5896 4353 5899
rect 4341 5868 6316 5896
rect 4341 5865 4353 5868
rect 4295 5859 4353 5865
rect 3697 5831 3755 5837
rect 3697 5828 3709 5831
rect 2700 5800 3709 5828
rect 2700 5769 2728 5800
rect 3697 5797 3709 5800
rect 3743 5797 3755 5831
rect 3697 5791 3755 5797
rect 3896 5800 4108 5828
rect 1112 5763 1170 5769
rect 1112 5729 1124 5763
rect 1158 5760 1170 5763
rect 2501 5763 2559 5769
rect 1158 5732 2084 5760
rect 1158 5729 1170 5732
rect 1112 5723 1170 5729
rect 842 5652 848 5704
rect 900 5652 906 5704
rect 2056 5624 2084 5732
rect 2501 5729 2513 5763
rect 2547 5729 2559 5763
rect 2501 5723 2559 5729
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5729 2743 5763
rect 2685 5723 2743 5729
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5760 2835 5763
rect 2823 5732 2857 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 2406 5652 2412 5704
rect 2464 5692 2470 5704
rect 2516 5692 2544 5723
rect 2792 5692 2820 5723
rect 3050 5720 3056 5772
rect 3108 5720 3114 5772
rect 3421 5763 3479 5769
rect 3421 5729 3433 5763
rect 3467 5729 3479 5763
rect 3421 5723 3479 5729
rect 2464 5664 3280 5692
rect 2464 5652 2470 5664
rect 3053 5627 3111 5633
rect 3053 5624 3065 5627
rect 2056 5596 3065 5624
rect 3053 5593 3065 5596
rect 3099 5593 3111 5627
rect 3053 5587 3111 5593
rect 3252 5568 3280 5664
rect 3436 5624 3464 5723
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 3896 5760 3924 5800
rect 3660 5732 3924 5760
rect 3660 5720 3666 5732
rect 3970 5720 3976 5772
rect 4028 5720 4034 5772
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 3694 5692 3700 5704
rect 3568 5664 3700 5692
rect 3568 5652 3574 5664
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 4080 5701 4108 5800
rect 5626 5788 5632 5840
rect 5684 5828 5690 5840
rect 6288 5828 6316 5868
rect 7098 5856 7104 5908
rect 7156 5896 7162 5908
rect 7282 5896 7288 5908
rect 7156 5868 7288 5896
rect 7156 5856 7162 5868
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 8386 5896 8392 5908
rect 7432 5868 8392 5896
rect 7432 5856 7438 5868
rect 8386 5856 8392 5868
rect 8444 5896 8450 5908
rect 15562 5896 15568 5908
rect 8444 5868 15568 5896
rect 8444 5856 8450 5868
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 16022 5856 16028 5908
rect 16080 5856 16086 5908
rect 16114 5856 16120 5908
rect 16172 5856 16178 5908
rect 16206 5856 16212 5908
rect 16264 5896 16270 5908
rect 16264 5868 16360 5896
rect 16264 5856 16270 5868
rect 9861 5831 9919 5837
rect 5684 5800 6132 5828
rect 6288 5800 9628 5828
rect 5684 5788 5690 5800
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5729 6055 5763
rect 6104 5760 6132 5800
rect 9600 5772 9628 5800
rect 9861 5797 9873 5831
rect 9907 5828 9919 5831
rect 15194 5828 15200 5840
rect 9907 5800 10364 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 6104 5732 6285 5760
rect 5997 5723 6055 5729
rect 6273 5729 6285 5732
rect 6319 5729 6331 5763
rect 6273 5723 6331 5729
rect 3881 5695 3939 5701
rect 3881 5661 3893 5695
rect 3927 5661 3939 5695
rect 3881 5655 3939 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4890 5692 4896 5704
rect 4111 5664 4896 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 3602 5624 3608 5636
rect 3436 5596 3608 5624
rect 3602 5584 3608 5596
rect 3660 5624 3666 5636
rect 3896 5624 3924 5655
rect 4890 5652 4896 5664
rect 4948 5692 4954 5704
rect 5534 5692 5540 5704
rect 4948 5664 5540 5692
rect 4948 5652 4954 5664
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 5258 5624 5264 5636
rect 3660 5596 5264 5624
rect 3660 5584 3666 5596
rect 5258 5584 5264 5596
rect 5316 5584 5322 5636
rect 6012 5624 6040 5723
rect 6362 5720 6368 5772
rect 6420 5720 6426 5772
rect 6546 5720 6552 5772
rect 6604 5720 6610 5772
rect 7006 5720 7012 5772
rect 7064 5760 7070 5772
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 7064 5732 7113 5760
rect 7064 5720 7070 5732
rect 7101 5729 7113 5732
rect 7147 5729 7159 5763
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 7101 5723 7159 5729
rect 7208 5732 9413 5760
rect 6178 5652 6184 5704
rect 6236 5652 6242 5704
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7208 5692 7236 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9582 5720 9588 5772
rect 9640 5720 9646 5772
rect 10336 5769 10364 5800
rect 12360 5800 13492 5828
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 6880 5664 7236 5692
rect 6880 5652 6886 5664
rect 7282 5652 7288 5704
rect 7340 5692 7346 5704
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 7340 5664 7389 5692
rect 7340 5652 7346 5664
rect 7377 5661 7389 5664
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8628 5664 9137 5692
rect 8628 5652 8634 5664
rect 9125 5661 9137 5664
rect 9171 5692 9183 5695
rect 10060 5692 10088 5723
rect 9171 5664 10088 5692
rect 10336 5692 10364 5723
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 11977 5763 12035 5769
rect 11977 5760 11989 5763
rect 11388 5732 11989 5760
rect 11388 5720 11394 5732
rect 11977 5729 11989 5732
rect 12023 5729 12035 5763
rect 11977 5723 12035 5729
rect 12161 5763 12219 5769
rect 12161 5729 12173 5763
rect 12207 5729 12219 5763
rect 12161 5723 12219 5729
rect 12176 5692 12204 5723
rect 12250 5720 12256 5772
rect 12308 5720 12314 5772
rect 12360 5769 12388 5800
rect 12345 5763 12403 5769
rect 12345 5729 12357 5763
rect 12391 5729 12403 5763
rect 12345 5723 12403 5729
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 12860 5732 12909 5760
rect 12860 5720 12866 5732
rect 12897 5729 12909 5732
rect 12943 5729 12955 5763
rect 12897 5723 12955 5729
rect 12989 5763 13047 5769
rect 12989 5729 13001 5763
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 10336 5664 11836 5692
rect 12176 5664 12725 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 9416 5636 9444 5664
rect 11808 5636 11836 5664
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 13004 5692 13032 5723
rect 13262 5720 13268 5772
rect 13320 5720 13326 5772
rect 12713 5655 12771 5661
rect 12820 5664 13032 5692
rect 13464 5692 13492 5800
rect 13556 5800 14596 5828
rect 13556 5769 13584 5800
rect 14568 5772 14596 5800
rect 15120 5800 15200 5828
rect 13541 5763 13599 5769
rect 13541 5729 13553 5763
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 13630 5720 13636 5772
rect 13688 5720 13694 5772
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 13909 5763 13967 5769
rect 13909 5760 13921 5763
rect 13872 5732 13921 5760
rect 13872 5720 13878 5732
rect 13909 5729 13921 5732
rect 13955 5729 13967 5763
rect 13909 5723 13967 5729
rect 13648 5692 13676 5720
rect 13464 5664 13676 5692
rect 8662 5624 8668 5636
rect 6012 5596 8668 5624
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 8938 5584 8944 5636
rect 8996 5584 9002 5636
rect 9398 5584 9404 5636
rect 9456 5584 9462 5636
rect 9585 5627 9643 5633
rect 9585 5593 9597 5627
rect 9631 5624 9643 5627
rect 10226 5624 10232 5636
rect 9631 5596 10232 5624
rect 9631 5593 9643 5596
rect 9585 5587 9643 5593
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 11790 5584 11796 5636
rect 11848 5624 11854 5636
rect 12820 5624 12848 5664
rect 11848 5596 12848 5624
rect 11848 5584 11854 5596
rect 12894 5584 12900 5636
rect 12952 5584 12958 5636
rect 13004 5624 13032 5664
rect 13538 5624 13544 5636
rect 13004 5596 13544 5624
rect 13538 5584 13544 5596
rect 13596 5584 13602 5636
rect 13924 5624 13952 5723
rect 14550 5720 14556 5772
rect 14608 5720 14614 5772
rect 15120 5769 15148 5800
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 15580 5769 15608 5856
rect 16040 5828 16068 5856
rect 15672 5800 16068 5828
rect 14829 5763 14887 5769
rect 14829 5729 14841 5763
rect 14875 5760 14887 5763
rect 15105 5763 15163 5769
rect 15105 5760 15117 5763
rect 14875 5732 15117 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 15105 5729 15117 5732
rect 15151 5729 15163 5763
rect 15105 5723 15163 5729
rect 15381 5763 15439 5769
rect 15381 5729 15393 5763
rect 15427 5729 15439 5763
rect 15381 5723 15439 5729
rect 15565 5763 15623 5769
rect 15565 5729 15577 5763
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 14645 5627 14703 5633
rect 14645 5624 14657 5627
rect 13924 5596 14657 5624
rect 14645 5593 14657 5596
rect 14691 5593 14703 5627
rect 15396 5624 15424 5723
rect 15672 5701 15700 5800
rect 15746 5720 15752 5772
rect 15804 5720 15810 5772
rect 15933 5763 15991 5769
rect 15933 5729 15945 5763
rect 15979 5760 15991 5763
rect 16132 5760 16160 5856
rect 16332 5828 16360 5868
rect 16332 5800 16712 5828
rect 16332 5769 16360 5800
rect 15979 5732 16160 5760
rect 16301 5763 16360 5769
rect 15979 5729 15991 5732
rect 15933 5723 15991 5729
rect 16301 5729 16313 5763
rect 16347 5732 16360 5763
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 16390 5720 16396 5772
rect 16448 5760 16454 5772
rect 16684 5769 16712 5800
rect 16485 5763 16543 5769
rect 16485 5760 16497 5763
rect 16448 5732 16497 5760
rect 16448 5720 16454 5732
rect 16485 5729 16497 5732
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 16945 5763 17003 5769
rect 16945 5729 16957 5763
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 16960 5692 16988 5723
rect 17126 5720 17132 5772
rect 17184 5720 17190 5772
rect 15657 5655 15715 5661
rect 16224 5664 16988 5692
rect 16224 5633 16252 5664
rect 16209 5627 16267 5633
rect 16209 5624 16221 5627
rect 15396 5596 16221 5624
rect 14645 5587 14703 5593
rect 16209 5593 16221 5596
rect 16255 5593 16267 5627
rect 16209 5587 16267 5593
rect 16758 5584 16764 5636
rect 16816 5584 16822 5636
rect 2222 5516 2228 5568
rect 2280 5516 2286 5568
rect 3234 5516 3240 5568
rect 3292 5516 3298 5568
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6178 5556 6184 5568
rect 5859 5528 6184 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 6917 5559 6975 5565
rect 6917 5556 6929 5559
rect 6512 5528 6929 5556
rect 6512 5516 6518 5528
rect 6917 5525 6929 5528
rect 6963 5525 6975 5559
rect 6917 5519 6975 5525
rect 7285 5559 7343 5565
rect 7285 5525 7297 5559
rect 7331 5556 7343 5559
rect 8956 5556 8984 5584
rect 7331 5528 8984 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 9214 5516 9220 5568
rect 9272 5516 9278 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9677 5559 9735 5565
rect 9677 5556 9689 5559
rect 9548 5528 9689 5556
rect 9548 5516 9554 5528
rect 9677 5525 9689 5528
rect 9723 5525 9735 5559
rect 9677 5519 9735 5525
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10137 5559 10195 5565
rect 10137 5556 10149 5559
rect 10100 5528 10149 5556
rect 10100 5516 10106 5528
rect 10137 5525 10149 5528
rect 10183 5525 10195 5559
rect 10137 5519 10195 5525
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 11238 5556 11244 5568
rect 10836 5528 11244 5556
rect 10836 5516 10842 5528
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 11974 5556 11980 5568
rect 11756 5528 11980 5556
rect 11756 5516 11762 5528
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 12621 5559 12679 5565
rect 12621 5556 12633 5559
rect 12584 5528 12633 5556
rect 12584 5516 12590 5528
rect 12621 5525 12633 5528
rect 12667 5525 12679 5559
rect 12912 5556 12940 5584
rect 13173 5559 13231 5565
rect 13173 5556 13185 5559
rect 12912 5528 13185 5556
rect 12621 5519 12679 5525
rect 13173 5525 13185 5528
rect 13219 5525 13231 5559
rect 13173 5519 13231 5525
rect 13262 5516 13268 5568
rect 13320 5556 13326 5568
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 13320 5528 13369 5556
rect 13320 5516 13326 5528
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 13357 5519 13415 5525
rect 13817 5559 13875 5565
rect 13817 5525 13829 5559
rect 13863 5556 13875 5559
rect 14090 5556 14096 5568
rect 13863 5528 14096 5556
rect 13863 5525 13875 5528
rect 13817 5519 13875 5525
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 14182 5516 14188 5568
rect 14240 5556 14246 5568
rect 14921 5559 14979 5565
rect 14921 5556 14933 5559
rect 14240 5528 14933 5556
rect 14240 5516 14246 5528
rect 14921 5525 14933 5528
rect 14967 5525 14979 5559
rect 14921 5519 14979 5525
rect 15194 5516 15200 5568
rect 15252 5516 15258 5568
rect 16942 5516 16948 5568
rect 17000 5516 17006 5568
rect 552 5466 17664 5488
rect 552 5414 1366 5466
rect 1418 5414 1430 5466
rect 1482 5414 1494 5466
rect 1546 5414 1558 5466
rect 1610 5414 1622 5466
rect 1674 5414 1686 5466
rect 1738 5414 7366 5466
rect 7418 5414 7430 5466
rect 7482 5414 7494 5466
rect 7546 5414 7558 5466
rect 7610 5414 7622 5466
rect 7674 5414 7686 5466
rect 7738 5414 13366 5466
rect 13418 5414 13430 5466
rect 13482 5414 13494 5466
rect 13546 5414 13558 5466
rect 13610 5414 13622 5466
rect 13674 5414 13686 5466
rect 13738 5414 17664 5466
rect 552 5392 17664 5414
rect 937 5355 995 5361
rect 937 5321 949 5355
rect 983 5352 995 5355
rect 2041 5355 2099 5361
rect 2041 5352 2053 5355
rect 983 5324 2053 5352
rect 983 5321 995 5324
rect 937 5315 995 5321
rect 2041 5321 2053 5324
rect 2087 5321 2099 5355
rect 2041 5315 2099 5321
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 3421 5355 3479 5361
rect 3421 5352 3433 5355
rect 2915 5324 3433 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 3421 5321 3433 5324
rect 3467 5321 3479 5355
rect 3421 5315 3479 5321
rect 5629 5355 5687 5361
rect 5629 5321 5641 5355
rect 5675 5352 5687 5355
rect 6822 5352 6828 5364
rect 5675 5324 6828 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7561 5355 7619 5361
rect 7561 5321 7573 5355
rect 7607 5352 7619 5355
rect 8110 5352 8116 5364
rect 7607 5324 8116 5352
rect 7607 5321 7619 5324
rect 7561 5315 7619 5321
rect 8110 5312 8116 5324
rect 8168 5352 8174 5364
rect 8570 5352 8576 5364
rect 8168 5324 8576 5352
rect 8168 5312 8174 5324
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 9766 5352 9772 5364
rect 8680 5324 9772 5352
rect 2409 5287 2467 5293
rect 2409 5284 2421 5287
rect 1412 5256 2421 5284
rect 1412 5216 1440 5256
rect 2409 5253 2421 5256
rect 2455 5253 2467 5287
rect 4249 5287 4307 5293
rect 4249 5284 4261 5287
rect 2409 5247 2467 5253
rect 3988 5256 4261 5284
rect 2038 5216 2044 5228
rect 860 5188 1440 5216
rect 860 5157 888 5188
rect 1412 5157 1440 5188
rect 1504 5188 2044 5216
rect 845 5151 903 5157
rect 845 5117 857 5151
rect 891 5117 903 5151
rect 845 5111 903 5117
rect 1029 5151 1087 5157
rect 1029 5117 1041 5151
rect 1075 5148 1087 5151
rect 1305 5151 1363 5157
rect 1075 5120 1256 5148
rect 1075 5117 1087 5120
rect 1029 5111 1087 5117
rect 1228 5021 1256 5120
rect 1305 5117 1317 5151
rect 1351 5117 1363 5151
rect 1305 5111 1363 5117
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 1320 5080 1348 5111
rect 1504 5092 1532 5188
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2424 5216 2452 5247
rect 2424 5188 2728 5216
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2406 5148 2412 5160
rect 2363 5120 2412 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 2590 5108 2596 5160
rect 2648 5108 2654 5160
rect 1486 5080 1492 5092
rect 1320 5052 1492 5080
rect 1486 5040 1492 5052
rect 1544 5040 1550 5092
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5049 1639 5083
rect 1581 5043 1639 5049
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5080 1823 5083
rect 2009 5083 2067 5089
rect 2009 5080 2021 5083
rect 1811 5052 2021 5080
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 2009 5049 2021 5052
rect 2055 5049 2067 5083
rect 2009 5043 2067 5049
rect 1213 5015 1271 5021
rect 1213 4981 1225 5015
rect 1259 5012 1271 5015
rect 1596 5012 1624 5043
rect 2130 5040 2136 5092
rect 2188 5080 2194 5092
rect 2225 5083 2283 5089
rect 2225 5080 2237 5083
rect 2188 5052 2237 5080
rect 2188 5040 2194 5052
rect 2225 5049 2237 5052
rect 2271 5049 2283 5083
rect 2225 5043 2283 5049
rect 2501 5083 2559 5089
rect 2501 5049 2513 5083
rect 2547 5080 2559 5083
rect 2700 5080 2728 5188
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3384 5188 3801 5216
rect 3384 5176 3390 5188
rect 3789 5185 3801 5188
rect 3835 5216 3847 5219
rect 3988 5216 4016 5256
rect 4249 5253 4261 5256
rect 4295 5284 4307 5287
rect 6546 5284 6552 5296
rect 4295 5256 6552 5284
rect 4295 5253 4307 5256
rect 4249 5247 4307 5253
rect 6546 5244 6552 5256
rect 6604 5244 6610 5296
rect 8680 5284 8708 5324
rect 9766 5312 9772 5324
rect 9824 5352 9830 5364
rect 9824 5324 12756 5352
rect 9824 5312 9830 5324
rect 7024 5256 8708 5284
rect 3835 5188 4016 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 5166 5176 5172 5228
rect 5224 5176 5230 5228
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5810 5216 5816 5228
rect 5307 5188 5816 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 6052 5188 6193 5216
rect 6052 5176 6058 5188
rect 6181 5185 6193 5188
rect 6227 5216 6239 5219
rect 6270 5216 6276 5228
rect 6227 5188 6276 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 6362 5176 6368 5228
rect 6420 5216 6426 5228
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6420 5188 6469 5216
rect 6420 5176 6426 5188
rect 6457 5185 6469 5188
rect 6503 5216 6515 5219
rect 7024 5216 7052 5256
rect 8754 5244 8760 5296
rect 8812 5284 8818 5296
rect 8849 5287 8907 5293
rect 8849 5284 8861 5287
rect 8812 5256 8861 5284
rect 8812 5244 8818 5256
rect 8849 5253 8861 5256
rect 8895 5253 8907 5287
rect 8849 5247 8907 5253
rect 9398 5244 9404 5296
rect 9456 5244 9462 5296
rect 9674 5284 9680 5296
rect 9646 5244 9680 5284
rect 9732 5244 9738 5296
rect 11333 5287 11391 5293
rect 11333 5284 11345 5287
rect 9876 5256 11345 5284
rect 6503 5188 7052 5216
rect 6503 5185 6515 5188
rect 6457 5179 6515 5185
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8772 5216 8800 5244
rect 9646 5216 9674 5244
rect 8076 5188 8800 5216
rect 8956 5188 9352 5216
rect 8076 5176 8082 5188
rect 3602 5108 3608 5160
rect 3660 5108 3666 5160
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5117 3755 5151
rect 3697 5111 3755 5117
rect 2837 5083 2895 5089
rect 2837 5080 2849 5083
rect 2547 5052 2636 5080
rect 2700 5052 2849 5080
rect 2547 5049 2559 5052
rect 2501 5043 2559 5049
rect 2608 5024 2636 5052
rect 2837 5049 2849 5052
rect 2883 5049 2895 5083
rect 2837 5043 2895 5049
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 3510 5080 3516 5092
rect 3099 5052 3516 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 3510 5040 3516 5052
rect 3568 5040 3574 5092
rect 3712 5080 3740 5111
rect 3878 5108 3884 5160
rect 3936 5108 3942 5160
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5117 4123 5151
rect 4065 5111 4123 5117
rect 3970 5080 3976 5092
rect 3712 5052 3976 5080
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 1259 4984 1624 5012
rect 1259 4981 1271 4984
rect 1213 4975 1271 4981
rect 1854 4972 1860 5024
rect 1912 4972 1918 5024
rect 2590 4972 2596 5024
rect 2648 4972 2654 5024
rect 2682 4972 2688 5024
rect 2740 4972 2746 5024
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3878 5012 3884 5024
rect 3016 4984 3884 5012
rect 3016 4972 3022 4984
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 4080 5012 4108 5111
rect 4890 5108 4896 5160
rect 4948 5108 4954 5160
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 5534 5148 5540 5160
rect 5491 5120 5540 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 5092 5080 5120 5111
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 7285 5151 7343 5157
rect 7285 5148 7297 5151
rect 5776 5120 7297 5148
rect 5776 5108 5782 5120
rect 7285 5117 7297 5120
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 7374 5108 7380 5160
rect 7432 5108 7438 5160
rect 7558 5108 7564 5160
rect 7616 5148 7622 5160
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7616 5120 7665 5148
rect 7616 5108 7622 5120
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 8386 5108 8392 5160
rect 8444 5108 8450 5160
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 8536 5120 8585 5148
rect 8536 5108 8542 5120
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8662 5108 8668 5160
rect 8720 5108 8726 5160
rect 8956 5157 8984 5188
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5117 8999 5151
rect 8941 5111 8999 5117
rect 9030 5108 9036 5160
rect 9088 5108 9094 5160
rect 9324 5157 9352 5188
rect 9508 5188 9674 5216
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 9508 5148 9536 5188
rect 9876 5160 9904 5256
rect 11333 5253 11345 5256
rect 11379 5284 11391 5287
rect 11379 5256 12388 5284
rect 11379 5253 11391 5256
rect 11333 5247 11391 5253
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 10060 5188 10609 5216
rect 10060 5160 10088 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10778 5176 10784 5228
rect 10836 5176 10842 5228
rect 11425 5219 11483 5225
rect 11425 5185 11437 5219
rect 11471 5216 11483 5219
rect 11514 5216 11520 5228
rect 11471 5188 11520 5216
rect 11471 5185 11483 5188
rect 11425 5179 11483 5185
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 11716 5188 12020 5216
rect 9355 5120 9536 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 9582 5108 9588 5160
rect 9640 5108 9646 5160
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5148 9735 5151
rect 9766 5148 9772 5160
rect 9723 5120 9772 5148
rect 9723 5117 9735 5120
rect 9677 5111 9735 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 9858 5108 9864 5160
rect 9916 5108 9922 5160
rect 10042 5108 10048 5160
rect 10100 5108 10106 5160
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 10192 5120 10333 5148
rect 10192 5108 10198 5120
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5117 10563 5151
rect 10505 5111 10563 5117
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 10796 5148 10824 5176
rect 10735 5120 10824 5148
rect 10873 5151 10931 5157
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 10873 5117 10885 5151
rect 10919 5148 10931 5151
rect 10965 5151 11023 5157
rect 10965 5148 10977 5151
rect 10919 5120 10977 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 10965 5117 10977 5120
rect 11011 5117 11023 5151
rect 10965 5111 11023 5117
rect 11149 5151 11207 5157
rect 11149 5117 11161 5151
rect 11195 5148 11207 5151
rect 11238 5148 11244 5160
rect 11195 5120 11244 5148
rect 11195 5117 11207 5120
rect 11149 5111 11207 5117
rect 5994 5080 6000 5092
rect 5092 5052 6000 5080
rect 5994 5040 6000 5052
rect 6052 5040 6058 5092
rect 7392 5080 7420 5108
rect 8110 5080 8116 5092
rect 6104 5052 7328 5080
rect 7392 5052 8116 5080
rect 4154 5012 4160 5024
rect 4080 4984 4160 5012
rect 4154 4972 4160 4984
rect 4212 5012 4218 5024
rect 6104 5012 6132 5052
rect 7300 5024 7328 5052
rect 8110 5040 8116 5052
rect 8168 5080 8174 5092
rect 10060 5080 10088 5108
rect 8168 5052 10088 5080
rect 10520 5080 10548 5111
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 10520 5052 10824 5080
rect 8168 5040 8174 5052
rect 10796 5024 10824 5052
rect 4212 4984 6132 5012
rect 4212 4972 4218 4984
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 6972 4984 7113 5012
rect 6972 4972 6978 4984
rect 7101 4981 7113 4984
rect 7147 4981 7159 5015
rect 7101 4975 7159 4981
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 8478 5012 8484 5024
rect 7340 4984 8484 5012
rect 7340 4972 7346 4984
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 9217 5015 9275 5021
rect 9217 4981 9229 5015
rect 9263 5012 9275 5015
rect 9674 5012 9680 5024
rect 9263 4984 9680 5012
rect 9263 4981 9275 4984
rect 9217 4975 9275 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 5012 9919 5015
rect 10042 5012 10048 5024
rect 9907 4984 10048 5012
rect 9907 4981 9919 4984
rect 9861 4975 9919 4981
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10134 4972 10140 5024
rect 10192 4972 10198 5024
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 11716 5012 11744 5188
rect 11882 5108 11888 5160
rect 11940 5108 11946 5160
rect 11992 5150 12020 5188
rect 12158 5176 12164 5228
rect 12216 5176 12222 5228
rect 12069 5151 12127 5157
rect 12069 5150 12081 5151
rect 11992 5122 12081 5150
rect 12069 5117 12081 5122
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12360 5148 12388 5256
rect 12728 5216 12756 5324
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 12860 5324 13645 5352
rect 12860 5312 12866 5324
rect 13633 5321 13645 5324
rect 13679 5321 13691 5355
rect 13633 5315 13691 5321
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 15746 5284 15752 5296
rect 12952 5256 15752 5284
rect 12952 5244 12958 5256
rect 15746 5244 15752 5256
rect 15804 5244 15810 5296
rect 12728 5188 13952 5216
rect 12299 5120 12388 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 12158 5040 12164 5092
rect 12216 5080 12222 5092
rect 12360 5080 12388 5120
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12483 5120 12848 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12216 5052 12388 5080
rect 12216 5040 12222 5052
rect 12618 5040 12624 5092
rect 12676 5040 12682 5092
rect 12820 5080 12848 5120
rect 12894 5108 12900 5160
rect 12952 5108 12958 5160
rect 13354 5108 13360 5160
rect 13412 5148 13418 5160
rect 13541 5151 13599 5157
rect 13541 5148 13553 5151
rect 13412 5120 13553 5148
rect 13412 5108 13418 5120
rect 13541 5117 13553 5120
rect 13587 5148 13599 5151
rect 13722 5148 13728 5160
rect 13587 5120 13728 5148
rect 13587 5117 13599 5120
rect 13541 5111 13599 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 13924 5157 13952 5188
rect 14090 5176 14096 5228
rect 14148 5176 14154 5228
rect 14550 5216 14556 5228
rect 14200 5188 14556 5216
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 13909 5151 13967 5157
rect 13909 5117 13921 5151
rect 13955 5148 13967 5151
rect 14200 5148 14228 5188
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 13955 5120 14228 5148
rect 13955 5117 13967 5120
rect 13909 5111 13967 5117
rect 13832 5080 13860 5111
rect 14274 5108 14280 5160
rect 14332 5108 14338 5160
rect 14292 5080 14320 5108
rect 12820 5052 14320 5080
rect 12713 5015 12771 5021
rect 12713 5012 12725 5015
rect 10836 4984 12725 5012
rect 10836 4972 10842 4984
rect 12713 4981 12725 4984
rect 12759 4981 12771 5015
rect 12713 4975 12771 4981
rect 552 4922 17664 4944
rect 552 4870 4366 4922
rect 4418 4870 4430 4922
rect 4482 4870 4494 4922
rect 4546 4870 4558 4922
rect 4610 4870 4622 4922
rect 4674 4870 4686 4922
rect 4738 4870 10366 4922
rect 10418 4870 10430 4922
rect 10482 4870 10494 4922
rect 10546 4870 10558 4922
rect 10610 4870 10622 4922
rect 10674 4870 10686 4922
rect 10738 4870 16366 4922
rect 16418 4870 16430 4922
rect 16482 4870 16494 4922
rect 16546 4870 16558 4922
rect 16610 4870 16622 4922
rect 16674 4870 16686 4922
rect 16738 4870 17664 4922
rect 552 4848 17664 4870
rect 1486 4768 1492 4820
rect 1544 4808 1550 4820
rect 1673 4811 1731 4817
rect 1673 4808 1685 4811
rect 1544 4780 1685 4808
rect 1544 4768 1550 4780
rect 1673 4777 1685 4780
rect 1719 4777 1731 4811
rect 1673 4771 1731 4777
rect 1854 4768 1860 4820
rect 1912 4768 1918 4820
rect 2682 4768 2688 4820
rect 2740 4768 2746 4820
rect 3050 4768 3056 4820
rect 3108 4768 3114 4820
rect 5810 4808 5816 4820
rect 5276 4780 5816 4808
rect 1872 4740 1900 4768
rect 1412 4712 1900 4740
rect 2700 4740 2728 4768
rect 2700 4712 3464 4740
rect 1412 4681 1440 4712
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 1762 4632 1768 4684
rect 1820 4632 1826 4684
rect 3326 4632 3332 4684
rect 3384 4632 3390 4684
rect 3436 4681 3464 4712
rect 5000 4712 5212 4740
rect 5000 4684 5028 4712
rect 3421 4675 3479 4681
rect 3421 4641 3433 4675
rect 3467 4641 3479 4675
rect 3421 4635 3479 4641
rect 4890 4632 4896 4684
rect 4948 4632 4954 4684
rect 4982 4632 4988 4684
rect 5040 4632 5046 4684
rect 5184 4681 5212 4712
rect 5276 4681 5304 4780
rect 5810 4768 5816 4780
rect 5868 4808 5874 4820
rect 5868 4780 6132 4808
rect 5868 4768 5874 4780
rect 5813 4685 5871 4691
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4641 5319 4675
rect 5261 4635 5319 4641
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 3068 4536 3096 4567
rect 3234 4564 3240 4616
rect 3292 4564 3298 4616
rect 3510 4604 3516 4616
rect 3344 4576 3516 4604
rect 3344 4536 3372 4576
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 5092 4604 5120 4635
rect 5442 4632 5448 4684
rect 5500 4632 5506 4684
rect 5813 4651 5825 4685
rect 5859 4651 5871 4685
rect 5813 4645 5871 4651
rect 5828 4616 5856 4645
rect 5994 4632 6000 4684
rect 6052 4632 6058 4684
rect 6104 4672 6132 4780
rect 7282 4768 7288 4820
rect 7340 4768 7346 4820
rect 7944 4780 8156 4808
rect 7300 4740 7328 4768
rect 7944 4740 7972 4780
rect 6380 4712 7328 4740
rect 7852 4712 7972 4740
rect 8128 4740 8156 4780
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 8662 4808 8668 4820
rect 8536 4780 8668 4808
rect 8536 4768 8542 4780
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 10060 4780 10200 4808
rect 8128 4712 8294 4740
rect 6380 4681 6408 4712
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 6104 4644 6193 4672
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 6365 4675 6423 4681
rect 6365 4641 6377 4675
rect 6411 4641 6423 4675
rect 6365 4635 6423 4641
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 6917 4675 6975 4681
rect 6917 4672 6929 4675
rect 6604 4644 6929 4672
rect 6604 4632 6610 4644
rect 6917 4641 6929 4644
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 7190 4632 7196 4684
rect 7248 4632 7254 4684
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 7558 4672 7564 4684
rect 7340 4644 7564 4672
rect 7340 4632 7346 4644
rect 7558 4632 7564 4644
rect 7616 4670 7622 4684
rect 7653 4675 7711 4681
rect 7653 4670 7665 4675
rect 7616 4642 7665 4670
rect 7616 4632 7622 4642
rect 7653 4641 7665 4642
rect 7699 4641 7711 4675
rect 7852 4672 7880 4712
rect 7653 4635 7711 4641
rect 7760 4644 7880 4672
rect 5092 4576 5212 4604
rect 4706 4536 4712 4548
rect 3068 4508 3372 4536
rect 3436 4508 4712 4536
rect 1210 4428 1216 4480
rect 1268 4428 1274 4480
rect 1670 4428 1676 4480
rect 1728 4468 1734 4480
rect 3436 4468 3464 4508
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 5184 4536 5212 4576
rect 5810 4564 5816 4616
rect 5868 4564 5874 4616
rect 6012 4536 6040 4632
rect 6086 4564 6092 4616
rect 6144 4564 6150 4616
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7760 4604 7788 4644
rect 8018 4632 8024 4684
rect 8076 4632 8082 4684
rect 8266 4681 8294 4712
rect 9490 4700 9496 4752
rect 9548 4740 9554 4752
rect 10060 4740 10088 4780
rect 9548 4712 10088 4740
rect 9548 4700 9554 4712
rect 8217 4675 8294 4681
rect 8217 4641 8229 4675
rect 8263 4644 8294 4675
rect 8263 4641 8275 4644
rect 8217 4635 8275 4641
rect 8478 4632 8484 4684
rect 8536 4632 8542 4684
rect 9048 4644 9536 4672
rect 7423 4576 7788 4604
rect 7837 4607 7895 4613
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4596 7987 4607
rect 8110 4596 8116 4616
rect 7975 4573 8116 4596
rect 7929 4568 8116 4573
rect 7929 4567 7987 4568
rect 5184 4508 6040 4536
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 7852 4536 7880 4567
rect 8110 4564 8116 4568
rect 8168 4564 8174 4616
rect 8496 4536 8524 4632
rect 9048 4616 9076 4644
rect 9030 4564 9036 4616
rect 9088 4564 9094 4616
rect 9398 4564 9404 4616
rect 9456 4564 9462 4616
rect 9508 4604 9536 4644
rect 9582 4632 9588 4684
rect 9640 4632 9646 4684
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 10172 4681 10200 4780
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11330 4808 11336 4820
rect 11112 4780 11336 4808
rect 11112 4768 11118 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 11977 4811 12035 4817
rect 11977 4808 11989 4811
rect 11940 4780 11989 4808
rect 11940 4768 11946 4780
rect 11977 4777 11989 4780
rect 12023 4777 12035 4811
rect 11977 4771 12035 4777
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 12158 4768 12164 4820
rect 12216 4768 12222 4820
rect 11609 4743 11667 4749
rect 11609 4709 11621 4743
rect 11655 4740 11667 4743
rect 11698 4740 11704 4752
rect 11655 4712 11704 4740
rect 11655 4709 11667 4712
rect 11609 4703 11667 4709
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 11790 4700 11796 4752
rect 11848 4700 11854 4752
rect 9861 4675 9919 4681
rect 9861 4674 9873 4675
rect 9784 4672 9873 4674
rect 9732 4646 9873 4672
rect 9732 4644 9812 4646
rect 9732 4632 9738 4644
rect 9861 4641 9873 4646
rect 9907 4641 9919 4675
rect 9861 4635 9919 4641
rect 9965 4675 10023 4681
rect 9965 4641 9977 4675
rect 10011 4641 10023 4675
rect 9965 4635 10023 4641
rect 10137 4675 10200 4681
rect 10137 4641 10149 4675
rect 10183 4644 10200 4675
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9508 4576 9781 4604
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 9968 4604 9996 4635
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 12084 4672 12112 4768
rect 11572 4644 12112 4672
rect 12176 4672 12204 4768
rect 14458 4700 14464 4752
rect 14516 4740 14522 4752
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 14516 4712 14657 4740
rect 14516 4700 14522 4712
rect 14645 4709 14657 4712
rect 14691 4740 14703 4743
rect 14691 4712 14964 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 12176 4644 12357 4672
rect 11572 4632 11578 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 13170 4632 13176 4684
rect 13228 4672 13234 4684
rect 14936 4681 14964 4712
rect 15654 4700 15660 4752
rect 15712 4700 15718 4752
rect 13725 4675 13783 4681
rect 13725 4672 13737 4675
rect 13228 4644 13737 4672
rect 13228 4632 13234 4644
rect 13725 4641 13737 4644
rect 13771 4641 13783 4675
rect 13725 4635 13783 4641
rect 14829 4675 14887 4681
rect 14829 4641 14841 4675
rect 14875 4641 14887 4675
rect 14829 4635 14887 4641
rect 14921 4675 14979 4681
rect 14921 4641 14933 4675
rect 14967 4641 14979 4675
rect 14921 4635 14979 4641
rect 10778 4604 10784 4616
rect 9968 4576 10784 4604
rect 9674 4536 9680 4548
rect 6696 4508 7512 4536
rect 7852 4508 8294 4536
rect 8496 4508 9680 4536
rect 6696 4496 6702 4508
rect 1728 4440 3464 4468
rect 1728 4428 1734 4440
rect 3510 4428 3516 4480
rect 3568 4468 3574 4480
rect 3605 4471 3663 4477
rect 3605 4468 3617 4471
rect 3568 4440 3617 4468
rect 3568 4428 3574 4440
rect 3605 4437 3617 4440
rect 3651 4437 3663 4471
rect 3605 4431 3663 4437
rect 5629 4471 5687 4477
rect 5629 4437 5641 4471
rect 5675 4468 5687 4471
rect 6270 4468 6276 4480
rect 5675 4440 6276 4468
rect 5675 4437 5687 4440
rect 5629 4431 5687 4437
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4468 6607 4471
rect 6914 4468 6920 4480
rect 6595 4440 6920 4468
rect 6595 4437 6607 4440
rect 6549 4431 6607 4437
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7484 4477 7512 4508
rect 7469 4471 7527 4477
rect 7469 4437 7481 4471
rect 7515 4437 7527 4471
rect 8266 4468 8294 4508
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 9784 4536 9812 4567
rect 9858 4536 9864 4548
rect 9784 4508 9864 4536
rect 9858 4496 9864 4508
rect 9916 4496 9922 4548
rect 9968 4468 9996 4576
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 12069 4607 12127 4613
rect 12069 4573 12081 4607
rect 12115 4604 12127 4607
rect 12250 4604 12256 4616
rect 12115 4576 12256 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 12250 4564 12256 4576
rect 12308 4564 12314 4616
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 13817 4607 13875 4613
rect 13817 4604 13829 4607
rect 12768 4576 13829 4604
rect 12768 4564 12774 4576
rect 13817 4573 13829 4576
rect 13863 4573 13875 4607
rect 13817 4567 13875 4573
rect 13906 4564 13912 4616
rect 13964 4564 13970 4616
rect 13998 4564 14004 4616
rect 14056 4564 14062 4616
rect 14844 4604 14872 4635
rect 15102 4632 15108 4684
rect 15160 4632 15166 4684
rect 15672 4604 15700 4700
rect 16577 4675 16635 4681
rect 16577 4641 16589 4675
rect 16623 4672 16635 4675
rect 16758 4672 16764 4684
rect 16623 4644 16764 4672
rect 16623 4641 16635 4644
rect 16577 4635 16635 4641
rect 16758 4632 16764 4644
rect 16816 4632 16822 4684
rect 14844 4576 15700 4604
rect 16669 4607 16727 4613
rect 16669 4573 16681 4607
rect 16715 4604 16727 4607
rect 16850 4604 16856 4616
rect 16715 4576 16856 4604
rect 16715 4573 16727 4576
rect 16669 4567 16727 4573
rect 16850 4564 16856 4576
rect 16908 4604 16914 4616
rect 17034 4604 17040 4616
rect 16908 4576 17040 4604
rect 16908 4564 16914 4576
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 8266 4440 9996 4468
rect 7469 4431 7527 4437
rect 14182 4428 14188 4480
rect 14240 4428 14246 4480
rect 14458 4428 14464 4480
rect 14516 4428 14522 4480
rect 14642 4428 14648 4480
rect 14700 4468 14706 4480
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14700 4440 15025 4468
rect 14700 4428 14706 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15013 4431 15071 4437
rect 16206 4428 16212 4480
rect 16264 4428 16270 4480
rect 552 4378 17664 4400
rect 552 4326 1366 4378
rect 1418 4326 1430 4378
rect 1482 4326 1494 4378
rect 1546 4326 1558 4378
rect 1610 4326 1622 4378
rect 1674 4326 1686 4378
rect 1738 4326 7366 4378
rect 7418 4326 7430 4378
rect 7482 4326 7494 4378
rect 7546 4326 7558 4378
rect 7610 4326 7622 4378
rect 7674 4326 7686 4378
rect 7738 4326 13366 4378
rect 13418 4326 13430 4378
rect 13482 4326 13494 4378
rect 13546 4326 13558 4378
rect 13610 4326 13622 4378
rect 13674 4326 13686 4378
rect 13738 4326 17664 4378
rect 552 4304 17664 4326
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 4212 4236 4629 4264
rect 4212 4224 4218 4236
rect 4617 4233 4629 4236
rect 4663 4264 4675 4267
rect 5442 4264 5448 4276
rect 4663 4236 5448 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 6181 4267 6239 4273
rect 6181 4233 6193 4267
rect 6227 4264 6239 4267
rect 6227 4236 7144 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 5166 4196 5172 4208
rect 4764 4168 5172 4196
rect 4764 4156 4770 4168
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 6546 4196 6552 4208
rect 5736 4168 6552 4196
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 1872 4100 3249 4128
rect 842 4020 848 4072
rect 900 4060 906 4072
rect 1872 4060 1900 4100
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 900 4032 1900 4060
rect 900 4020 906 4032
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 3510 4069 3516 4072
rect 2501 4063 2559 4069
rect 2501 4060 2513 4063
rect 2372 4032 2513 4060
rect 2372 4020 2378 4032
rect 2501 4029 2513 4032
rect 2547 4029 2559 4063
rect 2501 4023 2559 4029
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4029 2743 4063
rect 3504 4060 3516 4069
rect 3471 4032 3516 4060
rect 2685 4023 2743 4029
rect 3504 4023 3516 4032
rect 1112 3995 1170 4001
rect 1112 3961 1124 3995
rect 1158 3992 1170 3995
rect 1210 3992 1216 4004
rect 1158 3964 1216 3992
rect 1158 3961 1170 3964
rect 1112 3955 1170 3961
rect 1210 3952 1216 3964
rect 1268 3952 1274 4004
rect 2700 3936 2728 4023
rect 3510 4020 3516 4023
rect 3568 4020 3574 4072
rect 3878 4020 3884 4072
rect 3936 4060 3942 4072
rect 5626 4060 5632 4072
rect 3936 4032 5632 4060
rect 3936 4020 3942 4032
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 5736 4069 5764 4168
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 7116 4196 7144 4236
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 11238 4264 11244 4276
rect 7248 4236 11244 4264
rect 7248 4224 7254 4236
rect 11238 4224 11244 4236
rect 11296 4264 11302 4276
rect 11425 4267 11483 4273
rect 11425 4264 11437 4267
rect 11296 4236 11437 4264
rect 11296 4224 11302 4236
rect 7561 4199 7619 4205
rect 7561 4196 7573 4199
rect 7116 4168 7573 4196
rect 7561 4165 7573 4168
rect 7607 4165 7619 4199
rect 8018 4196 8024 4208
rect 7561 4159 7619 4165
rect 7668 4168 8024 4196
rect 6822 4128 6828 4140
rect 5828 4100 6828 4128
rect 5828 4069 5856 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4029 5871 4063
rect 5813 4023 5871 4029
rect 5994 4020 6000 4072
rect 6052 4020 6058 4072
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4029 6147 4063
rect 6089 4023 6147 4029
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3992 2927 3995
rect 5534 3992 5540 4004
rect 2915 3964 5540 3992
rect 2915 3961 2927 3964
rect 2869 3955 2927 3961
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 6104 3992 6132 4023
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 6328 4032 6377 4060
rect 6328 4020 6334 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 6972 4032 7389 4060
rect 6972 4020 6978 4032
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7377 4023 7435 4029
rect 5736 3964 6132 3992
rect 7576 3992 7604 4159
rect 7668 4137 7696 4168
rect 8018 4156 8024 4168
rect 8076 4156 8082 4208
rect 8478 4156 8484 4208
rect 8536 4196 8542 4208
rect 11054 4196 11060 4208
rect 8536 4168 11060 4196
rect 8536 4156 8542 4168
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 10962 4128 10968 4140
rect 8168 4100 10968 4128
rect 8168 4088 8174 4100
rect 10962 4088 10968 4100
rect 11020 4128 11026 4140
rect 11348 4137 11376 4236
rect 11425 4233 11437 4236
rect 11471 4233 11483 4267
rect 13541 4267 13599 4273
rect 13541 4264 13553 4267
rect 11425 4227 11483 4233
rect 13004 4236 13553 4264
rect 11333 4131 11391 4137
rect 11020 4100 11100 4128
rect 11020 4088 11026 4100
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 9030 4060 9036 4072
rect 7800 4032 9036 4060
rect 7800 4020 7806 4032
rect 9030 4020 9036 4032
rect 9088 4060 9094 4072
rect 9585 4063 9643 4069
rect 9585 4060 9597 4063
rect 9088 4032 9597 4060
rect 9088 4020 9094 4032
rect 9585 4029 9597 4032
rect 9631 4029 9643 4063
rect 9585 4023 9643 4029
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10042 4060 10048 4072
rect 9916 4032 10048 4060
rect 9916 4020 9922 4032
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 11072 4069 11100 4100
rect 11333 4097 11345 4131
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 12250 4088 12256 4140
rect 12308 4128 12314 4140
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12308 4100 12633 4128
rect 12308 4088 12314 4100
rect 12621 4097 12633 4100
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 12802 4088 12808 4140
rect 12860 4088 12866 4140
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13004 4128 13032 4236
rect 13541 4233 13553 4236
rect 13587 4233 13599 4267
rect 13541 4227 13599 4233
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14366 4264 14372 4276
rect 14056 4236 14372 4264
rect 14056 4224 14062 4236
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 14550 4224 14556 4276
rect 14608 4224 14614 4276
rect 15102 4224 15108 4276
rect 15160 4224 15166 4276
rect 15654 4224 15660 4276
rect 15712 4224 15718 4276
rect 14016 4196 14044 4224
rect 13556 4168 14044 4196
rect 13556 4128 13584 4168
rect 14461 4131 14519 4137
rect 14461 4128 14473 4131
rect 12943 4100 13032 4128
rect 13096 4100 13584 4128
rect 13648 4100 14473 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4029 11115 4063
rect 11057 4023 11115 4029
rect 11514 4020 11520 4072
rect 11572 4060 11578 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11572 4032 11621 4060
rect 11572 4020 11578 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 12345 4063 12403 4069
rect 12345 4029 12357 4063
rect 12391 4029 12403 4063
rect 12820 4060 12848 4088
rect 13096 4069 13124 4100
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12820 4032 13001 4060
rect 12345 4023 12403 4029
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 9214 3992 9220 4004
rect 7576 3964 9220 3992
rect 5736 3936 5764 3964
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 9674 3952 9680 4004
rect 9732 3992 9738 4004
rect 12360 3992 12388 4023
rect 13170 4020 13176 4072
rect 13228 4060 13234 4072
rect 13648 4060 13676 4100
rect 14461 4097 14473 4100
rect 14507 4097 14519 4131
rect 14568 4128 14596 4224
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14568 4100 14657 4128
rect 14461 4091 14519 4097
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4128 14795 4131
rect 14826 4128 14832 4140
rect 14783 4100 14832 4128
rect 14783 4097 14795 4100
rect 14737 4091 14795 4097
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 13228 4032 13676 4060
rect 13228 4020 13234 4032
rect 13814 4020 13820 4072
rect 13872 4020 13878 4072
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4029 13967 4063
rect 13909 4023 13967 4029
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14090 4060 14096 4072
rect 14047 4032 14096 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 13446 3992 13452 4004
rect 9732 3964 13452 3992
rect 9732 3952 9738 3964
rect 13446 3952 13452 3964
rect 13504 3992 13510 4004
rect 13924 3992 13952 4023
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 14553 4063 14611 4069
rect 14553 4029 14565 4063
rect 14599 4060 14611 4063
rect 15120 4060 15148 4224
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 15672 4128 15700 4224
rect 16117 4199 16175 4205
rect 16117 4165 16129 4199
rect 16163 4196 16175 4199
rect 16758 4196 16764 4208
rect 16163 4168 16764 4196
rect 16163 4165 16175 4168
rect 16117 4159 16175 4165
rect 16758 4156 16764 4168
rect 16816 4156 16822 4208
rect 16209 4131 16267 4137
rect 15252 4100 15424 4128
rect 15672 4100 16068 4128
rect 15252 4088 15258 4100
rect 15396 4069 15424 4100
rect 16040 4069 16068 4100
rect 16209 4097 16221 4131
rect 16255 4128 16267 4131
rect 16255 4100 16988 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 16960 4072 16988 4100
rect 14599 4032 15148 4060
rect 15289 4063 15347 4069
rect 14599 4029 14611 4032
rect 14553 4023 14611 4029
rect 15289 4029 15301 4063
rect 15335 4029 15347 4063
rect 15289 4023 15347 4029
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4029 15439 4063
rect 15381 4023 15439 4029
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15703 4032 15853 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 15841 4029 15853 4032
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 16025 4063 16083 4069
rect 16025 4029 16037 4063
rect 16071 4029 16083 4063
rect 16025 4023 16083 4029
rect 13504 3964 13952 3992
rect 13504 3952 13510 3964
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 1820 3896 2237 3924
rect 1820 3884 1826 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 2225 3887 2283 3893
rect 2314 3884 2320 3936
rect 2372 3884 2378 3936
rect 2682 3884 2688 3936
rect 2740 3884 2746 3936
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 3418 3924 3424 3936
rect 3007 3896 3424 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 3418 3884 3424 3896
rect 3476 3924 3482 3936
rect 4890 3924 4896 3936
rect 3476 3896 4896 3924
rect 3476 3884 3482 3896
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 5718 3884 5724 3936
rect 5776 3884 5782 3936
rect 6362 3884 6368 3936
rect 6420 3924 6426 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 6420 3896 6561 3924
rect 6420 3884 6426 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 7190 3884 7196 3936
rect 7248 3884 7254 3936
rect 9769 3927 9827 3933
rect 9769 3893 9781 3927
rect 9815 3924 9827 3927
rect 10042 3924 10048 3936
rect 9815 3896 10048 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 13354 3884 13360 3936
rect 13412 3884 13418 3936
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 14200 3924 14228 4023
rect 15304 3992 15332 4023
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 16172 4032 16313 4060
rect 16172 4020 16178 4032
rect 16301 4029 16313 4032
rect 16347 4029 16359 4063
rect 16301 4023 16359 4029
rect 16758 4020 16764 4072
rect 16816 4020 16822 4072
rect 16942 4020 16948 4072
rect 17000 4020 17006 4072
rect 17310 4020 17316 4072
rect 17368 4020 17374 4072
rect 14568 3964 15332 3992
rect 15749 3995 15807 4001
rect 14568 3936 14596 3964
rect 15749 3961 15761 3995
rect 15795 3992 15807 3995
rect 16850 3992 16856 4004
rect 15795 3964 16856 3992
rect 15795 3961 15807 3964
rect 15749 3955 15807 3961
rect 16850 3952 16856 3964
rect 16908 3992 16914 4004
rect 17221 3995 17279 4001
rect 17221 3992 17233 3995
rect 16908 3964 17233 3992
rect 16908 3952 16914 3964
rect 17221 3961 17233 3964
rect 17267 3961 17279 3995
rect 17221 3955 17279 3961
rect 13596 3896 14228 3924
rect 13596 3884 13602 3896
rect 14274 3884 14280 3936
rect 14332 3884 14338 3936
rect 14550 3884 14556 3936
rect 14608 3884 14614 3936
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 15105 3927 15163 3933
rect 15105 3924 15117 3927
rect 14884 3896 15117 3924
rect 14884 3884 14890 3896
rect 15105 3893 15117 3896
rect 15151 3893 15163 3927
rect 15105 3887 15163 3893
rect 552 3834 17664 3856
rect 552 3782 4366 3834
rect 4418 3782 4430 3834
rect 4482 3782 4494 3834
rect 4546 3782 4558 3834
rect 4610 3782 4622 3834
rect 4674 3782 4686 3834
rect 4738 3782 10366 3834
rect 10418 3782 10430 3834
rect 10482 3782 10494 3834
rect 10546 3782 10558 3834
rect 10610 3782 10622 3834
rect 10674 3782 10686 3834
rect 10738 3782 16366 3834
rect 16418 3782 16430 3834
rect 16482 3782 16494 3834
rect 16546 3782 16558 3834
rect 16610 3782 16622 3834
rect 16674 3782 16686 3834
rect 16738 3782 17664 3834
rect 552 3760 17664 3782
rect 2225 3723 2283 3729
rect 2225 3720 2237 3723
rect 1964 3692 2237 3720
rect 1964 3448 1992 3692
rect 2225 3689 2237 3692
rect 2271 3689 2283 3723
rect 2225 3683 2283 3689
rect 2314 3680 2320 3732
rect 2372 3680 2378 3732
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 2866 3720 2872 3732
rect 2823 3692 2872 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 2866 3680 2872 3692
rect 2924 3720 2930 3732
rect 5442 3720 5448 3732
rect 2924 3692 5448 3720
rect 2924 3680 2930 3692
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 8110 3720 8116 3732
rect 6052 3692 8116 3720
rect 6052 3680 6058 3692
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 9122 3720 9128 3732
rect 8956 3692 9128 3720
rect 2332 3652 2360 3680
rect 2682 3652 2688 3664
rect 2056 3624 2360 3652
rect 2608 3624 2688 3652
rect 2056 3593 2084 3624
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3553 2099 3587
rect 2041 3547 2099 3553
rect 2130 3544 2136 3596
rect 2188 3584 2194 3596
rect 2317 3587 2375 3593
rect 2317 3584 2329 3587
rect 2188 3556 2329 3584
rect 2188 3544 2194 3556
rect 2317 3553 2329 3556
rect 2363 3553 2375 3587
rect 2317 3547 2375 3553
rect 2406 3544 2412 3596
rect 2464 3544 2470 3596
rect 2608 3593 2636 3624
rect 2682 3612 2688 3624
rect 2740 3652 2746 3664
rect 2740 3624 3832 3652
rect 2740 3612 2746 3624
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3553 2651 3587
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 2593 3547 2651 3553
rect 2792 3556 2881 3584
rect 2792 3528 2820 3556
rect 2869 3553 2881 3556
rect 2915 3584 2927 3587
rect 3142 3584 3148 3596
rect 2915 3556 3148 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3804 3593 3832 3624
rect 4982 3612 4988 3664
rect 5040 3612 5046 3664
rect 5258 3612 5264 3664
rect 5316 3612 5322 3664
rect 5902 3612 5908 3664
rect 5960 3652 5966 3664
rect 6089 3655 6147 3661
rect 6089 3652 6101 3655
rect 5960 3624 6101 3652
rect 5960 3612 5966 3624
rect 6089 3621 6101 3624
rect 6135 3621 6147 3655
rect 6089 3615 6147 3621
rect 6273 3655 6331 3661
rect 6273 3621 6285 3655
rect 6319 3652 6331 3655
rect 8386 3652 8392 3664
rect 6319 3624 7972 3652
rect 6319 3621 6331 3624
rect 6273 3615 6331 3621
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3584 3847 3587
rect 4154 3584 4160 3596
rect 3835 3556 4160 3584
rect 3835 3553 3847 3556
rect 3789 3547 3847 3553
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 5000 3584 5028 3612
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5000 3556 5457 3584
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 6365 3587 6423 3593
rect 6365 3553 6377 3587
rect 6411 3553 6423 3587
rect 6546 3584 6552 3596
rect 6365 3547 6423 3553
rect 6472 3556 6552 3584
rect 2774 3476 2780 3528
rect 2832 3476 2838 3528
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 3878 3516 3884 3528
rect 3559 3488 3884 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6380 3516 6408 3547
rect 6144 3488 6408 3516
rect 6144 3476 6150 3488
rect 2866 3448 2872 3460
rect 1964 3420 2872 3448
rect 2866 3408 2872 3420
rect 2924 3408 2930 3460
rect 5629 3451 5687 3457
rect 5629 3417 5641 3451
rect 5675 3448 5687 3451
rect 6472 3448 6500 3556
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 7098 3544 7104 3596
rect 7156 3584 7162 3596
rect 7944 3593 7972 3624
rect 8036 3624 8392 3652
rect 8036 3593 8064 3624
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 8956 3661 8984 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9766 3680 9772 3732
rect 9824 3680 9830 3732
rect 9858 3680 9864 3732
rect 9916 3680 9922 3732
rect 10042 3680 10048 3732
rect 10100 3680 10106 3732
rect 10410 3680 10416 3732
rect 10468 3720 10474 3732
rect 11238 3720 11244 3732
rect 10468 3692 11244 3720
rect 10468 3680 10474 3692
rect 11238 3680 11244 3692
rect 11296 3720 11302 3732
rect 11606 3720 11612 3732
rect 11296 3692 11612 3720
rect 11296 3680 11302 3692
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 12434 3680 12440 3732
rect 12492 3680 12498 3732
rect 13262 3680 13268 3732
rect 13320 3680 13326 3732
rect 13446 3680 13452 3732
rect 13504 3680 13510 3732
rect 13814 3680 13820 3732
rect 13872 3680 13878 3732
rect 13906 3680 13912 3732
rect 13964 3680 13970 3732
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 15010 3720 15016 3732
rect 14240 3692 15016 3720
rect 14240 3680 14246 3692
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 8941 3655 8999 3661
rect 8941 3621 8953 3655
rect 8987 3621 8999 3655
rect 8941 3615 8999 3621
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 9493 3655 9551 3661
rect 9493 3652 9505 3655
rect 9272 3624 9505 3652
rect 9272 3612 9278 3624
rect 9493 3621 9505 3624
rect 9539 3621 9551 3655
rect 9493 3615 9551 3621
rect 9784 3593 9812 3680
rect 9876 3652 9904 3680
rect 10060 3652 10088 3680
rect 12069 3655 12127 3661
rect 9876 3624 9996 3652
rect 10060 3624 10548 3652
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 7156 3556 7849 3584
rect 7156 3544 7162 3556
rect 7837 3553 7849 3556
rect 7883 3553 7895 3587
rect 7837 3547 7895 3553
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3553 7987 3587
rect 7929 3547 7987 3553
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3553 8079 3587
rect 8021 3547 8079 3553
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8205 3547 8263 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 9171 3556 9781 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9769 3553 9781 3556
rect 9815 3553 9827 3587
rect 9769 3547 9827 3553
rect 7944 3516 7972 3547
rect 8220 3516 8248 3547
rect 9858 3544 9864 3596
rect 9916 3544 9922 3596
rect 9968 3593 9996 3624
rect 9953 3587 10011 3593
rect 9953 3553 9965 3587
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 10100 3556 10149 3584
rect 10100 3544 10106 3556
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 10520 3593 10548 3624
rect 12069 3621 12081 3655
rect 12115 3652 12127 3655
rect 12452 3652 12480 3680
rect 12115 3624 12480 3652
rect 12115 3621 12127 3624
rect 12069 3615 12127 3621
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 10284 3556 10333 3584
rect 10284 3544 10290 3556
rect 10321 3553 10333 3556
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11020 3556 12020 3584
rect 11020 3544 11026 3556
rect 10060 3516 10088 3544
rect 7944 3488 8064 3516
rect 8220 3488 10088 3516
rect 5675 3420 6500 3448
rect 6549 3451 6607 3457
rect 5675 3417 5687 3420
rect 5629 3411 5687 3417
rect 6549 3417 6561 3451
rect 6595 3448 6607 3451
rect 7098 3448 7104 3460
rect 6595 3420 7104 3448
rect 6595 3417 6607 3420
rect 6549 3411 6607 3417
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 8036 3448 8064 3488
rect 10410 3476 10416 3528
rect 10468 3476 10474 3528
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 11882 3516 11888 3528
rect 10827 3488 11888 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 8938 3448 8944 3460
rect 7208 3420 7972 3448
rect 8036 3420 8944 3448
rect 1854 3340 1860 3392
rect 1912 3340 1918 3392
rect 2406 3340 2412 3392
rect 2464 3340 2470 3392
rect 5905 3383 5963 3389
rect 5905 3349 5917 3383
rect 5951 3380 5963 3383
rect 5994 3380 6000 3392
rect 5951 3352 6000 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7208 3380 7236 3420
rect 6880 3352 7236 3380
rect 7561 3383 7619 3389
rect 6880 3340 6886 3352
rect 7561 3349 7573 3383
rect 7607 3380 7619 3383
rect 7834 3380 7840 3392
rect 7607 3352 7840 3380
rect 7607 3349 7619 3352
rect 7561 3343 7619 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 7944 3380 7972 3420
rect 8938 3408 8944 3420
rect 8996 3408 9002 3460
rect 9309 3451 9367 3457
rect 9309 3417 9321 3451
rect 9355 3448 9367 3451
rect 10612 3448 10640 3479
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 11992 3516 12020 3556
rect 12158 3544 12164 3596
rect 12216 3544 12222 3596
rect 12452 3593 12480 3624
rect 13280 3593 13308 3680
rect 13464 3652 13492 3680
rect 13372 3624 13492 3652
rect 13372 3593 13400 3624
rect 13832 3593 13860 3680
rect 14384 3624 14780 3652
rect 12429 3587 12487 3593
rect 12429 3553 12441 3587
rect 12475 3553 12487 3587
rect 12429 3547 12487 3553
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 13081 3587 13139 3593
rect 12667 3556 12701 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 13081 3553 13093 3587
rect 13127 3553 13139 3587
rect 13081 3547 13139 3553
rect 13265 3587 13323 3593
rect 13265 3553 13277 3587
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 13449 3587 13507 3593
rect 13449 3553 13461 3587
rect 13495 3584 13507 3587
rect 13817 3587 13875 3593
rect 13495 3556 13768 3584
rect 13495 3553 13507 3556
rect 13449 3547 13507 3553
rect 12636 3516 12664 3547
rect 12894 3516 12900 3528
rect 11992 3488 12900 3516
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13096 3516 13124 3547
rect 13538 3516 13544 3528
rect 13096 3488 13544 3516
rect 9355 3420 10640 3448
rect 9355 3417 9367 3420
rect 9309 3411 9367 3417
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 11701 3451 11759 3457
rect 11701 3448 11713 3451
rect 11572 3420 11713 3448
rect 11572 3408 11578 3420
rect 11701 3417 11713 3420
rect 11747 3417 11759 3451
rect 11701 3411 11759 3417
rect 11790 3408 11796 3460
rect 11848 3448 11854 3460
rect 12345 3451 12403 3457
rect 12345 3448 12357 3451
rect 11848 3420 12357 3448
rect 11848 3408 11854 3420
rect 12345 3417 12357 3420
rect 12391 3448 12403 3451
rect 13096 3448 13124 3488
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 13740 3516 13768 3556
rect 13817 3553 13829 3587
rect 13863 3553 13875 3587
rect 13817 3547 13875 3553
rect 13998 3544 14004 3596
rect 14056 3544 14062 3596
rect 14384 3584 14412 3624
rect 14752 3596 14780 3624
rect 16500 3624 16896 3652
rect 14108 3556 14412 3584
rect 14108 3516 14136 3556
rect 14458 3544 14464 3596
rect 14516 3544 14522 3596
rect 14734 3544 14740 3596
rect 14792 3544 14798 3596
rect 16500 3593 16528 3624
rect 16868 3596 16896 3624
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3553 16543 3587
rect 16485 3547 16543 3553
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3553 16819 3587
rect 16761 3547 16819 3553
rect 13740 3488 14136 3516
rect 14182 3476 14188 3528
rect 14240 3476 14246 3528
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14642 3516 14648 3528
rect 14415 3488 14648 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 14292 3448 14320 3479
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15378 3516 15384 3528
rect 15068 3488 15384 3516
rect 15068 3476 15074 3488
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 16206 3476 16212 3528
rect 16264 3516 16270 3528
rect 16393 3519 16451 3525
rect 16393 3516 16405 3519
rect 16264 3488 16405 3516
rect 16264 3476 16270 3488
rect 16393 3485 16405 3488
rect 16439 3485 16451 3519
rect 16776 3516 16804 3547
rect 16850 3544 16856 3596
rect 16908 3544 16914 3596
rect 17034 3516 17040 3528
rect 16776 3488 17040 3516
rect 16393 3479 16451 3485
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 12391 3420 13124 3448
rect 14016 3420 14320 3448
rect 12391 3417 12403 3420
rect 12345 3411 12403 3417
rect 14016 3392 14044 3420
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 16117 3451 16175 3457
rect 16117 3448 16129 3451
rect 14608 3420 16129 3448
rect 14608 3408 14614 3420
rect 16117 3417 16129 3420
rect 16163 3417 16175 3451
rect 16117 3411 16175 3417
rect 10410 3380 10416 3392
rect 7944 3352 10416 3380
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 11054 3340 11060 3392
rect 11112 3380 11118 3392
rect 11609 3383 11667 3389
rect 11609 3380 11621 3383
rect 11112 3352 11621 3380
rect 11112 3340 11118 3352
rect 11609 3349 11621 3352
rect 11655 3349 11667 3383
rect 11609 3343 11667 3349
rect 12250 3340 12256 3392
rect 12308 3380 12314 3392
rect 12529 3383 12587 3389
rect 12529 3380 12541 3383
rect 12308 3352 12541 3380
rect 12308 3340 12314 3352
rect 12529 3349 12541 3352
rect 12575 3349 12587 3383
rect 12529 3343 12587 3349
rect 13725 3383 13783 3389
rect 13725 3349 13737 3383
rect 13771 3380 13783 3383
rect 13906 3380 13912 3392
rect 13771 3352 13912 3380
rect 13771 3349 13783 3352
rect 13725 3343 13783 3349
rect 13906 3340 13912 3352
rect 13964 3340 13970 3392
rect 13998 3340 14004 3392
rect 14056 3340 14062 3392
rect 14642 3340 14648 3392
rect 14700 3340 14706 3392
rect 16758 3340 16764 3392
rect 16816 3380 16822 3392
rect 16853 3383 16911 3389
rect 16853 3380 16865 3383
rect 16816 3352 16865 3380
rect 16816 3340 16822 3352
rect 16853 3349 16865 3352
rect 16899 3349 16911 3383
rect 16853 3343 16911 3349
rect 17221 3383 17279 3389
rect 17221 3349 17233 3383
rect 17267 3380 17279 3383
rect 17267 3352 17724 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 552 3290 17664 3312
rect 552 3238 1366 3290
rect 1418 3238 1430 3290
rect 1482 3238 1494 3290
rect 1546 3238 1558 3290
rect 1610 3238 1622 3290
rect 1674 3238 1686 3290
rect 1738 3238 7366 3290
rect 7418 3238 7430 3290
rect 7482 3238 7494 3290
rect 7546 3238 7558 3290
rect 7610 3238 7622 3290
rect 7674 3238 7686 3290
rect 7738 3238 13366 3290
rect 13418 3238 13430 3290
rect 13482 3238 13494 3290
rect 13546 3238 13558 3290
rect 13610 3238 13622 3290
rect 13674 3238 13686 3290
rect 13738 3238 17664 3290
rect 552 3216 17664 3238
rect 2130 3136 2136 3188
rect 2188 3136 2194 3188
rect 2314 3136 2320 3188
rect 2372 3136 2378 3188
rect 2406 3136 2412 3188
rect 2464 3136 2470 3188
rect 4798 3136 4804 3188
rect 4856 3136 4862 3188
rect 6822 3176 6828 3188
rect 5276 3148 5856 3176
rect 2148 3108 2176 3136
rect 1780 3080 2176 3108
rect 1780 3049 1808 3080
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3009 1823 3043
rect 2332 3040 2360 3136
rect 1765 3003 1823 3009
rect 2148 3012 2360 3040
rect 2148 2981 2176 3012
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2941 2191 2975
rect 2133 2935 2191 2941
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2972 2375 2975
rect 2424 2972 2452 3136
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3712 3012 3985 3040
rect 3712 2981 3740 3012
rect 3973 3009 3985 3012
rect 4019 3040 4031 3043
rect 4246 3040 4252 3052
rect 4019 3012 4252 3040
rect 4019 3009 4031 3012
rect 3973 3003 4031 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4816 3040 4844 3136
rect 4632 3012 4844 3040
rect 2363 2944 2452 2972
rect 3697 2975 3755 2981
rect 2363 2941 2375 2944
rect 2317 2935 2375 2941
rect 3697 2941 3709 2975
rect 3743 2941 3755 2975
rect 3697 2935 3755 2941
rect 3881 2975 3939 2981
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 3927 2944 4169 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4157 2941 4169 2944
rect 4203 2972 4215 2975
rect 4430 2972 4436 2984
rect 4203 2944 4436 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 1688 2904 1716 2935
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 4632 2981 4660 3012
rect 5276 2984 5304 3148
rect 5718 3068 5724 3120
rect 5776 3068 5782 3120
rect 5736 3040 5764 3068
rect 5460 3012 5764 3040
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2941 4675 2975
rect 4617 2935 4675 2941
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 2774 2904 2780 2916
rect 1688 2876 2780 2904
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 4724 2904 4752 2935
rect 5258 2932 5264 2984
rect 5316 2932 5322 2984
rect 5460 2981 5488 3012
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 5718 2932 5724 2984
rect 5776 2932 5782 2984
rect 5828 2981 5856 3148
rect 6472 3148 6828 3176
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2941 5871 2975
rect 5813 2935 5871 2941
rect 5902 2932 5908 2984
rect 5960 2932 5966 2984
rect 5994 2932 6000 2984
rect 6052 2981 6058 2984
rect 6052 2975 6081 2981
rect 6069 2941 6081 2975
rect 6052 2935 6081 2941
rect 6181 2975 6239 2981
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 6270 2972 6276 2984
rect 6227 2944 6276 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 6052 2932 6058 2935
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 6362 2932 6368 2984
rect 6420 2932 6426 2984
rect 6472 2981 6500 3148
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 7282 3176 7288 3188
rect 7239 3148 7288 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 7834 3136 7840 3188
rect 7892 3136 7898 3188
rect 9030 3136 9036 3188
rect 9088 3136 9094 3188
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 9272 3148 9904 3176
rect 9272 3136 9278 3148
rect 6546 3068 6552 3120
rect 6604 3108 6610 3120
rect 6604 3080 6684 3108
rect 6604 3068 6610 3080
rect 6656 3049 6684 3080
rect 6649 3043 6707 3049
rect 6649 3009 6661 3043
rect 6695 3009 6707 3043
rect 7024 3040 7052 3136
rect 7300 3040 7328 3136
rect 7653 3043 7711 3049
rect 7024 3012 7236 3040
rect 7300 3012 7604 3040
rect 6649 3003 6707 3009
rect 6457 2975 6515 2981
rect 6457 2941 6469 2975
rect 6503 2941 6515 2975
rect 6457 2935 6515 2941
rect 6549 2975 6607 2981
rect 6549 2941 6561 2975
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7098 2972 7104 2984
rect 7055 2944 7104 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 4120 2876 4752 2904
rect 5353 2907 5411 2913
rect 4120 2864 4126 2876
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 5399 2876 6408 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 2038 2796 2044 2848
rect 2096 2796 2102 2848
rect 3786 2796 3792 2848
rect 3844 2796 3850 2848
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4341 2839 4399 2845
rect 4341 2836 4353 2839
rect 4304 2808 4353 2836
rect 4304 2796 4310 2808
rect 4341 2805 4353 2808
rect 4387 2805 4399 2839
rect 4341 2799 4399 2805
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2836 4491 2839
rect 4798 2836 4804 2848
rect 4479 2808 4804 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 6178 2836 6184 2848
rect 5583 2808 6184 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 6178 2796 6184 2808
rect 6236 2796 6242 2848
rect 6380 2836 6408 2876
rect 6564 2836 6592 2935
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 6380 2808 6592 2836
rect 6825 2839 6883 2845
rect 6825 2805 6837 2839
rect 6871 2836 6883 2839
rect 7006 2836 7012 2848
rect 6871 2808 7012 2836
rect 6871 2805 6883 2808
rect 6825 2799 6883 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7208 2836 7236 3012
rect 7282 2932 7288 2984
rect 7340 2972 7346 2984
rect 7576 2972 7604 3012
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7852 3040 7880 3136
rect 7699 3012 7880 3040
rect 7929 3043 7987 3049
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 9048 3040 9076 3136
rect 7975 3012 8064 3040
rect 9048 3012 9720 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8036 2984 8064 3012
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 7340 2944 7512 2972
rect 7576 2944 7757 2972
rect 7340 2932 7346 2944
rect 7484 2904 7512 2944
rect 7745 2941 7757 2944
rect 7791 2941 7803 2975
rect 7745 2935 7803 2941
rect 7834 2932 7840 2984
rect 7892 2932 7898 2984
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 9692 2981 9720 3012
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 9876 3049 9904 3148
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 11790 3176 11796 3188
rect 10100 3148 11796 3176
rect 10100 3136 10106 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 14550 3176 14556 3188
rect 12078 3148 14556 3176
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 12078 3040 12106 3148
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 16114 3136 16120 3188
rect 16172 3136 16178 3188
rect 16206 3136 16212 3188
rect 16264 3176 16270 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 16264 3148 16865 3176
rect 16264 3136 16270 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 13722 3108 13728 3120
rect 12952 3080 13728 3108
rect 12952 3068 12958 3080
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 13906 3068 13912 3120
rect 13964 3068 13970 3120
rect 15010 3108 15016 3120
rect 14292 3080 15016 3108
rect 12526 3040 12532 3052
rect 9861 3003 9919 3009
rect 11992 3012 12106 3040
rect 12268 3012 12532 3040
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 8076 2944 9597 2972
rect 8076 2932 8082 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2941 9735 2975
rect 9677 2935 9735 2941
rect 11054 2932 11060 2984
rect 11112 2932 11118 2984
rect 11790 2932 11796 2984
rect 11848 2932 11854 2984
rect 11992 2981 12020 3012
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12066 2932 12072 2984
rect 12124 2932 12130 2984
rect 12268 2981 12296 3012
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 13541 3043 13599 3049
rect 13541 3040 13553 3043
rect 13044 3012 13553 3040
rect 13044 3000 13050 3012
rect 13541 3009 13553 3012
rect 13587 3009 13599 3043
rect 13541 3003 13599 3009
rect 13814 3000 13820 3052
rect 13872 3000 13878 3052
rect 13924 3040 13952 3068
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13924 3012 14013 3040
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14292 3040 14320 3080
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 14001 3003 14059 3009
rect 14108 3012 14320 3040
rect 14384 3012 15577 3040
rect 12253 2975 12311 2981
rect 12253 2941 12265 2975
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2941 12403 2975
rect 12345 2935 12403 2941
rect 13173 2975 13231 2981
rect 13173 2941 13185 2975
rect 13219 2941 13231 2975
rect 13173 2935 13231 2941
rect 11072 2904 11100 2932
rect 12360 2904 12388 2935
rect 13188 2904 13216 2935
rect 13354 2932 13360 2984
rect 13412 2972 13418 2984
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13412 2944 13737 2972
rect 13412 2932 13418 2944
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 13725 2935 13783 2941
rect 13909 2975 13967 2981
rect 13909 2941 13921 2975
rect 13955 2972 13967 2975
rect 14108 2972 14136 3012
rect 14384 2972 14412 3012
rect 15565 3009 15577 3012
rect 15611 3040 15623 3043
rect 16132 3040 16160 3136
rect 15611 3012 16160 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 16850 3000 16856 3052
rect 16908 3000 16914 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17696 3040 17724 3352
rect 17083 3012 17724 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 14734 2972 14740 2984
rect 13955 2944 14136 2972
rect 14200 2944 14412 2972
rect 14476 2944 14740 2972
rect 13955 2941 13967 2944
rect 13909 2935 13967 2941
rect 14200 2904 14228 2944
rect 7484 2876 9674 2904
rect 11072 2876 12388 2904
rect 13096 2876 14228 2904
rect 14369 2907 14427 2913
rect 7469 2839 7527 2845
rect 7469 2836 7481 2839
rect 7208 2808 7481 2836
rect 7469 2805 7481 2808
rect 7515 2836 7527 2839
rect 8018 2836 8024 2848
rect 7515 2808 8024 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8110 2796 8116 2848
rect 8168 2796 8174 2848
rect 9398 2796 9404 2848
rect 9456 2796 9462 2848
rect 9646 2836 9674 2876
rect 13096 2836 13124 2876
rect 14369 2873 14381 2907
rect 14415 2904 14427 2907
rect 14476 2904 14504 2944
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 15286 2932 15292 2984
rect 15344 2932 15350 2984
rect 16114 2932 16120 2984
rect 16172 2972 16178 2984
rect 16393 2975 16451 2981
rect 16393 2972 16405 2975
rect 16172 2944 16405 2972
rect 16172 2932 16178 2944
rect 16393 2941 16405 2944
rect 16439 2941 16451 2975
rect 16393 2935 16451 2941
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2972 16819 2975
rect 16868 2972 16896 3000
rect 16807 2944 16896 2972
rect 16807 2941 16819 2944
rect 16761 2935 16819 2941
rect 17126 2932 17132 2984
rect 17184 2932 17190 2984
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 14415 2876 14504 2904
rect 14553 2907 14611 2913
rect 14415 2873 14427 2876
rect 14369 2867 14427 2873
rect 14553 2873 14565 2907
rect 14599 2873 14611 2907
rect 15304 2904 15332 2932
rect 16942 2904 16948 2916
rect 15304 2876 16948 2904
rect 14553 2867 14611 2873
rect 9646 2808 13124 2836
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 13354 2836 13360 2848
rect 13228 2808 13360 2836
rect 13228 2796 13234 2808
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 14182 2796 14188 2848
rect 14240 2796 14246 2848
rect 14274 2796 14280 2848
rect 14332 2836 14338 2848
rect 14568 2836 14596 2867
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 17037 2907 17095 2913
rect 17037 2873 17049 2907
rect 17083 2904 17095 2907
rect 17218 2904 17224 2916
rect 17083 2876 17224 2904
rect 17083 2873 17095 2876
rect 17037 2867 17095 2873
rect 17218 2864 17224 2876
rect 17276 2904 17282 2916
rect 17328 2904 17356 2935
rect 17276 2876 17356 2904
rect 17276 2864 17282 2876
rect 14918 2836 14924 2848
rect 14332 2808 14924 2836
rect 14332 2796 14338 2808
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 15562 2836 15568 2848
rect 15160 2808 15568 2836
rect 15160 2796 15166 2808
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 16577 2839 16635 2845
rect 16577 2805 16589 2839
rect 16623 2836 16635 2839
rect 16758 2836 16764 2848
rect 16623 2808 16764 2836
rect 16623 2805 16635 2808
rect 16577 2799 16635 2805
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 17310 2796 17316 2848
rect 17368 2796 17374 2848
rect 552 2746 17664 2768
rect 552 2694 4366 2746
rect 4418 2694 4430 2746
rect 4482 2694 4494 2746
rect 4546 2694 4558 2746
rect 4610 2694 4622 2746
rect 4674 2694 4686 2746
rect 4738 2694 10366 2746
rect 10418 2694 10430 2746
rect 10482 2694 10494 2746
rect 10546 2694 10558 2746
rect 10610 2694 10622 2746
rect 10674 2694 10686 2746
rect 10738 2694 16366 2746
rect 16418 2694 16430 2746
rect 16482 2694 16494 2746
rect 16546 2694 16558 2746
rect 16610 2694 16622 2746
rect 16674 2694 16686 2746
rect 16738 2694 17664 2746
rect 552 2672 17664 2694
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 3418 2632 3424 2644
rect 3283 2604 3424 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 3418 2592 3424 2604
rect 3476 2632 3482 2644
rect 4430 2632 4436 2644
rect 3476 2604 4436 2632
rect 3476 2592 3482 2604
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5810 2592 5816 2644
rect 5868 2592 5874 2644
rect 8662 2632 8668 2644
rect 6012 2604 8668 2632
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 3602 2564 3608 2576
rect 3191 2536 3608 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 3602 2524 3608 2536
rect 3660 2524 3666 2576
rect 6012 2508 6040 2604
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 11238 2632 11244 2644
rect 11195 2604 11244 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 14792 2604 16160 2632
rect 14792 2592 14798 2604
rect 7098 2524 7104 2576
rect 7156 2564 7162 2576
rect 7469 2567 7527 2573
rect 7469 2564 7481 2567
rect 7156 2536 7481 2564
rect 7156 2524 7162 2536
rect 7469 2533 7481 2536
rect 7515 2533 7527 2567
rect 7469 2527 7527 2533
rect 7650 2524 7656 2576
rect 7708 2564 7714 2576
rect 8202 2564 8208 2576
rect 7708 2536 8208 2564
rect 7708 2524 7714 2536
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 8294 2524 8300 2576
rect 8352 2524 8358 2576
rect 11057 2567 11115 2573
rect 11057 2564 11069 2567
rect 9140 2536 11069 2564
rect 1029 2499 1087 2505
rect 1029 2465 1041 2499
rect 1075 2496 1087 2499
rect 1762 2496 1768 2508
rect 1075 2468 1768 2496
rect 1075 2465 1087 2468
rect 1029 2459 1087 2465
rect 1762 2456 1768 2468
rect 1820 2456 1826 2508
rect 2958 2456 2964 2508
rect 3016 2496 3022 2508
rect 3053 2499 3111 2505
rect 3053 2496 3065 2499
rect 3016 2468 3065 2496
rect 3016 2456 3022 2468
rect 3053 2465 3065 2468
rect 3099 2465 3111 2499
rect 3053 2459 3111 2465
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 3694 2496 3700 2508
rect 3467 2468 3700 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3694 2456 3700 2468
rect 3752 2456 3758 2508
rect 3786 2456 3792 2508
rect 3844 2496 3850 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3844 2468 4077 2496
rect 3844 2456 3850 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4246 2456 4252 2508
rect 4304 2456 4310 2508
rect 5994 2456 6000 2508
rect 6052 2456 6058 2508
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 7282 2496 7288 2508
rect 6595 2468 7288 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 1121 2431 1179 2437
rect 1121 2397 1133 2431
rect 1167 2428 1179 2431
rect 3510 2428 3516 2440
rect 1167 2400 3516 2428
rect 1167 2397 1179 2400
rect 1121 2391 1179 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 6273 2431 6331 2437
rect 6273 2397 6285 2431
rect 6319 2428 6331 2431
rect 6822 2428 6828 2440
rect 6319 2400 6828 2428
rect 6319 2397 6331 2400
rect 6273 2391 6331 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 8312 2428 8340 2524
rect 9030 2456 9036 2508
rect 9088 2456 9094 2508
rect 9140 2505 9168 2536
rect 11057 2533 11069 2536
rect 11103 2564 11115 2567
rect 11103 2536 11376 2564
rect 11103 2533 11115 2536
rect 11057 2527 11115 2533
rect 9125 2499 9183 2505
rect 9125 2465 9137 2499
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 9306 2456 9312 2508
rect 9364 2456 9370 2508
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2496 9459 2499
rect 9447 2468 9674 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 9646 2428 9674 2468
rect 10594 2456 10600 2508
rect 10652 2496 10658 2508
rect 11238 2496 11244 2508
rect 10652 2468 11244 2496
rect 10652 2456 10658 2468
rect 11238 2456 11244 2468
rect 11296 2456 11302 2508
rect 11348 2505 11376 2536
rect 12342 2524 12348 2576
rect 12400 2564 12406 2576
rect 12710 2564 12716 2576
rect 12400 2536 12480 2564
rect 12400 2524 12406 2536
rect 12452 2505 12480 2536
rect 12636 2536 12716 2564
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 12428 2499 12486 2505
rect 12428 2465 12440 2499
rect 12474 2465 12486 2499
rect 12428 2459 12486 2465
rect 11054 2428 11060 2440
rect 6932 2400 8248 2428
rect 8312 2400 9076 2428
rect 9646 2400 11060 2428
rect 1397 2363 1455 2369
rect 1397 2329 1409 2363
rect 1443 2360 1455 2363
rect 1762 2360 1768 2372
rect 1443 2332 1768 2360
rect 1443 2329 1455 2332
rect 1397 2323 1455 2329
rect 1762 2320 1768 2332
rect 1820 2320 1826 2372
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 4338 2360 4344 2372
rect 3292 2332 4344 2360
rect 3292 2320 3298 2332
rect 4338 2320 4344 2332
rect 4396 2360 4402 2372
rect 5718 2360 5724 2372
rect 4396 2332 5724 2360
rect 4396 2320 4402 2332
rect 5718 2320 5724 2332
rect 5776 2360 5782 2372
rect 6365 2363 6423 2369
rect 6365 2360 6377 2363
rect 5776 2332 6377 2360
rect 5776 2320 5782 2332
rect 6365 2329 6377 2332
rect 6411 2329 6423 2363
rect 6365 2323 6423 2329
rect 3326 2252 3332 2304
rect 3384 2252 3390 2304
rect 4062 2252 4068 2304
rect 4120 2252 4126 2304
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 6932 2292 6960 2400
rect 7006 2320 7012 2372
rect 7064 2360 7070 2372
rect 8018 2360 8024 2372
rect 7064 2332 8024 2360
rect 7064 2320 7070 2332
rect 8018 2320 8024 2332
rect 8076 2320 8082 2372
rect 8220 2360 8248 2400
rect 9048 2372 9076 2400
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 8220 2332 8984 2360
rect 5592 2264 6960 2292
rect 5592 2252 5598 2264
rect 7282 2252 7288 2304
rect 7340 2252 7346 2304
rect 8846 2252 8852 2304
rect 8904 2252 8910 2304
rect 8956 2292 8984 2332
rect 9030 2320 9036 2372
rect 9088 2320 9094 2372
rect 10594 2360 10600 2372
rect 9646 2332 10600 2360
rect 9646 2292 9674 2332
rect 10594 2320 10600 2332
rect 10652 2320 10658 2372
rect 11348 2360 11376 2459
rect 12526 2456 12532 2508
rect 12584 2456 12590 2508
rect 12636 2428 12664 2536
rect 12710 2524 12716 2536
rect 12768 2564 12774 2576
rect 13998 2564 14004 2576
rect 12768 2536 14004 2564
rect 12768 2524 12774 2536
rect 13998 2524 14004 2536
rect 14056 2564 14062 2576
rect 15010 2564 15016 2576
rect 14056 2536 14412 2564
rect 14056 2524 14062 2536
rect 12805 2499 12863 2505
rect 12805 2494 12817 2499
rect 12360 2400 12664 2428
rect 12728 2466 12817 2494
rect 12066 2360 12072 2372
rect 11348 2332 12072 2360
rect 12066 2320 12072 2332
rect 12124 2360 12130 2372
rect 12253 2363 12311 2369
rect 12253 2360 12265 2363
rect 12124 2332 12265 2360
rect 12124 2320 12130 2332
rect 12253 2329 12265 2332
rect 12299 2329 12311 2363
rect 12253 2323 12311 2329
rect 8956 2264 9674 2292
rect 9766 2252 9772 2304
rect 9824 2292 9830 2304
rect 11517 2295 11575 2301
rect 11517 2292 11529 2295
rect 9824 2264 11529 2292
rect 9824 2252 9830 2264
rect 11517 2261 11529 2264
rect 11563 2292 11575 2295
rect 12360 2292 12388 2400
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12728 2360 12756 2466
rect 12805 2465 12817 2466
rect 12851 2465 12863 2499
rect 12805 2459 12863 2465
rect 14274 2456 14280 2508
rect 14332 2456 14338 2508
rect 14384 2496 14412 2536
rect 14752 2536 15016 2564
rect 14452 2499 14510 2505
rect 14452 2496 14464 2499
rect 14384 2468 14464 2496
rect 14452 2465 14464 2468
rect 14498 2465 14510 2499
rect 14452 2459 14510 2465
rect 14550 2456 14556 2508
rect 14608 2456 14614 2508
rect 14752 2505 14780 2536
rect 15010 2524 15016 2536
rect 15068 2524 15074 2576
rect 15194 2524 15200 2576
rect 15252 2564 15258 2576
rect 16132 2573 16160 2604
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 16317 2635 16375 2641
rect 16317 2632 16329 2635
rect 16264 2604 16329 2632
rect 16264 2592 16270 2604
rect 16317 2601 16329 2604
rect 16363 2601 16375 2635
rect 17126 2632 17132 2644
rect 16317 2595 16375 2601
rect 16408 2604 17132 2632
rect 16117 2567 16175 2573
rect 15252 2536 15700 2564
rect 15252 2524 15258 2536
rect 14737 2499 14795 2505
rect 14737 2465 14749 2499
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 14918 2456 14924 2508
rect 14976 2456 14982 2508
rect 15105 2499 15163 2505
rect 15105 2465 15117 2499
rect 15151 2465 15163 2499
rect 15105 2459 15163 2465
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14415 2400 14841 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 12492 2332 12756 2360
rect 12492 2320 12498 2332
rect 12802 2320 12808 2372
rect 12860 2360 12866 2372
rect 12989 2363 13047 2369
rect 12989 2360 13001 2363
rect 12860 2332 13001 2360
rect 12860 2320 12866 2332
rect 12989 2329 13001 2332
rect 13035 2329 13047 2363
rect 15120 2360 15148 2459
rect 15304 2428 15332 2459
rect 15378 2456 15384 2508
rect 15436 2456 15442 2508
rect 15562 2456 15568 2508
rect 15620 2456 15626 2508
rect 15672 2505 15700 2536
rect 16117 2533 16129 2567
rect 16163 2564 16175 2567
rect 16408 2564 16436 2604
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 16163 2536 16436 2564
rect 17037 2567 17095 2573
rect 16163 2533 16175 2536
rect 16117 2527 16175 2533
rect 17037 2533 17049 2567
rect 17083 2564 17095 2567
rect 17494 2564 17500 2576
rect 17083 2536 17500 2564
rect 17083 2533 17095 2536
rect 17037 2527 17095 2533
rect 17328 2505 17356 2536
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 17586 2524 17592 2576
rect 17644 2524 17650 2576
rect 15657 2499 15715 2505
rect 15657 2465 15669 2499
rect 15703 2465 15715 2499
rect 15657 2459 15715 2465
rect 16853 2499 16911 2505
rect 16853 2465 16865 2499
rect 16899 2496 16911 2499
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16899 2468 17141 2496
rect 16899 2465 16911 2468
rect 16853 2459 16911 2465
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 17313 2499 17371 2505
rect 17313 2465 17325 2499
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 15473 2431 15531 2437
rect 15473 2428 15485 2431
rect 15304 2400 15485 2428
rect 15473 2397 15485 2400
rect 15519 2397 15531 2431
rect 17144 2428 17172 2459
rect 17604 2428 17632 2524
rect 17144 2400 17632 2428
rect 15473 2391 15531 2397
rect 15120 2332 15424 2360
rect 12989 2323 13047 2329
rect 11563 2264 12388 2292
rect 12713 2295 12771 2301
rect 11563 2261 11575 2264
rect 11517 2255 11575 2261
rect 12713 2261 12725 2295
rect 12759 2292 12771 2295
rect 13998 2292 14004 2304
rect 12759 2264 14004 2292
rect 12759 2261 12771 2264
rect 12713 2255 12771 2261
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 14093 2295 14151 2301
rect 14093 2261 14105 2295
rect 14139 2292 14151 2295
rect 14274 2292 14280 2304
rect 14139 2264 14280 2292
rect 14139 2261 14151 2264
rect 14093 2255 14151 2261
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 14550 2252 14556 2304
rect 14608 2292 14614 2304
rect 14734 2292 14740 2304
rect 14608 2264 14740 2292
rect 14608 2252 14614 2264
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 15286 2252 15292 2304
rect 15344 2252 15350 2304
rect 15396 2292 15424 2332
rect 15562 2320 15568 2372
rect 15620 2360 15626 2372
rect 17494 2360 17500 2372
rect 15620 2332 17500 2360
rect 15620 2320 15626 2332
rect 17494 2320 17500 2332
rect 17552 2320 17558 2372
rect 15470 2292 15476 2304
rect 15396 2264 15476 2292
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 15838 2252 15844 2304
rect 15896 2252 15902 2304
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 16301 2295 16359 2301
rect 16301 2292 16313 2295
rect 16080 2264 16313 2292
rect 16080 2252 16086 2264
rect 16301 2261 16313 2264
rect 16347 2292 16359 2295
rect 16390 2292 16396 2304
rect 16347 2264 16396 2292
rect 16347 2261 16359 2264
rect 16301 2255 16359 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 16482 2252 16488 2304
rect 16540 2252 16546 2304
rect 16669 2295 16727 2301
rect 16669 2261 16681 2295
rect 16715 2292 16727 2295
rect 16850 2292 16856 2304
rect 16715 2264 16856 2292
rect 16715 2261 16727 2264
rect 16669 2255 16727 2261
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 552 2202 17664 2224
rect 552 2150 1366 2202
rect 1418 2150 1430 2202
rect 1482 2150 1494 2202
rect 1546 2150 1558 2202
rect 1610 2150 1622 2202
rect 1674 2150 1686 2202
rect 1738 2150 7366 2202
rect 7418 2150 7430 2202
rect 7482 2150 7494 2202
rect 7546 2150 7558 2202
rect 7610 2150 7622 2202
rect 7674 2150 7686 2202
rect 7738 2150 13366 2202
rect 13418 2150 13430 2202
rect 13482 2150 13494 2202
rect 13546 2150 13558 2202
rect 13610 2150 13622 2202
rect 13674 2150 13686 2202
rect 13738 2150 17664 2202
rect 552 2128 17664 2150
rect 1762 2048 1768 2100
rect 1820 2048 1826 2100
rect 3326 2048 3332 2100
rect 3384 2088 3390 2100
rect 3421 2091 3479 2097
rect 3421 2088 3433 2091
rect 3384 2060 3433 2088
rect 3384 2048 3390 2060
rect 3421 2057 3433 2060
rect 3467 2057 3479 2091
rect 3421 2051 3479 2057
rect 3528 2060 4660 2088
rect 1489 1955 1547 1961
rect 1489 1921 1501 1955
rect 1535 1952 1547 1955
rect 1780 1952 1808 2048
rect 3528 2032 3556 2060
rect 2038 1980 2044 2032
rect 2096 1980 2102 2032
rect 3510 1980 3516 2032
rect 3568 1980 3574 2032
rect 3605 2023 3663 2029
rect 3605 1989 3617 2023
rect 3651 2020 3663 2023
rect 4522 2020 4528 2032
rect 3651 1992 4528 2020
rect 3651 1989 3663 1992
rect 3605 1983 3663 1989
rect 4522 1980 4528 1992
rect 4580 1980 4586 2032
rect 1535 1924 1808 1952
rect 1535 1921 1547 1924
rect 1489 1915 1547 1921
rect 1397 1887 1455 1893
rect 1397 1853 1409 1887
rect 1443 1884 1455 1887
rect 1854 1884 1860 1896
rect 1443 1856 1860 1884
rect 1443 1853 1455 1856
rect 1397 1847 1455 1853
rect 1854 1844 1860 1856
rect 1912 1844 1918 1896
rect 1946 1844 1952 1896
rect 2004 1844 2010 1896
rect 2056 1884 2084 1980
rect 4246 1952 4252 1964
rect 2332 1924 3480 1952
rect 2332 1896 2360 1924
rect 2133 1887 2191 1893
rect 2133 1884 2145 1887
rect 2056 1856 2145 1884
rect 2133 1853 2145 1856
rect 2179 1853 2191 1887
rect 2133 1847 2191 1853
rect 2225 1887 2283 1893
rect 2225 1853 2237 1887
rect 2271 1884 2283 1887
rect 2314 1884 2320 1896
rect 2271 1856 2320 1884
rect 2271 1853 2283 1856
rect 2225 1847 2283 1853
rect 2314 1844 2320 1856
rect 2372 1844 2378 1896
rect 2501 1887 2559 1893
rect 2501 1853 2513 1887
rect 2547 1853 2559 1887
rect 2501 1847 2559 1853
rect 2516 1816 2544 1847
rect 2682 1844 2688 1896
rect 2740 1884 2746 1896
rect 2777 1887 2835 1893
rect 2777 1884 2789 1887
rect 2740 1856 2789 1884
rect 2740 1844 2746 1856
rect 2777 1853 2789 1856
rect 2823 1853 2835 1887
rect 2777 1847 2835 1853
rect 2961 1887 3019 1893
rect 2961 1853 2973 1887
rect 3007 1853 3019 1887
rect 2961 1847 3019 1853
rect 3452 1884 3480 1924
rect 3712 1924 4252 1952
rect 3510 1884 3516 1896
rect 3452 1853 3516 1884
rect 2976 1816 3004 1847
rect 1780 1788 2544 1816
rect 2608 1788 3004 1816
rect 1780 1757 1808 1788
rect 1765 1751 1823 1757
rect 1765 1717 1777 1751
rect 1811 1748 1823 1751
rect 1854 1748 1860 1760
rect 1811 1720 1860 1748
rect 1811 1717 1823 1720
rect 1765 1711 1823 1717
rect 1854 1708 1860 1720
rect 1912 1708 1918 1760
rect 2133 1751 2191 1757
rect 2133 1717 2145 1751
rect 2179 1748 2191 1751
rect 2317 1751 2375 1757
rect 2317 1748 2329 1751
rect 2179 1720 2329 1748
rect 2179 1717 2191 1720
rect 2133 1711 2191 1717
rect 2317 1717 2329 1720
rect 2363 1748 2375 1751
rect 2406 1748 2412 1760
rect 2363 1720 2412 1748
rect 2363 1717 2375 1720
rect 2317 1711 2375 1717
rect 2406 1708 2412 1720
rect 2464 1748 2470 1760
rect 2608 1748 2636 1788
rect 3234 1776 3240 1828
rect 3292 1776 3298 1828
rect 3452 1822 3479 1853
rect 3467 1819 3479 1822
rect 3513 1844 3516 1853
rect 3568 1844 3574 1896
rect 3712 1893 3740 1924
rect 4246 1912 4252 1924
rect 4304 1912 4310 1964
rect 4338 1912 4344 1964
rect 4396 1912 4402 1964
rect 4430 1912 4436 1964
rect 4488 1912 4494 1964
rect 4632 1952 4660 2060
rect 6086 2048 6092 2100
rect 6144 2048 6150 2100
rect 10686 2088 10692 2100
rect 6288 2060 8708 2088
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 5261 2023 5319 2029
rect 5261 2020 5273 2023
rect 4764 1992 5273 2020
rect 4764 1980 4770 1992
rect 5261 1989 5273 1992
rect 5307 1989 5319 2023
rect 5261 1983 5319 1989
rect 5350 1980 5356 2032
rect 5408 1980 5414 2032
rect 5902 1952 5908 1964
rect 4632 1924 4752 1952
rect 3697 1887 3755 1893
rect 3697 1853 3709 1887
rect 3743 1853 3755 1887
rect 3697 1847 3755 1853
rect 3786 1844 3792 1896
rect 3844 1844 3850 1896
rect 3878 1844 3884 1896
rect 3936 1884 3942 1896
rect 3973 1887 4031 1893
rect 3973 1884 3985 1887
rect 3936 1856 3985 1884
rect 3936 1844 3942 1856
rect 3973 1853 3985 1856
rect 4019 1853 4031 1887
rect 3973 1847 4031 1853
rect 4062 1844 4068 1896
rect 4120 1844 4126 1896
rect 4448 1884 4476 1912
rect 4724 1893 4752 1924
rect 5184 1924 5908 1952
rect 4617 1887 4675 1893
rect 4617 1884 4629 1887
rect 4172 1856 4404 1884
rect 4448 1856 4629 1884
rect 3513 1819 3525 1844
rect 3467 1813 3525 1819
rect 2464 1720 2636 1748
rect 2685 1751 2743 1757
rect 2464 1708 2470 1720
rect 2685 1717 2697 1751
rect 2731 1748 2743 1751
rect 2774 1748 2780 1760
rect 2731 1720 2780 1748
rect 2731 1717 2743 1720
rect 2685 1711 2743 1717
rect 2774 1708 2780 1720
rect 2832 1708 2838 1760
rect 2958 1708 2964 1760
rect 3016 1708 3022 1760
rect 3326 1708 3332 1760
rect 3384 1748 3390 1760
rect 4172 1748 4200 1856
rect 4376 1816 4404 1856
rect 4617 1853 4629 1856
rect 4663 1853 4675 1887
rect 4617 1847 4675 1853
rect 4709 1887 4767 1893
rect 4709 1853 4721 1887
rect 4755 1853 4767 1887
rect 4709 1847 4767 1853
rect 4982 1844 4988 1896
rect 5040 1844 5046 1896
rect 5184 1893 5212 1924
rect 5902 1912 5908 1924
rect 5960 1952 5966 1964
rect 6288 1952 6316 2060
rect 8680 2032 8708 2060
rect 9600 2060 10692 2088
rect 6454 1980 6460 2032
rect 6512 1980 6518 2032
rect 7558 2020 7564 2032
rect 6564 1992 7564 2020
rect 5960 1924 6316 1952
rect 5960 1912 5966 1924
rect 5169 1887 5227 1893
rect 5169 1853 5181 1887
rect 5215 1853 5227 1887
rect 5169 1847 5227 1853
rect 5445 1887 5503 1893
rect 5445 1853 5457 1887
rect 5491 1884 5503 1887
rect 5994 1884 6000 1896
rect 5491 1856 6000 1884
rect 5491 1853 5503 1856
rect 5445 1847 5503 1853
rect 5994 1844 6000 1856
rect 6052 1844 6058 1896
rect 6288 1893 6316 1924
rect 6564 1893 6592 1992
rect 7558 1980 7564 1992
rect 7616 2020 7622 2032
rect 8294 2020 8300 2032
rect 7616 1992 8300 2020
rect 7616 1980 7622 1992
rect 8294 1980 8300 1992
rect 8352 1980 8358 2032
rect 8662 1980 8668 2032
rect 8720 1980 8726 2032
rect 9122 1980 9128 2032
rect 9180 1980 9186 2032
rect 6730 1912 6736 1964
rect 6788 1952 6794 1964
rect 6917 1955 6975 1961
rect 6917 1952 6929 1955
rect 6788 1924 6929 1952
rect 6788 1912 6794 1924
rect 6917 1921 6929 1924
rect 6963 1921 6975 1955
rect 6917 1915 6975 1921
rect 7101 1955 7159 1961
rect 7101 1921 7113 1955
rect 7147 1952 7159 1955
rect 7282 1952 7288 1964
rect 7147 1924 7288 1952
rect 7147 1921 7159 1924
rect 7101 1915 7159 1921
rect 7282 1912 7288 1924
rect 7340 1912 7346 1964
rect 7377 1955 7435 1961
rect 7377 1921 7389 1955
rect 7423 1952 7435 1955
rect 8202 1952 8208 1964
rect 7423 1924 8208 1952
rect 7423 1921 7435 1924
rect 7377 1915 7435 1921
rect 8202 1912 8208 1924
rect 8260 1912 8266 1964
rect 8938 1912 8944 1964
rect 8996 1952 9002 1964
rect 9600 1961 9628 2060
rect 10686 2048 10692 2060
rect 10744 2088 10750 2100
rect 10781 2091 10839 2097
rect 10781 2088 10793 2091
rect 10744 2060 10793 2088
rect 10744 2048 10750 2060
rect 10781 2057 10793 2060
rect 10827 2088 10839 2091
rect 12066 2088 12072 2100
rect 10827 2060 12072 2088
rect 10827 2057 10839 2060
rect 10781 2051 10839 2057
rect 12066 2048 12072 2060
rect 12124 2048 12130 2100
rect 14182 2048 14188 2100
rect 14240 2088 14246 2100
rect 14826 2088 14832 2100
rect 14240 2060 14832 2088
rect 14240 2048 14246 2060
rect 14826 2048 14832 2060
rect 14884 2048 14890 2100
rect 15470 2048 15476 2100
rect 15528 2088 15534 2100
rect 15528 2060 16344 2088
rect 15528 2048 15534 2060
rect 10505 2023 10563 2029
rect 10505 2020 10517 2023
rect 9876 1992 10517 2020
rect 9585 1955 9643 1961
rect 8996 1924 9352 1952
rect 8996 1912 9002 1924
rect 6273 1887 6331 1893
rect 6273 1853 6285 1887
rect 6319 1853 6331 1887
rect 6273 1847 6331 1853
rect 6365 1887 6423 1893
rect 6365 1853 6377 1887
rect 6411 1853 6423 1887
rect 6365 1847 6423 1853
rect 6549 1887 6607 1893
rect 6549 1853 6561 1887
rect 6595 1853 6607 1887
rect 6549 1847 6607 1853
rect 6825 1887 6883 1893
rect 6825 1853 6837 1887
rect 6871 1853 6883 1887
rect 6825 1847 6883 1853
rect 6380 1816 6408 1847
rect 4376 1788 6408 1816
rect 6840 1816 6868 1847
rect 7006 1844 7012 1896
rect 7064 1844 7070 1896
rect 7650 1844 7656 1896
rect 7708 1884 7714 1896
rect 7834 1884 7840 1896
rect 7708 1856 7840 1884
rect 7708 1844 7714 1856
rect 7834 1844 7840 1856
rect 7892 1844 7898 1896
rect 8018 1844 8024 1896
rect 8076 1844 8082 1896
rect 8389 1887 8447 1893
rect 8389 1853 8401 1887
rect 8435 1884 8447 1887
rect 8665 1887 8723 1893
rect 8665 1884 8677 1887
rect 8435 1856 8677 1884
rect 8435 1853 8447 1856
rect 8389 1847 8447 1853
rect 8665 1853 8677 1856
rect 8711 1853 8723 1887
rect 8665 1847 8723 1853
rect 8846 1844 8852 1896
rect 8904 1844 8910 1896
rect 9030 1844 9036 1896
rect 9088 1844 9094 1896
rect 9324 1893 9352 1924
rect 9585 1921 9597 1955
rect 9631 1921 9643 1955
rect 9585 1915 9643 1921
rect 9876 1896 9904 1992
rect 10505 1989 10517 1992
rect 10551 1989 10563 2023
rect 11149 2023 11207 2029
rect 11149 2020 11161 2023
rect 10505 1983 10563 1989
rect 10704 1992 11161 2020
rect 9309 1887 9367 1893
rect 9309 1853 9321 1887
rect 9355 1853 9367 1887
rect 9309 1847 9367 1853
rect 9493 1887 9551 1893
rect 9493 1853 9505 1887
rect 9539 1853 9551 1887
rect 9493 1847 9551 1853
rect 7190 1816 7196 1828
rect 6840 1788 7196 1816
rect 7190 1776 7196 1788
rect 7248 1776 7254 1828
rect 8036 1816 8064 1844
rect 9508 1816 9536 1847
rect 9674 1844 9680 1896
rect 9732 1844 9738 1896
rect 9766 1844 9772 1896
rect 9824 1844 9830 1896
rect 9858 1844 9864 1896
rect 9916 1844 9922 1896
rect 10704 1893 10732 1992
rect 11149 1989 11161 1992
rect 11195 2020 11207 2023
rect 12434 2020 12440 2032
rect 11195 1992 12440 2020
rect 11195 1989 11207 1992
rect 11149 1983 11207 1989
rect 12434 1980 12440 1992
rect 12492 1980 12498 2032
rect 12529 2023 12587 2029
rect 12529 1989 12541 2023
rect 12575 2020 12587 2023
rect 13078 2020 13084 2032
rect 12575 1992 13084 2020
rect 12575 1989 12587 1992
rect 12529 1983 12587 1989
rect 13078 1980 13084 1992
rect 13136 1980 13142 2032
rect 14093 2023 14151 2029
rect 14093 2020 14105 2023
rect 13556 1992 14105 2020
rect 11054 1912 11060 1964
rect 11112 1912 11118 1964
rect 11974 1912 11980 1964
rect 12032 1912 12038 1964
rect 12253 1955 12311 1961
rect 12253 1921 12265 1955
rect 12299 1952 12311 1955
rect 12452 1952 12480 1980
rect 12299 1924 12480 1952
rect 12299 1921 12311 1924
rect 12253 1915 12311 1921
rect 12618 1912 12624 1964
rect 12676 1952 12682 1964
rect 13354 1952 13360 1964
rect 12676 1924 13032 1952
rect 12676 1912 12682 1924
rect 9953 1887 10011 1893
rect 9953 1853 9965 1887
rect 9999 1884 10011 1887
rect 10413 1887 10471 1893
rect 9999 1856 10364 1884
rect 9999 1853 10011 1856
rect 9953 1847 10011 1853
rect 10042 1816 10048 1828
rect 8036 1788 9536 1816
rect 9600 1788 10048 1816
rect 3384 1720 4200 1748
rect 4249 1751 4307 1757
rect 3384 1708 3390 1720
rect 4249 1717 4261 1751
rect 4295 1748 4307 1751
rect 4525 1751 4583 1757
rect 4525 1748 4537 1751
rect 4295 1720 4537 1748
rect 4295 1717 4307 1720
rect 4249 1711 4307 1717
rect 4525 1717 4537 1720
rect 4571 1717 4583 1751
rect 4525 1711 4583 1717
rect 4890 1708 4896 1760
rect 4948 1708 4954 1760
rect 7285 1751 7343 1757
rect 7285 1717 7297 1751
rect 7331 1748 7343 1751
rect 8478 1748 8484 1760
rect 7331 1720 8484 1748
rect 7331 1717 7343 1720
rect 7285 1711 7343 1717
rect 8478 1708 8484 1720
rect 8536 1708 8542 1760
rect 8570 1708 8576 1760
rect 8628 1708 8634 1760
rect 8662 1708 8668 1760
rect 8720 1748 8726 1760
rect 9600 1748 9628 1788
rect 10042 1776 10048 1788
rect 10100 1816 10106 1828
rect 10336 1816 10364 1856
rect 10413 1853 10425 1887
rect 10459 1884 10471 1887
rect 10689 1887 10747 1893
rect 10689 1884 10701 1887
rect 10459 1856 10701 1884
rect 10459 1853 10471 1856
rect 10413 1847 10471 1853
rect 10689 1853 10701 1856
rect 10735 1853 10747 1887
rect 10689 1847 10747 1853
rect 10965 1887 11023 1893
rect 10965 1853 10977 1887
rect 11011 1884 11023 1887
rect 11072 1884 11100 1912
rect 11333 1887 11391 1893
rect 11333 1884 11345 1887
rect 11011 1856 11345 1884
rect 11011 1853 11023 1856
rect 10965 1847 11023 1853
rect 11333 1853 11345 1856
rect 11379 1853 11391 1887
rect 11333 1847 11391 1853
rect 12342 1844 12348 1896
rect 12400 1844 12406 1896
rect 12434 1844 12440 1896
rect 12492 1884 12498 1896
rect 13004 1893 13032 1924
rect 13096 1924 13360 1952
rect 13096 1893 13124 1924
rect 13354 1912 13360 1924
rect 13412 1912 13418 1964
rect 12897 1887 12955 1893
rect 12897 1884 12909 1887
rect 12492 1856 12909 1884
rect 12492 1844 12498 1856
rect 12897 1853 12909 1856
rect 12943 1853 12955 1887
rect 12897 1847 12955 1853
rect 12989 1887 13047 1893
rect 12989 1853 13001 1887
rect 13035 1853 13047 1887
rect 12989 1847 13047 1853
rect 13081 1887 13139 1893
rect 13081 1853 13093 1887
rect 13127 1853 13139 1887
rect 13081 1847 13139 1853
rect 13265 1887 13323 1893
rect 13265 1853 13277 1887
rect 13311 1884 13323 1887
rect 13556 1884 13584 1992
rect 14093 1989 14105 1992
rect 14139 1989 14151 2023
rect 14093 1983 14151 1989
rect 14645 2023 14703 2029
rect 14645 1989 14657 2023
rect 14691 2020 14703 2023
rect 14691 1992 16160 2020
rect 14691 1989 14703 1992
rect 14645 1983 14703 1989
rect 13630 1912 13636 1964
rect 13688 1912 13694 1964
rect 13725 1955 13783 1961
rect 13725 1921 13737 1955
rect 13771 1921 13783 1955
rect 13725 1915 13783 1921
rect 13311 1856 13584 1884
rect 13311 1853 13323 1856
rect 13265 1847 13323 1853
rect 10870 1816 10876 1828
rect 10100 1788 10272 1816
rect 10336 1788 10876 1816
rect 10100 1776 10106 1788
rect 8720 1720 9628 1748
rect 8720 1708 8726 1720
rect 10134 1708 10140 1760
rect 10192 1708 10198 1760
rect 10244 1757 10272 1788
rect 10870 1776 10876 1788
rect 10928 1776 10934 1828
rect 12158 1776 12164 1828
rect 12216 1816 12222 1828
rect 12216 1788 12756 1816
rect 12216 1776 12222 1788
rect 10229 1751 10287 1757
rect 10229 1717 10241 1751
rect 10275 1717 10287 1751
rect 10229 1711 10287 1717
rect 10686 1708 10692 1760
rect 10744 1748 10750 1760
rect 10962 1748 10968 1760
rect 10744 1720 10968 1748
rect 10744 1708 10750 1720
rect 10962 1708 10968 1720
rect 11020 1708 11026 1760
rect 12618 1708 12624 1760
rect 12676 1708 12682 1760
rect 12728 1748 12756 1788
rect 13170 1776 13176 1828
rect 13228 1816 13234 1828
rect 13740 1816 13768 1915
rect 13906 1912 13912 1964
rect 13964 1912 13970 1964
rect 15102 1912 15108 1964
rect 15160 1912 15166 1964
rect 15654 1912 15660 1964
rect 15712 1912 15718 1964
rect 13814 1844 13820 1896
rect 13872 1844 13878 1896
rect 14369 1887 14427 1893
rect 14369 1853 14381 1887
rect 14415 1853 14427 1887
rect 14369 1847 14427 1853
rect 14461 1887 14519 1893
rect 14461 1853 14473 1887
rect 14507 1884 14519 1887
rect 14550 1884 14556 1896
rect 14507 1856 14556 1884
rect 14507 1853 14519 1856
rect 14461 1847 14519 1853
rect 13228 1788 13768 1816
rect 14384 1816 14412 1847
rect 14550 1844 14556 1856
rect 14608 1844 14614 1896
rect 14645 1887 14703 1893
rect 14645 1853 14657 1887
rect 14691 1884 14703 1887
rect 14918 1884 14924 1896
rect 14691 1856 14924 1884
rect 14691 1853 14703 1856
rect 14645 1847 14703 1853
rect 14918 1844 14924 1856
rect 14976 1844 14982 1896
rect 15010 1844 15016 1896
rect 15068 1844 15074 1896
rect 15289 1887 15347 1893
rect 15289 1853 15301 1887
rect 15335 1884 15347 1887
rect 15378 1884 15384 1896
rect 15335 1856 15384 1884
rect 15335 1853 15347 1856
rect 15289 1847 15347 1853
rect 15378 1844 15384 1856
rect 15436 1844 15442 1896
rect 15672 1884 15700 1912
rect 16132 1893 16160 1992
rect 16316 1893 16344 2060
rect 16482 2048 16488 2100
rect 16540 2048 16546 2100
rect 16945 2091 17003 2097
rect 16945 2057 16957 2091
rect 16991 2088 17003 2091
rect 17129 2091 17187 2097
rect 17129 2088 17141 2091
rect 16991 2060 17141 2088
rect 16991 2057 17003 2060
rect 16945 2051 17003 2057
rect 17129 2057 17141 2060
rect 17175 2057 17187 2091
rect 17129 2051 17187 2057
rect 15841 1887 15899 1893
rect 15841 1884 15853 1887
rect 15672 1856 15853 1884
rect 15841 1853 15853 1856
rect 15887 1853 15899 1887
rect 15841 1847 15899 1853
rect 16117 1887 16175 1893
rect 16117 1853 16129 1887
rect 16163 1853 16175 1887
rect 16117 1847 16175 1853
rect 16301 1887 16359 1893
rect 16301 1853 16313 1887
rect 16347 1853 16359 1887
rect 16500 1884 16528 2048
rect 16574 1980 16580 2032
rect 16632 1980 16638 2032
rect 16592 1952 16620 1980
rect 16592 1924 17264 1952
rect 16577 1887 16635 1893
rect 16577 1884 16589 1887
rect 16500 1856 16589 1884
rect 16301 1847 16359 1853
rect 16577 1853 16589 1856
rect 16623 1853 16635 1887
rect 16577 1847 16635 1853
rect 16669 1887 16727 1893
rect 16669 1853 16681 1887
rect 16715 1853 16727 1887
rect 16669 1847 16727 1853
rect 14384 1788 15792 1816
rect 13228 1776 13234 1788
rect 14277 1751 14335 1757
rect 14277 1748 14289 1751
rect 12728 1720 14289 1748
rect 14277 1717 14289 1720
rect 14323 1717 14335 1751
rect 14277 1711 14335 1717
rect 14829 1751 14887 1757
rect 14829 1717 14841 1751
rect 14875 1748 14887 1751
rect 15562 1748 15568 1760
rect 14875 1720 15568 1748
rect 14875 1717 14887 1720
rect 14829 1711 14887 1717
rect 15562 1708 15568 1720
rect 15620 1708 15626 1760
rect 15654 1708 15660 1760
rect 15712 1708 15718 1760
rect 15764 1748 15792 1788
rect 15930 1776 15936 1828
rect 15988 1776 15994 1828
rect 16022 1776 16028 1828
rect 16080 1776 16086 1828
rect 16132 1816 16160 1847
rect 16684 1816 16712 1847
rect 17034 1844 17040 1896
rect 17092 1844 17098 1896
rect 17129 1887 17187 1893
rect 17129 1853 17141 1887
rect 17175 1853 17187 1887
rect 17236 1884 17264 1924
rect 17310 1893 17316 1896
rect 17307 1884 17316 1893
rect 17236 1856 17316 1884
rect 17129 1847 17187 1853
rect 17307 1847 17316 1856
rect 16132 1788 16712 1816
rect 16393 1751 16451 1757
rect 16393 1748 16405 1751
rect 15764 1720 16405 1748
rect 16393 1717 16405 1720
rect 16439 1717 16451 1751
rect 16393 1711 16451 1717
rect 16482 1708 16488 1760
rect 16540 1748 16546 1760
rect 17144 1748 17172 1847
rect 17310 1844 17316 1847
rect 17368 1844 17374 1896
rect 16540 1720 17172 1748
rect 16540 1708 16546 1720
rect 552 1658 17664 1680
rect 552 1606 4366 1658
rect 4418 1606 4430 1658
rect 4482 1606 4494 1658
rect 4546 1606 4558 1658
rect 4610 1606 4622 1658
rect 4674 1606 4686 1658
rect 4738 1606 10366 1658
rect 10418 1606 10430 1658
rect 10482 1606 10494 1658
rect 10546 1606 10558 1658
rect 10610 1606 10622 1658
rect 10674 1606 10686 1658
rect 10738 1606 16366 1658
rect 16418 1606 16430 1658
rect 16482 1606 16494 1658
rect 16546 1606 16558 1658
rect 16610 1606 16622 1658
rect 16674 1606 16686 1658
rect 16738 1606 17664 1658
rect 552 1584 17664 1606
rect 1210 1504 1216 1556
rect 1268 1504 1274 1556
rect 1762 1504 1768 1556
rect 1820 1504 1826 1556
rect 2038 1504 2044 1556
rect 2096 1504 2102 1556
rect 2409 1547 2467 1553
rect 2409 1513 2421 1547
rect 2455 1544 2467 1547
rect 2682 1544 2688 1556
rect 2455 1516 2688 1544
rect 2455 1513 2467 1516
rect 2409 1507 2467 1513
rect 2682 1504 2688 1516
rect 2740 1504 2746 1556
rect 2961 1547 3019 1553
rect 2961 1513 2973 1547
rect 3007 1544 3019 1547
rect 3326 1544 3332 1556
rect 3007 1516 3332 1544
rect 3007 1513 3019 1516
rect 2961 1507 3019 1513
rect 3326 1504 3332 1516
rect 3384 1504 3390 1556
rect 3510 1504 3516 1556
rect 3568 1544 3574 1556
rect 3697 1547 3755 1553
rect 3697 1544 3709 1547
rect 3568 1516 3709 1544
rect 3568 1504 3574 1516
rect 3697 1513 3709 1516
rect 3743 1513 3755 1547
rect 3697 1507 3755 1513
rect 4798 1504 4804 1556
rect 4856 1504 4862 1556
rect 5810 1504 5816 1556
rect 5868 1504 5874 1556
rect 6914 1504 6920 1556
rect 6972 1504 6978 1556
rect 7006 1504 7012 1556
rect 7064 1504 7070 1556
rect 7650 1504 7656 1556
rect 7708 1504 7714 1556
rect 7834 1504 7840 1556
rect 7892 1504 7898 1556
rect 8110 1544 8116 1556
rect 7944 1516 8116 1544
rect 1228 1408 1256 1504
rect 1305 1411 1363 1417
rect 1305 1408 1317 1411
rect 1228 1380 1317 1408
rect 1305 1377 1317 1380
rect 1351 1377 1363 1411
rect 1305 1371 1363 1377
rect 1673 1411 1731 1417
rect 1673 1377 1685 1411
rect 1719 1408 1731 1411
rect 1780 1408 1808 1504
rect 1946 1436 1952 1488
rect 2004 1436 2010 1488
rect 2056 1476 2084 1504
rect 2225 1479 2283 1485
rect 2225 1476 2237 1479
rect 2056 1448 2237 1476
rect 2225 1445 2237 1448
rect 2271 1445 2283 1479
rect 2593 1479 2651 1485
rect 2593 1476 2605 1479
rect 2225 1439 2283 1445
rect 2424 1448 2605 1476
rect 1719 1380 1808 1408
rect 1964 1408 1992 1436
rect 2041 1411 2099 1417
rect 2041 1408 2053 1411
rect 1964 1380 2053 1408
rect 1719 1377 1731 1380
rect 1673 1371 1731 1377
rect 2041 1377 2053 1380
rect 2087 1377 2099 1411
rect 2041 1371 2099 1377
rect 2424 1272 2452 1448
rect 2593 1445 2605 1448
rect 2639 1445 2651 1479
rect 2793 1479 2851 1485
rect 2793 1476 2805 1479
rect 2593 1439 2651 1445
rect 2700 1448 2805 1476
rect 2498 1368 2504 1420
rect 2556 1408 2562 1420
rect 2700 1408 2728 1448
rect 2793 1445 2805 1448
rect 2839 1445 2851 1479
rect 2793 1439 2851 1445
rect 3786 1436 3792 1488
rect 3844 1476 3850 1488
rect 4816 1476 4844 1504
rect 3844 1448 4844 1476
rect 3844 1436 3850 1448
rect 2556 1380 2728 1408
rect 2556 1368 2562 1380
rect 2958 1368 2964 1420
rect 3016 1408 3022 1420
rect 3237 1411 3295 1417
rect 3237 1408 3249 1411
rect 3016 1380 3249 1408
rect 3016 1368 3022 1380
rect 3237 1377 3249 1380
rect 3283 1377 3295 1411
rect 3237 1371 3295 1377
rect 3329 1411 3387 1417
rect 3329 1377 3341 1411
rect 3375 1408 3387 1411
rect 3694 1408 3700 1420
rect 3375 1380 3700 1408
rect 3375 1377 3387 1380
rect 3329 1371 3387 1377
rect 3694 1368 3700 1380
rect 3752 1368 3758 1420
rect 3970 1368 3976 1420
rect 4028 1368 4034 1420
rect 4062 1368 4068 1420
rect 4120 1368 4126 1420
rect 4157 1411 4215 1417
rect 4157 1377 4169 1411
rect 4203 1406 4215 1411
rect 4246 1406 4252 1420
rect 4203 1378 4252 1406
rect 4203 1377 4215 1378
rect 4157 1371 4215 1377
rect 4246 1368 4252 1378
rect 4304 1368 4310 1420
rect 4376 1417 4404 1448
rect 4890 1436 4896 1488
rect 4948 1436 4954 1488
rect 5828 1476 5856 1504
rect 5828 1448 6500 1476
rect 4341 1411 4404 1417
rect 4341 1377 4353 1411
rect 4387 1378 4404 1411
rect 4387 1377 4399 1378
rect 4341 1371 4399 1377
rect 4798 1368 4804 1420
rect 4856 1368 4862 1420
rect 4908 1408 4936 1436
rect 4908 1380 5488 1408
rect 3418 1300 3424 1352
rect 3476 1300 3482 1352
rect 3513 1343 3571 1349
rect 3513 1309 3525 1343
rect 3559 1340 3571 1343
rect 3602 1340 3608 1352
rect 3559 1312 3608 1340
rect 3559 1309 3571 1312
rect 3513 1303 3571 1309
rect 3602 1300 3608 1312
rect 3660 1300 3666 1352
rect 3988 1340 4016 1368
rect 4709 1343 4767 1349
rect 4709 1340 4721 1343
rect 3988 1312 4721 1340
rect 4709 1309 4721 1312
rect 4755 1309 4767 1343
rect 4709 1303 4767 1309
rect 5169 1343 5227 1349
rect 5169 1309 5181 1343
rect 5215 1309 5227 1343
rect 5460 1340 5488 1380
rect 5534 1368 5540 1420
rect 5592 1368 5598 1420
rect 5902 1368 5908 1420
rect 5960 1408 5966 1420
rect 5997 1411 6055 1417
rect 5997 1408 6009 1411
rect 5960 1380 6009 1408
rect 5960 1368 5966 1380
rect 5997 1377 6009 1380
rect 6043 1377 6055 1411
rect 5997 1371 6055 1377
rect 6273 1411 6331 1417
rect 6273 1377 6285 1411
rect 6319 1408 6331 1411
rect 6362 1408 6368 1420
rect 6319 1380 6368 1408
rect 6319 1377 6331 1380
rect 6273 1371 6331 1377
rect 6362 1368 6368 1380
rect 6420 1368 6426 1420
rect 6472 1417 6500 1448
rect 6932 1417 6960 1504
rect 7668 1476 7696 1504
rect 7208 1448 7696 1476
rect 6457 1411 6515 1417
rect 6457 1377 6469 1411
rect 6503 1377 6515 1411
rect 6457 1371 6515 1377
rect 6917 1411 6975 1417
rect 6917 1377 6929 1411
rect 6963 1377 6975 1411
rect 6917 1371 6975 1377
rect 7009 1411 7067 1417
rect 7009 1377 7021 1411
rect 7055 1408 7067 1411
rect 7098 1408 7104 1420
rect 7055 1380 7104 1408
rect 7055 1377 7067 1380
rect 7009 1371 7067 1377
rect 6089 1343 6147 1349
rect 6089 1340 6101 1343
rect 5460 1312 6101 1340
rect 5169 1303 5227 1309
rect 6089 1309 6101 1312
rect 6135 1309 6147 1343
rect 6089 1303 6147 1309
rect 6181 1343 6239 1349
rect 6181 1309 6193 1343
rect 6227 1340 6239 1343
rect 6638 1340 6644 1352
rect 6227 1312 6644 1340
rect 6227 1309 6239 1312
rect 6181 1303 6239 1309
rect 3234 1272 3240 1284
rect 2424 1244 3240 1272
rect 3234 1232 3240 1244
rect 3292 1232 3298 1284
rect 3436 1272 3464 1300
rect 3881 1275 3939 1281
rect 3881 1272 3893 1275
rect 3436 1244 3893 1272
rect 3881 1241 3893 1244
rect 3927 1241 3939 1275
rect 5184 1272 5212 1303
rect 6638 1300 6644 1312
rect 6696 1300 6702 1352
rect 6932 1340 6960 1371
rect 7098 1368 7104 1380
rect 7156 1368 7162 1420
rect 7208 1417 7236 1448
rect 7193 1411 7251 1417
rect 7193 1377 7205 1411
rect 7239 1377 7251 1411
rect 7193 1371 7251 1377
rect 7469 1411 7527 1417
rect 7469 1377 7481 1411
rect 7515 1408 7527 1411
rect 7558 1408 7564 1420
rect 7515 1380 7564 1408
rect 7515 1377 7527 1380
rect 7469 1371 7527 1377
rect 7558 1368 7564 1380
rect 7616 1368 7622 1420
rect 7653 1411 7711 1417
rect 7653 1377 7665 1411
rect 7699 1408 7711 1411
rect 7852 1408 7880 1504
rect 7944 1417 7972 1516
rect 8110 1504 8116 1516
rect 8168 1504 8174 1556
rect 9766 1504 9772 1556
rect 9824 1504 9830 1556
rect 10042 1504 10048 1556
rect 10100 1544 10106 1556
rect 12434 1544 12440 1556
rect 10100 1516 10226 1544
rect 10100 1504 10106 1516
rect 8018 1436 8024 1488
rect 8076 1476 8082 1488
rect 8076 1448 8156 1476
rect 8076 1436 8082 1448
rect 8128 1417 8156 1448
rect 8478 1436 8484 1488
rect 8536 1476 8542 1488
rect 8938 1476 8944 1488
rect 8536 1448 8944 1476
rect 8536 1436 8542 1448
rect 8938 1436 8944 1448
rect 8996 1436 9002 1488
rect 9784 1476 9812 1504
rect 10198 1476 10226 1516
rect 10520 1516 12440 1544
rect 9048 1448 9904 1476
rect 10198 1448 10364 1476
rect 9048 1417 9076 1448
rect 7699 1380 7880 1408
rect 7929 1411 7987 1417
rect 7699 1377 7711 1380
rect 7653 1371 7711 1377
rect 7929 1377 7941 1411
rect 7975 1377 7987 1411
rect 7929 1371 7987 1377
rect 8113 1411 8171 1417
rect 8113 1377 8125 1411
rect 8159 1377 8171 1411
rect 9033 1411 9091 1417
rect 8113 1371 8171 1377
rect 8220 1380 8984 1408
rect 7285 1343 7343 1349
rect 7285 1340 7297 1343
rect 6932 1312 7297 1340
rect 7285 1309 7297 1312
rect 7331 1309 7343 1343
rect 7285 1303 7343 1309
rect 7742 1300 7748 1352
rect 7800 1300 7806 1352
rect 7837 1343 7895 1349
rect 7837 1309 7849 1343
rect 7883 1309 7895 1343
rect 7837 1303 7895 1309
rect 5184 1244 6408 1272
rect 3881 1235 3939 1241
rect 6380 1216 6408 1244
rect 1118 1164 1124 1216
rect 1176 1164 1182 1216
rect 1489 1207 1547 1213
rect 1489 1173 1501 1207
rect 1535 1204 1547 1207
rect 1762 1204 1768 1216
rect 1535 1176 1768 1204
rect 1535 1173 1547 1176
rect 1489 1167 1547 1173
rect 1762 1164 1768 1176
rect 1820 1164 1826 1216
rect 2774 1164 2780 1216
rect 2832 1164 2838 1216
rect 3602 1164 3608 1216
rect 3660 1204 3666 1216
rect 4249 1207 4307 1213
rect 4249 1204 4261 1207
rect 3660 1176 4261 1204
rect 3660 1164 3666 1176
rect 4249 1173 4261 1176
rect 4295 1173 4307 1207
rect 4249 1167 4307 1173
rect 5350 1164 5356 1216
rect 5408 1164 5414 1216
rect 5810 1164 5816 1216
rect 5868 1164 5874 1216
rect 6362 1164 6368 1216
rect 6420 1164 6426 1216
rect 6638 1164 6644 1216
rect 6696 1164 6702 1216
rect 6730 1164 6736 1216
rect 6788 1164 6794 1216
rect 6822 1164 6828 1216
rect 6880 1204 6886 1216
rect 7852 1204 7880 1303
rect 8220 1204 8248 1380
rect 8297 1343 8355 1349
rect 8297 1309 8309 1343
rect 8343 1340 8355 1343
rect 8478 1340 8484 1352
rect 8343 1312 8484 1340
rect 8343 1309 8355 1312
rect 8297 1303 8355 1309
rect 8478 1300 8484 1312
rect 8536 1300 8542 1352
rect 8956 1340 8984 1380
rect 9033 1377 9045 1411
rect 9079 1377 9091 1411
rect 9033 1371 9091 1377
rect 9214 1368 9220 1420
rect 9272 1368 9278 1420
rect 9677 1411 9735 1417
rect 9677 1377 9689 1411
rect 9723 1377 9735 1411
rect 9677 1371 9735 1377
rect 9306 1340 9312 1352
rect 8956 1312 9312 1340
rect 9306 1300 9312 1312
rect 9364 1300 9370 1352
rect 9692 1340 9720 1371
rect 9766 1368 9772 1420
rect 9824 1368 9830 1420
rect 9876 1417 9904 1448
rect 9861 1411 9919 1417
rect 9861 1377 9873 1411
rect 9907 1377 9919 1411
rect 9861 1371 9919 1377
rect 10042 1368 10048 1420
rect 10100 1368 10106 1420
rect 10336 1417 10364 1448
rect 10321 1411 10379 1417
rect 10321 1377 10333 1411
rect 10367 1377 10379 1411
rect 10520 1408 10548 1516
rect 12434 1504 12440 1516
rect 12492 1504 12498 1556
rect 12526 1504 12532 1556
rect 12584 1544 12590 1556
rect 12621 1547 12679 1553
rect 12621 1544 12633 1547
rect 12584 1516 12633 1544
rect 12584 1504 12590 1516
rect 12621 1513 12633 1516
rect 12667 1513 12679 1547
rect 12621 1507 12679 1513
rect 13446 1504 13452 1556
rect 13504 1544 13510 1556
rect 15013 1547 15071 1553
rect 13504 1516 14596 1544
rect 13504 1504 13510 1516
rect 10686 1436 10692 1488
rect 10744 1476 10750 1488
rect 11422 1476 11428 1488
rect 10744 1448 11192 1476
rect 10744 1436 10750 1448
rect 10321 1371 10379 1377
rect 10428 1380 10548 1408
rect 10597 1411 10655 1417
rect 10428 1340 10456 1380
rect 10597 1377 10609 1411
rect 10643 1408 10655 1411
rect 10643 1380 11100 1408
rect 10643 1377 10655 1380
rect 10597 1371 10655 1377
rect 11072 1352 11100 1380
rect 9692 1312 10456 1340
rect 10502 1300 10508 1352
rect 10560 1300 10566 1352
rect 10962 1300 10968 1352
rect 11020 1300 11026 1352
rect 11054 1300 11060 1352
rect 11112 1300 11118 1352
rect 11164 1340 11192 1448
rect 11256 1448 11428 1476
rect 11256 1417 11284 1448
rect 11422 1436 11428 1448
rect 11480 1436 11486 1488
rect 11885 1479 11943 1485
rect 11885 1445 11897 1479
rect 11931 1476 11943 1479
rect 11931 1448 12580 1476
rect 11931 1445 11943 1448
rect 11885 1439 11943 1445
rect 11241 1411 11299 1417
rect 11241 1377 11253 1411
rect 11287 1377 11299 1411
rect 12345 1411 12403 1417
rect 12345 1408 12357 1411
rect 11241 1371 11299 1377
rect 11348 1380 12357 1408
rect 11348 1340 11376 1380
rect 12345 1377 12357 1380
rect 12391 1377 12403 1411
rect 12345 1371 12403 1377
rect 11164 1312 11376 1340
rect 12066 1300 12072 1352
rect 12124 1300 12130 1352
rect 12158 1300 12164 1352
rect 12216 1300 12222 1352
rect 8846 1232 8852 1284
rect 8904 1232 8910 1284
rect 8938 1232 8944 1284
rect 8996 1272 9002 1284
rect 8996 1244 9996 1272
rect 8996 1232 9002 1244
rect 6880 1176 8248 1204
rect 6880 1164 6886 1176
rect 8386 1164 8392 1216
rect 8444 1204 8450 1216
rect 9401 1207 9459 1213
rect 9401 1204 9413 1207
rect 8444 1176 9413 1204
rect 8444 1164 8450 1176
rect 9401 1173 9413 1176
rect 9447 1173 9459 1207
rect 9968 1204 9996 1244
rect 10042 1232 10048 1284
rect 10100 1272 10106 1284
rect 10137 1275 10195 1281
rect 10137 1272 10149 1275
rect 10100 1244 10149 1272
rect 10100 1232 10106 1244
rect 10137 1241 10149 1244
rect 10183 1241 10195 1275
rect 10137 1235 10195 1241
rect 10413 1275 10471 1281
rect 10413 1241 10425 1275
rect 10459 1272 10471 1275
rect 12176 1272 12204 1300
rect 10459 1244 12204 1272
rect 12552 1272 12580 1448
rect 13170 1436 13176 1488
rect 13228 1436 13234 1488
rect 13262 1436 13268 1488
rect 13320 1476 13326 1488
rect 13320 1448 13584 1476
rect 13320 1436 13326 1448
rect 12710 1368 12716 1420
rect 12768 1368 12774 1420
rect 12805 1411 12863 1417
rect 12805 1377 12817 1411
rect 12851 1408 12863 1411
rect 12894 1408 12900 1420
rect 12851 1380 12900 1408
rect 12851 1377 12863 1380
rect 12805 1371 12863 1377
rect 12894 1368 12900 1380
rect 12952 1368 12958 1420
rect 12986 1368 12992 1420
rect 13044 1368 13050 1420
rect 13354 1368 13360 1420
rect 13412 1368 13418 1420
rect 13556 1417 13584 1448
rect 13541 1411 13599 1417
rect 13541 1377 13553 1411
rect 13587 1377 13599 1411
rect 13541 1371 13599 1377
rect 13906 1368 13912 1420
rect 13964 1368 13970 1420
rect 14090 1368 14096 1420
rect 14148 1368 14154 1420
rect 14366 1368 14372 1420
rect 14424 1368 14430 1420
rect 14568 1417 14596 1516
rect 15013 1513 15025 1547
rect 15059 1544 15071 1547
rect 15286 1544 15292 1556
rect 15059 1516 15292 1544
rect 15059 1513 15071 1516
rect 15013 1507 15071 1513
rect 15286 1504 15292 1516
rect 15344 1504 15350 1556
rect 15470 1504 15476 1556
rect 15528 1544 15534 1556
rect 15749 1547 15807 1553
rect 15749 1544 15761 1547
rect 15528 1516 15761 1544
rect 15528 1504 15534 1516
rect 15749 1513 15761 1516
rect 15795 1513 15807 1547
rect 15749 1507 15807 1513
rect 16022 1504 16028 1556
rect 16080 1544 16086 1556
rect 16080 1516 16896 1544
rect 16080 1504 16086 1516
rect 16868 1485 16896 1516
rect 16209 1479 16267 1485
rect 16209 1476 16221 1479
rect 15028 1448 16221 1476
rect 14553 1411 14611 1417
rect 14553 1377 14565 1411
rect 14599 1377 14611 1411
rect 14553 1371 14611 1377
rect 14734 1368 14740 1420
rect 14792 1408 14798 1420
rect 14829 1411 14887 1417
rect 14829 1408 14841 1411
rect 14792 1380 14841 1408
rect 14792 1368 14798 1380
rect 14829 1377 14841 1380
rect 14875 1377 14887 1411
rect 14829 1371 14887 1377
rect 12728 1340 12756 1368
rect 13081 1343 13139 1349
rect 13081 1340 13093 1343
rect 12728 1312 13093 1340
rect 13081 1309 13093 1312
rect 13127 1340 13139 1343
rect 13633 1343 13691 1349
rect 13633 1340 13645 1343
rect 13127 1312 13645 1340
rect 13127 1309 13139 1312
rect 13081 1303 13139 1309
rect 13633 1309 13645 1312
rect 13679 1340 13691 1343
rect 14185 1343 14243 1349
rect 14185 1340 14197 1343
rect 13679 1312 14197 1340
rect 13679 1309 13691 1312
rect 13633 1303 13691 1309
rect 14185 1309 14197 1312
rect 14231 1309 14243 1343
rect 14185 1303 14243 1309
rect 14277 1343 14335 1349
rect 14277 1309 14289 1343
rect 14323 1309 14335 1343
rect 15028 1340 15056 1448
rect 16209 1445 16221 1448
rect 16255 1445 16267 1479
rect 16209 1439 16267 1445
rect 16853 1479 16911 1485
rect 16853 1445 16865 1479
rect 16899 1476 16911 1479
rect 17218 1476 17224 1488
rect 16899 1448 17224 1476
rect 16899 1445 16911 1448
rect 16853 1439 16911 1445
rect 17218 1436 17224 1448
rect 17276 1436 17282 1488
rect 17402 1436 17408 1488
rect 17460 1436 17466 1488
rect 15102 1368 15108 1420
rect 15160 1408 15166 1420
rect 15381 1411 15439 1417
rect 15381 1408 15393 1411
rect 15160 1380 15393 1408
rect 15160 1368 15166 1380
rect 15381 1377 15393 1380
rect 15427 1377 15439 1411
rect 15381 1371 15439 1377
rect 15746 1368 15752 1420
rect 15804 1368 15810 1420
rect 15930 1368 15936 1420
rect 15988 1408 15994 1420
rect 17034 1408 17040 1420
rect 15988 1380 17040 1408
rect 15988 1368 15994 1380
rect 17034 1368 17040 1380
rect 17092 1408 17098 1420
rect 17420 1408 17448 1436
rect 17092 1380 17448 1408
rect 17092 1368 17098 1380
rect 14277 1303 14335 1309
rect 14660 1312 15056 1340
rect 15289 1343 15347 1349
rect 13725 1275 13783 1281
rect 13725 1272 13737 1275
rect 12552 1244 13737 1272
rect 10459 1241 10471 1244
rect 10413 1235 10471 1241
rect 13725 1241 13737 1244
rect 13771 1241 13783 1275
rect 13725 1235 13783 1241
rect 14090 1232 14096 1284
rect 14148 1272 14154 1284
rect 14292 1272 14320 1303
rect 14148 1244 14320 1272
rect 14148 1232 14154 1244
rect 11057 1207 11115 1213
rect 11057 1204 11069 1207
rect 9968 1176 11069 1204
rect 9401 1167 9459 1173
rect 11057 1173 11069 1176
rect 11103 1173 11115 1207
rect 11057 1167 11115 1173
rect 11425 1207 11483 1213
rect 11425 1173 11437 1207
rect 11471 1204 11483 1207
rect 11514 1204 11520 1216
rect 11471 1176 11520 1204
rect 11471 1173 11483 1176
rect 11425 1167 11483 1173
rect 11514 1164 11520 1176
rect 11572 1164 11578 1216
rect 11606 1164 11612 1216
rect 11664 1164 11670 1216
rect 11882 1164 11888 1216
rect 11940 1204 11946 1216
rect 12161 1207 12219 1213
rect 12161 1204 12173 1207
rect 11940 1176 12173 1204
rect 11940 1164 11946 1176
rect 12161 1173 12173 1176
rect 12207 1173 12219 1207
rect 12161 1167 12219 1173
rect 12529 1207 12587 1213
rect 12529 1173 12541 1207
rect 12575 1204 12587 1207
rect 14660 1204 14688 1312
rect 15289 1309 15301 1343
rect 15335 1340 15347 1343
rect 15764 1340 15792 1368
rect 16669 1343 16727 1349
rect 16669 1340 16681 1343
rect 15335 1312 15424 1340
rect 15764 1312 16681 1340
rect 15335 1309 15347 1312
rect 15289 1303 15347 1309
rect 15396 1284 15424 1312
rect 16669 1309 16681 1312
rect 16715 1309 16727 1343
rect 16669 1303 16727 1309
rect 14737 1275 14795 1281
rect 14737 1241 14749 1275
rect 14783 1272 14795 1275
rect 15194 1272 15200 1284
rect 14783 1244 15200 1272
rect 14783 1241 14795 1244
rect 14737 1235 14795 1241
rect 15194 1232 15200 1244
rect 15252 1232 15258 1284
rect 15378 1232 15384 1284
rect 15436 1232 15442 1284
rect 15580 1244 16344 1272
rect 12575 1176 14688 1204
rect 12575 1173 12587 1176
rect 12529 1167 12587 1173
rect 14918 1164 14924 1216
rect 14976 1204 14982 1216
rect 15580 1204 15608 1244
rect 16316 1213 16344 1244
rect 14976 1176 15608 1204
rect 16301 1207 16359 1213
rect 14976 1164 14982 1176
rect 16301 1173 16313 1207
rect 16347 1173 16359 1207
rect 16301 1167 16359 1173
rect 552 1114 17664 1136
rect 552 1062 1366 1114
rect 1418 1062 1430 1114
rect 1482 1062 1494 1114
rect 1546 1062 1558 1114
rect 1610 1062 1622 1114
rect 1674 1062 1686 1114
rect 1738 1062 7366 1114
rect 7418 1062 7430 1114
rect 7482 1062 7494 1114
rect 7546 1062 7558 1114
rect 7610 1062 7622 1114
rect 7674 1062 7686 1114
rect 7738 1062 13366 1114
rect 13418 1062 13430 1114
rect 13482 1062 13494 1114
rect 13546 1062 13558 1114
rect 13610 1062 13622 1114
rect 13674 1062 13686 1114
rect 13738 1062 17664 1114
rect 552 1040 17664 1062
rect 2498 960 2504 1012
rect 2556 960 2562 1012
rect 5810 960 5816 1012
rect 5868 960 5874 1012
rect 8846 960 8852 1012
rect 8904 960 8910 1012
rect 9306 960 9312 1012
rect 9364 960 9370 1012
rect 9861 1003 9919 1009
rect 9861 969 9873 1003
rect 9907 1000 9919 1003
rect 9950 1000 9956 1012
rect 9907 972 9956 1000
rect 9907 969 9919 972
rect 9861 963 9919 969
rect 9950 960 9956 972
rect 10008 960 10014 1012
rect 10505 1003 10563 1009
rect 10505 969 10517 1003
rect 10551 969 10563 1003
rect 10505 963 10563 969
rect 11057 1003 11115 1009
rect 11057 969 11069 1003
rect 11103 1000 11115 1003
rect 11146 1000 11152 1012
rect 11103 972 11152 1000
rect 11103 969 11115 972
rect 11057 963 11115 969
rect 2038 892 2044 944
rect 2096 932 2102 944
rect 2685 935 2743 941
rect 2685 932 2697 935
rect 2096 904 2697 932
rect 2096 892 2102 904
rect 2685 901 2697 904
rect 2731 901 2743 935
rect 2685 895 2743 901
rect 2406 824 2412 876
rect 2464 864 2470 876
rect 5828 864 5856 960
rect 8110 864 8116 876
rect 2464 836 2544 864
rect 2464 824 2470 836
rect 1118 756 1124 808
rect 1176 756 1182 808
rect 1581 799 1639 805
rect 1581 765 1593 799
rect 1627 796 1639 799
rect 1762 796 1768 808
rect 1627 768 1768 796
rect 1627 765 1639 768
rect 1581 759 1639 765
rect 1762 756 1768 768
rect 1820 756 1826 808
rect 1854 756 1860 808
rect 1912 796 1918 808
rect 2225 799 2283 805
rect 2225 796 2237 799
rect 1912 768 2237 796
rect 1912 756 1918 768
rect 2225 765 2237 768
rect 2271 765 2283 799
rect 2225 759 2283 765
rect 2314 756 2320 808
rect 2372 756 2378 808
rect 2516 805 2544 836
rect 2884 836 5856 864
rect 6012 836 8116 864
rect 2884 805 2912 836
rect 2501 799 2559 805
rect 2501 765 2513 799
rect 2547 765 2559 799
rect 2501 759 2559 765
rect 2869 799 2927 805
rect 2869 765 2881 799
rect 2915 765 2927 799
rect 2869 759 2927 765
rect 3513 799 3571 805
rect 3513 765 3525 799
rect 3559 765 3571 799
rect 3513 759 3571 765
rect 3881 799 3939 805
rect 3881 765 3893 799
rect 3927 796 3939 799
rect 4154 796 4160 808
rect 3927 768 4160 796
rect 3927 765 3939 768
rect 3881 759 3939 765
rect 2332 728 2360 756
rect 2409 731 2467 737
rect 2409 728 2421 731
rect 2332 700 2421 728
rect 2409 697 2421 700
rect 2455 697 2467 731
rect 3528 728 3556 759
rect 4154 756 4160 768
rect 4212 756 4218 808
rect 4617 799 4675 805
rect 4617 765 4629 799
rect 4663 796 4675 799
rect 5258 796 5264 808
rect 4663 768 5264 796
rect 4663 765 4675 768
rect 4617 759 4675 765
rect 5258 756 5264 768
rect 5316 756 5322 808
rect 5350 756 5356 808
rect 5408 756 5414 808
rect 6012 728 6040 836
rect 8110 824 8116 836
rect 8168 824 8174 876
rect 8864 864 8892 960
rect 8220 836 8892 864
rect 6086 756 6092 808
rect 6144 756 6150 808
rect 6638 756 6644 808
rect 6696 756 6702 808
rect 6730 756 6736 808
rect 6788 796 6794 808
rect 8220 805 8248 836
rect 6825 799 6883 805
rect 6825 796 6837 799
rect 6788 768 6837 796
rect 6788 756 6794 768
rect 6825 765 6837 768
rect 6871 765 6883 799
rect 6825 759 6883 765
rect 7285 799 7343 805
rect 7285 765 7297 799
rect 7331 765 7343 799
rect 7285 759 7343 765
rect 8205 799 8263 805
rect 8205 765 8217 799
rect 8251 765 8263 799
rect 8205 759 8263 765
rect 3528 700 6040 728
rect 6656 728 6684 756
rect 7300 728 7328 759
rect 8478 756 8484 808
rect 8536 756 8542 808
rect 6656 700 7328 728
rect 2409 691 2467 697
rect 8110 688 8116 740
rect 8168 728 8174 740
rect 9324 728 9352 960
rect 9398 892 9404 944
rect 9456 932 9462 944
rect 10520 932 10548 963
rect 11146 960 11152 972
rect 11204 960 11210 1012
rect 11238 960 11244 1012
rect 11296 1000 11302 1012
rect 11609 1003 11667 1009
rect 11609 1000 11621 1003
rect 11296 972 11621 1000
rect 11296 960 11302 972
rect 11609 969 11621 972
rect 11655 969 11667 1003
rect 11609 963 11667 969
rect 12713 1003 12771 1009
rect 12713 969 12725 1003
rect 12759 1000 12771 1003
rect 12802 1000 12808 1012
rect 12759 972 12808 1000
rect 12759 969 12771 972
rect 12713 963 12771 969
rect 12802 960 12808 972
rect 12860 960 12866 1012
rect 13170 1000 13176 1012
rect 12912 972 13176 1000
rect 12912 932 12940 972
rect 13170 960 13176 972
rect 13228 960 13234 1012
rect 14182 1000 14188 1012
rect 13924 972 14188 1000
rect 9456 904 10548 932
rect 12406 904 12940 932
rect 13081 935 13139 941
rect 9456 892 9462 904
rect 12406 864 12434 904
rect 13081 901 13093 935
rect 13127 932 13139 935
rect 13924 932 13952 972
rect 14182 960 14188 972
rect 14240 960 14246 1012
rect 14274 960 14280 1012
rect 14332 1000 14338 1012
rect 14369 1003 14427 1009
rect 14369 1000 14381 1003
rect 14332 972 14381 1000
rect 14332 960 14338 972
rect 14369 969 14381 972
rect 14415 969 14427 1003
rect 14369 963 14427 969
rect 14642 960 14648 1012
rect 14700 1000 14706 1012
rect 14921 1003 14979 1009
rect 14921 1000 14933 1003
rect 14700 972 14933 1000
rect 14700 960 14706 972
rect 14921 969 14933 972
rect 14967 969 14979 1003
rect 14921 963 14979 969
rect 15010 960 15016 1012
rect 15068 1000 15074 1012
rect 15289 1003 15347 1009
rect 15289 1000 15301 1003
rect 15068 972 15301 1000
rect 15068 960 15074 972
rect 15289 969 15301 972
rect 15335 969 15347 1003
rect 15289 963 15347 969
rect 16301 1003 16359 1009
rect 16301 969 16313 1003
rect 16347 969 16359 1003
rect 16301 963 16359 969
rect 13127 904 13952 932
rect 13127 901 13139 904
rect 13081 895 13139 901
rect 13998 892 14004 944
rect 14056 932 14062 944
rect 16316 932 16344 963
rect 17034 960 17040 1012
rect 17092 960 17098 1012
rect 14056 904 16344 932
rect 14056 892 14062 904
rect 9600 836 12434 864
rect 9600 805 9628 836
rect 12710 824 12716 876
rect 12768 864 12774 876
rect 13173 867 13231 873
rect 13173 864 13185 867
rect 12768 836 13185 864
rect 12768 824 12774 836
rect 13173 833 13185 836
rect 13219 833 13231 867
rect 13173 827 13231 833
rect 13354 824 13360 876
rect 13412 864 13418 876
rect 15749 867 15807 873
rect 15749 864 15761 867
rect 13412 836 15761 864
rect 13412 824 13418 836
rect 15749 833 15761 836
rect 15795 833 15807 867
rect 15749 827 15807 833
rect 16669 867 16727 873
rect 16669 833 16681 867
rect 16715 864 16727 867
rect 17126 864 17132 876
rect 16715 836 17132 864
rect 16715 833 16727 836
rect 16669 827 16727 833
rect 17126 824 17132 836
rect 17184 824 17190 876
rect 9585 799 9643 805
rect 9585 765 9597 799
rect 9631 765 9643 799
rect 9585 759 9643 765
rect 9769 799 9827 805
rect 9769 765 9781 799
rect 9815 796 9827 799
rect 9858 796 9864 808
rect 9815 768 9864 796
rect 9815 765 9827 768
rect 9769 759 9827 765
rect 9784 728 9812 759
rect 9858 756 9864 768
rect 9916 756 9922 808
rect 10045 799 10103 805
rect 10045 765 10057 799
rect 10091 796 10103 799
rect 10091 768 10824 796
rect 10091 765 10103 768
rect 10045 759 10103 765
rect 8168 700 8616 728
rect 9324 700 9812 728
rect 10229 731 10287 737
rect 8168 688 8174 700
rect 566 620 572 672
rect 624 660 630 672
rect 937 663 995 669
rect 937 660 949 663
rect 624 632 949 660
rect 624 620 630 632
rect 937 629 949 632
rect 983 629 995 663
rect 937 623 995 629
rect 1302 620 1308 672
rect 1360 620 1366 672
rect 2774 620 2780 672
rect 2832 660 2838 672
rect 3329 663 3387 669
rect 3329 660 3341 663
rect 2832 632 3341 660
rect 2832 620 2838 632
rect 3329 629 3341 632
rect 3375 629 3387 663
rect 3329 623 3387 629
rect 3694 620 3700 672
rect 3752 620 3758 672
rect 4246 620 4252 672
rect 4304 660 4310 672
rect 4433 663 4491 669
rect 4433 660 4445 663
rect 4304 632 4445 660
rect 4304 620 4310 632
rect 4433 629 4445 632
rect 4479 629 4491 663
rect 4433 623 4491 629
rect 5166 620 5172 672
rect 5224 620 5230 672
rect 5902 620 5908 672
rect 5960 620 5966 672
rect 6638 620 6644 672
rect 6696 620 6702 672
rect 7190 620 7196 672
rect 7248 660 7254 672
rect 7469 663 7527 669
rect 7469 660 7481 663
rect 7248 632 7481 660
rect 7248 620 7254 632
rect 7469 629 7481 632
rect 7515 629 7527 663
rect 7469 623 7527 629
rect 8021 663 8079 669
rect 8021 629 8033 663
rect 8067 660 8079 663
rect 8386 660 8392 672
rect 8067 632 8392 660
rect 8067 629 8079 632
rect 8021 623 8079 629
rect 8386 620 8392 632
rect 8444 620 8450 672
rect 8588 669 8616 700
rect 10229 697 10241 731
rect 10275 728 10287 731
rect 10413 731 10471 737
rect 10413 728 10425 731
rect 10275 700 10425 728
rect 10275 697 10287 700
rect 10229 691 10287 697
rect 10413 697 10425 700
rect 10459 697 10471 731
rect 10796 728 10824 768
rect 10962 756 10968 808
rect 11020 756 11026 808
rect 11241 799 11299 805
rect 11241 796 11253 799
rect 11072 768 11253 796
rect 11072 740 11100 768
rect 11241 765 11253 768
rect 11287 765 11299 799
rect 11241 759 11299 765
rect 11790 756 11796 808
rect 11848 756 11854 808
rect 11977 799 12035 805
rect 11977 765 11989 799
rect 12023 765 12035 799
rect 11977 759 12035 765
rect 11054 728 11060 740
rect 10796 700 11060 728
rect 10413 691 10471 697
rect 11054 688 11060 700
rect 11112 688 11118 740
rect 11146 688 11152 740
rect 11204 728 11210 740
rect 11992 728 12020 759
rect 12434 756 12440 808
rect 12492 756 12498 808
rect 12897 799 12955 805
rect 12897 765 12909 799
rect 12943 796 12955 799
rect 12943 768 13124 796
rect 12943 765 12955 768
rect 12897 759 12955 765
rect 11204 700 11560 728
rect 11992 700 12296 728
rect 11204 688 11210 700
rect 8573 663 8631 669
rect 8573 629 8585 663
rect 8619 629 8631 663
rect 8573 623 8631 629
rect 9493 663 9551 669
rect 9493 629 9505 663
rect 9539 660 9551 663
rect 10134 660 10140 672
rect 9539 632 10140 660
rect 9539 629 9551 632
rect 9493 623 9551 629
rect 10134 620 10140 632
rect 10192 620 10198 672
rect 11422 620 11428 672
rect 11480 620 11486 672
rect 11532 660 11560 700
rect 12161 663 12219 669
rect 12161 660 12173 663
rect 11532 632 12173 660
rect 12161 629 12173 632
rect 12207 629 12219 663
rect 12268 660 12296 700
rect 12342 688 12348 740
rect 12400 728 12406 740
rect 13096 728 13124 768
rect 13262 756 13268 808
rect 13320 796 13326 808
rect 13633 799 13691 805
rect 13633 796 13645 799
rect 13320 768 13645 796
rect 13320 756 13326 768
rect 13633 765 13645 768
rect 13679 765 13691 799
rect 13633 759 13691 765
rect 13906 756 13912 808
rect 13964 756 13970 808
rect 14090 756 14096 808
rect 14148 796 14154 808
rect 14277 799 14335 805
rect 14277 796 14289 799
rect 14148 768 14289 796
rect 14148 756 14154 768
rect 14277 765 14289 768
rect 14323 765 14335 799
rect 14277 759 14335 765
rect 13924 728 13952 756
rect 12400 700 13032 728
rect 13096 700 13952 728
rect 14292 728 14320 759
rect 14366 756 14372 808
rect 14424 796 14430 808
rect 14553 799 14611 805
rect 14553 796 14565 799
rect 14424 768 14565 796
rect 14424 756 14430 768
rect 14553 765 14565 768
rect 14599 765 14611 799
rect 14829 799 14887 805
rect 14829 796 14841 799
rect 14553 759 14611 765
rect 14660 768 14841 796
rect 14660 728 14688 768
rect 14829 765 14841 768
rect 14875 765 14887 799
rect 14829 759 14887 765
rect 15102 756 15108 808
rect 15160 756 15166 808
rect 15194 756 15200 808
rect 15252 796 15258 808
rect 15252 768 15516 796
rect 15252 756 15258 768
rect 15488 737 15516 768
rect 16850 756 16856 808
rect 16908 756 16914 808
rect 14292 700 14688 728
rect 14737 731 14795 737
rect 12400 688 12406 700
rect 12894 660 12900 672
rect 12268 632 12900 660
rect 12161 623 12219 629
rect 12894 620 12900 632
rect 12952 620 12958 672
rect 13004 660 13032 700
rect 14737 697 14749 731
rect 14783 697 14795 731
rect 14737 691 14795 697
rect 15473 731 15531 737
rect 15473 697 15485 731
rect 15519 697 15531 731
rect 15473 691 15531 697
rect 13725 663 13783 669
rect 13725 660 13737 663
rect 13004 632 13737 660
rect 13725 629 13737 632
rect 13771 629 13783 663
rect 14752 660 14780 691
rect 16206 688 16212 740
rect 16264 688 16270 740
rect 16114 660 16120 672
rect 14752 632 16120 660
rect 13725 623 13783 629
rect 16114 620 16120 632
rect 16172 620 16178 672
rect 552 570 17664 592
rect 552 518 4366 570
rect 4418 518 4430 570
rect 4482 518 4494 570
rect 4546 518 4558 570
rect 4610 518 4622 570
rect 4674 518 4686 570
rect 4738 518 10366 570
rect 10418 518 10430 570
rect 10482 518 10494 570
rect 10546 518 10558 570
rect 10610 518 10622 570
rect 10674 518 10686 570
rect 10738 518 16366 570
rect 16418 518 16430 570
rect 16482 518 16494 570
rect 16546 518 16558 570
rect 16610 518 16622 570
rect 16674 518 16686 570
rect 16738 518 17664 570
rect 552 496 17664 518
rect 5258 416 5264 468
rect 5316 416 5322 468
rect 6086 416 6092 468
rect 6144 456 6150 468
rect 12802 456 12808 468
rect 6144 428 12808 456
rect 6144 416 6150 428
rect 12802 416 12808 428
rect 12860 416 12866 468
rect 12894 416 12900 468
rect 12952 456 12958 468
rect 14366 456 14372 468
rect 12952 428 14372 456
rect 12952 416 12958 428
rect 14366 416 14372 428
rect 14424 416 14430 468
rect 14734 416 14740 468
rect 14792 416 14798 468
rect 16206 416 16212 468
rect 16264 416 16270 468
rect 5276 320 5304 416
rect 6362 348 6368 400
rect 6420 388 6426 400
rect 9674 388 9680 400
rect 6420 360 9680 388
rect 6420 348 6426 360
rect 9674 348 9680 360
rect 9732 348 9738 400
rect 11422 348 11428 400
rect 11480 388 11486 400
rect 14752 388 14780 416
rect 11480 360 14780 388
rect 11480 348 11486 360
rect 12526 320 12532 332
rect 5276 292 12532 320
rect 12526 280 12532 292
rect 12584 280 12590 332
rect 7834 212 7840 264
rect 7892 252 7898 264
rect 11974 252 11980 264
rect 7892 224 11980 252
rect 7892 212 7898 224
rect 11974 212 11980 224
rect 12032 252 12038 264
rect 14090 252 14096 264
rect 12032 224 14096 252
rect 12032 212 12038 224
rect 14090 212 14096 224
rect 14148 212 14154 264
rect 4154 144 4160 196
rect 4212 184 4218 196
rect 10042 184 10048 196
rect 4212 156 10048 184
rect 4212 144 4218 156
rect 10042 144 10048 156
rect 10100 144 10106 196
rect 11514 144 11520 196
rect 11572 184 11578 196
rect 16224 184 16252 416
rect 11572 156 16252 184
rect 11572 144 11578 156
<< via1 >>
rect 12808 17620 12860 17672
rect 14096 17620 14148 17672
rect 7288 17552 7340 17604
rect 11796 17552 11848 17604
rect 14832 17552 14884 17604
rect 2964 17484 3016 17536
rect 7196 17484 7248 17536
rect 11428 17484 11480 17536
rect 12992 17484 13044 17536
rect 13636 17484 13688 17536
rect 14556 17484 14608 17536
rect 1366 17382 1418 17434
rect 1430 17382 1482 17434
rect 1494 17382 1546 17434
rect 1558 17382 1610 17434
rect 1622 17382 1674 17434
rect 1686 17382 1738 17434
rect 7366 17382 7418 17434
rect 7430 17382 7482 17434
rect 7494 17382 7546 17434
rect 7558 17382 7610 17434
rect 7622 17382 7674 17434
rect 7686 17382 7738 17434
rect 13366 17382 13418 17434
rect 13430 17382 13482 17434
rect 13494 17382 13546 17434
rect 13558 17382 13610 17434
rect 13622 17382 13674 17434
rect 13686 17382 13738 17434
rect 1216 17323 1268 17332
rect 1216 17289 1225 17323
rect 1225 17289 1259 17323
rect 1259 17289 1268 17323
rect 1216 17280 1268 17289
rect 2044 17323 2096 17332
rect 2044 17289 2053 17323
rect 2053 17289 2087 17323
rect 2087 17289 2096 17323
rect 2044 17280 2096 17289
rect 2872 17280 2924 17332
rect 3700 17280 3752 17332
rect 4528 17280 4580 17332
rect 5356 17280 5408 17332
rect 6184 17280 6236 17332
rect 6736 17212 6788 17264
rect 7012 17280 7064 17332
rect 7840 17280 7892 17332
rect 8668 17280 8720 17332
rect 11152 17280 11204 17332
rect 2780 17076 2832 17128
rect 2964 17187 3016 17196
rect 2964 17153 2973 17187
rect 2973 17153 3007 17187
rect 3007 17153 3016 17187
rect 2964 17144 3016 17153
rect 3056 17144 3108 17196
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 7288 17144 7340 17196
rect 12992 17212 13044 17264
rect 4252 17119 4304 17128
rect 4252 17085 4261 17119
rect 4261 17085 4295 17119
rect 4295 17085 4304 17119
rect 4252 17076 4304 17085
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 7104 17119 7156 17128
rect 7104 17085 7113 17119
rect 7113 17085 7147 17119
rect 7147 17085 7156 17119
rect 7104 17076 7156 17085
rect 6460 17008 6512 17060
rect 6552 17051 6604 17060
rect 6552 17017 6561 17051
rect 6561 17017 6595 17051
rect 6595 17017 6604 17051
rect 6552 17008 6604 17017
rect 11612 17187 11664 17196
rect 11612 17153 11621 17187
rect 11621 17153 11655 17187
rect 11655 17153 11664 17187
rect 11612 17144 11664 17153
rect 3792 16940 3844 16992
rect 4252 16940 4304 16992
rect 5448 16940 5500 16992
rect 6368 16940 6420 16992
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 9036 17119 9088 17128
rect 9036 17085 9045 17119
rect 9045 17085 9079 17119
rect 9079 17085 9088 17119
rect 9036 17076 9088 17085
rect 9496 17076 9548 17128
rect 10324 17076 10376 17128
rect 10784 17119 10836 17128
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 10784 17076 10836 17085
rect 11428 17119 11480 17128
rect 11428 17085 11437 17119
rect 11437 17085 11471 17119
rect 11471 17085 11480 17119
rect 11428 17076 11480 17085
rect 11980 17076 12032 17128
rect 8576 16940 8628 16992
rect 9312 16983 9364 16992
rect 9312 16949 9321 16983
rect 9321 16949 9355 16983
rect 9355 16949 9364 16983
rect 9312 16940 9364 16949
rect 9404 16940 9456 16992
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 10140 16983 10192 16992
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 12716 17008 12768 17060
rect 13452 17076 13504 17128
rect 15292 17280 15344 17332
rect 16212 17280 16264 17332
rect 13820 17255 13872 17264
rect 13820 17221 13829 17255
rect 13829 17221 13863 17255
rect 13863 17221 13872 17255
rect 13820 17212 13872 17221
rect 16120 17144 16172 17196
rect 14096 17076 14148 17128
rect 14372 17076 14424 17128
rect 15384 17076 15436 17128
rect 12072 16940 12124 16992
rect 15108 17008 15160 17060
rect 15844 16940 15896 16992
rect 4366 16838 4418 16890
rect 4430 16838 4482 16890
rect 4494 16838 4546 16890
rect 4558 16838 4610 16890
rect 4622 16838 4674 16890
rect 4686 16838 4738 16890
rect 10366 16838 10418 16890
rect 10430 16838 10482 16890
rect 10494 16838 10546 16890
rect 10558 16838 10610 16890
rect 10622 16838 10674 16890
rect 10686 16838 10738 16890
rect 16366 16838 16418 16890
rect 16430 16838 16482 16890
rect 16494 16838 16546 16890
rect 16558 16838 16610 16890
rect 16622 16838 16674 16890
rect 16686 16838 16738 16890
rect 1676 16736 1728 16788
rect 3792 16736 3844 16788
rect 5540 16736 5592 16788
rect 6368 16779 6420 16788
rect 6368 16745 6377 16779
rect 6377 16745 6411 16779
rect 6411 16745 6420 16779
rect 6368 16736 6420 16745
rect 6552 16779 6604 16788
rect 6552 16745 6561 16779
rect 6561 16745 6595 16779
rect 6595 16745 6604 16779
rect 6552 16736 6604 16745
rect 9312 16736 9364 16788
rect 10140 16736 10192 16788
rect 12808 16736 12860 16788
rect 13728 16736 13780 16788
rect 14464 16736 14516 16788
rect 2780 16600 2832 16652
rect 2964 16600 3016 16652
rect 3056 16643 3108 16652
rect 3056 16609 3065 16643
rect 3065 16609 3099 16643
rect 3099 16609 3108 16643
rect 3056 16600 3108 16609
rect 3240 16600 3292 16652
rect 848 16532 900 16584
rect 4252 16532 4304 16584
rect 5908 16600 5960 16652
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 6276 16600 6328 16652
rect 9220 16668 9272 16720
rect 6184 16532 6236 16584
rect 2780 16396 2832 16448
rect 6368 16464 6420 16516
rect 4252 16396 4304 16448
rect 4620 16439 4672 16448
rect 4620 16405 4629 16439
rect 4629 16405 4663 16439
rect 4663 16405 4672 16439
rect 4620 16396 4672 16405
rect 5356 16439 5408 16448
rect 5356 16405 5365 16439
rect 5365 16405 5399 16439
rect 5399 16405 5408 16439
rect 5356 16396 5408 16405
rect 7012 16532 7064 16584
rect 7380 16464 7432 16516
rect 7012 16396 7064 16448
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 10048 16600 10100 16652
rect 11060 16600 11112 16652
rect 13176 16600 13228 16652
rect 13360 16600 13412 16652
rect 14372 16668 14424 16720
rect 8576 16396 8628 16448
rect 9220 16396 9272 16448
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 11520 16464 11572 16516
rect 13452 16532 13504 16584
rect 14556 16600 14608 16652
rect 16212 16736 16264 16788
rect 16028 16600 16080 16652
rect 14832 16532 14884 16584
rect 15844 16532 15896 16584
rect 12532 16396 12584 16448
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 14188 16396 14240 16448
rect 15016 16464 15068 16516
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 15568 16439 15620 16448
rect 15568 16405 15577 16439
rect 15577 16405 15611 16439
rect 15611 16405 15620 16439
rect 15568 16396 15620 16405
rect 16120 16439 16172 16448
rect 16120 16405 16129 16439
rect 16129 16405 16163 16439
rect 16163 16405 16172 16439
rect 16120 16396 16172 16405
rect 1366 16294 1418 16346
rect 1430 16294 1482 16346
rect 1494 16294 1546 16346
rect 1558 16294 1610 16346
rect 1622 16294 1674 16346
rect 1686 16294 1738 16346
rect 7366 16294 7418 16346
rect 7430 16294 7482 16346
rect 7494 16294 7546 16346
rect 7558 16294 7610 16346
rect 7622 16294 7674 16346
rect 7686 16294 7738 16346
rect 13366 16294 13418 16346
rect 13430 16294 13482 16346
rect 13494 16294 13546 16346
rect 13558 16294 13610 16346
rect 13622 16294 13674 16346
rect 13686 16294 13738 16346
rect 6736 16192 6788 16244
rect 6828 16192 6880 16244
rect 7196 16192 7248 16244
rect 7288 16235 7340 16244
rect 7288 16201 7297 16235
rect 7297 16201 7331 16235
rect 7331 16201 7340 16235
rect 7288 16192 7340 16201
rect 3240 16124 3292 16176
rect 848 15988 900 16040
rect 2780 16056 2832 16108
rect 3056 15988 3108 16040
rect 6460 16099 6512 16108
rect 6460 16065 6469 16099
rect 6469 16065 6503 16099
rect 6503 16065 6512 16099
rect 6460 16056 6512 16065
rect 9588 16192 9640 16244
rect 10784 16192 10836 16244
rect 11520 16192 11572 16244
rect 11152 16167 11204 16176
rect 11152 16133 11161 16167
rect 11161 16133 11195 16167
rect 11195 16133 11204 16167
rect 12348 16192 12400 16244
rect 13268 16192 13320 16244
rect 11152 16124 11204 16133
rect 12624 16167 12676 16176
rect 12624 16133 12633 16167
rect 12633 16133 12667 16167
rect 12667 16133 12676 16167
rect 12624 16124 12676 16133
rect 13084 16124 13136 16176
rect 5356 15988 5408 16040
rect 1492 15963 1544 15972
rect 1492 15929 1526 15963
rect 1526 15929 1544 15963
rect 1492 15920 1544 15929
rect 2596 15895 2648 15904
rect 2596 15861 2605 15895
rect 2605 15861 2639 15895
rect 2639 15861 2648 15895
rect 2596 15852 2648 15861
rect 3240 15895 3292 15904
rect 3240 15861 3249 15895
rect 3249 15861 3283 15895
rect 3283 15861 3292 15895
rect 3240 15852 3292 15861
rect 4620 15920 4672 15972
rect 5540 15920 5592 15972
rect 5632 15920 5684 15972
rect 7840 15988 7892 16040
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 11428 16056 11480 16108
rect 11612 16099 11664 16108
rect 11612 16065 11621 16099
rect 11621 16065 11655 16099
rect 11655 16065 11664 16099
rect 11612 16056 11664 16065
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 8208 15988 8260 16040
rect 8852 15920 8904 15972
rect 9404 15988 9456 16040
rect 10968 16031 11020 16040
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 10968 15988 11020 15997
rect 12716 16031 12768 16040
rect 12716 15997 12725 16031
rect 12725 15997 12759 16031
rect 12759 15997 12768 16031
rect 12716 15988 12768 15997
rect 9312 15920 9364 15972
rect 9680 15920 9732 15972
rect 11704 15963 11756 15972
rect 11704 15929 11713 15963
rect 11713 15929 11747 15963
rect 11747 15929 11756 15963
rect 11704 15920 11756 15929
rect 12808 15920 12860 15972
rect 13820 16056 13872 16108
rect 14464 16124 14516 16176
rect 15016 16099 15068 16108
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 15292 15988 15344 16040
rect 15568 15988 15620 16040
rect 14832 15920 14884 15972
rect 15200 15963 15252 15972
rect 15200 15929 15209 15963
rect 15209 15929 15243 15963
rect 15243 15929 15252 15963
rect 15200 15920 15252 15929
rect 15752 15920 15804 15972
rect 5724 15852 5776 15904
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 7472 15852 7524 15904
rect 8484 15852 8536 15904
rect 8944 15852 8996 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 13084 15852 13136 15904
rect 13912 15852 13964 15904
rect 14280 15852 14332 15904
rect 15476 15852 15528 15904
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 17040 15895 17092 15904
rect 17040 15861 17049 15895
rect 17049 15861 17083 15895
rect 17083 15861 17092 15895
rect 17040 15852 17092 15861
rect 4366 15750 4418 15802
rect 4430 15750 4482 15802
rect 4494 15750 4546 15802
rect 4558 15750 4610 15802
rect 4622 15750 4674 15802
rect 4686 15750 4738 15802
rect 10366 15750 10418 15802
rect 10430 15750 10482 15802
rect 10494 15750 10546 15802
rect 10558 15750 10610 15802
rect 10622 15750 10674 15802
rect 10686 15750 10738 15802
rect 16366 15750 16418 15802
rect 16430 15750 16482 15802
rect 16494 15750 16546 15802
rect 16558 15750 16610 15802
rect 16622 15750 16674 15802
rect 16686 15750 16738 15802
rect 1492 15648 1544 15700
rect 2044 15691 2096 15700
rect 2044 15657 2053 15691
rect 2053 15657 2087 15691
rect 2087 15657 2096 15691
rect 2044 15648 2096 15657
rect 2596 15648 2648 15700
rect 2044 15512 2096 15564
rect 2780 15580 2832 15632
rect 3056 15580 3108 15632
rect 2688 15376 2740 15428
rect 3240 15648 3292 15700
rect 3976 15648 4028 15700
rect 4896 15648 4948 15700
rect 4620 15623 4672 15632
rect 4620 15589 4629 15623
rect 4629 15589 4663 15623
rect 4663 15589 4672 15623
rect 4620 15580 4672 15589
rect 4988 15580 5040 15632
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 4160 15512 4212 15564
rect 4252 15512 4304 15564
rect 5264 15580 5316 15632
rect 5816 15648 5868 15700
rect 6276 15648 6328 15700
rect 6368 15648 6420 15700
rect 3884 15444 3936 15496
rect 5356 15512 5408 15564
rect 5724 15512 5776 15564
rect 6460 15580 6512 15632
rect 3792 15376 3844 15428
rect 6276 15555 6328 15564
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 6276 15512 6328 15521
rect 7472 15580 7524 15632
rect 7932 15648 7984 15700
rect 9312 15648 9364 15700
rect 10968 15648 11020 15700
rect 6644 15444 6696 15496
rect 7196 15444 7248 15496
rect 7288 15444 7340 15496
rect 8760 15512 8812 15564
rect 9128 15444 9180 15496
rect 10048 15512 10100 15564
rect 10232 15512 10284 15564
rect 13084 15648 13136 15700
rect 13176 15648 13228 15700
rect 15016 15691 15068 15700
rect 15016 15657 15025 15691
rect 15025 15657 15059 15691
rect 15059 15657 15068 15691
rect 15016 15648 15068 15657
rect 15568 15648 15620 15700
rect 15752 15648 15804 15700
rect 16120 15648 16172 15700
rect 17040 15648 17092 15700
rect 11980 15580 12032 15632
rect 12164 15580 12216 15632
rect 11520 15512 11572 15564
rect 12348 15512 12400 15564
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 12716 15512 12768 15564
rect 9956 15376 10008 15428
rect 11152 15376 11204 15428
rect 11612 15376 11664 15428
rect 13084 15512 13136 15564
rect 13912 15555 13964 15564
rect 13912 15521 13921 15555
rect 13921 15521 13955 15555
rect 13955 15521 13964 15555
rect 13912 15512 13964 15521
rect 14280 15512 14332 15564
rect 15200 15512 15252 15564
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 14556 15444 14608 15496
rect 16028 15444 16080 15496
rect 12808 15376 12860 15428
rect 13268 15376 13320 15428
rect 13452 15376 13504 15428
rect 13912 15376 13964 15428
rect 14188 15376 14240 15428
rect 15476 15376 15528 15428
rect 2872 15351 2924 15360
rect 2872 15317 2881 15351
rect 2881 15317 2915 15351
rect 2915 15317 2924 15351
rect 2872 15308 2924 15317
rect 3516 15308 3568 15360
rect 4160 15351 4212 15360
rect 4160 15317 4169 15351
rect 4169 15317 4203 15351
rect 4203 15317 4212 15351
rect 4160 15308 4212 15317
rect 4252 15308 4304 15360
rect 4804 15351 4856 15360
rect 4804 15317 4813 15351
rect 4813 15317 4847 15351
rect 4847 15317 4856 15351
rect 4804 15308 4856 15317
rect 4988 15308 5040 15360
rect 5172 15308 5224 15360
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 7932 15308 7984 15360
rect 8576 15308 8628 15360
rect 8852 15308 8904 15360
rect 10140 15308 10192 15360
rect 12716 15308 12768 15360
rect 12992 15308 13044 15360
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 15108 15308 15160 15360
rect 15936 15308 15988 15360
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 1366 15206 1418 15258
rect 1430 15206 1482 15258
rect 1494 15206 1546 15258
rect 1558 15206 1610 15258
rect 1622 15206 1674 15258
rect 1686 15206 1738 15258
rect 7366 15206 7418 15258
rect 7430 15206 7482 15258
rect 7494 15206 7546 15258
rect 7558 15206 7610 15258
rect 7622 15206 7674 15258
rect 7686 15206 7738 15258
rect 13366 15206 13418 15258
rect 13430 15206 13482 15258
rect 13494 15206 13546 15258
rect 13558 15206 13610 15258
rect 13622 15206 13674 15258
rect 13686 15206 13738 15258
rect 2688 15147 2740 15156
rect 2688 15113 2697 15147
rect 2697 15113 2731 15147
rect 2731 15113 2740 15147
rect 2688 15104 2740 15113
rect 2964 15104 3016 15156
rect 3516 15104 3568 15156
rect 848 14943 900 14952
rect 848 14909 857 14943
rect 857 14909 891 14943
rect 891 14909 900 14943
rect 848 14900 900 14909
rect 1400 14832 1452 14884
rect 2044 14764 2096 14816
rect 3148 15036 3200 15088
rect 3516 15011 3568 15020
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 3516 14968 3568 14977
rect 5172 15104 5224 15156
rect 6000 15104 6052 15156
rect 6552 15104 6604 15156
rect 7656 15104 7708 15156
rect 4252 15036 4304 15088
rect 3424 14943 3476 14952
rect 3424 14909 3433 14943
rect 3433 14909 3467 14943
rect 3467 14909 3476 14943
rect 3424 14900 3476 14909
rect 3976 14900 4028 14952
rect 4160 14900 4212 14952
rect 4896 15011 4948 15020
rect 4896 14977 4905 15011
rect 4905 14977 4939 15011
rect 4939 14977 4948 15011
rect 4896 14968 4948 14977
rect 5540 14968 5592 15020
rect 6092 14968 6144 15020
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 6644 15036 6696 15088
rect 7380 14968 7432 15020
rect 3792 14832 3844 14884
rect 5264 14900 5316 14952
rect 5816 14900 5868 14952
rect 6276 14900 6328 14952
rect 6552 14900 6604 14952
rect 6736 14900 6788 14952
rect 6920 14900 6972 14952
rect 8024 15036 8076 15088
rect 7748 14900 7800 14952
rect 8576 15147 8628 15156
rect 8576 15113 8585 15147
rect 8585 15113 8619 15147
rect 8619 15113 8628 15147
rect 8576 15104 8628 15113
rect 8760 15147 8812 15156
rect 8760 15113 8769 15147
rect 8769 15113 8803 15147
rect 8803 15113 8812 15147
rect 8760 15104 8812 15113
rect 8392 15036 8444 15088
rect 13452 15104 13504 15156
rect 13912 15104 13964 15156
rect 15016 15104 15068 15156
rect 15384 15104 15436 15156
rect 11796 15036 11848 15088
rect 12900 15036 12952 15088
rect 10048 14968 10100 15020
rect 8576 14943 8628 14952
rect 8576 14909 8585 14943
rect 8585 14909 8619 14943
rect 8619 14909 8628 14943
rect 8576 14900 8628 14909
rect 8852 14900 8904 14952
rect 9588 14900 9640 14952
rect 6368 14832 6420 14884
rect 8208 14832 8260 14884
rect 3700 14764 3752 14816
rect 4620 14764 4672 14816
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 6000 14764 6052 14816
rect 6552 14764 6604 14816
rect 7104 14764 7156 14816
rect 7380 14807 7432 14816
rect 7380 14773 7389 14807
rect 7389 14773 7423 14807
rect 7423 14773 7432 14807
rect 7380 14764 7432 14773
rect 9864 14764 9916 14816
rect 14556 15036 14608 15088
rect 14740 15036 14792 15088
rect 13268 14968 13320 15020
rect 14188 14968 14240 15020
rect 14372 14968 14424 15020
rect 11888 14900 11940 14952
rect 12256 14900 12308 14952
rect 11428 14764 11480 14816
rect 12348 14832 12400 14884
rect 12624 14875 12676 14884
rect 12624 14841 12642 14875
rect 12642 14841 12676 14875
rect 12624 14832 12676 14841
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 13452 14832 13504 14884
rect 14004 14900 14056 14952
rect 14556 14900 14608 14952
rect 13912 14832 13964 14884
rect 11704 14764 11756 14816
rect 13084 14764 13136 14816
rect 14096 14764 14148 14816
rect 17040 14764 17092 14816
rect 4366 14662 4418 14714
rect 4430 14662 4482 14714
rect 4494 14662 4546 14714
rect 4558 14662 4610 14714
rect 4622 14662 4674 14714
rect 4686 14662 4738 14714
rect 10366 14662 10418 14714
rect 10430 14662 10482 14714
rect 10494 14662 10546 14714
rect 10558 14662 10610 14714
rect 10622 14662 10674 14714
rect 10686 14662 10738 14714
rect 16366 14662 16418 14714
rect 16430 14662 16482 14714
rect 16494 14662 16546 14714
rect 16558 14662 16610 14714
rect 16622 14662 16674 14714
rect 16686 14662 16738 14714
rect 1400 14560 1452 14612
rect 2872 14560 2924 14612
rect 3516 14560 3568 14612
rect 2044 14467 2096 14476
rect 2044 14433 2053 14467
rect 2053 14433 2087 14467
rect 2087 14433 2096 14467
rect 2044 14424 2096 14433
rect 2504 14424 2556 14476
rect 2688 14467 2740 14476
rect 2688 14433 2697 14467
rect 2697 14433 2731 14467
rect 2731 14433 2740 14467
rect 2688 14424 2740 14433
rect 1768 14356 1820 14408
rect 2596 14399 2648 14408
rect 2596 14365 2605 14399
rect 2605 14365 2639 14399
rect 2639 14365 2648 14399
rect 2596 14356 2648 14365
rect 2964 14424 3016 14476
rect 3792 14424 3844 14476
rect 5080 14560 5132 14612
rect 5264 14560 5316 14612
rect 4528 14535 4580 14544
rect 4528 14501 4537 14535
rect 4537 14501 4571 14535
rect 4571 14501 4580 14535
rect 4528 14492 4580 14501
rect 5540 14492 5592 14544
rect 5632 14492 5684 14544
rect 6276 14492 6328 14544
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 5080 14424 5132 14476
rect 4896 14356 4948 14408
rect 5816 14424 5868 14476
rect 7380 14560 7432 14612
rect 7656 14560 7708 14612
rect 7932 14492 7984 14544
rect 8576 14560 8628 14612
rect 8760 14560 8812 14612
rect 9220 14560 9272 14612
rect 12164 14560 12216 14612
rect 12348 14560 12400 14612
rect 6368 14356 6420 14408
rect 6828 14356 6880 14408
rect 8300 14424 8352 14476
rect 8392 14424 8444 14476
rect 9128 14424 9180 14476
rect 8668 14356 8720 14408
rect 8852 14356 8904 14408
rect 9496 14467 9548 14476
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 9956 14424 10008 14476
rect 10600 14467 10652 14476
rect 10600 14433 10609 14467
rect 10609 14433 10643 14467
rect 10643 14433 10652 14467
rect 10600 14424 10652 14433
rect 11888 14492 11940 14544
rect 11336 14424 11388 14476
rect 12348 14424 12400 14476
rect 10876 14356 10928 14408
rect 9772 14288 9824 14340
rect 9864 14288 9916 14340
rect 11612 14356 11664 14408
rect 1860 14220 1912 14272
rect 2964 14220 3016 14272
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 5816 14263 5868 14272
rect 5816 14229 5825 14263
rect 5825 14229 5859 14263
rect 5859 14229 5868 14263
rect 5816 14220 5868 14229
rect 7840 14220 7892 14272
rect 12532 14356 12584 14408
rect 13820 14424 13872 14476
rect 13912 14467 13964 14476
rect 13912 14433 13921 14467
rect 13921 14433 13955 14467
rect 13955 14433 13964 14467
rect 13912 14424 13964 14433
rect 14004 14467 14056 14476
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 12900 14356 12952 14408
rect 14372 14424 14424 14476
rect 15936 14467 15988 14476
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 11060 14220 11112 14272
rect 11152 14263 11204 14272
rect 11152 14229 11161 14263
rect 11161 14229 11195 14263
rect 11195 14229 11204 14263
rect 11152 14220 11204 14229
rect 11520 14220 11572 14272
rect 11704 14263 11756 14272
rect 11704 14229 11713 14263
rect 11713 14229 11747 14263
rect 11747 14229 11756 14263
rect 11704 14220 11756 14229
rect 11796 14220 11848 14272
rect 14004 14288 14056 14340
rect 15936 14433 15945 14467
rect 15945 14433 15979 14467
rect 15979 14433 15988 14467
rect 15936 14424 15988 14433
rect 15752 14331 15804 14340
rect 15752 14297 15761 14331
rect 15761 14297 15795 14331
rect 15795 14297 15804 14331
rect 15752 14288 15804 14297
rect 16028 14288 16080 14340
rect 12440 14220 12492 14272
rect 12716 14263 12768 14272
rect 12716 14229 12725 14263
rect 12725 14229 12759 14263
rect 12759 14229 12768 14263
rect 12716 14220 12768 14229
rect 1366 14118 1418 14170
rect 1430 14118 1482 14170
rect 1494 14118 1546 14170
rect 1558 14118 1610 14170
rect 1622 14118 1674 14170
rect 1686 14118 1738 14170
rect 7366 14118 7418 14170
rect 7430 14118 7482 14170
rect 7494 14118 7546 14170
rect 7558 14118 7610 14170
rect 7622 14118 7674 14170
rect 7686 14118 7738 14170
rect 13366 14118 13418 14170
rect 13430 14118 13482 14170
rect 13494 14118 13546 14170
rect 13558 14118 13610 14170
rect 13622 14118 13674 14170
rect 13686 14118 13738 14170
rect 3424 14016 3476 14068
rect 4988 14016 5040 14068
rect 5356 14016 5408 14068
rect 1860 13948 1912 14000
rect 2504 13880 2556 13932
rect 3608 13880 3660 13932
rect 4344 13880 4396 13932
rect 2596 13812 2648 13864
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 3884 13812 3936 13864
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 4068 13855 4120 13864
rect 4068 13821 4077 13855
rect 4077 13821 4111 13855
rect 4111 13821 4120 13855
rect 4068 13812 4120 13821
rect 4252 13855 4304 13864
rect 4252 13821 4262 13855
rect 4262 13821 4296 13855
rect 4296 13821 4304 13855
rect 4252 13812 4304 13821
rect 4804 13812 4856 13864
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 5816 14016 5868 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 6828 14016 6880 14068
rect 7196 14059 7248 14068
rect 7196 14025 7205 14059
rect 7205 14025 7239 14059
rect 7239 14025 7248 14059
rect 7196 14016 7248 14025
rect 6460 13948 6512 14000
rect 8024 14016 8076 14068
rect 6092 13880 6144 13932
rect 6276 13855 6328 13864
rect 6276 13821 6285 13855
rect 6285 13821 6319 13855
rect 6319 13821 6328 13855
rect 6276 13812 6328 13821
rect 7288 13880 7340 13932
rect 8208 13880 8260 13932
rect 8300 13880 8352 13932
rect 8760 13880 8812 13932
rect 4252 13676 4304 13728
rect 6000 13676 6052 13728
rect 6368 13744 6420 13796
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 7748 13855 7800 13864
rect 7748 13821 7757 13855
rect 7757 13821 7791 13855
rect 7791 13821 7800 13855
rect 7748 13812 7800 13821
rect 7932 13812 7984 13864
rect 9220 14016 9272 14068
rect 10600 14016 10652 14068
rect 11796 14016 11848 14068
rect 10968 13948 11020 14000
rect 11244 13948 11296 14000
rect 12164 13948 12216 14000
rect 12256 13948 12308 14000
rect 9496 13812 9548 13864
rect 9588 13812 9640 13864
rect 9128 13744 9180 13796
rect 9680 13787 9732 13796
rect 9680 13753 9689 13787
rect 9689 13753 9723 13787
rect 9723 13753 9732 13787
rect 9680 13744 9732 13753
rect 10048 13744 10100 13796
rect 12072 13880 12124 13932
rect 11060 13787 11112 13796
rect 8392 13676 8444 13728
rect 8760 13676 8812 13728
rect 9864 13676 9916 13728
rect 10232 13676 10284 13728
rect 11060 13753 11087 13787
rect 11087 13753 11112 13787
rect 11060 13744 11112 13753
rect 11336 13744 11388 13796
rect 11612 13744 11664 13796
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 13728 14016 13780 14068
rect 14096 14016 14148 14068
rect 14004 13948 14056 14000
rect 13912 13880 13964 13932
rect 12532 13855 12584 13864
rect 12532 13821 12541 13855
rect 12541 13821 12575 13855
rect 12575 13821 12584 13855
rect 12532 13812 12584 13821
rect 12624 13812 12676 13864
rect 14372 13855 14424 13864
rect 14372 13821 14381 13855
rect 14381 13821 14415 13855
rect 14415 13821 14424 13855
rect 14372 13812 14424 13821
rect 10600 13676 10652 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 13820 13676 13872 13728
rect 14096 13787 14148 13796
rect 14096 13753 14105 13787
rect 14105 13753 14139 13787
rect 14139 13753 14148 13787
rect 14096 13744 14148 13753
rect 15752 13812 15804 13864
rect 15936 13948 15988 14000
rect 17132 13948 17184 14000
rect 16212 13880 16264 13932
rect 16396 13923 16448 13932
rect 16396 13889 16405 13923
rect 16405 13889 16439 13923
rect 16439 13889 16448 13923
rect 16396 13880 16448 13889
rect 16764 13812 16816 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 14740 13744 14792 13796
rect 17040 13744 17092 13796
rect 17408 13676 17460 13728
rect 4366 13574 4418 13626
rect 4430 13574 4482 13626
rect 4494 13574 4546 13626
rect 4558 13574 4610 13626
rect 4622 13574 4674 13626
rect 4686 13574 4738 13626
rect 10366 13574 10418 13626
rect 10430 13574 10482 13626
rect 10494 13574 10546 13626
rect 10558 13574 10610 13626
rect 10622 13574 10674 13626
rect 10686 13574 10738 13626
rect 16366 13574 16418 13626
rect 16430 13574 16482 13626
rect 16494 13574 16546 13626
rect 16558 13574 16610 13626
rect 16622 13574 16674 13626
rect 16686 13574 16738 13626
rect 2136 13472 2188 13524
rect 2596 13404 2648 13456
rect 3516 13472 3568 13524
rect 3608 13515 3660 13524
rect 3608 13481 3617 13515
rect 3617 13481 3651 13515
rect 3651 13481 3660 13515
rect 3608 13472 3660 13481
rect 3976 13472 4028 13524
rect 4344 13472 4396 13524
rect 1216 13379 1268 13388
rect 1216 13345 1250 13379
rect 1250 13345 1268 13379
rect 1216 13336 1268 13345
rect 848 13268 900 13320
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 2504 13132 2556 13184
rect 3240 13132 3292 13184
rect 6368 13404 6420 13456
rect 6920 13472 6972 13524
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 9128 13472 9180 13524
rect 10048 13472 10100 13524
rect 10876 13472 10928 13524
rect 12072 13472 12124 13524
rect 6828 13447 6880 13456
rect 6828 13413 6837 13447
rect 6837 13413 6871 13447
rect 6871 13413 6880 13447
rect 6828 13404 6880 13413
rect 7380 13404 7432 13456
rect 7932 13404 7984 13456
rect 4344 13336 4396 13388
rect 4620 13336 4672 13388
rect 4896 13336 4948 13388
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 5632 13379 5684 13388
rect 5632 13345 5641 13379
rect 5641 13345 5675 13379
rect 5675 13345 5684 13379
rect 5632 13336 5684 13345
rect 6092 13336 6144 13388
rect 6920 13379 6972 13388
rect 6920 13345 6929 13379
rect 6929 13345 6963 13379
rect 6963 13345 6972 13379
rect 6920 13336 6972 13345
rect 8392 13404 8444 13456
rect 9588 13404 9640 13456
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 8668 13336 8720 13388
rect 9404 13336 9456 13388
rect 7840 13268 7892 13320
rect 9772 13268 9824 13320
rect 4988 13200 5040 13252
rect 5724 13200 5776 13252
rect 9680 13200 9732 13252
rect 10232 13404 10284 13456
rect 12624 13404 12676 13456
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 12900 13472 12952 13524
rect 13084 13472 13136 13524
rect 13360 13447 13412 13456
rect 13360 13413 13369 13447
rect 13369 13413 13403 13447
rect 13403 13413 13412 13447
rect 13360 13404 13412 13413
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 14004 13404 14056 13456
rect 17132 13472 17184 13524
rect 10600 13336 10652 13388
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 11520 13336 11572 13388
rect 12164 13336 12216 13388
rect 13820 13336 13872 13388
rect 14924 13336 14976 13388
rect 15568 13336 15620 13388
rect 15936 13379 15988 13388
rect 15936 13345 15945 13379
rect 15945 13345 15979 13379
rect 15979 13345 15988 13379
rect 15936 13336 15988 13345
rect 16028 13336 16080 13388
rect 16396 13336 16448 13388
rect 10232 13200 10284 13252
rect 10324 13200 10376 13252
rect 5172 13132 5224 13184
rect 7932 13132 7984 13184
rect 9864 13132 9916 13184
rect 10600 13132 10652 13184
rect 10692 13132 10744 13184
rect 11428 13268 11480 13320
rect 14556 13268 14608 13320
rect 16764 13379 16816 13388
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 16764 13336 16816 13345
rect 14740 13200 14792 13252
rect 15292 13200 15344 13252
rect 13176 13132 13228 13184
rect 15384 13132 15436 13184
rect 15752 13132 15804 13184
rect 17132 13175 17184 13184
rect 17132 13141 17141 13175
rect 17141 13141 17175 13175
rect 17175 13141 17184 13175
rect 17132 13132 17184 13141
rect 1366 13030 1418 13082
rect 1430 13030 1482 13082
rect 1494 13030 1546 13082
rect 1558 13030 1610 13082
rect 1622 13030 1674 13082
rect 1686 13030 1738 13082
rect 7366 13030 7418 13082
rect 7430 13030 7482 13082
rect 7494 13030 7546 13082
rect 7558 13030 7610 13082
rect 7622 13030 7674 13082
rect 7686 13030 7738 13082
rect 13366 13030 13418 13082
rect 13430 13030 13482 13082
rect 13494 13030 13546 13082
rect 13558 13030 13610 13082
rect 13622 13030 13674 13082
rect 13686 13030 13738 13082
rect 1216 12928 1268 12980
rect 1768 12928 1820 12980
rect 2872 12971 2924 12980
rect 2872 12937 2881 12971
rect 2881 12937 2915 12971
rect 2915 12937 2924 12971
rect 2872 12928 2924 12937
rect 1676 12860 1728 12912
rect 5356 12928 5408 12980
rect 5908 12928 5960 12980
rect 7012 12928 7064 12980
rect 8392 12928 8444 12980
rect 9496 12928 9548 12980
rect 9680 12928 9732 12980
rect 4620 12903 4672 12912
rect 4620 12869 4629 12903
rect 4629 12869 4663 12903
rect 4663 12869 4672 12903
rect 4620 12860 4672 12869
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 11796 12860 11848 12912
rect 9772 12792 9824 12844
rect 11428 12792 11480 12844
rect 1952 12724 2004 12776
rect 2412 12724 2464 12776
rect 5080 12767 5132 12776
rect 5080 12733 5089 12767
rect 5089 12733 5123 12767
rect 5123 12733 5132 12767
rect 5080 12724 5132 12733
rect 2596 12656 2648 12708
rect 2780 12588 2832 12640
rect 2964 12588 3016 12640
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 3516 12699 3568 12708
rect 3516 12665 3550 12699
rect 3550 12665 3568 12699
rect 3516 12656 3568 12665
rect 3608 12656 3660 12708
rect 4160 12656 4212 12708
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 6276 12724 6328 12776
rect 6184 12656 6236 12708
rect 7104 12724 7156 12776
rect 8392 12724 8444 12776
rect 9588 12724 9640 12776
rect 10692 12767 10744 12776
rect 6736 12656 6788 12708
rect 6828 12656 6880 12708
rect 8300 12656 8352 12708
rect 7012 12588 7064 12640
rect 7840 12588 7892 12640
rect 9404 12656 9456 12708
rect 10692 12733 10701 12767
rect 10701 12733 10735 12767
rect 10735 12733 10744 12767
rect 10692 12724 10744 12733
rect 11980 12792 12032 12844
rect 12164 12792 12216 12844
rect 12532 12792 12584 12844
rect 9956 12699 10008 12708
rect 9956 12665 9965 12699
rect 9965 12665 9999 12699
rect 9999 12665 10008 12699
rect 9956 12656 10008 12665
rect 8668 12588 8720 12640
rect 9128 12588 9180 12640
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 10324 12699 10376 12708
rect 10324 12665 10333 12699
rect 10333 12665 10367 12699
rect 10367 12665 10376 12699
rect 10324 12656 10376 12665
rect 10876 12656 10928 12708
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 13268 12928 13320 12980
rect 14556 12928 14608 12980
rect 16856 12928 16908 12980
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 12624 12767 12676 12776
rect 12624 12733 12633 12767
rect 12633 12733 12667 12767
rect 12667 12733 12676 12767
rect 12624 12724 12676 12733
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 14004 12724 14056 12776
rect 14280 12724 14332 12776
rect 14924 12724 14976 12776
rect 15200 12724 15252 12776
rect 17132 12724 17184 12776
rect 13084 12656 13136 12708
rect 14188 12656 14240 12708
rect 15292 12656 15344 12708
rect 15476 12656 15528 12708
rect 16396 12656 16448 12708
rect 9496 12588 9548 12597
rect 11796 12588 11848 12640
rect 12624 12588 12676 12640
rect 12808 12588 12860 12640
rect 13636 12588 13688 12640
rect 14832 12588 14884 12640
rect 15936 12588 15988 12640
rect 4366 12486 4418 12538
rect 4430 12486 4482 12538
rect 4494 12486 4546 12538
rect 4558 12486 4610 12538
rect 4622 12486 4674 12538
rect 4686 12486 4738 12538
rect 10366 12486 10418 12538
rect 10430 12486 10482 12538
rect 10494 12486 10546 12538
rect 10558 12486 10610 12538
rect 10622 12486 10674 12538
rect 10686 12486 10738 12538
rect 16366 12486 16418 12538
rect 16430 12486 16482 12538
rect 16494 12486 16546 12538
rect 16558 12486 16610 12538
rect 16622 12486 16674 12538
rect 16686 12486 16738 12538
rect 2964 12384 3016 12436
rect 3516 12384 3568 12436
rect 4160 12384 4212 12436
rect 6828 12384 6880 12436
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 8392 12427 8444 12436
rect 8392 12393 8401 12427
rect 8401 12393 8435 12427
rect 8435 12393 8444 12427
rect 8392 12384 8444 12393
rect 12532 12384 12584 12436
rect 13268 12384 13320 12436
rect 1124 12291 1176 12300
rect 1124 12257 1158 12291
rect 1158 12257 1176 12291
rect 1124 12248 1176 12257
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 2964 12248 3016 12257
rect 5724 12316 5776 12368
rect 848 12223 900 12232
rect 848 12189 857 12223
rect 857 12189 891 12223
rect 891 12189 900 12223
rect 848 12180 900 12189
rect 2228 12180 2280 12232
rect 4252 12180 4304 12232
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 6460 12316 6512 12368
rect 6736 12248 6788 12300
rect 7288 12248 7340 12300
rect 2136 12044 2188 12096
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 4988 12112 5040 12164
rect 6644 12180 6696 12232
rect 7104 12112 7156 12164
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 8300 12316 8352 12368
rect 11244 12316 11296 12368
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 9312 12248 9364 12300
rect 10968 12248 11020 12300
rect 11704 12291 11756 12300
rect 11704 12257 11738 12291
rect 11738 12257 11756 12291
rect 11704 12248 11756 12257
rect 8116 12112 8168 12164
rect 8576 12112 8628 12164
rect 8944 12112 8996 12164
rect 9404 12112 9456 12164
rect 4896 12044 4948 12096
rect 6552 12044 6604 12096
rect 7196 12044 7248 12096
rect 7748 12044 7800 12096
rect 7932 12044 7984 12096
rect 8484 12044 8536 12096
rect 11336 12044 11388 12096
rect 12532 12044 12584 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 13636 12316 13688 12368
rect 14556 12316 14608 12368
rect 15476 12384 15528 12436
rect 16948 12384 17000 12436
rect 17224 12384 17276 12436
rect 13820 12248 13872 12300
rect 13912 12291 13964 12300
rect 13912 12257 13921 12291
rect 13921 12257 13955 12291
rect 13955 12257 13964 12291
rect 13912 12248 13964 12257
rect 14280 12155 14332 12164
rect 14280 12121 14289 12155
rect 14289 12121 14323 12155
rect 14323 12121 14332 12155
rect 14280 12112 14332 12121
rect 14924 12044 14976 12096
rect 15200 12044 15252 12096
rect 17040 12180 17092 12232
rect 17408 12180 17460 12232
rect 16212 12044 16264 12096
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 1366 11942 1418 11994
rect 1430 11942 1482 11994
rect 1494 11942 1546 11994
rect 1558 11942 1610 11994
rect 1622 11942 1674 11994
rect 1686 11942 1738 11994
rect 7366 11942 7418 11994
rect 7430 11942 7482 11994
rect 7494 11942 7546 11994
rect 7558 11942 7610 11994
rect 7622 11942 7674 11994
rect 7686 11942 7738 11994
rect 13366 11942 13418 11994
rect 13430 11942 13482 11994
rect 13494 11942 13546 11994
rect 13558 11942 13610 11994
rect 13622 11942 13674 11994
rect 13686 11942 13738 11994
rect 1124 11840 1176 11892
rect 1768 11883 1820 11892
rect 1768 11849 1777 11883
rect 1777 11849 1811 11883
rect 1811 11849 1820 11883
rect 1768 11840 1820 11849
rect 2688 11840 2740 11892
rect 3148 11840 3200 11892
rect 7288 11840 7340 11892
rect 7840 11840 7892 11892
rect 2596 11772 2648 11824
rect 3332 11772 3384 11824
rect 2044 11636 2096 11688
rect 2412 11679 2464 11688
rect 2412 11645 2421 11679
rect 2421 11645 2455 11679
rect 2455 11645 2464 11679
rect 2412 11636 2464 11645
rect 6184 11772 6236 11824
rect 9404 11883 9456 11892
rect 9404 11849 9413 11883
rect 9413 11849 9447 11883
rect 9447 11849 9456 11883
rect 9404 11840 9456 11849
rect 11704 11840 11756 11892
rect 13084 11840 13136 11892
rect 3608 11704 3660 11756
rect 5908 11704 5960 11756
rect 6368 11704 6420 11756
rect 6644 11704 6696 11756
rect 9312 11772 9364 11824
rect 1952 11543 2004 11552
rect 1952 11509 1979 11543
rect 1979 11509 2004 11543
rect 1952 11500 2004 11509
rect 3976 11636 4028 11688
rect 4344 11679 4396 11688
rect 4344 11645 4353 11679
rect 4353 11645 4387 11679
rect 4387 11645 4396 11679
rect 4344 11636 4396 11645
rect 4804 11636 4856 11688
rect 3424 11568 3476 11620
rect 6460 11636 6512 11688
rect 7012 11636 7064 11688
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 7748 11679 7800 11688
rect 7748 11645 7757 11679
rect 7757 11645 7791 11679
rect 7791 11645 7800 11679
rect 7748 11636 7800 11645
rect 8024 11636 8076 11688
rect 6184 11568 6236 11620
rect 4160 11500 4212 11552
rect 4988 11500 5040 11552
rect 5356 11500 5408 11552
rect 7380 11500 7432 11552
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 9128 11568 9180 11620
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 9496 11636 9548 11688
rect 9588 11611 9640 11620
rect 9588 11577 9597 11611
rect 9597 11577 9631 11611
rect 9631 11577 9640 11611
rect 9588 11568 9640 11577
rect 9956 11636 10008 11688
rect 10232 11704 10284 11756
rect 11244 11679 11296 11688
rect 11244 11645 11253 11679
rect 11253 11645 11287 11679
rect 11287 11645 11296 11679
rect 13176 11772 13228 11824
rect 15568 11840 15620 11892
rect 14832 11772 14884 11824
rect 11244 11636 11296 11645
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 12808 11704 12860 11756
rect 12072 11568 12124 11620
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 10140 11500 10192 11552
rect 11060 11500 11112 11552
rect 11520 11500 11572 11552
rect 13084 11636 13136 11688
rect 13820 11704 13872 11756
rect 12348 11500 12400 11552
rect 12716 11500 12768 11552
rect 13728 11500 13780 11552
rect 14740 11636 14792 11688
rect 14924 11636 14976 11688
rect 14372 11543 14424 11552
rect 14372 11509 14394 11543
rect 14394 11509 14424 11543
rect 14372 11500 14424 11509
rect 15108 11568 15160 11620
rect 16120 11568 16172 11620
rect 4366 11398 4418 11450
rect 4430 11398 4482 11450
rect 4494 11398 4546 11450
rect 4558 11398 4610 11450
rect 4622 11398 4674 11450
rect 4686 11398 4738 11450
rect 10366 11398 10418 11450
rect 10430 11398 10482 11450
rect 10494 11398 10546 11450
rect 10558 11398 10610 11450
rect 10622 11398 10674 11450
rect 10686 11398 10738 11450
rect 16366 11398 16418 11450
rect 16430 11398 16482 11450
rect 16494 11398 16546 11450
rect 16558 11398 16610 11450
rect 16622 11398 16674 11450
rect 16686 11398 16738 11450
rect 1768 11296 1820 11348
rect 2412 11296 2464 11348
rect 4344 11296 4396 11348
rect 848 11228 900 11280
rect 1952 11160 2004 11212
rect 4068 11228 4120 11280
rect 4160 11228 4212 11280
rect 4804 11296 4856 11348
rect 6920 11296 6972 11348
rect 7932 11296 7984 11348
rect 8024 11339 8076 11348
rect 8024 11305 8033 11339
rect 8033 11305 8067 11339
rect 8067 11305 8076 11339
rect 8024 11296 8076 11305
rect 8392 11296 8444 11348
rect 8576 11296 8628 11348
rect 9036 11296 9088 11348
rect 9588 11296 9640 11348
rect 10232 11296 10284 11348
rect 11244 11296 11296 11348
rect 11704 11296 11756 11348
rect 12348 11296 12400 11348
rect 12900 11296 12952 11348
rect 13084 11296 13136 11348
rect 13912 11296 13964 11348
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 16212 11296 16264 11348
rect 16948 11296 17000 11348
rect 2320 11092 2372 11144
rect 2320 10999 2372 11008
rect 2320 10965 2329 10999
rect 2329 10965 2363 10999
rect 2363 10965 2372 10999
rect 2320 10956 2372 10965
rect 3608 11160 3660 11212
rect 4160 11092 4212 11144
rect 4804 11160 4856 11212
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 5080 11160 5132 11212
rect 5816 11203 5868 11212
rect 5172 11024 5224 11076
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 5724 11092 5776 11144
rect 6368 11092 6420 11144
rect 6644 11160 6696 11212
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 6828 11160 6880 11212
rect 7380 11203 7432 11212
rect 7380 11169 7389 11203
rect 7389 11169 7423 11203
rect 7423 11169 7432 11203
rect 7380 11160 7432 11169
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 9220 11160 9272 11212
rect 11336 11228 11388 11280
rect 14740 11228 14792 11280
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 12716 11160 12768 11212
rect 14096 11160 14148 11212
rect 14924 11160 14976 11212
rect 15108 11160 15160 11212
rect 8116 11092 8168 11144
rect 3332 10956 3384 11008
rect 3700 10956 3752 11008
rect 5356 10956 5408 11008
rect 5540 10956 5592 11008
rect 6460 10956 6512 11008
rect 6736 10956 6788 11008
rect 8576 11024 8628 11076
rect 9312 11092 9364 11144
rect 9956 11092 10008 11144
rect 11060 11092 11112 11144
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 14556 11092 14608 11144
rect 15016 11092 15068 11144
rect 13636 11024 13688 11076
rect 14280 11024 14332 11076
rect 9588 10999 9640 11008
rect 9588 10965 9597 10999
rect 9597 10965 9631 10999
rect 9631 10965 9640 10999
rect 9588 10956 9640 10965
rect 10140 10956 10192 11008
rect 11152 10956 11204 11008
rect 12072 10956 12124 11008
rect 14556 10956 14608 11008
rect 16304 11203 16356 11212
rect 16304 11169 16313 11203
rect 16313 11169 16347 11203
rect 16347 11169 16356 11203
rect 16304 11160 16356 11169
rect 16580 11203 16632 11212
rect 16580 11169 16589 11203
rect 16589 11169 16623 11203
rect 16623 11169 16632 11203
rect 16580 11160 16632 11169
rect 17500 11024 17552 11076
rect 15844 10999 15896 11008
rect 15844 10965 15853 10999
rect 15853 10965 15887 10999
rect 15887 10965 15896 10999
rect 15844 10956 15896 10965
rect 1366 10854 1418 10906
rect 1430 10854 1482 10906
rect 1494 10854 1546 10906
rect 1558 10854 1610 10906
rect 1622 10854 1674 10906
rect 1686 10854 1738 10906
rect 7366 10854 7418 10906
rect 7430 10854 7482 10906
rect 7494 10854 7546 10906
rect 7558 10854 7610 10906
rect 7622 10854 7674 10906
rect 7686 10854 7738 10906
rect 13366 10854 13418 10906
rect 13430 10854 13482 10906
rect 13494 10854 13546 10906
rect 13558 10854 13610 10906
rect 13622 10854 13674 10906
rect 13686 10854 13738 10906
rect 4252 10752 4304 10804
rect 5816 10752 5868 10804
rect 6920 10752 6972 10804
rect 7012 10795 7064 10804
rect 7012 10761 7021 10795
rect 7021 10761 7055 10795
rect 7055 10761 7064 10795
rect 7012 10752 7064 10761
rect 4344 10684 4396 10736
rect 6460 10684 6512 10736
rect 6552 10684 6604 10736
rect 8024 10752 8076 10804
rect 9404 10752 9456 10804
rect 9588 10752 9640 10804
rect 12808 10752 12860 10804
rect 13176 10752 13228 10804
rect 13912 10752 13964 10804
rect 14832 10752 14884 10804
rect 16304 10752 16356 10804
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 5264 10616 5316 10668
rect 1768 10548 1820 10600
rect 2320 10548 2372 10600
rect 4620 10548 4672 10600
rect 5080 10548 5132 10600
rect 5264 10480 5316 10532
rect 6368 10616 6420 10668
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 4252 10412 4304 10464
rect 5356 10412 5408 10464
rect 6368 10523 6420 10532
rect 6368 10489 6377 10523
rect 6377 10489 6411 10523
rect 6411 10489 6420 10523
rect 6368 10480 6420 10489
rect 6460 10523 6512 10532
rect 6460 10489 6469 10523
rect 6469 10489 6503 10523
rect 6503 10489 6512 10523
rect 6460 10480 6512 10489
rect 6828 10548 6880 10600
rect 7104 10616 7156 10668
rect 7932 10684 7984 10736
rect 8576 10684 8628 10736
rect 9036 10684 9088 10736
rect 11244 10684 11296 10736
rect 11336 10684 11388 10736
rect 7472 10548 7524 10600
rect 8116 10616 8168 10668
rect 6736 10480 6788 10532
rect 7380 10523 7432 10532
rect 7380 10489 7389 10523
rect 7389 10489 7423 10523
rect 7423 10489 7432 10523
rect 7380 10480 7432 10489
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6276 10412 6328 10464
rect 7104 10412 7156 10464
rect 7656 10412 7708 10464
rect 10876 10548 10928 10600
rect 12716 10616 12768 10668
rect 11704 10548 11756 10600
rect 14004 10616 14056 10668
rect 15200 10684 15252 10736
rect 15844 10684 15896 10736
rect 15292 10616 15344 10668
rect 15568 10616 15620 10668
rect 16212 10616 16264 10668
rect 9036 10480 9088 10532
rect 13360 10548 13412 10600
rect 13820 10548 13872 10600
rect 14096 10548 14148 10600
rect 8484 10412 8536 10464
rect 8576 10412 8628 10464
rect 10232 10412 10284 10464
rect 14372 10480 14424 10532
rect 15844 10548 15896 10600
rect 13544 10412 13596 10464
rect 15108 10480 15160 10532
rect 16212 10412 16264 10464
rect 16948 10412 17000 10464
rect 4366 10310 4418 10362
rect 4430 10310 4482 10362
rect 4494 10310 4546 10362
rect 4558 10310 4610 10362
rect 4622 10310 4674 10362
rect 4686 10310 4738 10362
rect 10366 10310 10418 10362
rect 10430 10310 10482 10362
rect 10494 10310 10546 10362
rect 10558 10310 10610 10362
rect 10622 10310 10674 10362
rect 10686 10310 10738 10362
rect 16366 10310 16418 10362
rect 16430 10310 16482 10362
rect 16494 10310 16546 10362
rect 16558 10310 16610 10362
rect 16622 10310 16674 10362
rect 16686 10310 16738 10362
rect 3976 10208 4028 10260
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 4712 10208 4764 10260
rect 4988 10208 5040 10260
rect 5080 10208 5132 10260
rect 5356 10208 5408 10260
rect 5908 10208 5960 10260
rect 6368 10208 6420 10260
rect 1584 10072 1636 10124
rect 3884 10072 3936 10124
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 4804 10072 4856 10124
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 848 10047 900 10056
rect 848 10013 857 10047
rect 857 10013 891 10047
rect 891 10013 900 10047
rect 848 10004 900 10013
rect 4344 10004 4396 10056
rect 9128 10208 9180 10260
rect 10416 10208 10468 10260
rect 11336 10208 11388 10260
rect 12348 10251 12400 10260
rect 12348 10217 12357 10251
rect 12357 10217 12391 10251
rect 12391 10217 12400 10251
rect 12348 10208 12400 10217
rect 12532 10208 12584 10260
rect 12808 10208 12860 10260
rect 13820 10208 13872 10260
rect 15200 10208 15252 10260
rect 15292 10208 15344 10260
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 5724 10072 5776 10124
rect 7472 10140 7524 10192
rect 6828 10072 6880 10124
rect 7196 10072 7248 10124
rect 4252 9936 4304 9988
rect 6092 10004 6144 10056
rect 6276 10004 6328 10056
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 5172 9936 5224 9988
rect 2688 9868 2740 9920
rect 4160 9868 4212 9920
rect 4804 9868 4856 9920
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9220 10115 9272 10124
rect 9220 10081 9229 10115
rect 9229 10081 9263 10115
rect 9263 10081 9272 10115
rect 9220 10072 9272 10081
rect 10784 10140 10836 10192
rect 11612 10140 11664 10192
rect 17592 10208 17644 10260
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 9956 10072 10008 10124
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 10416 10072 10468 10124
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 13544 10072 13596 10124
rect 14464 10072 14516 10124
rect 15292 10072 15344 10124
rect 15752 10072 15804 10124
rect 13912 10004 13964 10056
rect 14740 10004 14792 10056
rect 15108 10004 15160 10056
rect 16764 10115 16816 10124
rect 16764 10081 16773 10115
rect 16773 10081 16807 10115
rect 16807 10081 16816 10115
rect 16764 10072 16816 10081
rect 7104 9868 7156 9920
rect 7932 9868 7984 9920
rect 9680 9868 9732 9920
rect 9956 9868 10008 9920
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 10416 9868 10468 9920
rect 10784 9868 10836 9920
rect 12348 9936 12400 9988
rect 16028 10004 16080 10056
rect 17040 10115 17092 10124
rect 17040 10081 17049 10115
rect 17049 10081 17083 10115
rect 17083 10081 17092 10115
rect 17040 10072 17092 10081
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 15476 9911 15528 9920
rect 15476 9877 15485 9911
rect 15485 9877 15519 9911
rect 15519 9877 15528 9911
rect 15476 9868 15528 9877
rect 17132 9911 17184 9920
rect 17132 9877 17141 9911
rect 17141 9877 17175 9911
rect 17175 9877 17184 9911
rect 17132 9868 17184 9877
rect 1366 9766 1418 9818
rect 1430 9766 1482 9818
rect 1494 9766 1546 9818
rect 1558 9766 1610 9818
rect 1622 9766 1674 9818
rect 1686 9766 1738 9818
rect 7366 9766 7418 9818
rect 7430 9766 7482 9818
rect 7494 9766 7546 9818
rect 7558 9766 7610 9818
rect 7622 9766 7674 9818
rect 7686 9766 7738 9818
rect 13366 9766 13418 9818
rect 13430 9766 13482 9818
rect 13494 9766 13546 9818
rect 13558 9766 13610 9818
rect 13622 9766 13674 9818
rect 13686 9766 13738 9818
rect 4160 9664 4212 9716
rect 5264 9664 5316 9716
rect 5816 9664 5868 9716
rect 9772 9664 9824 9716
rect 11612 9664 11664 9716
rect 12348 9664 12400 9716
rect 3884 9596 3936 9648
rect 5724 9596 5776 9648
rect 6644 9596 6696 9648
rect 6828 9596 6880 9648
rect 7196 9596 7248 9648
rect 9128 9596 9180 9648
rect 10232 9596 10284 9648
rect 10416 9639 10468 9648
rect 10416 9605 10425 9639
rect 10425 9605 10459 9639
rect 10459 9605 10468 9639
rect 10416 9596 10468 9605
rect 13912 9664 13964 9716
rect 1952 9528 2004 9580
rect 2228 9528 2280 9580
rect 3516 9528 3568 9580
rect 5172 9528 5224 9580
rect 9312 9528 9364 9580
rect 9956 9528 10008 9580
rect 14280 9596 14332 9648
rect 17040 9596 17092 9648
rect 848 9503 900 9512
rect 848 9469 857 9503
rect 857 9469 891 9503
rect 891 9469 900 9503
rect 848 9460 900 9469
rect 1860 9392 1912 9444
rect 3792 9503 3844 9512
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 4160 9460 4212 9512
rect 4528 9460 4580 9512
rect 3884 9392 3936 9444
rect 4620 9392 4672 9444
rect 5264 9460 5316 9512
rect 6184 9503 6236 9512
rect 6184 9469 6193 9503
rect 6193 9469 6227 9503
rect 6227 9469 6236 9503
rect 6184 9460 6236 9469
rect 6368 9460 6420 9512
rect 6460 9503 6512 9512
rect 6460 9469 6469 9503
rect 6469 9469 6503 9503
rect 6503 9469 6512 9503
rect 6460 9460 6512 9469
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 9036 9460 9088 9512
rect 9772 9503 9824 9512
rect 9772 9469 9781 9503
rect 9781 9469 9815 9503
rect 9815 9469 9824 9503
rect 9772 9460 9824 9469
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 10324 9460 10376 9512
rect 11060 9460 11112 9512
rect 11704 9460 11756 9512
rect 12256 9503 12308 9512
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 12256 9460 12308 9469
rect 13268 9528 13320 9580
rect 6736 9435 6788 9444
rect 6736 9401 6771 9435
rect 6771 9401 6788 9435
rect 6736 9392 6788 9401
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 6184 9324 6236 9376
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 6644 9324 6696 9376
rect 6920 9324 6972 9376
rect 7288 9324 7340 9376
rect 9312 9367 9364 9376
rect 9312 9333 9321 9367
rect 9321 9333 9355 9367
rect 9355 9333 9364 9367
rect 9312 9324 9364 9333
rect 10232 9324 10284 9376
rect 12808 9460 12860 9512
rect 17408 9528 17460 9580
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 14372 9503 14424 9512
rect 14372 9469 14381 9503
rect 14381 9469 14415 9503
rect 14415 9469 14424 9503
rect 14372 9460 14424 9469
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 14924 9460 14976 9512
rect 16212 9460 16264 9512
rect 11060 9324 11112 9376
rect 11152 9324 11204 9376
rect 12348 9324 12400 9376
rect 12440 9324 12492 9376
rect 12624 9392 12676 9444
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 14004 9324 14056 9376
rect 14372 9324 14424 9376
rect 14556 9324 14608 9376
rect 16856 9324 16908 9376
rect 4366 9222 4418 9274
rect 4430 9222 4482 9274
rect 4494 9222 4546 9274
rect 4558 9222 4610 9274
rect 4622 9222 4674 9274
rect 4686 9222 4738 9274
rect 10366 9222 10418 9274
rect 10430 9222 10482 9274
rect 10494 9222 10546 9274
rect 10558 9222 10610 9274
rect 10622 9222 10674 9274
rect 10686 9222 10738 9274
rect 16366 9222 16418 9274
rect 16430 9222 16482 9274
rect 16494 9222 16546 9274
rect 16558 9222 16610 9274
rect 16622 9222 16674 9274
rect 16686 9222 16738 9274
rect 4160 9120 4212 9172
rect 4896 9120 4948 9172
rect 6184 9163 6236 9172
rect 6184 9129 6193 9163
rect 6193 9129 6227 9163
rect 6227 9129 6236 9163
rect 6184 9120 6236 9129
rect 6460 9120 6512 9172
rect 9956 9120 10008 9172
rect 10140 9120 10192 9172
rect 848 8984 900 9036
rect 2596 8984 2648 9036
rect 3792 8984 3844 9036
rect 5540 8984 5592 9036
rect 7288 9052 7340 9104
rect 8944 9095 8996 9104
rect 8944 9061 8953 9095
rect 8953 9061 8987 9095
rect 8987 9061 8996 9095
rect 8944 9052 8996 9061
rect 9128 9052 9180 9104
rect 11060 9120 11112 9172
rect 13820 9120 13872 9172
rect 4804 8916 4856 8968
rect 5172 8916 5224 8968
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 6736 8984 6788 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 6920 9027 6972 9036
rect 6920 8993 6929 9027
rect 6929 8993 6963 9027
rect 6963 8993 6972 9027
rect 6920 8984 6972 8993
rect 6276 8848 6328 8900
rect 6644 8916 6696 8968
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 6092 8823 6144 8832
rect 6092 8789 6101 8823
rect 6101 8789 6135 8823
rect 6135 8789 6144 8823
rect 6092 8780 6144 8789
rect 6460 8780 6512 8832
rect 7104 8848 7156 8900
rect 7840 8984 7892 9036
rect 9312 9027 9364 9036
rect 9312 8993 9321 9027
rect 9321 8993 9355 9027
rect 9355 8993 9364 9027
rect 9312 8984 9364 8993
rect 8484 8848 8536 8900
rect 9772 8916 9824 8968
rect 10048 8984 10100 9036
rect 10416 9027 10468 9036
rect 10416 8993 10425 9027
rect 10425 8993 10459 9027
rect 10459 8993 10468 9027
rect 10416 8984 10468 8993
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 10784 8984 10836 9036
rect 11336 9095 11388 9104
rect 11336 9061 11345 9095
rect 11345 9061 11379 9095
rect 11379 9061 11388 9095
rect 11336 9052 11388 9061
rect 11704 9052 11756 9104
rect 12072 8984 12124 9036
rect 12440 9052 12492 9104
rect 12716 8984 12768 9036
rect 12808 9008 12860 9060
rect 13176 9052 13228 9104
rect 13912 9052 13964 9104
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 13820 8984 13872 8993
rect 14280 9120 14332 9172
rect 16764 9120 16816 9172
rect 17040 9120 17092 9172
rect 14556 8984 14608 9036
rect 12808 8916 12860 8968
rect 12256 8848 12308 8900
rect 9680 8780 9732 8832
rect 12624 8780 12676 8832
rect 14464 8848 14516 8900
rect 15752 8984 15804 9036
rect 16856 8984 16908 9036
rect 16028 8916 16080 8968
rect 17132 8916 17184 8968
rect 15200 8780 15252 8832
rect 17132 8780 17184 8832
rect 17408 8780 17460 8832
rect 1366 8678 1418 8730
rect 1430 8678 1482 8730
rect 1494 8678 1546 8730
rect 1558 8678 1610 8730
rect 1622 8678 1674 8730
rect 1686 8678 1738 8730
rect 7366 8678 7418 8730
rect 7430 8678 7482 8730
rect 7494 8678 7546 8730
rect 7558 8678 7610 8730
rect 7622 8678 7674 8730
rect 7686 8678 7738 8730
rect 13366 8678 13418 8730
rect 13430 8678 13482 8730
rect 13494 8678 13546 8730
rect 13558 8678 13610 8730
rect 13622 8678 13674 8730
rect 13686 8678 13738 8730
rect 3148 8576 3200 8628
rect 5540 8619 5592 8628
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 6092 8576 6144 8628
rect 6828 8576 6880 8628
rect 6920 8576 6972 8628
rect 7840 8576 7892 8628
rect 9312 8576 9364 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 12348 8576 12400 8628
rect 13176 8576 13228 8628
rect 16856 8576 16908 8628
rect 848 8440 900 8492
rect 3976 8440 4028 8492
rect 5908 8508 5960 8560
rect 3884 8372 3936 8424
rect 3792 8347 3844 8356
rect 3792 8313 3801 8347
rect 3801 8313 3835 8347
rect 3835 8313 3844 8347
rect 3792 8304 3844 8313
rect 5632 8372 5684 8424
rect 5908 8372 5960 8424
rect 6552 8304 6604 8356
rect 6736 8440 6788 8492
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 10784 8508 10836 8560
rect 11428 8508 11480 8560
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 7840 8415 7892 8424
rect 5172 8236 5224 8288
rect 7380 8304 7432 8356
rect 7840 8381 7849 8415
rect 7849 8381 7883 8415
rect 7883 8381 7892 8415
rect 7840 8372 7892 8381
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 9128 8372 9180 8424
rect 9680 8440 9732 8492
rect 10324 8440 10376 8492
rect 8024 8347 8076 8356
rect 8024 8313 8033 8347
rect 8033 8313 8067 8347
rect 8067 8313 8076 8347
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 10048 8415 10100 8424
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 12256 8440 12308 8492
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 14924 8440 14976 8492
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 8024 8304 8076 8313
rect 10232 8304 10284 8356
rect 10968 8236 11020 8288
rect 11060 8279 11112 8288
rect 11060 8245 11069 8279
rect 11069 8245 11103 8279
rect 11103 8245 11112 8279
rect 11060 8236 11112 8245
rect 11428 8347 11480 8356
rect 11428 8313 11437 8347
rect 11437 8313 11471 8347
rect 11471 8313 11480 8347
rect 11428 8304 11480 8313
rect 11888 8304 11940 8356
rect 14188 8372 14240 8424
rect 16764 8304 16816 8356
rect 12164 8236 12216 8288
rect 13544 8236 13596 8288
rect 13636 8236 13688 8288
rect 13820 8236 13872 8288
rect 14188 8236 14240 8288
rect 14280 8279 14332 8288
rect 14280 8245 14289 8279
rect 14289 8245 14323 8279
rect 14323 8245 14332 8279
rect 14280 8236 14332 8245
rect 14372 8236 14424 8288
rect 4366 8134 4418 8186
rect 4430 8134 4482 8186
rect 4494 8134 4546 8186
rect 4558 8134 4610 8186
rect 4622 8134 4674 8186
rect 4686 8134 4738 8186
rect 10366 8134 10418 8186
rect 10430 8134 10482 8186
rect 10494 8134 10546 8186
rect 10558 8134 10610 8186
rect 10622 8134 10674 8186
rect 10686 8134 10738 8186
rect 16366 8134 16418 8186
rect 16430 8134 16482 8186
rect 16494 8134 16546 8186
rect 16558 8134 16610 8186
rect 16622 8134 16674 8186
rect 16686 8134 16738 8186
rect 2228 8032 2280 8084
rect 2688 8032 2740 8084
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 4252 8032 4304 8084
rect 7012 8032 7064 8084
rect 10140 8032 10192 8084
rect 1952 7896 2004 7948
rect 2228 7896 2280 7948
rect 2320 7896 2372 7948
rect 2596 7896 2648 7948
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 3148 7896 3200 7948
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 5172 7964 5224 8016
rect 5908 8007 5960 8016
rect 5908 7973 5917 8007
rect 5917 7973 5951 8007
rect 5951 7973 5960 8007
rect 5908 7964 5960 7973
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 4896 7896 4948 7948
rect 5264 7896 5316 7948
rect 5540 7896 5592 7948
rect 1952 7760 2004 7812
rect 3516 7760 3568 7812
rect 3976 7760 4028 7812
rect 8116 7964 8168 8016
rect 8300 7964 8352 8016
rect 9220 7964 9272 8016
rect 13820 8032 13872 8084
rect 8024 7896 8076 7948
rect 6092 7828 6144 7880
rect 11244 7896 11296 7948
rect 1768 7735 1820 7744
rect 1768 7701 1777 7735
rect 1777 7701 1811 7735
rect 1811 7701 1820 7735
rect 1768 7692 1820 7701
rect 2596 7735 2648 7744
rect 2596 7701 2605 7735
rect 2605 7701 2639 7735
rect 2639 7701 2648 7735
rect 2596 7692 2648 7701
rect 4988 7692 5040 7744
rect 7104 7760 7156 7812
rect 11520 7828 11572 7880
rect 12164 7939 12216 7948
rect 12164 7905 12173 7939
rect 12173 7905 12207 7939
rect 12207 7905 12216 7939
rect 12164 7896 12216 7905
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 13176 7896 13228 7948
rect 13544 7896 13596 7948
rect 13636 7939 13688 7948
rect 13636 7905 13649 7939
rect 13649 7905 13683 7939
rect 13683 7905 13688 7939
rect 13636 7896 13688 7905
rect 13820 7939 13872 7948
rect 13820 7905 13829 7939
rect 13829 7905 13863 7939
rect 13863 7905 13872 7939
rect 13820 7896 13872 7905
rect 14188 7896 14240 7948
rect 10784 7760 10836 7812
rect 5264 7735 5316 7744
rect 5264 7701 5273 7735
rect 5273 7701 5307 7735
rect 5307 7701 5316 7735
rect 5264 7692 5316 7701
rect 5448 7692 5500 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 8484 7692 8536 7744
rect 10048 7692 10100 7744
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 10692 7692 10744 7744
rect 11704 7760 11756 7812
rect 11612 7735 11664 7744
rect 11612 7701 11621 7735
rect 11621 7701 11655 7735
rect 11655 7701 11664 7735
rect 11612 7692 11664 7701
rect 13544 7760 13596 7812
rect 14556 7939 14608 7948
rect 14556 7905 14565 7939
rect 14565 7905 14599 7939
rect 14599 7905 14608 7939
rect 14556 7896 14608 7905
rect 15200 8032 15252 8084
rect 16764 8032 16816 8084
rect 14740 7896 14792 7948
rect 14924 7896 14976 7948
rect 15200 7939 15252 7948
rect 15200 7905 15209 7939
rect 15209 7905 15243 7939
rect 15243 7905 15252 7939
rect 15200 7896 15252 7905
rect 15752 7964 15804 8016
rect 14648 7760 14700 7812
rect 12348 7692 12400 7744
rect 13820 7692 13872 7744
rect 14924 7692 14976 7744
rect 15016 7735 15068 7744
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 1366 7590 1418 7642
rect 1430 7590 1482 7642
rect 1494 7590 1546 7642
rect 1558 7590 1610 7642
rect 1622 7590 1674 7642
rect 1686 7590 1738 7642
rect 7366 7590 7418 7642
rect 7430 7590 7482 7642
rect 7494 7590 7546 7642
rect 7558 7590 7610 7642
rect 7622 7590 7674 7642
rect 7686 7590 7738 7642
rect 13366 7590 13418 7642
rect 13430 7590 13482 7642
rect 13494 7590 13546 7642
rect 13558 7590 13610 7642
rect 13622 7590 13674 7642
rect 13686 7590 13738 7642
rect 1860 7488 1912 7540
rect 1952 7488 2004 7540
rect 2596 7488 2648 7540
rect 4252 7488 4304 7540
rect 4160 7463 4212 7472
rect 4160 7429 4169 7463
rect 4169 7429 4203 7463
rect 4203 7429 4212 7463
rect 4160 7420 4212 7429
rect 4988 7488 5040 7540
rect 5448 7488 5500 7540
rect 5816 7488 5868 7540
rect 5908 7488 5960 7540
rect 6460 7488 6512 7540
rect 9496 7488 9548 7540
rect 9680 7488 9732 7540
rect 5264 7420 5316 7472
rect 7932 7420 7984 7472
rect 5172 7352 5224 7404
rect 2320 7284 2372 7336
rect 1768 7148 1820 7200
rect 2044 7148 2096 7200
rect 2228 7148 2280 7200
rect 2504 7327 2556 7336
rect 2504 7293 2513 7327
rect 2513 7293 2547 7327
rect 2547 7293 2556 7327
rect 2504 7284 2556 7293
rect 2688 7327 2740 7336
rect 2688 7293 2697 7327
rect 2697 7293 2731 7327
rect 2731 7293 2740 7327
rect 2688 7284 2740 7293
rect 3240 7216 3292 7268
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 3884 7216 3936 7268
rect 4344 7216 4396 7268
rect 4896 7284 4948 7336
rect 5540 7284 5592 7336
rect 6000 7352 6052 7404
rect 6552 7352 6604 7404
rect 6828 7284 6880 7336
rect 8116 7284 8168 7336
rect 9772 7420 9824 7472
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 10416 7488 10468 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 11612 7488 11664 7540
rect 11704 7488 11756 7540
rect 12164 7488 12216 7540
rect 12348 7531 12400 7540
rect 12348 7497 12357 7531
rect 12357 7497 12391 7531
rect 12391 7497 12400 7531
rect 12348 7488 12400 7497
rect 12440 7488 12492 7540
rect 12900 7488 12952 7540
rect 13820 7488 13872 7540
rect 14740 7488 14792 7540
rect 10324 7420 10376 7472
rect 4896 7148 4948 7200
rect 5172 7148 5224 7200
rect 6368 7148 6420 7200
rect 7104 7148 7156 7200
rect 8576 7148 8628 7200
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 11060 7352 11112 7404
rect 15568 7420 15620 7472
rect 15752 7420 15804 7472
rect 11980 7352 12032 7404
rect 14372 7352 14424 7404
rect 14924 7352 14976 7404
rect 15016 7352 15068 7404
rect 10508 7327 10560 7336
rect 10508 7293 10517 7327
rect 10517 7293 10551 7327
rect 10551 7293 10560 7327
rect 10508 7284 10560 7293
rect 11612 7284 11664 7336
rect 12348 7284 12400 7336
rect 12900 7284 12952 7336
rect 14280 7284 14332 7336
rect 15384 7284 15436 7336
rect 15568 7284 15620 7336
rect 15660 7284 15712 7336
rect 16212 7284 16264 7336
rect 17224 7284 17276 7336
rect 9036 7148 9088 7200
rect 9128 7148 9180 7200
rect 9312 7148 9364 7200
rect 10140 7148 10192 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 13176 7148 13228 7200
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 4366 7046 4418 7098
rect 4430 7046 4482 7098
rect 4494 7046 4546 7098
rect 4558 7046 4610 7098
rect 4622 7046 4674 7098
rect 4686 7046 4738 7098
rect 10366 7046 10418 7098
rect 10430 7046 10482 7098
rect 10494 7046 10546 7098
rect 10558 7046 10610 7098
rect 10622 7046 10674 7098
rect 10686 7046 10738 7098
rect 16366 7046 16418 7098
rect 16430 7046 16482 7098
rect 16494 7046 16546 7098
rect 16558 7046 16610 7098
rect 16622 7046 16674 7098
rect 16686 7046 16738 7098
rect 3884 6944 3936 6996
rect 4344 6944 4396 6996
rect 6000 6944 6052 6996
rect 3516 6876 3568 6928
rect 1860 6808 1912 6860
rect 848 6783 900 6792
rect 848 6749 857 6783
rect 857 6749 891 6783
rect 891 6749 900 6783
rect 848 6740 900 6749
rect 2504 6808 2556 6860
rect 3884 6808 3936 6860
rect 4160 6876 4212 6928
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 5264 6876 5316 6928
rect 7012 6876 7064 6928
rect 7196 6876 7248 6928
rect 8116 6876 8168 6928
rect 7288 6851 7340 6860
rect 7288 6817 7297 6851
rect 7297 6817 7331 6851
rect 7331 6817 7340 6851
rect 7288 6808 7340 6817
rect 9036 6944 9088 6996
rect 10968 6944 11020 6996
rect 15200 6944 15252 6996
rect 15384 6944 15436 6996
rect 8576 6876 8628 6928
rect 9496 6876 9548 6928
rect 4068 6672 4120 6724
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 7472 6740 7524 6792
rect 7748 6740 7800 6792
rect 4804 6672 4856 6724
rect 7932 6740 7984 6792
rect 3608 6604 3660 6656
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 4344 6604 4396 6656
rect 6552 6604 6604 6656
rect 7932 6604 7984 6656
rect 9128 6808 9180 6860
rect 10048 6808 10100 6860
rect 10140 6808 10192 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11888 6876 11940 6928
rect 13268 6876 13320 6928
rect 14096 6876 14148 6928
rect 14372 6876 14424 6928
rect 14648 6876 14700 6928
rect 16212 6876 16264 6928
rect 16488 6876 16540 6928
rect 11336 6808 11388 6860
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 9220 6740 9272 6792
rect 9496 6740 9548 6792
rect 10324 6740 10376 6792
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11060 6740 11112 6792
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 9772 6672 9824 6724
rect 8484 6604 8536 6656
rect 15936 6808 15988 6860
rect 16120 6808 16172 6860
rect 11704 6672 11756 6724
rect 14924 6740 14976 6792
rect 14372 6672 14424 6724
rect 14832 6672 14884 6724
rect 12164 6604 12216 6656
rect 12532 6604 12584 6656
rect 13084 6604 13136 6656
rect 1366 6502 1418 6554
rect 1430 6502 1482 6554
rect 1494 6502 1546 6554
rect 1558 6502 1610 6554
rect 1622 6502 1674 6554
rect 1686 6502 1738 6554
rect 7366 6502 7418 6554
rect 7430 6502 7482 6554
rect 7494 6502 7546 6554
rect 7558 6502 7610 6554
rect 7622 6502 7674 6554
rect 7686 6502 7738 6554
rect 13366 6502 13418 6554
rect 13430 6502 13482 6554
rect 13494 6502 13546 6554
rect 13558 6502 13610 6554
rect 13622 6502 13674 6554
rect 13686 6502 13738 6554
rect 3700 6400 3752 6452
rect 6460 6400 6512 6452
rect 7012 6400 7064 6452
rect 8576 6400 8628 6452
rect 5816 6375 5868 6384
rect 5816 6341 5825 6375
rect 5825 6341 5859 6375
rect 5859 6341 5868 6375
rect 5816 6332 5868 6341
rect 6276 6332 6328 6384
rect 2596 6196 2648 6248
rect 6828 6264 6880 6316
rect 7104 6264 7156 6316
rect 7196 6239 7248 6248
rect 2228 6128 2280 6180
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 2044 6060 2096 6112
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 2504 6060 2556 6112
rect 5724 6060 5776 6112
rect 6184 6060 6236 6112
rect 7196 6060 7248 6112
rect 8116 6196 8168 6248
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 9404 6400 9456 6452
rect 9772 6400 9824 6452
rect 11060 6443 11112 6452
rect 11060 6409 11069 6443
rect 11069 6409 11103 6443
rect 11103 6409 11112 6443
rect 11060 6400 11112 6409
rect 11244 6400 11296 6452
rect 8944 6332 8996 6384
rect 11336 6332 11388 6384
rect 12256 6400 12308 6452
rect 15568 6400 15620 6452
rect 15844 6400 15896 6452
rect 16212 6400 16264 6452
rect 8668 6196 8720 6248
rect 11428 6264 11480 6316
rect 9956 6196 10008 6248
rect 10324 6196 10376 6248
rect 10968 6196 11020 6248
rect 11796 6196 11848 6248
rect 8024 6060 8076 6112
rect 11704 6060 11756 6112
rect 12256 6196 12308 6248
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 12164 6128 12216 6180
rect 12256 6060 12308 6112
rect 14188 6196 14240 6248
rect 14556 6196 14608 6248
rect 14832 6264 14884 6316
rect 15200 6128 15252 6180
rect 15568 6196 15620 6248
rect 16120 6196 16172 6248
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 17224 6196 17276 6248
rect 14832 6103 14884 6112
rect 14832 6069 14841 6103
rect 14841 6069 14875 6103
rect 14875 6069 14884 6103
rect 14832 6060 14884 6069
rect 15568 6060 15620 6112
rect 16120 6103 16172 6112
rect 16120 6069 16129 6103
rect 16129 6069 16163 6103
rect 16163 6069 16172 6103
rect 16120 6060 16172 6069
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 4366 5958 4418 6010
rect 4430 5958 4482 6010
rect 4494 5958 4546 6010
rect 4558 5958 4610 6010
rect 4622 5958 4674 6010
rect 4686 5958 4738 6010
rect 10366 5958 10418 6010
rect 10430 5958 10482 6010
rect 10494 5958 10546 6010
rect 10558 5958 10610 6010
rect 10622 5958 10674 6010
rect 10686 5958 10738 6010
rect 16366 5958 16418 6010
rect 16430 5958 16482 6010
rect 16494 5958 16546 6010
rect 16558 5958 16610 6010
rect 16622 5958 16674 6010
rect 16686 5958 16738 6010
rect 1860 5856 1912 5908
rect 3332 5856 3384 5908
rect 3976 5856 4028 5908
rect 848 5695 900 5704
rect 848 5661 857 5695
rect 857 5661 891 5695
rect 891 5661 900 5695
rect 848 5652 900 5661
rect 2412 5652 2464 5704
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 3056 5720 3108 5729
rect 3608 5763 3660 5772
rect 3608 5729 3617 5763
rect 3617 5729 3651 5763
rect 3651 5729 3660 5763
rect 3608 5720 3660 5729
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 3516 5652 3568 5704
rect 3700 5695 3752 5704
rect 3700 5661 3709 5695
rect 3709 5661 3743 5695
rect 3743 5661 3752 5695
rect 3700 5652 3752 5661
rect 5632 5788 5684 5840
rect 7104 5856 7156 5908
rect 7288 5856 7340 5908
rect 7380 5856 7432 5908
rect 8392 5856 8444 5908
rect 15568 5856 15620 5908
rect 16028 5856 16080 5908
rect 16120 5856 16172 5908
rect 16212 5856 16264 5908
rect 3608 5584 3660 5636
rect 4896 5652 4948 5704
rect 5540 5652 5592 5704
rect 5264 5584 5316 5636
rect 6368 5763 6420 5772
rect 6368 5729 6377 5763
rect 6377 5729 6411 5763
rect 6411 5729 6420 5763
rect 6368 5720 6420 5729
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 7012 5720 7064 5772
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 6828 5652 6880 5704
rect 9588 5720 9640 5772
rect 7288 5652 7340 5704
rect 8576 5652 8628 5704
rect 11336 5720 11388 5772
rect 12256 5763 12308 5772
rect 12256 5729 12265 5763
rect 12265 5729 12299 5763
rect 12299 5729 12308 5763
rect 12256 5720 12308 5729
rect 12808 5720 12860 5772
rect 13268 5763 13320 5772
rect 13268 5729 13277 5763
rect 13277 5729 13311 5763
rect 13311 5729 13320 5763
rect 13268 5720 13320 5729
rect 13636 5763 13688 5772
rect 13636 5729 13645 5763
rect 13645 5729 13679 5763
rect 13679 5729 13688 5763
rect 13636 5720 13688 5729
rect 13820 5720 13872 5772
rect 8668 5584 8720 5636
rect 8944 5584 8996 5636
rect 9404 5584 9456 5636
rect 10232 5584 10284 5636
rect 11796 5584 11848 5636
rect 12900 5584 12952 5636
rect 13544 5584 13596 5636
rect 14556 5720 14608 5772
rect 15200 5788 15252 5840
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 16396 5720 16448 5772
rect 17132 5763 17184 5772
rect 17132 5729 17141 5763
rect 17141 5729 17175 5763
rect 17175 5729 17184 5763
rect 17132 5720 17184 5729
rect 16764 5627 16816 5636
rect 16764 5593 16773 5627
rect 16773 5593 16807 5627
rect 16807 5593 16816 5627
rect 16764 5584 16816 5593
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 3240 5559 3292 5568
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 6184 5516 6236 5568
rect 6460 5516 6512 5568
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 9496 5516 9548 5568
rect 10048 5516 10100 5568
rect 10784 5516 10836 5568
rect 11244 5516 11296 5568
rect 11704 5516 11756 5568
rect 11980 5516 12032 5568
rect 12532 5516 12584 5568
rect 13268 5516 13320 5568
rect 14096 5516 14148 5568
rect 14188 5516 14240 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 16948 5559 17000 5568
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 1366 5414 1418 5466
rect 1430 5414 1482 5466
rect 1494 5414 1546 5466
rect 1558 5414 1610 5466
rect 1622 5414 1674 5466
rect 1686 5414 1738 5466
rect 7366 5414 7418 5466
rect 7430 5414 7482 5466
rect 7494 5414 7546 5466
rect 7558 5414 7610 5466
rect 7622 5414 7674 5466
rect 7686 5414 7738 5466
rect 13366 5414 13418 5466
rect 13430 5414 13482 5466
rect 13494 5414 13546 5466
rect 13558 5414 13610 5466
rect 13622 5414 13674 5466
rect 13686 5414 13738 5466
rect 6828 5312 6880 5364
rect 8116 5312 8168 5364
rect 8576 5312 8628 5364
rect 2044 5176 2096 5228
rect 2412 5108 2464 5160
rect 2596 5151 2648 5160
rect 2596 5117 2605 5151
rect 2605 5117 2639 5151
rect 2639 5117 2648 5151
rect 2596 5108 2648 5117
rect 1492 5040 1544 5092
rect 2136 5040 2188 5092
rect 3332 5176 3384 5228
rect 6552 5244 6604 5296
rect 9772 5312 9824 5364
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 5816 5176 5868 5228
rect 6000 5176 6052 5228
rect 6276 5176 6328 5228
rect 6368 5176 6420 5228
rect 8760 5244 8812 5296
rect 9404 5287 9456 5296
rect 9404 5253 9413 5287
rect 9413 5253 9447 5287
rect 9447 5253 9456 5287
rect 9404 5244 9456 5253
rect 9680 5244 9732 5296
rect 8024 5176 8076 5228
rect 3608 5151 3660 5160
rect 3608 5117 3617 5151
rect 3617 5117 3651 5151
rect 3651 5117 3660 5151
rect 3608 5108 3660 5117
rect 3516 5040 3568 5092
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 3976 5040 4028 5092
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 2596 4972 2648 5024
rect 2688 5015 2740 5024
rect 2688 4981 2697 5015
rect 2697 4981 2731 5015
rect 2731 4981 2740 5015
rect 2688 4972 2740 4981
rect 2964 4972 3016 5024
rect 3884 4972 3936 5024
rect 4896 5151 4948 5160
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 5540 5108 5592 5160
rect 5724 5108 5776 5160
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 7564 5108 7616 5160
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 8484 5108 8536 5160
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 10784 5176 10836 5228
rect 11520 5176 11572 5228
rect 9588 5151 9640 5160
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 9772 5108 9824 5160
rect 9864 5108 9916 5160
rect 10048 5108 10100 5160
rect 10140 5108 10192 5160
rect 6000 5040 6052 5092
rect 4160 4972 4212 5024
rect 8116 5040 8168 5092
rect 11244 5108 11296 5160
rect 6920 4972 6972 5024
rect 7288 4972 7340 5024
rect 8484 4972 8536 5024
rect 9680 4972 9732 5024
rect 10048 4972 10100 5024
rect 10140 5015 10192 5024
rect 10140 4981 10149 5015
rect 10149 4981 10183 5015
rect 10183 4981 10192 5015
rect 10140 4972 10192 4981
rect 10784 4972 10836 5024
rect 11888 5151 11940 5160
rect 11888 5117 11897 5151
rect 11897 5117 11931 5151
rect 11931 5117 11940 5151
rect 11888 5108 11940 5117
rect 12164 5219 12216 5228
rect 12164 5185 12173 5219
rect 12173 5185 12207 5219
rect 12207 5185 12216 5219
rect 12164 5176 12216 5185
rect 12808 5312 12860 5364
rect 12900 5244 12952 5296
rect 15752 5244 15804 5296
rect 12164 5040 12216 5092
rect 12624 5083 12676 5092
rect 12624 5049 12633 5083
rect 12633 5049 12667 5083
rect 12667 5049 12676 5083
rect 12624 5040 12676 5049
rect 12900 5151 12952 5160
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 13360 5108 13412 5160
rect 13728 5108 13780 5160
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 14556 5176 14608 5228
rect 14280 5108 14332 5160
rect 4366 4870 4418 4922
rect 4430 4870 4482 4922
rect 4494 4870 4546 4922
rect 4558 4870 4610 4922
rect 4622 4870 4674 4922
rect 4686 4870 4738 4922
rect 10366 4870 10418 4922
rect 10430 4870 10482 4922
rect 10494 4870 10546 4922
rect 10558 4870 10610 4922
rect 10622 4870 10674 4922
rect 10686 4870 10738 4922
rect 16366 4870 16418 4922
rect 16430 4870 16482 4922
rect 16494 4870 16546 4922
rect 16558 4870 16610 4922
rect 16622 4870 16674 4922
rect 16686 4870 16738 4922
rect 1492 4768 1544 4820
rect 1860 4768 1912 4820
rect 2688 4768 2740 4820
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 4988 4632 5040 4684
rect 5816 4768 5868 4820
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 3516 4564 3568 4616
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 7288 4768 7340 4820
rect 8484 4768 8536 4820
rect 8668 4768 8720 4820
rect 6552 4632 6604 4684
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 7288 4632 7340 4684
rect 7564 4632 7616 4684
rect 1216 4471 1268 4480
rect 1216 4437 1225 4471
rect 1225 4437 1259 4471
rect 1259 4437 1268 4471
rect 1216 4428 1268 4437
rect 1676 4428 1728 4480
rect 4712 4496 4764 4548
rect 5816 4564 5868 4616
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 8024 4675 8076 4684
rect 8024 4641 8033 4675
rect 8033 4641 8067 4675
rect 8067 4641 8076 4675
rect 8024 4632 8076 4641
rect 9496 4700 9548 4752
rect 8484 4632 8536 4684
rect 6644 4496 6696 4548
rect 8116 4564 8168 4616
rect 9036 4564 9088 4616
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 9588 4675 9640 4684
rect 9588 4641 9597 4675
rect 9597 4641 9631 4675
rect 9631 4641 9640 4675
rect 9588 4632 9640 4641
rect 9680 4632 9732 4684
rect 11060 4768 11112 4820
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 11888 4768 11940 4820
rect 12072 4768 12124 4820
rect 12164 4768 12216 4820
rect 11704 4700 11756 4752
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 14464 4700 14516 4752
rect 11520 4632 11572 4641
rect 13176 4632 13228 4684
rect 15660 4700 15712 4752
rect 3516 4428 3568 4480
rect 6276 4428 6328 4480
rect 6920 4428 6972 4480
rect 9680 4496 9732 4548
rect 9864 4496 9916 4548
rect 10784 4564 10836 4616
rect 12256 4564 12308 4616
rect 12716 4564 12768 4616
rect 13912 4607 13964 4616
rect 13912 4573 13921 4607
rect 13921 4573 13955 4607
rect 13955 4573 13964 4607
rect 13912 4564 13964 4573
rect 14004 4607 14056 4616
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 16764 4632 16816 4684
rect 16856 4564 16908 4616
rect 17040 4564 17092 4616
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 14464 4471 14516 4480
rect 14464 4437 14473 4471
rect 14473 4437 14507 4471
rect 14507 4437 14516 4471
rect 14464 4428 14516 4437
rect 14648 4428 14700 4480
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 1366 4326 1418 4378
rect 1430 4326 1482 4378
rect 1494 4326 1546 4378
rect 1558 4326 1610 4378
rect 1622 4326 1674 4378
rect 1686 4326 1738 4378
rect 7366 4326 7418 4378
rect 7430 4326 7482 4378
rect 7494 4326 7546 4378
rect 7558 4326 7610 4378
rect 7622 4326 7674 4378
rect 7686 4326 7738 4378
rect 13366 4326 13418 4378
rect 13430 4326 13482 4378
rect 13494 4326 13546 4378
rect 13558 4326 13610 4378
rect 13622 4326 13674 4378
rect 13686 4326 13738 4378
rect 4160 4224 4212 4276
rect 5448 4224 5500 4276
rect 4712 4156 4764 4208
rect 5172 4156 5224 4208
rect 848 4063 900 4072
rect 848 4029 857 4063
rect 857 4029 891 4063
rect 891 4029 900 4063
rect 848 4020 900 4029
rect 2320 4020 2372 4072
rect 3516 4063 3568 4072
rect 3516 4029 3550 4063
rect 3550 4029 3568 4063
rect 1216 3952 1268 4004
rect 3516 4020 3568 4029
rect 3884 4020 3936 4072
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 6552 4156 6604 4208
rect 7196 4224 7248 4276
rect 11244 4224 11296 4276
rect 6828 4088 6880 4140
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 5540 3952 5592 4004
rect 6276 4020 6328 4072
rect 6920 4020 6972 4072
rect 8024 4156 8076 4208
rect 8484 4156 8536 4208
rect 11060 4156 11112 4208
rect 8116 4088 8168 4140
rect 10968 4088 11020 4140
rect 7748 4020 7800 4072
rect 9036 4020 9088 4072
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 9864 4020 9916 4072
rect 10048 4020 10100 4072
rect 12256 4088 12308 4140
rect 12808 4088 12860 4140
rect 14004 4224 14056 4276
rect 14372 4224 14424 4276
rect 14556 4224 14608 4276
rect 15108 4224 15160 4276
rect 15660 4224 15712 4276
rect 11520 4020 11572 4072
rect 9220 3952 9272 4004
rect 9680 3952 9732 4004
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 14832 4088 14884 4140
rect 13176 4020 13228 4029
rect 13820 4063 13872 4072
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 13820 4020 13872 4029
rect 13452 3952 13504 4004
rect 14096 4020 14148 4072
rect 15200 4088 15252 4140
rect 16764 4156 16816 4208
rect 1768 3884 1820 3936
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 2688 3884 2740 3936
rect 3424 3884 3476 3936
rect 4896 3884 4948 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 5724 3884 5776 3936
rect 6368 3884 6420 3936
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 10048 3884 10100 3936
rect 13360 3927 13412 3936
rect 13360 3893 13369 3927
rect 13369 3893 13403 3927
rect 13403 3893 13412 3927
rect 13360 3884 13412 3893
rect 13544 3884 13596 3936
rect 16120 4020 16172 4072
rect 16764 4063 16816 4072
rect 16764 4029 16773 4063
rect 16773 4029 16807 4063
rect 16807 4029 16816 4063
rect 16764 4020 16816 4029
rect 16948 4063 17000 4072
rect 16948 4029 16957 4063
rect 16957 4029 16991 4063
rect 16991 4029 17000 4063
rect 16948 4020 17000 4029
rect 17316 4063 17368 4072
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 16856 3952 16908 4004
rect 14280 3927 14332 3936
rect 14280 3893 14289 3927
rect 14289 3893 14323 3927
rect 14323 3893 14332 3927
rect 14280 3884 14332 3893
rect 14556 3884 14608 3936
rect 14832 3884 14884 3936
rect 4366 3782 4418 3834
rect 4430 3782 4482 3834
rect 4494 3782 4546 3834
rect 4558 3782 4610 3834
rect 4622 3782 4674 3834
rect 4686 3782 4738 3834
rect 10366 3782 10418 3834
rect 10430 3782 10482 3834
rect 10494 3782 10546 3834
rect 10558 3782 10610 3834
rect 10622 3782 10674 3834
rect 10686 3782 10738 3834
rect 16366 3782 16418 3834
rect 16430 3782 16482 3834
rect 16494 3782 16546 3834
rect 16558 3782 16610 3834
rect 16622 3782 16674 3834
rect 16686 3782 16738 3834
rect 2320 3680 2372 3732
rect 2872 3680 2924 3732
rect 5448 3680 5500 3732
rect 6000 3680 6052 3732
rect 8116 3680 8168 3732
rect 2136 3544 2188 3596
rect 2412 3587 2464 3596
rect 2412 3553 2421 3587
rect 2421 3553 2455 3587
rect 2455 3553 2464 3587
rect 2412 3544 2464 3553
rect 2688 3612 2740 3664
rect 3148 3544 3200 3596
rect 4988 3612 5040 3664
rect 5264 3655 5316 3664
rect 5264 3621 5273 3655
rect 5273 3621 5307 3655
rect 5307 3621 5316 3655
rect 5264 3612 5316 3621
rect 5908 3612 5960 3664
rect 4160 3544 4212 3596
rect 2780 3476 2832 3528
rect 3884 3476 3936 3528
rect 6092 3476 6144 3528
rect 2872 3408 2924 3460
rect 6552 3544 6604 3596
rect 7104 3544 7156 3596
rect 8392 3612 8444 3664
rect 9128 3680 9180 3732
rect 9772 3680 9824 3732
rect 9864 3680 9916 3732
rect 10048 3680 10100 3732
rect 10416 3680 10468 3732
rect 11244 3680 11296 3732
rect 11612 3680 11664 3732
rect 12440 3680 12492 3732
rect 13268 3680 13320 3732
rect 13452 3680 13504 3732
rect 13820 3680 13872 3732
rect 13912 3723 13964 3732
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 14188 3680 14240 3732
rect 15016 3680 15068 3732
rect 9220 3612 9272 3664
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 10048 3544 10100 3596
rect 10232 3544 10284 3596
rect 10968 3544 11020 3596
rect 7104 3408 7156 3460
rect 10416 3519 10468 3528
rect 10416 3485 10425 3519
rect 10425 3485 10459 3519
rect 10459 3485 10468 3519
rect 10416 3476 10468 3485
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2412 3383 2464 3392
rect 2412 3349 2421 3383
rect 2421 3349 2455 3383
rect 2455 3349 2464 3383
rect 2412 3340 2464 3349
rect 6000 3340 6052 3392
rect 6828 3340 6880 3392
rect 7840 3340 7892 3392
rect 8944 3408 8996 3460
rect 11888 3476 11940 3528
rect 12164 3587 12216 3596
rect 12164 3553 12173 3587
rect 12173 3553 12207 3587
rect 12207 3553 12216 3587
rect 12164 3544 12216 3553
rect 12900 3476 12952 3528
rect 11520 3408 11572 3460
rect 11796 3408 11848 3460
rect 13544 3476 13596 3528
rect 14004 3587 14056 3596
rect 14004 3553 14013 3587
rect 14013 3553 14047 3587
rect 14047 3553 14056 3587
rect 14004 3544 14056 3553
rect 14464 3587 14516 3596
rect 14464 3553 14473 3587
rect 14473 3553 14507 3587
rect 14507 3553 14516 3587
rect 14464 3544 14516 3553
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 14188 3476 14240 3485
rect 14648 3476 14700 3528
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 15384 3476 15436 3528
rect 16212 3476 16264 3528
rect 16856 3544 16908 3596
rect 17040 3476 17092 3528
rect 14556 3408 14608 3460
rect 10416 3340 10468 3392
rect 11060 3340 11112 3392
rect 12256 3340 12308 3392
rect 13912 3340 13964 3392
rect 14004 3340 14056 3392
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 16764 3340 16816 3392
rect 1366 3238 1418 3290
rect 1430 3238 1482 3290
rect 1494 3238 1546 3290
rect 1558 3238 1610 3290
rect 1622 3238 1674 3290
rect 1686 3238 1738 3290
rect 7366 3238 7418 3290
rect 7430 3238 7482 3290
rect 7494 3238 7546 3290
rect 7558 3238 7610 3290
rect 7622 3238 7674 3290
rect 7686 3238 7738 3290
rect 13366 3238 13418 3290
rect 13430 3238 13482 3290
rect 13494 3238 13546 3290
rect 13558 3238 13610 3290
rect 13622 3238 13674 3290
rect 13686 3238 13738 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 2320 3136 2372 3188
rect 2412 3136 2464 3188
rect 4804 3136 4856 3188
rect 4252 3000 4304 3052
rect 4436 2932 4488 2984
rect 5724 3068 5776 3120
rect 2780 2864 2832 2916
rect 4068 2864 4120 2916
rect 5264 2975 5316 2984
rect 5264 2941 5273 2975
rect 5273 2941 5307 2975
rect 5307 2941 5316 2975
rect 5264 2932 5316 2941
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 6000 2975 6052 2984
rect 6000 2941 6035 2975
rect 6035 2941 6052 2975
rect 6000 2932 6052 2941
rect 6276 2932 6328 2984
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 6828 3136 6880 3188
rect 7012 3136 7064 3188
rect 7288 3136 7340 3188
rect 7840 3136 7892 3188
rect 9036 3136 9088 3188
rect 9220 3136 9272 3188
rect 6552 3068 6604 3120
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 3792 2839 3844 2848
rect 3792 2805 3801 2839
rect 3801 2805 3835 2839
rect 3835 2805 3844 2839
rect 3792 2796 3844 2805
rect 4252 2796 4304 2848
rect 4804 2796 4856 2848
rect 6184 2796 6236 2848
rect 7104 2932 7156 2984
rect 7012 2796 7064 2848
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 7840 2975 7892 2984
rect 7840 2941 7849 2975
rect 7849 2941 7883 2975
rect 7883 2941 7892 2975
rect 7840 2932 7892 2941
rect 8024 2932 8076 2984
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10048 3136 10100 3188
rect 11796 3136 11848 3188
rect 14556 3136 14608 3188
rect 16120 3136 16172 3188
rect 16212 3136 16264 3188
rect 12900 3068 12952 3120
rect 13728 3068 13780 3120
rect 13912 3068 13964 3120
rect 11060 2932 11112 2984
rect 11796 2975 11848 2984
rect 11796 2941 11805 2975
rect 11805 2941 11839 2975
rect 11839 2941 11848 2975
rect 11796 2932 11848 2941
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 12532 3000 12584 3052
rect 12992 3000 13044 3052
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 15016 3068 15068 3120
rect 13360 2932 13412 2984
rect 16856 3000 16908 3052
rect 8024 2796 8076 2848
rect 8116 2839 8168 2848
rect 8116 2805 8125 2839
rect 8125 2805 8159 2839
rect 8159 2805 8168 2839
rect 8116 2796 8168 2805
rect 9404 2839 9456 2848
rect 9404 2805 9413 2839
rect 9413 2805 9447 2839
rect 9447 2805 9456 2839
rect 9404 2796 9456 2805
rect 14740 2932 14792 2984
rect 15292 2975 15344 2984
rect 15292 2941 15301 2975
rect 15301 2941 15335 2975
rect 15335 2941 15344 2975
rect 15292 2932 15344 2941
rect 16120 2932 16172 2984
rect 17132 2975 17184 2984
rect 17132 2941 17141 2975
rect 17141 2941 17175 2975
rect 17175 2941 17184 2975
rect 17132 2932 17184 2941
rect 13176 2796 13228 2848
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 14188 2839 14240 2848
rect 14188 2805 14197 2839
rect 14197 2805 14231 2839
rect 14231 2805 14240 2839
rect 14188 2796 14240 2805
rect 14280 2796 14332 2848
rect 16948 2864 17000 2916
rect 17224 2864 17276 2916
rect 14924 2796 14976 2848
rect 15108 2796 15160 2848
rect 15568 2796 15620 2848
rect 16764 2796 16816 2848
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 4366 2694 4418 2746
rect 4430 2694 4482 2746
rect 4494 2694 4546 2746
rect 4558 2694 4610 2746
rect 4622 2694 4674 2746
rect 4686 2694 4738 2746
rect 10366 2694 10418 2746
rect 10430 2694 10482 2746
rect 10494 2694 10546 2746
rect 10558 2694 10610 2746
rect 10622 2694 10674 2746
rect 10686 2694 10738 2746
rect 16366 2694 16418 2746
rect 16430 2694 16482 2746
rect 16494 2694 16546 2746
rect 16558 2694 16610 2746
rect 16622 2694 16674 2746
rect 16686 2694 16738 2746
rect 3424 2592 3476 2644
rect 4436 2592 4488 2644
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 3608 2524 3660 2576
rect 8668 2592 8720 2644
rect 11244 2592 11296 2644
rect 14740 2592 14792 2644
rect 7104 2524 7156 2576
rect 7656 2567 7708 2576
rect 7656 2533 7665 2567
rect 7665 2533 7699 2567
rect 7699 2533 7708 2567
rect 7656 2524 7708 2533
rect 8208 2524 8260 2576
rect 8300 2524 8352 2576
rect 1768 2456 1820 2508
rect 2964 2456 3016 2508
rect 3700 2456 3752 2508
rect 3792 2456 3844 2508
rect 4252 2499 4304 2508
rect 4252 2465 4261 2499
rect 4261 2465 4295 2499
rect 4295 2465 4304 2499
rect 4252 2456 4304 2465
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 7288 2456 7340 2508
rect 3516 2388 3568 2440
rect 6828 2388 6880 2440
rect 9036 2499 9088 2508
rect 9036 2465 9045 2499
rect 9045 2465 9079 2499
rect 9079 2465 9088 2499
rect 9036 2456 9088 2465
rect 9312 2499 9364 2508
rect 9312 2465 9321 2499
rect 9321 2465 9355 2499
rect 9355 2465 9364 2499
rect 9312 2456 9364 2465
rect 10600 2456 10652 2508
rect 11244 2456 11296 2508
rect 12348 2524 12400 2576
rect 1768 2320 1820 2372
rect 3240 2320 3292 2372
rect 4344 2320 4396 2372
rect 5724 2320 5776 2372
rect 3332 2295 3384 2304
rect 3332 2261 3341 2295
rect 3341 2261 3375 2295
rect 3375 2261 3384 2295
rect 3332 2252 3384 2261
rect 4068 2295 4120 2304
rect 4068 2261 4077 2295
rect 4077 2261 4111 2295
rect 4111 2261 4120 2295
rect 4068 2252 4120 2261
rect 5540 2252 5592 2304
rect 7012 2320 7064 2372
rect 8024 2320 8076 2372
rect 11060 2388 11112 2440
rect 7288 2295 7340 2304
rect 7288 2261 7297 2295
rect 7297 2261 7331 2295
rect 7331 2261 7340 2295
rect 7288 2252 7340 2261
rect 8852 2295 8904 2304
rect 8852 2261 8861 2295
rect 8861 2261 8895 2295
rect 8895 2261 8904 2295
rect 8852 2252 8904 2261
rect 9036 2320 9088 2372
rect 10600 2320 10652 2372
rect 12532 2499 12584 2508
rect 12532 2465 12541 2499
rect 12541 2465 12575 2499
rect 12575 2465 12584 2499
rect 12532 2456 12584 2465
rect 12716 2524 12768 2576
rect 14004 2524 14056 2576
rect 12072 2320 12124 2372
rect 9772 2252 9824 2304
rect 12440 2320 12492 2372
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 14556 2499 14608 2508
rect 14556 2465 14565 2499
rect 14565 2465 14599 2499
rect 14599 2465 14608 2499
rect 14556 2456 14608 2465
rect 15016 2524 15068 2576
rect 15200 2524 15252 2576
rect 16212 2592 16264 2644
rect 17132 2635 17184 2644
rect 14924 2499 14976 2508
rect 14924 2465 14933 2499
rect 14933 2465 14967 2499
rect 14967 2465 14976 2499
rect 14924 2456 14976 2465
rect 12808 2320 12860 2372
rect 15384 2499 15436 2508
rect 15384 2465 15393 2499
rect 15393 2465 15427 2499
rect 15427 2465 15436 2499
rect 15384 2456 15436 2465
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 15568 2456 15620 2465
rect 17132 2601 17141 2635
rect 17141 2601 17175 2635
rect 17175 2601 17184 2635
rect 17132 2592 17184 2601
rect 17500 2524 17552 2576
rect 17592 2524 17644 2576
rect 14004 2252 14056 2304
rect 14280 2252 14332 2304
rect 14556 2252 14608 2304
rect 14740 2252 14792 2304
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 15568 2320 15620 2372
rect 17500 2320 17552 2372
rect 15476 2252 15528 2304
rect 15844 2295 15896 2304
rect 15844 2261 15853 2295
rect 15853 2261 15887 2295
rect 15887 2261 15896 2295
rect 15844 2252 15896 2261
rect 16028 2252 16080 2304
rect 16396 2252 16448 2304
rect 16488 2295 16540 2304
rect 16488 2261 16497 2295
rect 16497 2261 16531 2295
rect 16531 2261 16540 2295
rect 16488 2252 16540 2261
rect 16856 2252 16908 2304
rect 1366 2150 1418 2202
rect 1430 2150 1482 2202
rect 1494 2150 1546 2202
rect 1558 2150 1610 2202
rect 1622 2150 1674 2202
rect 1686 2150 1738 2202
rect 7366 2150 7418 2202
rect 7430 2150 7482 2202
rect 7494 2150 7546 2202
rect 7558 2150 7610 2202
rect 7622 2150 7674 2202
rect 7686 2150 7738 2202
rect 13366 2150 13418 2202
rect 13430 2150 13482 2202
rect 13494 2150 13546 2202
rect 13558 2150 13610 2202
rect 13622 2150 13674 2202
rect 13686 2150 13738 2202
rect 1768 2048 1820 2100
rect 3332 2048 3384 2100
rect 2044 1980 2096 2032
rect 3516 1980 3568 2032
rect 4528 1980 4580 2032
rect 1860 1844 1912 1896
rect 1952 1887 2004 1896
rect 1952 1853 1961 1887
rect 1961 1853 1995 1887
rect 1995 1853 2004 1887
rect 1952 1844 2004 1853
rect 2320 1844 2372 1896
rect 2688 1844 2740 1896
rect 1860 1708 1912 1760
rect 2412 1708 2464 1760
rect 3240 1819 3292 1828
rect 3240 1785 3249 1819
rect 3249 1785 3283 1819
rect 3283 1785 3292 1819
rect 3240 1776 3292 1785
rect 3516 1844 3568 1896
rect 4252 1912 4304 1964
rect 4344 1955 4396 1964
rect 4344 1921 4353 1955
rect 4353 1921 4387 1955
rect 4387 1921 4396 1955
rect 4344 1912 4396 1921
rect 4436 1912 4488 1964
rect 6092 2091 6144 2100
rect 6092 2057 6101 2091
rect 6101 2057 6135 2091
rect 6135 2057 6144 2091
rect 6092 2048 6144 2057
rect 4712 1980 4764 2032
rect 5356 2023 5408 2032
rect 5356 1989 5365 2023
rect 5365 1989 5399 2023
rect 5399 1989 5408 2023
rect 5356 1980 5408 1989
rect 3792 1887 3844 1896
rect 3792 1853 3801 1887
rect 3801 1853 3835 1887
rect 3835 1853 3844 1887
rect 3792 1844 3844 1853
rect 3884 1844 3936 1896
rect 4068 1887 4120 1896
rect 4068 1853 4077 1887
rect 4077 1853 4111 1887
rect 4111 1853 4120 1887
rect 4068 1844 4120 1853
rect 2780 1708 2832 1760
rect 2964 1751 3016 1760
rect 2964 1717 2973 1751
rect 2973 1717 3007 1751
rect 3007 1717 3016 1751
rect 2964 1708 3016 1717
rect 3332 1708 3384 1760
rect 4988 1887 5040 1896
rect 4988 1853 4997 1887
rect 4997 1853 5031 1887
rect 5031 1853 5040 1887
rect 4988 1844 5040 1853
rect 5908 1912 5960 1964
rect 6460 2023 6512 2032
rect 6460 1989 6469 2023
rect 6469 1989 6503 2023
rect 6503 1989 6512 2023
rect 6460 1980 6512 1989
rect 6000 1844 6052 1896
rect 7564 1980 7616 2032
rect 8300 1980 8352 2032
rect 8668 1980 8720 2032
rect 9128 2023 9180 2032
rect 9128 1989 9137 2023
rect 9137 1989 9171 2023
rect 9171 1989 9180 2023
rect 9128 1980 9180 1989
rect 6736 1912 6788 1964
rect 7288 1912 7340 1964
rect 8208 1912 8260 1964
rect 8944 1912 8996 1964
rect 10692 2048 10744 2100
rect 12072 2048 12124 2100
rect 14188 2048 14240 2100
rect 14832 2048 14884 2100
rect 15476 2091 15528 2100
rect 15476 2057 15485 2091
rect 15485 2057 15519 2091
rect 15519 2057 15528 2091
rect 15476 2048 15528 2057
rect 7012 1887 7064 1896
rect 7012 1853 7021 1887
rect 7021 1853 7055 1887
rect 7055 1853 7064 1887
rect 7012 1844 7064 1853
rect 7656 1887 7708 1896
rect 7656 1853 7665 1887
rect 7665 1853 7699 1887
rect 7699 1853 7708 1887
rect 7656 1844 7708 1853
rect 7840 1844 7892 1896
rect 8024 1844 8076 1896
rect 8852 1887 8904 1896
rect 8852 1853 8861 1887
rect 8861 1853 8895 1887
rect 8895 1853 8904 1887
rect 8852 1844 8904 1853
rect 9036 1887 9088 1896
rect 9036 1853 9045 1887
rect 9045 1853 9079 1887
rect 9079 1853 9088 1887
rect 9036 1844 9088 1853
rect 7196 1776 7248 1828
rect 9680 1887 9732 1896
rect 9680 1853 9689 1887
rect 9689 1853 9723 1887
rect 9723 1853 9732 1887
rect 9680 1844 9732 1853
rect 9772 1887 9824 1896
rect 9772 1853 9781 1887
rect 9781 1853 9815 1887
rect 9815 1853 9824 1887
rect 9772 1844 9824 1853
rect 9864 1844 9916 1896
rect 12440 1980 12492 2032
rect 13084 1980 13136 2032
rect 11060 1912 11112 1964
rect 11980 1955 12032 1964
rect 11980 1921 11989 1955
rect 11989 1921 12023 1955
rect 12023 1921 12032 1955
rect 11980 1912 12032 1921
rect 12624 1912 12676 1964
rect 4896 1751 4948 1760
rect 4896 1717 4905 1751
rect 4905 1717 4939 1751
rect 4939 1717 4948 1751
rect 4896 1708 4948 1717
rect 8484 1708 8536 1760
rect 8576 1751 8628 1760
rect 8576 1717 8585 1751
rect 8585 1717 8619 1751
rect 8619 1717 8628 1751
rect 8576 1708 8628 1717
rect 8668 1708 8720 1760
rect 10048 1776 10100 1828
rect 12348 1887 12400 1896
rect 12348 1853 12357 1887
rect 12357 1853 12391 1887
rect 12391 1853 12400 1887
rect 12348 1844 12400 1853
rect 12440 1844 12492 1896
rect 13360 1912 13412 1964
rect 13636 1955 13688 1964
rect 13636 1921 13645 1955
rect 13645 1921 13679 1955
rect 13679 1921 13688 1955
rect 13636 1912 13688 1921
rect 10140 1751 10192 1760
rect 10140 1717 10149 1751
rect 10149 1717 10183 1751
rect 10183 1717 10192 1751
rect 10140 1708 10192 1717
rect 10876 1776 10928 1828
rect 12164 1776 12216 1828
rect 10692 1708 10744 1760
rect 10968 1708 11020 1760
rect 12624 1751 12676 1760
rect 12624 1717 12633 1751
rect 12633 1717 12667 1751
rect 12667 1717 12676 1751
rect 12624 1708 12676 1717
rect 13176 1776 13228 1828
rect 13912 1955 13964 1964
rect 13912 1921 13921 1955
rect 13921 1921 13955 1955
rect 13955 1921 13964 1955
rect 13912 1912 13964 1921
rect 15108 1955 15160 1964
rect 15108 1921 15117 1955
rect 15117 1921 15151 1955
rect 15151 1921 15160 1955
rect 15108 1912 15160 1921
rect 15660 1912 15712 1964
rect 13820 1887 13872 1896
rect 13820 1853 13829 1887
rect 13829 1853 13863 1887
rect 13863 1853 13872 1887
rect 13820 1844 13872 1853
rect 14556 1844 14608 1896
rect 14924 1844 14976 1896
rect 15016 1887 15068 1896
rect 15016 1853 15025 1887
rect 15025 1853 15059 1887
rect 15059 1853 15068 1887
rect 15016 1844 15068 1853
rect 15384 1844 15436 1896
rect 16488 2048 16540 2100
rect 16580 1980 16632 2032
rect 15568 1708 15620 1760
rect 15660 1751 15712 1760
rect 15660 1717 15669 1751
rect 15669 1717 15703 1751
rect 15703 1717 15712 1751
rect 15660 1708 15712 1717
rect 15936 1819 15988 1828
rect 15936 1785 15945 1819
rect 15945 1785 15979 1819
rect 15979 1785 15988 1819
rect 15936 1776 15988 1785
rect 16028 1819 16080 1828
rect 16028 1785 16037 1819
rect 16037 1785 16071 1819
rect 16071 1785 16080 1819
rect 16028 1776 16080 1785
rect 17040 1887 17092 1896
rect 17040 1853 17049 1887
rect 17049 1853 17083 1887
rect 17083 1853 17092 1887
rect 17040 1844 17092 1853
rect 17316 1887 17368 1896
rect 17316 1853 17319 1887
rect 17319 1853 17353 1887
rect 17353 1853 17368 1887
rect 16488 1708 16540 1760
rect 17316 1844 17368 1853
rect 4366 1606 4418 1658
rect 4430 1606 4482 1658
rect 4494 1606 4546 1658
rect 4558 1606 4610 1658
rect 4622 1606 4674 1658
rect 4686 1606 4738 1658
rect 10366 1606 10418 1658
rect 10430 1606 10482 1658
rect 10494 1606 10546 1658
rect 10558 1606 10610 1658
rect 10622 1606 10674 1658
rect 10686 1606 10738 1658
rect 16366 1606 16418 1658
rect 16430 1606 16482 1658
rect 16494 1606 16546 1658
rect 16558 1606 16610 1658
rect 16622 1606 16674 1658
rect 16686 1606 16738 1658
rect 1216 1504 1268 1556
rect 1768 1504 1820 1556
rect 2044 1504 2096 1556
rect 2688 1504 2740 1556
rect 3332 1504 3384 1556
rect 3516 1504 3568 1556
rect 4804 1504 4856 1556
rect 5816 1504 5868 1556
rect 6920 1504 6972 1556
rect 7012 1547 7064 1556
rect 7012 1513 7021 1547
rect 7021 1513 7055 1547
rect 7055 1513 7064 1547
rect 7012 1504 7064 1513
rect 7656 1504 7708 1556
rect 7840 1504 7892 1556
rect 1952 1436 2004 1488
rect 2504 1368 2556 1420
rect 3792 1479 3844 1488
rect 3792 1445 3801 1479
rect 3801 1445 3835 1479
rect 3835 1445 3844 1479
rect 3792 1436 3844 1445
rect 2964 1368 3016 1420
rect 3700 1368 3752 1420
rect 3976 1411 4028 1420
rect 3976 1377 3985 1411
rect 3985 1377 4019 1411
rect 4019 1377 4028 1411
rect 3976 1368 4028 1377
rect 4068 1411 4120 1420
rect 4068 1377 4077 1411
rect 4077 1377 4111 1411
rect 4111 1377 4120 1411
rect 4068 1368 4120 1377
rect 4252 1368 4304 1420
rect 4896 1436 4948 1488
rect 4804 1411 4856 1420
rect 4804 1377 4813 1411
rect 4813 1377 4847 1411
rect 4847 1377 4856 1411
rect 4804 1368 4856 1377
rect 3424 1343 3476 1352
rect 3424 1309 3433 1343
rect 3433 1309 3467 1343
rect 3467 1309 3476 1343
rect 3424 1300 3476 1309
rect 3608 1300 3660 1352
rect 5540 1411 5592 1420
rect 5540 1377 5549 1411
rect 5549 1377 5583 1411
rect 5583 1377 5592 1411
rect 5540 1368 5592 1377
rect 5908 1368 5960 1420
rect 6368 1368 6420 1420
rect 3240 1232 3292 1284
rect 6644 1300 6696 1352
rect 7104 1368 7156 1420
rect 7564 1368 7616 1420
rect 8116 1504 8168 1556
rect 9772 1504 9824 1556
rect 10048 1504 10100 1556
rect 8024 1436 8076 1488
rect 8484 1436 8536 1488
rect 8944 1436 8996 1488
rect 7748 1343 7800 1352
rect 7748 1309 7757 1343
rect 7757 1309 7791 1343
rect 7791 1309 7800 1343
rect 7748 1300 7800 1309
rect 1124 1207 1176 1216
rect 1124 1173 1133 1207
rect 1133 1173 1167 1207
rect 1167 1173 1176 1207
rect 1124 1164 1176 1173
rect 1768 1164 1820 1216
rect 2780 1207 2832 1216
rect 2780 1173 2789 1207
rect 2789 1173 2823 1207
rect 2823 1173 2832 1207
rect 2780 1164 2832 1173
rect 3608 1164 3660 1216
rect 5356 1207 5408 1216
rect 5356 1173 5365 1207
rect 5365 1173 5399 1207
rect 5399 1173 5408 1207
rect 5356 1164 5408 1173
rect 5816 1207 5868 1216
rect 5816 1173 5825 1207
rect 5825 1173 5859 1207
rect 5859 1173 5868 1207
rect 5816 1164 5868 1173
rect 6368 1164 6420 1216
rect 6644 1207 6696 1216
rect 6644 1173 6653 1207
rect 6653 1173 6687 1207
rect 6687 1173 6696 1207
rect 6644 1164 6696 1173
rect 6736 1207 6788 1216
rect 6736 1173 6745 1207
rect 6745 1173 6779 1207
rect 6779 1173 6788 1207
rect 6736 1164 6788 1173
rect 6828 1164 6880 1216
rect 8484 1300 8536 1352
rect 9220 1411 9272 1420
rect 9220 1377 9229 1411
rect 9229 1377 9263 1411
rect 9263 1377 9272 1411
rect 9220 1368 9272 1377
rect 9312 1343 9364 1352
rect 9312 1309 9321 1343
rect 9321 1309 9355 1343
rect 9355 1309 9364 1343
rect 9312 1300 9364 1309
rect 9772 1411 9824 1420
rect 9772 1377 9781 1411
rect 9781 1377 9815 1411
rect 9815 1377 9824 1411
rect 9772 1368 9824 1377
rect 10048 1411 10100 1420
rect 10048 1377 10057 1411
rect 10057 1377 10091 1411
rect 10091 1377 10100 1411
rect 10048 1368 10100 1377
rect 12440 1504 12492 1556
rect 12532 1504 12584 1556
rect 13452 1504 13504 1556
rect 10692 1436 10744 1488
rect 10508 1343 10560 1352
rect 10508 1309 10517 1343
rect 10517 1309 10551 1343
rect 10551 1309 10560 1343
rect 10508 1300 10560 1309
rect 10968 1343 11020 1352
rect 10968 1309 10977 1343
rect 10977 1309 11011 1343
rect 11011 1309 11020 1343
rect 10968 1300 11020 1309
rect 11060 1300 11112 1352
rect 11428 1436 11480 1488
rect 12072 1343 12124 1352
rect 12072 1309 12081 1343
rect 12081 1309 12115 1343
rect 12115 1309 12124 1343
rect 12072 1300 12124 1309
rect 12164 1300 12216 1352
rect 8852 1275 8904 1284
rect 8852 1241 8861 1275
rect 8861 1241 8895 1275
rect 8895 1241 8904 1275
rect 8852 1232 8904 1241
rect 8944 1232 8996 1284
rect 8392 1164 8444 1216
rect 10048 1232 10100 1284
rect 13176 1479 13228 1488
rect 13176 1445 13185 1479
rect 13185 1445 13219 1479
rect 13219 1445 13228 1479
rect 13176 1436 13228 1445
rect 13268 1436 13320 1488
rect 12716 1368 12768 1420
rect 12900 1368 12952 1420
rect 12992 1411 13044 1420
rect 12992 1377 13001 1411
rect 13001 1377 13035 1411
rect 13035 1377 13044 1411
rect 12992 1368 13044 1377
rect 13360 1411 13412 1420
rect 13360 1377 13369 1411
rect 13369 1377 13403 1411
rect 13403 1377 13412 1411
rect 13360 1368 13412 1377
rect 13912 1411 13964 1420
rect 13912 1377 13921 1411
rect 13921 1377 13955 1411
rect 13955 1377 13964 1411
rect 13912 1368 13964 1377
rect 14096 1411 14148 1420
rect 14096 1377 14105 1411
rect 14105 1377 14139 1411
rect 14139 1377 14148 1411
rect 14096 1368 14148 1377
rect 14372 1411 14424 1420
rect 14372 1377 14381 1411
rect 14381 1377 14415 1411
rect 14415 1377 14424 1411
rect 14372 1368 14424 1377
rect 15292 1504 15344 1556
rect 15476 1504 15528 1556
rect 16028 1504 16080 1556
rect 14740 1368 14792 1420
rect 17224 1436 17276 1488
rect 17408 1436 17460 1488
rect 15108 1368 15160 1420
rect 15752 1368 15804 1420
rect 15936 1368 15988 1420
rect 17040 1411 17092 1420
rect 17040 1377 17049 1411
rect 17049 1377 17083 1411
rect 17083 1377 17092 1411
rect 17040 1368 17092 1377
rect 14096 1232 14148 1284
rect 11520 1164 11572 1216
rect 11612 1207 11664 1216
rect 11612 1173 11621 1207
rect 11621 1173 11655 1207
rect 11655 1173 11664 1207
rect 11612 1164 11664 1173
rect 11888 1164 11940 1216
rect 15200 1232 15252 1284
rect 15384 1232 15436 1284
rect 14924 1164 14976 1216
rect 1366 1062 1418 1114
rect 1430 1062 1482 1114
rect 1494 1062 1546 1114
rect 1558 1062 1610 1114
rect 1622 1062 1674 1114
rect 1686 1062 1738 1114
rect 7366 1062 7418 1114
rect 7430 1062 7482 1114
rect 7494 1062 7546 1114
rect 7558 1062 7610 1114
rect 7622 1062 7674 1114
rect 7686 1062 7738 1114
rect 13366 1062 13418 1114
rect 13430 1062 13482 1114
rect 13494 1062 13546 1114
rect 13558 1062 13610 1114
rect 13622 1062 13674 1114
rect 13686 1062 13738 1114
rect 2504 1003 2556 1012
rect 2504 969 2513 1003
rect 2513 969 2547 1003
rect 2547 969 2556 1003
rect 2504 960 2556 969
rect 5816 960 5868 1012
rect 8852 960 8904 1012
rect 9312 960 9364 1012
rect 9956 960 10008 1012
rect 2044 892 2096 944
rect 2412 824 2464 876
rect 1124 799 1176 808
rect 1124 765 1133 799
rect 1133 765 1167 799
rect 1167 765 1176 799
rect 1124 756 1176 765
rect 1768 756 1820 808
rect 1860 756 1912 808
rect 2320 756 2372 808
rect 4160 756 4212 808
rect 5264 756 5316 808
rect 5356 799 5408 808
rect 5356 765 5365 799
rect 5365 765 5399 799
rect 5399 765 5408 799
rect 5356 756 5408 765
rect 8116 824 8168 876
rect 6092 799 6144 808
rect 6092 765 6101 799
rect 6101 765 6135 799
rect 6135 765 6144 799
rect 6092 756 6144 765
rect 6644 756 6696 808
rect 6736 756 6788 808
rect 8484 799 8536 808
rect 8484 765 8493 799
rect 8493 765 8527 799
rect 8527 765 8536 799
rect 8484 756 8536 765
rect 8116 688 8168 740
rect 9404 892 9456 944
rect 11152 960 11204 1012
rect 11244 960 11296 1012
rect 12808 960 12860 1012
rect 13176 960 13228 1012
rect 14188 960 14240 1012
rect 14280 960 14332 1012
rect 14648 960 14700 1012
rect 15016 960 15068 1012
rect 14004 892 14056 944
rect 17040 1003 17092 1012
rect 17040 969 17049 1003
rect 17049 969 17083 1003
rect 17083 969 17092 1003
rect 17040 960 17092 969
rect 12716 824 12768 876
rect 13360 824 13412 876
rect 17132 824 17184 876
rect 9864 756 9916 808
rect 572 620 624 672
rect 1308 663 1360 672
rect 1308 629 1317 663
rect 1317 629 1351 663
rect 1351 629 1360 663
rect 1308 620 1360 629
rect 2780 620 2832 672
rect 3700 663 3752 672
rect 3700 629 3709 663
rect 3709 629 3743 663
rect 3743 629 3752 663
rect 3700 620 3752 629
rect 4252 620 4304 672
rect 5172 663 5224 672
rect 5172 629 5181 663
rect 5181 629 5215 663
rect 5215 629 5224 663
rect 5172 620 5224 629
rect 5908 663 5960 672
rect 5908 629 5917 663
rect 5917 629 5951 663
rect 5951 629 5960 663
rect 5908 620 5960 629
rect 6644 663 6696 672
rect 6644 629 6653 663
rect 6653 629 6687 663
rect 6687 629 6696 663
rect 6644 620 6696 629
rect 7196 620 7248 672
rect 8392 620 8444 672
rect 10968 799 11020 808
rect 10968 765 10977 799
rect 10977 765 11011 799
rect 11011 765 11020 799
rect 10968 756 11020 765
rect 11796 799 11848 808
rect 11796 765 11805 799
rect 11805 765 11839 799
rect 11839 765 11848 799
rect 11796 756 11848 765
rect 11060 688 11112 740
rect 11152 688 11204 740
rect 12440 799 12492 808
rect 12440 765 12449 799
rect 12449 765 12483 799
rect 12483 765 12492 799
rect 12440 756 12492 765
rect 10140 620 10192 672
rect 11428 663 11480 672
rect 11428 629 11437 663
rect 11437 629 11471 663
rect 11471 629 11480 663
rect 11428 620 11480 629
rect 12348 688 12400 740
rect 13268 756 13320 808
rect 13912 756 13964 808
rect 14096 756 14148 808
rect 14372 756 14424 808
rect 15108 799 15160 808
rect 15108 765 15117 799
rect 15117 765 15151 799
rect 15151 765 15160 799
rect 15108 756 15160 765
rect 15200 756 15252 808
rect 16856 799 16908 808
rect 16856 765 16865 799
rect 16865 765 16899 799
rect 16899 765 16908 799
rect 16856 756 16908 765
rect 12900 620 12952 672
rect 16212 731 16264 740
rect 16212 697 16221 731
rect 16221 697 16255 731
rect 16255 697 16264 731
rect 16212 688 16264 697
rect 16120 620 16172 672
rect 4366 518 4418 570
rect 4430 518 4482 570
rect 4494 518 4546 570
rect 4558 518 4610 570
rect 4622 518 4674 570
rect 4686 518 4738 570
rect 10366 518 10418 570
rect 10430 518 10482 570
rect 10494 518 10546 570
rect 10558 518 10610 570
rect 10622 518 10674 570
rect 10686 518 10738 570
rect 16366 518 16418 570
rect 16430 518 16482 570
rect 16494 518 16546 570
rect 16558 518 16610 570
rect 16622 518 16674 570
rect 16686 518 16738 570
rect 5264 416 5316 468
rect 6092 416 6144 468
rect 12808 416 12860 468
rect 12900 416 12952 468
rect 14372 416 14424 468
rect 14740 416 14792 468
rect 16212 416 16264 468
rect 6368 348 6420 400
rect 9680 348 9732 400
rect 11428 348 11480 400
rect 12532 280 12584 332
rect 7840 212 7892 264
rect 11980 212 12032 264
rect 14096 212 14148 264
rect 4160 144 4212 196
rect 10048 144 10100 196
rect 11520 144 11572 196
<< metal2 >>
rect 1214 17845 1270 18245
rect 2042 17845 2098 18245
rect 2870 17845 2926 18245
rect 3698 17845 3754 18245
rect 4526 17845 4582 18245
rect 5354 17845 5410 18245
rect 6182 17845 6238 18245
rect 7010 17845 7066 18245
rect 7838 17845 7894 18245
rect 8666 17845 8722 18245
rect 9494 17845 9550 18245
rect 10322 17845 10378 18245
rect 11150 17845 11206 18245
rect 11978 17845 12034 18245
rect 12806 17845 12862 18245
rect 13634 17845 13690 18245
rect 14462 17845 14518 18245
rect 15290 17845 15346 18245
rect 16118 17845 16174 18245
rect 16946 17845 17002 18245
rect 1228 17338 1256 17845
rect 1364 17436 1740 17445
rect 1420 17434 1444 17436
rect 1500 17434 1524 17436
rect 1580 17434 1604 17436
rect 1660 17434 1684 17436
rect 1420 17382 1430 17434
rect 1674 17382 1684 17434
rect 1420 17380 1444 17382
rect 1500 17380 1524 17382
rect 1580 17380 1604 17382
rect 1660 17380 1684 17382
rect 1364 17371 1740 17380
rect 2056 17338 2084 17845
rect 2884 17338 2912 17845
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 1216 17332 1268 17338
rect 1216 17274 1268 17280
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2976 17202 3004 17478
rect 3712 17338 3740 17845
rect 4540 17338 4568 17845
rect 5368 17338 5396 17845
rect 6196 17338 6224 17845
rect 7024 17338 7052 17845
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16794 1716 16934
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 2792 16658 2820 17070
rect 3068 16658 3096 17138
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4264 16998 4292 17070
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 3804 16794 3832 16934
rect 4364 16892 4740 16901
rect 4420 16890 4444 16892
rect 4500 16890 4524 16892
rect 4580 16890 4604 16892
rect 4660 16890 4684 16892
rect 4420 16838 4430 16890
rect 4674 16838 4684 16890
rect 4420 16836 4444 16838
rect 4500 16836 4524 16838
rect 4580 16836 4604 16838
rect 4660 16836 4684 16838
rect 4364 16827 4740 16836
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 4908 16697 4936 17070
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 4894 16688 4950 16697
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 3240 16652 3292 16658
rect 4894 16623 4950 16632
rect 3240 16594 3292 16600
rect 848 16584 900 16590
rect 848 16526 900 16532
rect 860 16046 888 16526
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 1364 16348 1740 16357
rect 1420 16346 1444 16348
rect 1500 16346 1524 16348
rect 1580 16346 1604 16348
rect 1660 16346 1684 16348
rect 1420 16294 1430 16346
rect 1674 16294 1684 16346
rect 1420 16292 1444 16294
rect 1500 16292 1524 16294
rect 1580 16292 1604 16294
rect 1660 16292 1684 16294
rect 1364 16283 1740 16292
rect 2792 16114 2820 16390
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 848 16040 900 16046
rect 848 15982 900 15988
rect 860 14958 888 15982
rect 1492 15972 1544 15978
rect 1492 15914 1544 15920
rect 1504 15706 1532 15914
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2042 15736 2098 15745
rect 1492 15700 1544 15706
rect 2608 15706 2636 15846
rect 2042 15671 2044 15680
rect 1492 15642 1544 15648
rect 2096 15671 2098 15680
rect 2596 15700 2648 15706
rect 2044 15642 2096 15648
rect 2596 15642 2648 15648
rect 2056 15570 2084 15642
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 1364 15260 1740 15269
rect 1420 15258 1444 15260
rect 1500 15258 1524 15260
rect 1580 15258 1604 15260
rect 1660 15258 1684 15260
rect 1420 15206 1430 15258
rect 1674 15206 1684 15258
rect 1420 15204 1444 15206
rect 1500 15204 1524 15206
rect 1580 15204 1604 15206
rect 1660 15204 1684 15206
rect 1364 15195 1740 15204
rect 2700 15162 2728 15370
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 848 14952 900 14958
rect 848 14894 900 14900
rect 2686 14920 2742 14929
rect 860 13326 888 14894
rect 1400 14884 1452 14890
rect 2686 14855 2742 14864
rect 1400 14826 1452 14832
rect 1412 14618 1440 14826
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 2056 14482 2084 14758
rect 2700 14482 2728 14855
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1364 14172 1740 14181
rect 1420 14170 1444 14172
rect 1500 14170 1524 14172
rect 1580 14170 1604 14172
rect 1660 14170 1684 14172
rect 1420 14118 1430 14170
rect 1674 14118 1684 14170
rect 1420 14116 1444 14118
rect 1500 14116 1524 14118
rect 1580 14116 1604 14118
rect 1660 14116 1684 14118
rect 1364 14107 1740 14116
rect 1216 13388 1268 13394
rect 1216 13330 1268 13336
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 12238 888 13262
rect 1228 12986 1256 13330
rect 1364 13084 1740 13093
rect 1420 13082 1444 13084
rect 1500 13082 1524 13084
rect 1580 13082 1604 13084
rect 1660 13082 1684 13084
rect 1420 13030 1430 13082
rect 1674 13030 1684 13082
rect 1420 13028 1444 13030
rect 1500 13028 1524 13030
rect 1580 13028 1604 13030
rect 1660 13028 1684 13030
rect 1364 13019 1740 13028
rect 1780 12986 1808 14350
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1872 14006 1900 14214
rect 1860 14000 1912 14006
rect 1860 13942 1912 13948
rect 1216 12980 1268 12986
rect 1216 12922 1268 12928
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1676 12912 1728 12918
rect 1872 12866 1900 13942
rect 2516 13938 2544 14418
rect 2596 14408 2648 14414
rect 2686 14376 2742 14385
rect 2648 14356 2686 14362
rect 2596 14350 2686 14356
rect 2608 14334 2686 14350
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 1728 12860 1900 12866
rect 1676 12854 1900 12860
rect 1688 12838 1900 12854
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1124 12300 1176 12306
rect 1124 12242 1176 12248
rect 848 12232 900 12238
rect 848 12174 900 12180
rect 860 11286 888 12174
rect 1136 11898 1164 12242
rect 1364 11996 1740 12005
rect 1420 11994 1444 11996
rect 1500 11994 1524 11996
rect 1580 11994 1604 11996
rect 1660 11994 1684 11996
rect 1420 11942 1430 11994
rect 1674 11942 1684 11994
rect 1420 11940 1444 11942
rect 1500 11940 1524 11942
rect 1580 11940 1604 11942
rect 1660 11940 1684 11942
rect 1364 11931 1740 11940
rect 1780 11898 1808 12718
rect 1124 11892 1176 11898
rect 1124 11834 1176 11840
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1964 11558 1992 12718
rect 2148 12102 2176 13466
rect 2516 13190 2544 13874
rect 2608 13870 2636 14334
rect 2686 14311 2742 14320
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2608 13462 2636 13806
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 848 11280 900 11286
rect 848 11222 900 11228
rect 1364 10908 1740 10917
rect 1420 10906 1444 10908
rect 1500 10906 1524 10908
rect 1580 10906 1604 10908
rect 1660 10906 1684 10908
rect 1420 10854 1430 10906
rect 1674 10854 1684 10906
rect 1420 10852 1444 10854
rect 1500 10852 1524 10854
rect 1580 10852 1604 10854
rect 1660 10852 1684 10854
rect 1364 10843 1740 10852
rect 1780 10606 1808 11290
rect 1964 11218 1992 11494
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10130 1624 10406
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 848 10056 900 10062
rect 848 9998 900 10004
rect 860 9518 888 9998
rect 1364 9820 1740 9829
rect 1420 9818 1444 9820
rect 1500 9818 1524 9820
rect 1580 9818 1604 9820
rect 1660 9818 1684 9820
rect 1420 9766 1430 9818
rect 1674 9766 1684 9818
rect 1420 9764 1444 9766
rect 1500 9764 1524 9766
rect 1580 9764 1604 9766
rect 1660 9764 1684 9766
rect 1364 9755 1740 9764
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 848 9512 900 9518
rect 848 9454 900 9460
rect 860 9042 888 9454
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 848 9036 900 9042
rect 848 8978 900 8984
rect 860 8498 888 8978
rect 1872 8945 1900 9386
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 1364 8732 1740 8741
rect 1420 8730 1444 8732
rect 1500 8730 1524 8732
rect 1580 8730 1604 8732
rect 1660 8730 1684 8732
rect 1420 8678 1430 8730
rect 1674 8678 1684 8730
rect 1420 8676 1444 8678
rect 1500 8676 1524 8678
rect 1580 8676 1604 8678
rect 1660 8676 1684 8678
rect 1364 8667 1740 8676
rect 848 8492 900 8498
rect 848 8434 900 8440
rect 860 6798 888 8434
rect 1964 7954 1992 9522
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1364 7644 1740 7653
rect 1420 7642 1444 7644
rect 1500 7642 1524 7644
rect 1580 7642 1604 7644
rect 1660 7642 1684 7644
rect 1420 7590 1430 7642
rect 1674 7590 1684 7642
rect 1420 7588 1444 7590
rect 1500 7588 1524 7590
rect 1580 7588 1604 7590
rect 1660 7588 1684 7590
rect 1364 7579 1740 7588
rect 1780 7290 1808 7686
rect 1872 7546 1900 7822
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1964 7546 1992 7754
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1780 7262 1992 7290
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 5710 888 6734
rect 1364 6556 1740 6565
rect 1420 6554 1444 6556
rect 1500 6554 1524 6556
rect 1580 6554 1604 6556
rect 1660 6554 1684 6556
rect 1420 6502 1430 6554
rect 1674 6502 1684 6554
rect 1420 6500 1444 6502
rect 1500 6500 1524 6502
rect 1580 6500 1604 6502
rect 1660 6500 1684 6502
rect 1364 6491 1740 6500
rect 848 5704 900 5710
rect 848 5646 900 5652
rect 860 4078 888 5646
rect 1364 5468 1740 5477
rect 1420 5466 1444 5468
rect 1500 5466 1524 5468
rect 1580 5466 1604 5468
rect 1660 5466 1684 5468
rect 1420 5414 1430 5466
rect 1674 5414 1684 5466
rect 1420 5412 1444 5414
rect 1500 5412 1524 5414
rect 1580 5412 1604 5414
rect 1660 5412 1684 5414
rect 1364 5403 1740 5412
rect 1492 5092 1544 5098
rect 1492 5034 1544 5040
rect 1504 4826 1532 5034
rect 1780 4978 1808 7142
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1872 5914 1900 6802
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1688 4950 1808 4978
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 1688 4486 1716 4950
rect 1872 4826 1900 4966
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1216 4480 1268 4486
rect 1216 4422 1268 4428
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 848 4072 900 4078
rect 848 4014 900 4020
rect 1228 4010 1256 4422
rect 1364 4380 1740 4389
rect 1420 4378 1444 4380
rect 1500 4378 1524 4380
rect 1580 4378 1604 4380
rect 1660 4378 1684 4380
rect 1420 4326 1430 4378
rect 1674 4326 1684 4378
rect 1420 4324 1444 4326
rect 1500 4324 1524 4326
rect 1580 4324 1604 4326
rect 1660 4324 1684 4326
rect 1364 4315 1740 4324
rect 1216 4004 1268 4010
rect 1216 3946 1268 3952
rect 1780 3942 1808 4626
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1364 3292 1740 3301
rect 1420 3290 1444 3292
rect 1500 3290 1524 3292
rect 1580 3290 1604 3292
rect 1660 3290 1684 3292
rect 1420 3238 1430 3290
rect 1674 3238 1684 3290
rect 1420 3236 1444 3238
rect 1500 3236 1524 3238
rect 1580 3236 1604 3238
rect 1660 3236 1684 3238
rect 1364 3227 1740 3236
rect 1306 2544 1362 2553
rect 1228 2502 1306 2530
rect 1228 1562 1256 2502
rect 1780 2514 1808 3878
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1306 2479 1362 2488
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 1364 2204 1740 2213
rect 1420 2202 1444 2204
rect 1500 2202 1524 2204
rect 1580 2202 1604 2204
rect 1660 2202 1684 2204
rect 1420 2150 1430 2202
rect 1674 2150 1684 2202
rect 1420 2148 1444 2150
rect 1500 2148 1524 2150
rect 1580 2148 1604 2150
rect 1660 2148 1684 2150
rect 1364 2139 1740 2148
rect 1780 2106 1808 2314
rect 1768 2100 1820 2106
rect 1768 2042 1820 2048
rect 1872 1902 1900 3334
rect 1964 1902 1992 7262
rect 2056 7206 2084 11630
rect 2148 7970 2176 12038
rect 2240 11132 2268 12174
rect 2332 11234 2360 13126
rect 2424 12782 2452 13126
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2686 12744 2742 12753
rect 2596 12708 2648 12714
rect 2686 12679 2742 12688
rect 2596 12650 2648 12656
rect 2608 11830 2636 12650
rect 2700 11898 2728 12679
rect 2792 12646 2820 15574
rect 2976 15450 3004 16594
rect 3068 16130 3096 16594
rect 3252 16182 3280 16594
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4264 16454 4292 16526
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 3240 16176 3292 16182
rect 3068 16102 3188 16130
rect 3240 16118 3292 16124
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3068 15638 3096 15982
rect 3056 15632 3108 15638
rect 3056 15574 3108 15580
rect 2976 15422 3096 15450
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2884 14618 2912 15302
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2976 14482 3004 15098
rect 3068 14940 3096 15422
rect 3160 15094 3188 16102
rect 3240 15904 3292 15910
rect 3292 15864 3372 15892
rect 3240 15846 3292 15852
rect 3238 15736 3294 15745
rect 3238 15671 3240 15680
rect 3292 15671 3294 15680
rect 3240 15642 3292 15648
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3068 14912 3188 14940
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2884 12889 2912 12922
rect 2870 12880 2926 12889
rect 2870 12815 2926 12824
rect 2976 12764 3004 14214
rect 2884 12736 3004 12764
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2424 11354 2452 11630
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2332 11206 2452 11234
rect 2320 11144 2372 11150
rect 2240 11104 2320 11132
rect 2320 11086 2372 11092
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2332 10606 2360 10950
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2240 8090 2268 9522
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2148 7954 2268 7970
rect 2148 7948 2280 7954
rect 2148 7942 2228 7948
rect 2228 7890 2280 7896
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2134 7848 2190 7857
rect 2134 7783 2190 7792
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5234 2084 6054
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2148 5098 2176 7783
rect 2240 7206 2268 7890
rect 2332 7342 2360 7890
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2424 6914 2452 11206
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2594 9072 2650 9081
rect 2594 9007 2596 9016
rect 2648 9007 2650 9016
rect 2596 8978 2648 8984
rect 2700 8090 2728 9862
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2608 7834 2636 7890
rect 2516 7806 2636 7834
rect 2516 7426 2544 7806
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2608 7546 2636 7686
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2516 7398 2636 7426
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2332 6886 2452 6914
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2240 5574 2268 6122
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2136 5092 2188 5098
rect 2136 5034 2188 5040
rect 2332 4078 2360 6886
rect 2516 6866 2544 7278
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2608 6254 2636 7398
rect 2700 7342 2728 8026
rect 2688 7336 2740 7342
rect 2884 7313 2912 12736
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2976 12442 3004 12582
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 3068 12322 3096 12582
rect 2976 12306 3096 12322
rect 2964 12300 3096 12306
rect 3016 12294 3096 12300
rect 2964 12242 3016 12248
rect 3160 11898 3188 14912
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3160 7954 3188 8570
rect 3252 8090 3280 13126
rect 3344 11830 3372 15864
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 15162 3556 15302
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3528 15026 3556 15098
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3436 14074 3464 14894
rect 3528 14618 3556 14962
rect 3804 14890 3832 15370
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3514 13968 3570 13977
rect 3514 13903 3570 13912
rect 3608 13932 3660 13938
rect 3528 13530 3556 13903
rect 3608 13874 3660 13880
rect 3620 13530 3648 13874
rect 3712 13870 3740 14758
rect 3804 14482 3832 14826
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3896 13870 3924 15438
rect 3988 14958 4016 15642
rect 4264 15570 4292 16390
rect 4632 15978 4660 16390
rect 5368 16046 5396 16390
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4364 15804 4740 15813
rect 4420 15802 4444 15804
rect 4500 15802 4524 15804
rect 4580 15802 4604 15804
rect 4660 15802 4684 15804
rect 4420 15750 4430 15802
rect 4674 15750 4684 15802
rect 4420 15748 4444 15750
rect 4500 15748 4524 15750
rect 4580 15748 4604 15750
rect 4660 15748 4684 15750
rect 4364 15739 4740 15748
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 5092 15694 5396 15722
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4080 15348 4108 15506
rect 4172 15450 4200 15506
rect 4172 15422 4292 15450
rect 4264 15366 4292 15422
rect 4160 15360 4212 15366
rect 4080 15320 4160 15348
rect 4160 15302 4212 15308
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4172 14958 4200 15302
rect 4264 15094 4292 15302
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 3988 14498 4016 14894
rect 4264 14804 4292 15030
rect 4632 14822 4660 15574
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4172 14776 4292 14804
rect 4620 14816 4672 14822
rect 4066 14512 4122 14521
rect 3988 14470 4066 14498
rect 4066 14447 4122 14456
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4172 13852 4200 14776
rect 4620 14758 4672 14764
rect 4364 14716 4740 14725
rect 4420 14714 4444 14716
rect 4500 14714 4524 14716
rect 4580 14714 4604 14716
rect 4660 14714 4684 14716
rect 4420 14662 4430 14714
rect 4674 14662 4684 14714
rect 4420 14660 4444 14662
rect 4500 14660 4524 14662
rect 4580 14660 4604 14662
rect 4660 14660 4684 14662
rect 4364 14651 4740 14660
rect 4528 14544 4580 14550
rect 4526 14512 4528 14521
rect 4580 14512 4582 14521
rect 4526 14447 4582 14456
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4632 14113 4660 14418
rect 4618 14104 4674 14113
rect 4618 14039 4674 14048
rect 4342 13968 4398 13977
rect 4342 13903 4344 13912
rect 4396 13903 4398 13912
rect 4344 13874 4396 13880
rect 4816 13870 4844 15302
rect 4908 15026 4936 15642
rect 4988 15632 5040 15638
rect 5092 15620 5120 15694
rect 5040 15592 5120 15620
rect 5264 15632 5316 15638
rect 4988 15574 5040 15580
rect 5264 15574 5316 15580
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4908 14929 4936 14962
rect 4894 14920 4950 14929
rect 4894 14855 4950 14864
rect 5000 14822 5028 15302
rect 5184 15162 5212 15302
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 5078 15056 5134 15065
rect 5078 14991 5134 15000
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14464 5028 14758
rect 5092 14618 5120 14991
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 5080 14476 5132 14482
rect 5000 14436 5080 14464
rect 5080 14418 5132 14424
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4252 13864 4304 13870
rect 4172 13824 4252 13852
rect 3988 13530 4016 13806
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4080 13433 4108 13806
rect 4066 13424 4122 13433
rect 4066 13359 4122 13368
rect 4172 13308 4200 13824
rect 4252 13806 4304 13812
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4264 13512 4292 13670
rect 4364 13628 4740 13637
rect 4420 13626 4444 13628
rect 4500 13626 4524 13628
rect 4580 13626 4604 13628
rect 4660 13626 4684 13628
rect 4420 13574 4430 13626
rect 4674 13574 4684 13626
rect 4420 13572 4444 13574
rect 4500 13572 4524 13574
rect 4580 13572 4604 13574
rect 4660 13572 4684 13574
rect 4364 13563 4740 13572
rect 4344 13524 4396 13530
rect 4264 13484 4344 13512
rect 4344 13466 4396 13472
rect 3804 13280 4200 13308
rect 4264 13394 4384 13410
rect 4908 13394 4936 14350
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4264 13388 4396 13394
rect 4264 13382 4344 13388
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3528 12442 3556 12650
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3436 11626 3464 12038
rect 3620 11762 3648 12650
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3620 11218 3648 11698
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3332 11008 3384 11014
rect 3700 11008 3752 11014
rect 3384 10968 3464 10996
rect 3332 10950 3384 10956
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2688 7278 2740 7284
rect 2870 7304 2926 7313
rect 2870 7239 2926 7248
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2424 5166 2452 5646
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2516 5012 2544 6054
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2596 5160 2648 5166
rect 2746 5120 3004 5148
rect 2746 5114 2774 5120
rect 2648 5108 2774 5114
rect 2596 5102 2774 5108
rect 2608 5086 2774 5102
rect 2976 5030 3004 5120
rect 2596 5024 2648 5030
rect 2516 4992 2596 5012
rect 2688 5024 2740 5030
rect 2648 4992 2650 5001
rect 2516 4984 2594 4992
rect 2688 4966 2740 4972
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2594 4927 2650 4936
rect 2700 4826 2728 4966
rect 3068 4826 3096 5714
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 2320 4072 2372 4078
rect 2372 4032 2452 4060
rect 2320 4014 2372 4020
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2332 3738 2360 3878
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 2148 3194 2176 3538
rect 2332 3194 2360 3674
rect 2424 3602 2452 4032
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3670 2728 3878
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2424 3194 2452 3334
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2792 2922 2820 3470
rect 2884 3466 2912 3674
rect 3160 3602 3188 7890
rect 3252 7274 3280 8026
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 4622 3280 5510
rect 3344 5234 3372 5850
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3344 4690 3372 5170
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3436 3942 3464 10968
rect 3700 10950 3752 10956
rect 3712 9897 3740 10950
rect 3804 10033 3832 13280
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4172 12442 4200 12650
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4264 12238 4292 13382
rect 4344 13330 4396 13336
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4632 12918 4660 13330
rect 5000 13258 5028 14010
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 5184 13190 5212 15098
rect 5276 14958 5304 15574
rect 5368 15570 5396 15694
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5276 14618 5304 14758
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5368 14074 5396 14758
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5264 13864 5316 13870
rect 5262 13832 5264 13841
rect 5316 13832 5318 13841
rect 5262 13767 5318 13776
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 5184 12850 5212 13126
rect 5368 12986 5396 13262
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5080 12776 5132 12782
rect 5368 12730 5396 12922
rect 5080 12718 5132 12724
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4364 12540 4740 12549
rect 4420 12538 4444 12540
rect 4500 12538 4524 12540
rect 4580 12538 4604 12540
rect 4660 12538 4684 12540
rect 4420 12486 4430 12538
rect 4674 12486 4684 12538
rect 4420 12484 4444 12486
rect 4500 12484 4524 12486
rect 4580 12484 4604 12486
rect 4660 12484 4684 12486
rect 4364 12475 4740 12484
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4264 11744 4292 12174
rect 4908 12102 4936 12582
rect 5092 12434 5120 12718
rect 5000 12406 5120 12434
rect 5184 12702 5396 12730
rect 5184 12434 5212 12702
rect 5460 12594 5488 16934
rect 6380 16794 6408 16934
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 5552 15978 5580 16730
rect 6472 16674 6500 17002
rect 6564 16794 6592 17002
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6276 16652 6328 16658
rect 6472 16646 6592 16674
rect 6276 16594 6328 16600
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5552 15026 5580 15914
rect 5644 15366 5672 15914
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5736 15570 5764 15846
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5644 14550 5672 15302
rect 5828 14958 5856 15642
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5552 14362 5580 14486
rect 5828 14482 5856 14894
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5552 14334 5672 14362
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5368 12566 5488 12594
rect 5184 12406 5304 12434
rect 5000 12170 5028 12406
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4172 11716 4292 11744
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3882 10976 3938 10985
rect 3882 10911 3938 10920
rect 3896 10130 3924 10911
rect 3988 10266 4016 11630
rect 4172 11558 4200 11716
rect 4344 11688 4396 11694
rect 4264 11648 4344 11676
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4172 11286 4200 11494
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4080 10849 4108 11222
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4066 10840 4122 10849
rect 4066 10775 4122 10784
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4080 10130 4108 10610
rect 4172 10266 4200 11086
rect 4264 10810 4292 11648
rect 4344 11630 4396 11636
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4364 11452 4740 11461
rect 4420 11450 4444 11452
rect 4500 11450 4524 11452
rect 4580 11450 4604 11452
rect 4660 11450 4684 11452
rect 4420 11398 4430 11450
rect 4674 11398 4684 11450
rect 4420 11396 4444 11398
rect 4500 11396 4524 11398
rect 4580 11396 4604 11398
rect 4660 11396 4684 11398
rect 4364 11387 4740 11396
rect 4816 11354 4844 11630
rect 4988 11552 5040 11558
rect 4908 11512 4988 11540
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4356 10742 4384 11290
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4620 10600 4672 10606
rect 4618 10568 4620 10577
rect 4672 10568 4674 10577
rect 4618 10503 4674 10512
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3790 10024 3846 10033
rect 3790 9959 3846 9968
rect 4172 9926 4200 10202
rect 4264 9994 4292 10406
rect 4364 10364 4740 10373
rect 4420 10362 4444 10364
rect 4500 10362 4524 10364
rect 4580 10362 4604 10364
rect 4660 10362 4684 10364
rect 4420 10310 4430 10362
rect 4674 10310 4684 10362
rect 4420 10308 4444 10310
rect 4500 10308 4524 10310
rect 4580 10308 4604 10310
rect 4660 10308 4684 10310
rect 4364 10299 4740 10308
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4342 10160 4398 10169
rect 4342 10095 4398 10104
rect 4356 10062 4384 10095
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4618 10024 4674 10033
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4160 9920 4212 9926
rect 3698 9888 3754 9897
rect 4160 9862 4212 9868
rect 3698 9823 3754 9832
rect 4172 9722 4200 9862
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 3884 9648 3936 9654
rect 3514 9616 3570 9625
rect 4356 9602 4384 9998
rect 4724 10010 4752 10202
rect 4816 10130 4844 11154
rect 4908 10146 4936 11512
rect 4988 11494 5040 11500
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5000 10266 5028 11154
rect 5092 11121 5120 11154
rect 5078 11112 5134 11121
rect 5276 11098 5304 12406
rect 5368 11558 5396 12566
rect 5552 12434 5580 14214
rect 5644 13394 5672 14334
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 14074 5856 14214
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5552 12406 5672 12434
rect 5644 11880 5672 12406
rect 5736 12374 5764 13194
rect 5920 12986 5948 16594
rect 6012 15162 6040 16594
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 15910 6224 16526
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6196 15026 6224 15846
rect 6288 15706 6316 16594
rect 6458 16552 6514 16561
rect 6368 16516 6420 16522
rect 6458 16487 6514 16496
rect 6368 16458 6420 16464
rect 6380 15706 6408 16458
rect 6472 16114 6500 16487
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6288 15065 6316 15506
rect 6274 15056 6330 15065
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 6184 15020 6236 15026
rect 6274 14991 6330 15000
rect 6184 14962 6236 14968
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 13734 6040 14758
rect 6104 13938 6132 14962
rect 6276 14952 6328 14958
rect 6196 14900 6276 14906
rect 6196 14894 6328 14900
rect 6366 14920 6422 14929
rect 6196 14878 6316 14894
rect 6196 13977 6224 14878
rect 6366 14855 6368 14864
rect 6420 14855 6422 14864
rect 6368 14826 6420 14832
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6182 13968 6238 13977
rect 6092 13932 6144 13938
rect 6182 13903 6238 13912
rect 6092 13874 6144 13880
rect 6000 13728 6052 13734
rect 5998 13696 6000 13705
rect 6052 13696 6054 13705
rect 5998 13631 6054 13640
rect 6196 13546 6224 13903
rect 6288 13870 6316 14486
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6380 13802 6408 14350
rect 6472 14006 6500 15574
rect 6564 15473 6592 16646
rect 6748 16250 6776 17206
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 6840 16250 6868 17070
rect 7012 16584 7064 16590
rect 6932 16532 7012 16538
rect 6932 16526 7064 16532
rect 6932 16510 7052 16526
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6644 15496 6696 15502
rect 6550 15464 6606 15473
rect 6644 15438 6696 15444
rect 6550 15399 6606 15408
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6564 14958 6592 15098
rect 6656 15094 6684 15438
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6366 13560 6422 13569
rect 6196 13518 6366 13546
rect 6366 13495 6422 13504
rect 6368 13456 6420 13462
rect 6090 13424 6146 13433
rect 6368 13398 6420 13404
rect 6090 13359 6092 13368
rect 6144 13359 6146 13368
rect 6092 13330 6144 13336
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6276 12776 6328 12782
rect 6380 12753 6408 13398
rect 6276 12718 6328 12724
rect 6366 12744 6422 12753
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 6196 12306 6224 12650
rect 6288 12481 6316 12718
rect 6366 12679 6422 12688
rect 6274 12472 6330 12481
rect 6274 12407 6330 12416
rect 6472 12374 6500 13942
rect 6564 12850 6592 14758
rect 6656 14074 6684 15030
rect 6932 14958 6960 16510
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6656 12322 6684 12786
rect 6748 12714 6776 14894
rect 6828 14408 6880 14414
rect 6880 14368 6960 14396
rect 6828 14350 6880 14356
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6840 13462 6868 14010
rect 6932 13530 6960 14368
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6932 13297 6960 13330
rect 6918 13288 6974 13297
rect 6918 13223 6974 13232
rect 7024 12986 7052 16390
rect 7116 15337 7144 17070
rect 7208 16250 7236 17478
rect 7300 17320 7328 17546
rect 7364 17436 7740 17445
rect 7420 17434 7444 17436
rect 7500 17434 7524 17436
rect 7580 17434 7604 17436
rect 7660 17434 7684 17436
rect 7420 17382 7430 17434
rect 7674 17382 7684 17434
rect 7420 17380 7444 17382
rect 7500 17380 7524 17382
rect 7580 17380 7604 17382
rect 7660 17380 7684 17382
rect 7364 17371 7740 17380
rect 7852 17338 7880 17845
rect 8680 17338 8708 17845
rect 7840 17332 7892 17338
rect 7300 17292 7420 17320
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7300 16250 7328 17138
rect 7392 16561 7420 17292
rect 7840 17274 7892 17280
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 9508 17134 9536 17845
rect 10336 17134 10364 17845
rect 11164 17338 11192 17845
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11440 17134 11468 17478
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 7378 16552 7434 16561
rect 7378 16487 7380 16496
rect 7432 16487 7434 16496
rect 7380 16458 7432 16464
rect 7364 16348 7740 16357
rect 7420 16346 7444 16348
rect 7500 16346 7524 16348
rect 7580 16346 7604 16348
rect 7660 16346 7684 16348
rect 7420 16294 7430 16346
rect 7674 16294 7684 16346
rect 7420 16292 7444 16294
rect 7500 16292 7524 16294
rect 7580 16292 7604 16294
rect 7660 16292 7684 16294
rect 7364 16283 7740 16292
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7944 16130 7972 17070
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8588 16454 8616 16934
rect 9048 16697 9076 17070
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 9324 16794 9352 16934
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9220 16720 9272 16726
rect 9034 16688 9090 16697
rect 9416 16674 9444 16934
rect 9272 16668 9444 16674
rect 9220 16662 9444 16668
rect 9232 16646 9444 16662
rect 10060 16658 10088 16934
rect 10152 16794 10180 16934
rect 10364 16892 10740 16901
rect 10420 16890 10444 16892
rect 10500 16890 10524 16892
rect 10580 16890 10604 16892
rect 10660 16890 10684 16892
rect 10420 16838 10430 16890
rect 10674 16838 10684 16890
rect 10420 16836 10444 16838
rect 10500 16836 10524 16838
rect 10580 16836 10604 16838
rect 10660 16836 10684 16838
rect 10364 16827 10740 16836
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 9034 16623 9090 16632
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 7944 16102 8156 16130
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 15638 7512 15846
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7102 15328 7158 15337
rect 7102 15263 7158 15272
rect 7102 15056 7158 15065
rect 7208 15042 7236 15438
rect 7158 15014 7236 15042
rect 7102 14991 7158 15000
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7012 12980 7064 12986
rect 6932 12940 7012 12968
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6840 12442 6868 12650
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5644 11852 6040 11880
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5814 11248 5870 11257
rect 5814 11183 5816 11192
rect 5868 11183 5870 11192
rect 5816 11154 5868 11160
rect 5724 11144 5776 11150
rect 5078 11047 5134 11056
rect 5172 11076 5224 11082
rect 5276 11070 5488 11098
rect 5724 11086 5776 11092
rect 5172 11018 5224 11024
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 10266 5120 10542
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4804 10124 4856 10130
rect 4908 10118 5028 10146
rect 4804 10066 4856 10072
rect 4724 9982 4936 10010
rect 4618 9959 4674 9968
rect 4526 9888 4582 9897
rect 4526 9823 4582 9832
rect 3936 9596 4384 9602
rect 3884 9590 4384 9596
rect 3896 9574 4384 9590
rect 3514 9551 3516 9560
rect 3568 9551 3570 9560
rect 3516 9522 3568 9528
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3804 9042 3832 9454
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3896 8430 3924 9386
rect 3988 8498 4016 9574
rect 4540 9518 4568 9823
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3516 7812 3568 7818
rect 3516 7754 3568 7760
rect 3528 6934 3556 7754
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 5778 3648 6598
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3712 5710 3740 6394
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3528 5098 3556 5646
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3620 5166 3648 5578
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3516 5092 3568 5098
rect 3516 5034 3568 5040
rect 3528 4622 3556 5034
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3528 4078 3556 4422
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3804 3652 3832 8298
rect 4080 7954 4108 9454
rect 4172 9178 4200 9454
rect 4632 9450 4660 9959
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4364 9276 4740 9285
rect 4420 9274 4444 9276
rect 4500 9274 4524 9276
rect 4580 9274 4604 9276
rect 4660 9274 4684 9276
rect 4420 9222 4430 9274
rect 4674 9222 4684 9274
rect 4420 9220 4444 9222
rect 4500 9220 4524 9222
rect 4580 9220 4604 9222
rect 4660 9220 4684 9222
rect 4364 9211 4740 9220
rect 4160 9172 4212 9178
rect 4212 9132 4292 9160
rect 4160 9114 4212 9120
rect 4264 8090 4292 9132
rect 4816 8974 4844 9862
rect 4908 9466 4936 9982
rect 5000 9602 5028 10118
rect 5080 10124 5132 10130
rect 5184 10112 5212 11018
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5262 10704 5318 10713
rect 5262 10639 5264 10648
rect 5316 10639 5318 10648
rect 5264 10610 5316 10616
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5276 10130 5304 10474
rect 5368 10470 5396 10950
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10266 5396 10406
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5132 10084 5212 10112
rect 5264 10124 5316 10130
rect 5080 10066 5132 10072
rect 5264 10066 5316 10072
rect 5172 9988 5224 9994
rect 5172 9930 5224 9936
rect 5000 9574 5120 9602
rect 5184 9586 5212 9930
rect 5276 9722 5304 10066
rect 5460 10010 5488 11070
rect 5540 11008 5592 11014
rect 5538 10976 5540 10985
rect 5592 10976 5594 10985
rect 5538 10911 5594 10920
rect 5736 10690 5764 11086
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5368 9982 5488 10010
rect 5552 10662 5764 10690
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 4908 9438 5028 9466
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 9178 4936 9318
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4364 8188 4740 8197
rect 4420 8186 4444 8188
rect 4500 8186 4524 8188
rect 4580 8186 4604 8188
rect 4660 8186 4684 8188
rect 4420 8134 4430 8186
rect 4674 8134 4684 8186
rect 4420 8132 4444 8134
rect 4500 8132 4524 8134
rect 4580 8132 4604 8134
rect 4660 8132 4684 8134
rect 4364 8123 4740 8132
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4896 7948 4948 7954
rect 5000 7936 5028 9438
rect 4948 7908 5028 7936
rect 4896 7890 4948 7896
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7342 4016 7754
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3896 7002 3924 7210
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3896 6866 3924 6938
rect 4172 6934 4200 7414
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3988 5778 4016 5850
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3896 5030 3924 5102
rect 3988 5098 4016 5714
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4078 3924 4966
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3528 3624 3832 3652
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2038 2084 2790
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2044 2032 2096 2038
rect 2044 1974 2096 1980
rect 1860 1896 1912 1902
rect 1766 1864 1822 1873
rect 1860 1838 1912 1844
rect 1952 1896 2004 1902
rect 1952 1838 2004 1844
rect 1766 1799 1822 1808
rect 1780 1562 1808 1799
rect 1860 1760 1912 1766
rect 1860 1702 1912 1708
rect 1216 1556 1268 1562
rect 1216 1498 1268 1504
rect 1768 1556 1820 1562
rect 1768 1498 1820 1504
rect 1124 1216 1176 1222
rect 1124 1158 1176 1164
rect 1768 1216 1820 1222
rect 1768 1158 1820 1164
rect 1136 814 1164 1158
rect 1364 1116 1740 1125
rect 1420 1114 1444 1116
rect 1500 1114 1524 1116
rect 1580 1114 1604 1116
rect 1660 1114 1684 1116
rect 1420 1062 1430 1114
rect 1674 1062 1684 1114
rect 1420 1060 1444 1062
rect 1500 1060 1524 1062
rect 1580 1060 1604 1062
rect 1660 1060 1684 1062
rect 1364 1051 1740 1060
rect 1780 814 1808 1158
rect 1872 814 1900 1702
rect 1964 1494 1992 1838
rect 2056 1562 2084 1974
rect 2320 1896 2372 1902
rect 2320 1838 2372 1844
rect 2688 1896 2740 1902
rect 2688 1838 2740 1844
rect 2044 1556 2096 1562
rect 2044 1498 2096 1504
rect 1952 1488 2004 1494
rect 1952 1430 2004 1436
rect 2044 944 2096 950
rect 2044 886 2096 892
rect 1124 808 1176 814
rect 1124 750 1176 756
rect 1768 808 1820 814
rect 1768 750 1820 756
rect 1860 808 1912 814
rect 1860 750 1912 756
rect 572 672 624 678
rect 572 614 624 620
rect 1308 672 1360 678
rect 1308 614 1360 620
rect 584 400 612 614
rect 1320 400 1348 614
rect 2056 400 2084 886
rect 2332 814 2360 1838
rect 2412 1760 2464 1766
rect 2412 1702 2464 1708
rect 2424 882 2452 1702
rect 2700 1562 2728 1838
rect 2976 1766 3004 2450
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3252 1834 3280 2314
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 2106 3372 2246
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 3240 1828 3292 1834
rect 3240 1770 3292 1776
rect 2780 1760 2832 1766
rect 2780 1702 2832 1708
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 2688 1556 2740 1562
rect 2688 1498 2740 1504
rect 2504 1420 2556 1426
rect 2504 1362 2556 1368
rect 2516 1018 2544 1362
rect 2792 1222 2820 1702
rect 2976 1426 3004 1702
rect 2964 1420 3016 1426
rect 2964 1362 3016 1368
rect 3252 1290 3280 1770
rect 3332 1760 3384 1766
rect 3332 1702 3384 1708
rect 3344 1562 3372 1702
rect 3332 1556 3384 1562
rect 3332 1498 3384 1504
rect 3436 1358 3464 2586
rect 3528 2553 3556 3624
rect 3896 3534 3924 4014
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 4080 2938 4108 6666
rect 4264 6662 4292 7482
rect 4356 7274 4384 7890
rect 4908 7342 4936 7890
rect 5000 7750 5028 7908
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4364 7100 4740 7109
rect 4420 7098 4444 7100
rect 4500 7098 4524 7100
rect 4580 7098 4604 7100
rect 4660 7098 4684 7100
rect 4420 7046 4430 7098
rect 4674 7046 4684 7098
rect 4420 7044 4444 7046
rect 4500 7044 4524 7046
rect 4580 7044 4604 7046
rect 4660 7044 4684 7046
rect 4364 7035 4740 7044
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4356 6866 4384 6938
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 6100 4384 6598
rect 4264 6072 4384 6100
rect 4160 5024 4212 5030
rect 4158 4992 4160 5001
rect 4212 4992 4214 5001
rect 4158 4927 4214 4936
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4172 3602 4200 4218
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4264 3058 4292 6072
rect 4364 6012 4740 6021
rect 4420 6010 4444 6012
rect 4500 6010 4524 6012
rect 4580 6010 4604 6012
rect 4660 6010 4684 6012
rect 4420 5958 4430 6010
rect 4674 5958 4684 6010
rect 4420 5956 4444 5958
rect 4500 5956 4524 5958
rect 4580 5956 4604 5958
rect 4660 5956 4684 5958
rect 4364 5947 4740 5956
rect 4364 4924 4740 4933
rect 4420 4922 4444 4924
rect 4500 4922 4524 4924
rect 4580 4922 4604 4924
rect 4660 4922 4684 4924
rect 4420 4870 4430 4922
rect 4674 4870 4684 4922
rect 4420 4868 4444 4870
rect 4500 4868 4524 4870
rect 4580 4868 4604 4870
rect 4660 4868 4684 4870
rect 4364 4859 4740 4868
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4724 4214 4752 4490
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4364 3836 4740 3845
rect 4420 3834 4444 3836
rect 4500 3834 4524 3836
rect 4580 3834 4604 3836
rect 4660 3834 4684 3836
rect 4420 3782 4430 3834
rect 4674 3782 4684 3834
rect 4420 3780 4444 3782
rect 4500 3780 4524 3782
rect 4580 3780 4604 3782
rect 4660 3780 4684 3782
rect 4364 3771 4740 3780
rect 4434 3360 4490 3369
rect 4434 3295 4490 3304
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4448 2990 4476 3295
rect 4816 3194 4844 6666
rect 4908 5710 4936 7142
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4896 5160 4948 5166
rect 5000 5137 5028 7482
rect 4896 5102 4948 5108
rect 4986 5128 5042 5137
rect 4908 4690 4936 5102
rect 4986 5063 5042 5072
rect 5000 4690 5028 5063
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4908 4593 4936 4626
rect 4894 4584 4950 4593
rect 4894 4519 4950 4528
rect 4894 4040 4950 4049
rect 4894 3975 4950 3984
rect 4908 3942 4936 3975
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 5000 3670 5028 4626
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 3712 2922 4108 2938
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 3712 2916 4120 2922
rect 3712 2910 4068 2916
rect 3608 2576 3660 2582
rect 3514 2544 3570 2553
rect 3608 2518 3660 2524
rect 3514 2479 3570 2488
rect 3528 2446 3556 2479
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3516 2032 3568 2038
rect 3620 2020 3648 2518
rect 3712 2514 3740 2910
rect 4068 2858 4120 2864
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 3804 2514 3832 2790
rect 4264 2514 4292 2790
rect 4364 2748 4740 2757
rect 4420 2746 4444 2748
rect 4500 2746 4524 2748
rect 4580 2746 4604 2748
rect 4660 2746 4684 2748
rect 4420 2694 4430 2746
rect 4674 2694 4684 2746
rect 4420 2692 4444 2694
rect 4500 2692 4524 2694
rect 4580 2692 4604 2694
rect 4660 2692 4684 2694
rect 4364 2683 4740 2692
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 3568 1992 3648 2020
rect 3516 1974 3568 1980
rect 3516 1896 3568 1902
rect 3516 1838 3568 1844
rect 3528 1562 3556 1838
rect 3516 1556 3568 1562
rect 3516 1498 3568 1504
rect 3620 1358 3648 1992
rect 3712 1426 3740 2450
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4080 1902 4108 2246
rect 4264 1970 4292 2450
rect 4344 2372 4396 2378
rect 4344 2314 4396 2320
rect 4356 1970 4384 2314
rect 4448 1970 4476 2586
rect 4528 2032 4580 2038
rect 4712 2032 4764 2038
rect 4580 1992 4712 2020
rect 4528 1974 4580 1980
rect 4712 1974 4764 1980
rect 4252 1964 4304 1970
rect 4252 1906 4304 1912
rect 4344 1964 4396 1970
rect 4344 1906 4396 1912
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 3884 1896 3936 1902
rect 4068 1896 4120 1902
rect 3884 1838 3936 1844
rect 3988 1856 4068 1884
rect 3804 1494 3832 1838
rect 3792 1488 3844 1494
rect 3792 1430 3844 1436
rect 3700 1420 3752 1426
rect 3700 1362 3752 1368
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 3608 1352 3660 1358
rect 3608 1294 3660 1300
rect 3896 1306 3924 1838
rect 3988 1426 4016 1856
rect 4068 1838 4120 1844
rect 4066 1456 4122 1465
rect 3976 1420 4028 1426
rect 4264 1426 4292 1906
rect 4364 1660 4740 1669
rect 4420 1658 4444 1660
rect 4500 1658 4524 1660
rect 4580 1658 4604 1660
rect 4660 1658 4684 1660
rect 4420 1606 4430 1658
rect 4674 1606 4684 1658
rect 4420 1604 4444 1606
rect 4500 1604 4524 1606
rect 4580 1604 4604 1606
rect 4660 1604 4684 1606
rect 4364 1595 4740 1604
rect 4816 1562 4844 2790
rect 5092 2774 5120 9574
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5184 8294 5212 8910
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 8022 5212 8230
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5184 7410 5212 7958
rect 5276 7954 5304 9454
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5276 7478 5304 7686
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 5234 5212 7142
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5276 5642 5304 6870
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5368 5522 5396 9982
rect 5552 9042 5580 10662
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10130 5764 10406
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5828 9722 5856 10746
rect 5920 10266 5948 11698
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5736 8634 5764 9590
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5552 7954 5580 8570
rect 5908 8560 5960 8566
rect 5828 8508 5908 8514
rect 5828 8502 5960 8508
rect 5828 8486 5948 8502
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7546 5488 7686
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5552 7342 5580 7890
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5644 7154 5672 8366
rect 5828 7546 5856 8486
rect 5908 8424 5960 8430
rect 5906 8392 5908 8401
rect 5960 8392 5962 8401
rect 5906 8327 5962 8336
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 6012 7970 6040 11852
rect 6196 11830 6224 12242
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6090 11520 6146 11529
rect 6090 11455 6146 11464
rect 6104 10062 6132 11455
rect 6196 10441 6224 11562
rect 6380 11150 6408 11698
rect 6472 11694 6500 12310
rect 6656 12306 6776 12322
rect 6656 12300 6788 12306
rect 6656 12294 6736 12300
rect 6736 12242 6788 12248
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10742 6500 10950
rect 6564 10742 6592 12038
rect 6656 11762 6684 12174
rect 6932 11801 6960 12940
rect 7012 12922 7064 12928
rect 7116 12782 7144 14758
rect 7300 14634 7328 15438
rect 7364 15260 7740 15269
rect 7420 15258 7444 15260
rect 7500 15258 7524 15260
rect 7580 15258 7604 15260
rect 7660 15258 7684 15260
rect 7420 15206 7430 15258
rect 7674 15206 7684 15258
rect 7420 15204 7444 15206
rect 7500 15204 7524 15206
rect 7580 15204 7604 15206
rect 7660 15204 7684 15206
rect 7364 15195 7740 15204
rect 7656 15156 7708 15162
rect 7852 15144 7880 15982
rect 7944 15706 7972 15982
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7708 15116 7880 15144
rect 7656 15098 7708 15104
rect 7944 15076 7972 15302
rect 7852 15048 7972 15076
rect 8024 15088 8076 15094
rect 7380 15020 7432 15026
rect 7432 14980 7696 15008
rect 7380 14962 7432 14968
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7208 14606 7328 14634
rect 7392 14618 7420 14758
rect 7668 14618 7696 14980
rect 7748 14952 7800 14958
rect 7746 14920 7748 14929
rect 7800 14920 7802 14929
rect 7746 14855 7802 14864
rect 7380 14612 7432 14618
rect 7208 14074 7236 14606
rect 7380 14554 7432 14560
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7286 14376 7342 14385
rect 7286 14311 7342 14320
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7300 13938 7328 14311
rect 7852 14278 7880 15048
rect 8024 15030 8076 15036
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7364 14172 7740 14181
rect 7420 14170 7444 14172
rect 7500 14170 7524 14172
rect 7580 14170 7604 14172
rect 7660 14170 7684 14172
rect 7420 14118 7430 14170
rect 7674 14118 7684 14170
rect 7420 14116 7444 14118
rect 7500 14116 7524 14118
rect 7580 14116 7604 14118
rect 7660 14116 7684 14118
rect 7364 14107 7740 14116
rect 7838 14104 7894 14113
rect 7484 14048 7838 14056
rect 7484 14039 7894 14048
rect 7484 14028 7880 14039
rect 7484 13977 7512 14028
rect 7470 13968 7526 13977
rect 7288 13932 7340 13938
rect 7470 13903 7526 13912
rect 7654 13968 7710 13977
rect 7654 13903 7710 13912
rect 7288 13874 7340 13880
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7392 13462 7420 13806
rect 7668 13530 7696 13903
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 7760 13172 7788 13806
rect 7852 13326 7880 14028
rect 7944 13870 7972 14486
rect 8036 14074 8064 15030
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7944 13462 7972 13806
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7932 13184 7984 13190
rect 7760 13144 7880 13172
rect 7364 13084 7740 13093
rect 7420 13082 7444 13084
rect 7500 13082 7524 13084
rect 7580 13082 7604 13084
rect 7660 13082 7684 13084
rect 7420 13030 7430 13082
rect 7674 13030 7684 13082
rect 7420 13028 7444 13030
rect 7500 13028 7524 13030
rect 7580 13028 7604 13030
rect 7660 13028 7684 13030
rect 7364 13019 7740 13028
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7852 12646 7880 13144
rect 8128 13172 8156 16102
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8220 14890 8248 15982
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8404 14929 8432 15030
rect 8390 14920 8446 14929
rect 8208 14884 8260 14890
rect 8390 14855 8446 14864
rect 8208 14826 8260 14832
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8312 13938 8340 14418
rect 8404 14249 8432 14418
rect 8390 14240 8446 14249
rect 8390 14175 8446 14184
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 7932 13126 7984 13132
rect 8036 13144 8156 13172
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7840 12640 7892 12646
rect 7944 12617 7972 13126
rect 7840 12582 7892 12588
rect 7930 12608 7986 12617
rect 6918 11792 6974 11801
rect 6644 11756 6696 11762
rect 6918 11727 6974 11736
rect 6644 11698 6696 11704
rect 7024 11694 7052 12582
rect 7930 12543 7986 12552
rect 7930 12472 7986 12481
rect 7930 12407 7932 12416
rect 7984 12407 7986 12416
rect 7932 12378 7984 12384
rect 8036 12322 8064 13144
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7760 12294 8064 12322
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6460 10736 6512 10742
rect 6366 10704 6422 10713
rect 6460 10678 6512 10684
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6366 10639 6368 10648
rect 6420 10639 6422 10648
rect 6368 10610 6420 10616
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6460 10532 6512 10538
rect 6460 10474 6512 10480
rect 6276 10464 6328 10470
rect 6182 10432 6238 10441
rect 6276 10406 6328 10412
rect 6182 10367 6238 10376
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6196 9518 6224 10367
rect 6288 10062 6316 10406
rect 6380 10266 6408 10474
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6472 10010 6500 10474
rect 6472 9982 6592 10010
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6460 9512 6512 9518
rect 6564 9500 6592 9982
rect 6656 9654 6684 11154
rect 6748 11121 6776 11154
rect 6734 11112 6790 11121
rect 6734 11047 6790 11056
rect 6736 11008 6788 11014
rect 6840 10996 6868 11154
rect 6788 10968 6868 10996
rect 6736 10950 6788 10956
rect 6840 10606 6868 10968
rect 6932 10810 6960 11290
rect 7010 10840 7066 10849
rect 6920 10804 6972 10810
rect 7010 10775 7012 10784
rect 6920 10746 6972 10752
rect 7064 10775 7066 10784
rect 7012 10746 7064 10752
rect 7116 10674 7144 12106
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7104 10668 7156 10674
rect 6932 10628 7104 10656
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6644 9512 6696 9518
rect 6564 9472 6644 9500
rect 6460 9454 6512 9460
rect 6644 9454 6696 9460
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6196 9178 6224 9318
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6288 8906 6316 9318
rect 6380 9042 6408 9454
rect 6472 9178 6500 9454
rect 6748 9450 6776 10474
rect 6840 10130 6868 10542
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6826 10024 6882 10033
rect 6826 9959 6882 9968
rect 6840 9654 6868 9959
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6644 9376 6696 9382
rect 6564 9336 6644 9364
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6104 8634 6132 8774
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5920 7546 5948 7958
rect 6012 7942 6224 7970
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5908 7540 5960 7546
rect 5960 7500 6040 7528
rect 5908 7482 5960 7488
rect 5276 5494 5396 5522
rect 5460 7126 5672 7154
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5184 3097 5212 4150
rect 5276 3670 5304 5494
rect 5460 5114 5488 7126
rect 5828 6474 5856 7482
rect 6012 7410 6040 7500
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6012 7002 6040 7346
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5828 6446 5948 6474
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5166 5580 5646
rect 5368 5086 5488 5114
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5368 4026 5396 5086
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5460 4282 5488 4626
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5644 4078 5672 5782
rect 5736 5166 5764 6054
rect 5828 5234 5856 6326
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4072 5684 4078
rect 5368 3998 5488 4026
rect 5632 4014 5684 4020
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5170 3088 5226 3097
rect 5170 3023 5226 3032
rect 5276 2990 5304 3606
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5000 2746 5120 2774
rect 5000 1902 5028 2746
rect 5368 2038 5396 3878
rect 5460 3738 5488 3998
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5552 3890 5580 3946
rect 5736 3942 5764 5102
rect 5828 4826 5856 5170
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5816 4616 5868 4622
rect 5814 4584 5816 4593
rect 5868 4584 5870 4593
rect 5814 4519 5870 4528
rect 5724 3936 5776 3942
rect 5630 3904 5686 3913
rect 5552 3862 5630 3890
rect 5724 3878 5776 3884
rect 5630 3839 5686 3848
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5920 3670 5948 6446
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6012 5098 6040 5170
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 6012 4690 6040 5034
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6104 4622 6132 7822
rect 6196 6118 6224 7942
rect 6380 7206 6408 8978
rect 6458 8936 6514 8945
rect 6458 8871 6514 8880
rect 6472 8838 6500 8871
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6564 8362 6592 9336
rect 6644 9318 6696 9324
rect 6748 9160 6776 9386
rect 6932 9382 6960 10628
rect 7104 10610 7156 10616
rect 7208 10554 7236 12038
rect 7300 11898 7328 12242
rect 7760 12102 7788 12294
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7364 11996 7740 12005
rect 7420 11994 7444 11996
rect 7500 11994 7524 11996
rect 7580 11994 7604 11996
rect 7660 11994 7684 11996
rect 7420 11942 7430 11994
rect 7674 11942 7684 11994
rect 7420 11940 7444 11942
rect 7500 11940 7524 11942
rect 7580 11940 7604 11942
rect 7660 11940 7684 11942
rect 7364 11931 7740 11940
rect 7852 11898 7880 12174
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7286 11792 7342 11801
rect 7286 11727 7342 11736
rect 7654 11792 7710 11801
rect 7654 11727 7710 11736
rect 7300 10690 7328 11727
rect 7668 11694 7696 11727
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7392 11218 7420 11494
rect 7380 11212 7432 11218
rect 7760 11200 7788 11630
rect 7944 11354 7972 12038
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8036 11354 8064 11630
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 8022 11248 8078 11257
rect 7760 11172 7972 11200
rect 8022 11183 8024 11192
rect 7380 11154 7432 11160
rect 7944 11098 7972 11172
rect 8076 11183 8078 11192
rect 8024 11154 8076 11160
rect 8128 11150 8156 12106
rect 8116 11144 8168 11150
rect 7944 11070 8064 11098
rect 8116 11086 8168 11092
rect 7364 10908 7740 10917
rect 7420 10906 7444 10908
rect 7500 10906 7524 10908
rect 7580 10906 7604 10908
rect 7660 10906 7684 10908
rect 7420 10854 7430 10906
rect 7674 10854 7684 10906
rect 7420 10852 7444 10854
rect 7500 10852 7524 10854
rect 7580 10852 7604 10854
rect 7660 10852 7684 10854
rect 7364 10843 7740 10852
rect 8036 10810 8064 11070
rect 8114 10976 8170 10985
rect 8114 10911 8170 10920
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7932 10736 7984 10742
rect 7300 10662 7788 10690
rect 7932 10678 7984 10684
rect 7024 10526 7236 10554
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7380 10532 7432 10538
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6656 9132 6776 9160
rect 6656 8974 6684 9132
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6748 8537 6776 8978
rect 6840 8634 6868 8978
rect 6932 8634 6960 8978
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6734 8528 6790 8537
rect 7024 8514 7052 10526
rect 7380 10474 7432 10480
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 9926 7144 10406
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7208 9738 7236 10066
rect 7392 9908 7420 10474
rect 7484 10198 7512 10542
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7668 10033 7696 10406
rect 7760 10044 7788 10662
rect 7654 10024 7710 10033
rect 7760 10016 7880 10044
rect 7654 9959 7710 9968
rect 7116 9710 7236 9738
rect 7300 9880 7420 9908
rect 7116 8906 7144 9710
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 6734 8463 6736 8472
rect 6788 8463 6790 8472
rect 6932 8486 7052 8514
rect 6736 8434 6788 8440
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6472 6458 6500 7482
rect 6564 7410 6592 7686
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5710 6224 6054
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6012 3738 6040 4014
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5908 3664 5960 3670
rect 5828 3624 5908 3652
rect 5724 3120 5776 3126
rect 5828 3074 5856 3624
rect 5908 3606 5960 3612
rect 6104 3534 6132 4558
rect 6196 3584 6224 5510
rect 6288 5234 6316 6326
rect 6564 5778 6592 6598
rect 6840 6322 6868 7278
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6932 6202 6960 8486
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 7024 8090 7052 8366
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7116 7818 7144 8842
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7208 7290 7236 9590
rect 7300 9382 7328 9880
rect 7364 9820 7740 9829
rect 7420 9818 7444 9820
rect 7500 9818 7524 9820
rect 7580 9818 7604 9820
rect 7660 9818 7684 9820
rect 7420 9766 7430 9818
rect 7674 9766 7684 9818
rect 7420 9764 7444 9766
rect 7500 9764 7524 9766
rect 7580 9764 7604 9766
rect 7660 9764 7684 9766
rect 7364 9755 7740 9764
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9110 7328 9318
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7852 9042 7880 10016
rect 7944 9926 7972 10678
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 8036 9674 8064 10746
rect 8128 10674 8156 10911
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7944 9646 8064 9674
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7300 8344 7328 8910
rect 7364 8732 7740 8741
rect 7420 8730 7444 8732
rect 7500 8730 7524 8732
rect 7580 8730 7604 8732
rect 7660 8730 7684 8732
rect 7420 8678 7430 8730
rect 7674 8678 7684 8730
rect 7420 8676 7444 8678
rect 7500 8676 7524 8678
rect 7580 8676 7604 8678
rect 7660 8676 7684 8678
rect 7364 8667 7740 8676
rect 7852 8634 7880 8978
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7378 8528 7434 8537
rect 7378 8463 7380 8472
rect 7432 8463 7434 8472
rect 7380 8434 7432 8440
rect 7472 8424 7524 8430
rect 7470 8392 7472 8401
rect 7840 8424 7892 8430
rect 7524 8392 7526 8401
rect 7380 8356 7432 8362
rect 7300 8316 7380 8344
rect 7840 8366 7892 8372
rect 7470 8327 7526 8336
rect 7380 8298 7432 8304
rect 7364 7644 7740 7653
rect 7420 7642 7444 7644
rect 7500 7642 7524 7644
rect 7580 7642 7604 7644
rect 7660 7642 7684 7644
rect 7420 7590 7430 7642
rect 7674 7590 7684 7642
rect 7420 7588 7444 7590
rect 7500 7588 7524 7590
rect 7580 7588 7604 7590
rect 7660 7588 7684 7590
rect 7364 7579 7740 7588
rect 7024 7262 7236 7290
rect 7470 7304 7526 7313
rect 7024 6934 7052 7262
rect 7470 7239 7526 7248
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7116 6798 7144 7142
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7024 6458 7052 6734
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7116 6322 7144 6734
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7208 6254 7236 6870
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 6840 6174 6960 6202
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7012 6180 7064 6186
rect 6840 5794 6868 6174
rect 7012 6122 7064 6128
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6748 5766 6868 5794
rect 7024 5778 7052 6122
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7012 5772 7064 5778
rect 6380 5234 6408 5714
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6288 4078 6316 4422
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6196 3556 6316 3584
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5776 3068 5948 3074
rect 5724 3062 5948 3068
rect 5736 3046 5948 3062
rect 5920 2990 5948 3046
rect 6012 2990 6040 3334
rect 6288 2990 6316 3556
rect 6380 2990 6408 3878
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 5736 2378 5764 2926
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 5814 2680 5870 2689
rect 5814 2615 5816 2624
rect 5868 2615 5870 2624
rect 5816 2586 5868 2592
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5356 2032 5408 2038
rect 5356 1974 5408 1980
rect 4988 1896 5040 1902
rect 4986 1864 4988 1873
rect 5040 1864 5042 1873
rect 4986 1799 5042 1808
rect 4896 1760 4948 1766
rect 4896 1702 4948 1708
rect 4804 1556 4856 1562
rect 4804 1498 4856 1504
rect 4908 1494 4936 1702
rect 4896 1488 4948 1494
rect 4802 1456 4858 1465
rect 4066 1391 4068 1400
rect 3976 1362 4028 1368
rect 4120 1391 4122 1400
rect 4252 1420 4304 1426
rect 4068 1362 4120 1368
rect 4896 1430 4948 1436
rect 5552 1426 5580 2246
rect 5828 1562 5856 2586
rect 6196 2514 6224 2790
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 5816 1556 5868 1562
rect 5816 1498 5868 1504
rect 5920 1426 5948 1906
rect 6012 1902 6040 2450
rect 6090 2408 6146 2417
rect 6090 2343 6146 2352
rect 6104 2106 6132 2343
rect 6092 2100 6144 2106
rect 6092 2042 6144 2048
rect 6472 2038 6500 5510
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 6564 4690 6592 5238
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6552 4208 6604 4214
rect 6550 4176 6552 4185
rect 6604 4176 6606 4185
rect 6550 4111 6606 4120
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6564 3126 6592 3538
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6460 2032 6512 2038
rect 6460 1974 6512 1980
rect 6000 1896 6052 1902
rect 6000 1838 6052 1844
rect 6366 1592 6422 1601
rect 6366 1527 6422 1536
rect 6380 1426 6408 1527
rect 4802 1391 4804 1400
rect 4252 1362 4304 1368
rect 4856 1391 4858 1400
rect 5540 1420 5592 1426
rect 4804 1362 4856 1368
rect 5540 1362 5592 1368
rect 5908 1420 5960 1426
rect 5908 1362 5960 1368
rect 6368 1420 6420 1426
rect 6368 1362 6420 1368
rect 4080 1306 4108 1362
rect 6656 1358 6684 4490
rect 6748 3924 6776 5766
rect 7012 5714 7064 5720
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5370 6868 5646
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4570 6960 4966
rect 7010 4720 7066 4729
rect 7010 4655 7066 4664
rect 7024 4622 7052 4655
rect 6840 4542 6960 4570
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6840 4146 6868 4542
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6932 4078 6960 4422
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6748 3896 6960 3924
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3194 6868 3334
rect 6828 3188 6880 3194
rect 6748 3148 6828 3176
rect 6748 1970 6776 3148
rect 6828 3130 6880 3136
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 3240 1284 3292 1290
rect 3240 1226 3292 1232
rect 3620 1222 3648 1294
rect 3896 1278 4108 1306
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6840 1222 6868 2382
rect 6932 1562 6960 3896
rect 7116 3720 7144 5850
rect 7208 4690 7236 6054
rect 7300 5914 7328 6802
rect 7484 6798 7512 7239
rect 7472 6792 7524 6798
rect 7748 6792 7800 6798
rect 7472 6734 7524 6740
rect 7746 6760 7748 6769
rect 7800 6760 7802 6769
rect 7746 6695 7802 6704
rect 7364 6556 7740 6565
rect 7420 6554 7444 6556
rect 7500 6554 7524 6556
rect 7580 6554 7604 6556
rect 7660 6554 7684 6556
rect 7420 6502 7430 6554
rect 7674 6502 7684 6554
rect 7420 6500 7444 6502
rect 7500 6500 7524 6502
rect 7580 6500 7604 6502
rect 7660 6500 7684 6502
rect 7364 6491 7740 6500
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5914 7420 6190
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7300 5148 7328 5646
rect 7364 5468 7740 5477
rect 7420 5466 7444 5468
rect 7500 5466 7524 5468
rect 7580 5466 7604 5468
rect 7660 5466 7684 5468
rect 7420 5414 7430 5466
rect 7674 5414 7684 5466
rect 7420 5412 7444 5414
rect 7500 5412 7524 5414
rect 7580 5412 7604 5414
rect 7660 5412 7684 5414
rect 7364 5403 7740 5412
rect 7380 5160 7432 5166
rect 7300 5120 7380 5148
rect 7564 5160 7616 5166
rect 7380 5102 7432 5108
rect 7562 5128 7564 5137
rect 7616 5128 7618 5137
rect 7562 5063 7618 5072
rect 7288 5024 7340 5030
rect 7852 4978 7880 8366
rect 7944 7478 7972 9646
rect 8128 9625 8156 9998
rect 8114 9616 8170 9625
rect 8114 9551 8170 9560
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 8036 7954 8064 8298
rect 8128 8022 8156 8366
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8128 6934 8156 7278
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 7932 6792 7984 6798
rect 7984 6740 8064 6746
rect 7932 6734 8064 6740
rect 7944 6718 8064 6734
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 5137 7972 6598
rect 8036 6118 8064 6718
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8128 5370 8156 6190
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7930 5128 7986 5137
rect 7930 5063 7986 5072
rect 7288 4966 7340 4972
rect 7300 4826 7328 4966
rect 7576 4950 7880 4978
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7576 4690 7604 4950
rect 7930 4856 7986 4865
rect 7930 4791 7986 4800
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7208 4282 7236 4626
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7024 3692 7144 3720
rect 7024 3194 7052 3692
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7116 3466 7144 3538
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7116 2990 7144 3402
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7024 2378 7052 2790
rect 7116 2582 7144 2926
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 7012 1896 7064 1902
rect 7012 1838 7064 1844
rect 7024 1562 7052 1838
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 7012 1556 7064 1562
rect 7012 1498 7064 1504
rect 7116 1426 7144 2518
rect 7208 1834 7236 3878
rect 7300 3194 7328 4626
rect 7364 4380 7740 4389
rect 7420 4378 7444 4380
rect 7500 4378 7524 4380
rect 7580 4378 7604 4380
rect 7660 4378 7684 4380
rect 7420 4326 7430 4378
rect 7674 4326 7684 4378
rect 7420 4324 7444 4326
rect 7500 4324 7524 4326
rect 7580 4324 7604 4326
rect 7660 4324 7684 4326
rect 7364 4315 7740 4324
rect 7748 4072 7800 4078
rect 7746 4040 7748 4049
rect 7800 4040 7802 4049
rect 7746 3975 7802 3984
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7364 3292 7740 3301
rect 7420 3290 7444 3292
rect 7500 3290 7524 3292
rect 7580 3290 7604 3292
rect 7660 3290 7684 3292
rect 7420 3238 7430 3290
rect 7674 3238 7684 3290
rect 7420 3236 7444 3238
rect 7500 3236 7524 3238
rect 7580 3236 7604 3238
rect 7660 3236 7684 3238
rect 7364 3227 7740 3236
rect 7852 3194 7880 3334
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7838 3088 7894 3097
rect 7838 3023 7894 3032
rect 7852 2990 7880 3023
rect 7288 2984 7340 2990
rect 7840 2984 7892 2990
rect 7288 2926 7340 2932
rect 7654 2952 7710 2961
rect 7300 2514 7328 2926
rect 7840 2926 7892 2932
rect 7654 2887 7710 2896
rect 7668 2582 7696 2887
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7300 1970 7328 2246
rect 7364 2204 7740 2213
rect 7420 2202 7444 2204
rect 7500 2202 7524 2204
rect 7580 2202 7604 2204
rect 7660 2202 7684 2204
rect 7420 2150 7430 2202
rect 7674 2150 7684 2202
rect 7420 2148 7444 2150
rect 7500 2148 7524 2150
rect 7580 2148 7604 2150
rect 7660 2148 7684 2150
rect 7364 2139 7740 2148
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 7288 1964 7340 1970
rect 7288 1906 7340 1912
rect 7196 1828 7248 1834
rect 7196 1770 7248 1776
rect 7576 1426 7604 1974
rect 7852 1902 7880 2926
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 7840 1896 7892 1902
rect 7840 1838 7892 1844
rect 7668 1562 7696 1838
rect 7656 1556 7708 1562
rect 7656 1498 7708 1504
rect 7840 1556 7892 1562
rect 7944 1544 7972 4791
rect 8036 4690 8064 5170
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8036 4214 8064 4626
rect 8128 4622 8156 5034
rect 8220 5001 8248 13874
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13462 8432 13670
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8404 12986 8432 13398
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8312 12374 8340 12650
rect 8404 12442 8432 12718
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8300 12232 8352 12238
rect 8496 12220 8524 15846
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8588 15162 8616 15302
rect 8772 15162 8800 15506
rect 8864 15366 8892 15914
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8588 14618 8616 14894
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8668 14408 8720 14414
rect 8588 14368 8668 14396
rect 8588 13394 8616 14368
rect 8668 14350 8720 14356
rect 8666 14240 8722 14249
rect 8666 14175 8722 14184
rect 8680 13433 8708 14175
rect 8772 14056 8800 14554
rect 8864 14414 8892 14894
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8772 14028 8892 14056
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13734 8800 13874
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8666 13424 8722 13433
rect 8576 13388 8628 13394
rect 8864 13410 8892 14028
rect 8666 13359 8668 13368
rect 8576 13330 8628 13336
rect 8720 13359 8722 13368
rect 8772 13382 8892 13410
rect 8668 13330 8720 13336
rect 8666 13152 8722 13161
rect 8588 13110 8666 13138
rect 8588 12288 8616 13110
rect 8666 13087 8722 13096
rect 8666 12744 8722 12753
rect 8666 12679 8722 12688
rect 8680 12646 8708 12679
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8588 12260 8708 12288
rect 8300 12174 8352 12180
rect 8404 12192 8524 12220
rect 8312 12073 8340 12174
rect 8298 12064 8354 12073
rect 8298 11999 8354 12008
rect 8404 11540 8432 12192
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8312 11512 8432 11540
rect 8312 8022 8340 11512
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8404 6848 8432 11290
rect 8496 10470 8524 12038
rect 8588 11354 8616 12106
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8588 10742 8616 11018
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8484 10464 8536 10470
rect 8482 10432 8484 10441
rect 8576 10464 8628 10470
rect 8536 10432 8538 10441
rect 8576 10406 8628 10412
rect 8482 10367 8538 10376
rect 8588 10062 8616 10406
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8496 8537 8524 8842
rect 8482 8528 8538 8537
rect 8482 8463 8538 8472
rect 8496 7857 8524 8463
rect 8482 7848 8538 7857
rect 8482 7783 8538 7792
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8312 6820 8432 6848
rect 8206 4992 8262 5001
rect 8206 4927 8262 4936
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8128 3738 8156 4082
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8036 2854 8064 2926
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 8036 1902 8064 2314
rect 8024 1896 8076 1902
rect 8024 1838 8076 1844
rect 7892 1516 7972 1544
rect 8022 1592 8078 1601
rect 8128 1562 8156 2790
rect 8312 2582 8340 6820
rect 8496 6746 8524 7686
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8588 6934 8616 7142
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8404 6718 8524 6746
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8404 6225 8432 6718
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8390 6216 8446 6225
rect 8390 6151 8446 6160
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8404 5545 8432 5850
rect 8496 5556 8524 6598
rect 8588 6458 8616 6734
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8680 6338 8708 12260
rect 8588 6310 8708 6338
rect 8588 5710 8616 6310
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8680 5642 8708 6190
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8390 5536 8446 5545
rect 8496 5528 8616 5556
rect 8588 5522 8616 5528
rect 8588 5494 8708 5522
rect 8390 5471 8446 5480
rect 8574 5400 8630 5409
rect 8574 5335 8576 5344
rect 8628 5335 8630 5344
rect 8576 5306 8628 5312
rect 8680 5273 8708 5494
rect 8772 5302 8800 13382
rect 8956 12170 8984 15846
rect 9232 15586 9260 16390
rect 9416 16046 9444 16646
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9600 16250 9628 16594
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9692 15978 9720 16390
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9324 15706 9352 15914
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9232 15558 9536 15586
rect 10060 15570 10088 16594
rect 10796 16250 10824 17070
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16658 11100 16934
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10364 15804 10740 15813
rect 10420 15802 10444 15804
rect 10500 15802 10524 15804
rect 10580 15802 10604 15804
rect 10660 15802 10684 15804
rect 10420 15750 10430 15802
rect 10674 15750 10684 15802
rect 10420 15748 10444 15750
rect 10500 15748 10524 15750
rect 10580 15748 10604 15750
rect 10660 15748 10684 15750
rect 10364 15739 10740 15748
rect 9128 15496 9180 15502
rect 9048 15456 9128 15484
rect 8944 12164 8996 12170
rect 8944 12106 8996 12112
rect 9048 12050 9076 15456
rect 9128 15438 9180 15444
rect 9310 15056 9366 15065
rect 9310 14991 9366 15000
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9140 13802 9168 14418
rect 9232 14074 9260 14554
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9140 13161 9168 13466
rect 9126 13152 9182 13161
rect 9126 13087 9182 13096
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8864 12022 9076 12050
rect 8760 5296 8812 5302
rect 8666 5264 8722 5273
rect 8760 5238 8812 5244
rect 8666 5199 8722 5208
rect 8392 5160 8444 5166
rect 8484 5160 8536 5166
rect 8392 5102 8444 5108
rect 8482 5128 8484 5137
rect 8668 5160 8720 5166
rect 8536 5128 8538 5137
rect 8404 3670 8432 5102
rect 8668 5102 8720 5108
rect 8482 5063 8538 5072
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 4826 8524 4966
rect 8680 4826 8708 5102
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8482 4720 8538 4729
rect 8482 4655 8484 4664
rect 8536 4655 8538 4664
rect 8484 4626 8536 4632
rect 8482 4584 8538 4593
rect 8482 4519 8538 4528
rect 8496 4214 8524 4519
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8864 2774 8892 12022
rect 9140 11914 9168 12582
rect 9324 12306 9352 14991
rect 9508 14482 9536 15558
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10244 15450 10272 15506
rect 9956 15428 10008 15434
rect 10060 15422 10272 15450
rect 10060 15416 10088 15422
rect 10008 15388 10088 15416
rect 9956 15370 10008 15376
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9508 13870 9536 14418
rect 9600 13870 9628 14894
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 14346 9904 14758
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9692 13705 9720 13738
rect 9678 13696 9734 13705
rect 9678 13631 9734 13640
rect 9586 13560 9642 13569
rect 9586 13495 9642 13504
rect 9600 13462 9628 13495
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9416 12714 9444 13330
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9508 12646 9536 12922
rect 9600 12782 9628 13398
rect 9784 13326 9812 14282
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9692 12986 9720 13194
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9784 12850 9812 13262
rect 9876 13190 9904 13670
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9968 12714 9996 14418
rect 10060 13802 10088 14962
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10060 13530 10088 13738
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10060 13433 10088 13466
rect 10046 13424 10102 13433
rect 10046 13359 10102 13368
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 10152 12434 10180 15302
rect 10364 14716 10740 14725
rect 10420 14714 10444 14716
rect 10500 14714 10524 14716
rect 10580 14714 10604 14716
rect 10660 14714 10684 14716
rect 10420 14662 10430 14714
rect 10674 14662 10684 14714
rect 10420 14660 10444 14662
rect 10500 14660 10524 14662
rect 10580 14660 10604 14662
rect 10660 14660 10684 14662
rect 10364 14651 10740 14660
rect 10506 14512 10562 14521
rect 10506 14447 10562 14456
rect 10600 14476 10652 14482
rect 10232 13728 10284 13734
rect 10520 13716 10548 14447
rect 10600 14418 10652 14424
rect 10612 14385 10640 14418
rect 10598 14376 10654 14385
rect 10598 14311 10654 14320
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 14074 10640 14214
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10600 13728 10652 13734
rect 10520 13688 10600 13716
rect 10232 13670 10284 13676
rect 10600 13670 10652 13676
rect 10244 13462 10272 13670
rect 10364 13628 10740 13637
rect 10420 13626 10444 13628
rect 10500 13626 10524 13628
rect 10580 13626 10604 13628
rect 10660 13626 10684 13628
rect 10420 13574 10430 13626
rect 10674 13574 10684 13626
rect 10420 13572 10444 13574
rect 10500 13572 10524 13574
rect 10580 13572 10604 13574
rect 10660 13572 10684 13574
rect 10364 13563 10740 13572
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10322 13288 10378 13297
rect 10232 13252 10284 13258
rect 10322 13223 10324 13232
rect 10232 13194 10284 13200
rect 10376 13223 10378 13232
rect 10324 13194 10376 13200
rect 9876 12406 10180 12434
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9310 12064 9366 12073
rect 9310 11999 9366 12008
rect 8956 11886 9168 11914
rect 8956 9194 8984 11886
rect 9324 11830 9352 11999
rect 9416 11898 9444 12106
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 9402 11792 9458 11801
rect 9458 11750 9536 11778
rect 9402 11727 9458 11736
rect 9508 11694 9536 11750
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9048 11354 9076 11630
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9034 10976 9090 10985
rect 9034 10911 9090 10920
rect 9048 10742 9076 10911
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9048 9518 9076 10474
rect 9140 10266 9168 11562
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9232 10130 9260 11154
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9128 10056 9180 10062
rect 9324 10010 9352 11086
rect 9416 10810 9444 11630
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11354 9628 11562
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10810 9628 10950
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9692 10441 9720 11494
rect 9770 11248 9826 11257
rect 9770 11183 9826 11192
rect 9678 10432 9734 10441
rect 9678 10367 9734 10376
rect 9784 10282 9812 11183
rect 9600 10254 9812 10282
rect 9600 10146 9628 10254
rect 9180 10004 9352 10010
rect 9128 9998 9352 10004
rect 9140 9982 9352 9998
rect 9508 10118 9628 10146
rect 9678 10160 9734 10169
rect 9140 9654 9168 9982
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9324 9382 9352 9522
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 8956 9166 9076 9194
rect 8944 9104 8996 9110
rect 8942 9072 8944 9081
rect 8996 9072 8998 9081
rect 8942 9007 8998 9016
rect 9048 7970 9076 9166
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9140 8430 9168 9046
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9324 8634 9352 8978
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8956 7942 9076 7970
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 8956 6497 8984 7942
rect 9232 7342 9260 7958
rect 9508 7546 9536 10118
rect 9678 10095 9734 10104
rect 9772 10124 9824 10130
rect 9692 10010 9720 10095
rect 9772 10066 9824 10072
rect 9600 9982 9720 10010
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9600 7449 9628 9982
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 8838 9720 9862
rect 9784 9722 9812 10066
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9784 9081 9812 9454
rect 9770 9072 9826 9081
rect 9770 9007 9826 9016
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8498 9720 8774
rect 9784 8634 9812 8910
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9586 7440 9642 7449
rect 9586 7375 9642 7384
rect 9128 7336 9180 7342
rect 9126 7304 9128 7313
rect 9220 7336 9272 7342
rect 9180 7304 9182 7313
rect 9496 7336 9548 7342
rect 9272 7296 9444 7324
rect 9220 7278 9272 7284
rect 9126 7239 9182 7248
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9048 7002 9076 7142
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9140 6866 9168 7142
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 8942 6488 8998 6497
rect 9140 6458 9168 6802
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 8942 6423 8998 6432
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 9126 6352 9182 6361
rect 8956 5642 8984 6326
rect 9126 6287 9182 6296
rect 9034 6216 9090 6225
rect 9034 6151 9090 6160
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 8942 5536 8998 5545
rect 8942 5471 8998 5480
rect 8956 3466 8984 5471
rect 9048 5166 9076 6151
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9048 4185 9076 4558
rect 9034 4176 9090 4185
rect 9034 4111 9090 4120
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 9048 3194 9076 4014
rect 9140 3913 9168 6287
rect 9232 5574 9260 6734
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 4010 9260 5510
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9126 3904 9182 3913
rect 9126 3839 9182 3848
rect 9140 3738 9168 3839
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9232 3194 9260 3606
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8680 2746 8984 2774
rect 8680 2650 8708 2746
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8220 1970 8248 2518
rect 8312 2038 8340 2518
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8300 2032 8352 2038
rect 8300 1974 8352 1980
rect 8668 2032 8720 2038
rect 8668 1974 8720 1980
rect 8208 1964 8260 1970
rect 8208 1906 8260 1912
rect 8574 1864 8630 1873
rect 8574 1799 8630 1808
rect 8588 1766 8616 1799
rect 8680 1766 8708 1974
rect 8864 1902 8892 2246
rect 8956 1970 8984 2746
rect 9034 2544 9090 2553
rect 9324 2514 9352 7142
rect 9416 6458 9444 7296
rect 9496 7278 9548 7284
rect 9508 6934 9536 7278
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9496 6792 9548 6798
rect 9692 6746 9720 7482
rect 9772 7472 9824 7478
rect 9770 7440 9772 7449
rect 9824 7440 9826 7449
rect 9770 7375 9826 7384
rect 9548 6740 9720 6746
rect 9496 6734 9720 6740
rect 9508 6718 9720 6734
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9784 6458 9812 6666
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9416 5302 9444 5578
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9508 4758 9536 5510
rect 9600 5166 9628 5714
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9588 5160 9640 5166
rect 9692 5137 9720 5238
rect 9784 5166 9812 5306
rect 9876 5273 9904 12406
rect 10244 11762 10272 13194
rect 10336 12714 10364 13194
rect 10612 13190 10640 13330
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12782 10732 13126
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10364 12540 10740 12549
rect 10420 12538 10444 12540
rect 10500 12538 10524 12540
rect 10580 12538 10604 12540
rect 10660 12538 10684 12540
rect 10420 12486 10430 12538
rect 10674 12486 10684 12538
rect 10420 12484 10444 12486
rect 10500 12484 10524 12486
rect 10580 12484 10604 12486
rect 10660 12484 10684 12486
rect 10364 12475 10740 12484
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9968 11150 9996 11630
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 10152 11014 10180 11494
rect 10244 11354 10272 11698
rect 10364 11452 10740 11461
rect 10420 11450 10444 11452
rect 10500 11450 10524 11452
rect 10580 11450 10604 11452
rect 10660 11450 10684 11452
rect 10420 11398 10430 11450
rect 10674 11398 10684 11450
rect 10420 11396 10444 11398
rect 10500 11396 10524 11398
rect 10580 11396 10604 11398
rect 10660 11396 10684 11398
rect 10364 11387 10740 11396
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10248 10272 10406
rect 10364 10364 10740 10373
rect 10420 10362 10444 10364
rect 10500 10362 10524 10364
rect 10580 10362 10604 10364
rect 10660 10362 10684 10364
rect 10420 10310 10430 10362
rect 10674 10310 10684 10362
rect 10420 10308 10444 10310
rect 10500 10308 10524 10310
rect 10580 10308 10604 10310
rect 10660 10308 10684 10310
rect 10364 10299 10740 10308
rect 10796 10282 10824 15846
rect 10980 15706 11008 15982
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11164 15434 11192 16118
rect 11440 16114 11468 17070
rect 11624 16538 11652 17138
rect 11532 16522 11652 16538
rect 11520 16516 11652 16522
rect 11572 16510 11652 16516
rect 11520 16458 11572 16464
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11334 15600 11390 15609
rect 11532 15570 11560 16186
rect 11624 16114 11652 16510
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11334 15535 11390 15544
rect 11520 15564 11572 15570
rect 11348 15502 11376 15535
rect 11520 15506 11572 15512
rect 11336 15496 11388 15502
rect 11532 15473 11560 15506
rect 11336 15438 11388 15444
rect 11518 15464 11574 15473
rect 11152 15428 11204 15434
rect 11624 15434 11652 16050
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11518 15399 11574 15408
rect 11612 15428 11664 15434
rect 11152 15370 11204 15376
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10888 13530 10916 14350
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10980 12753 11008 13942
rect 11072 13802 11100 14214
rect 11164 13977 11192 14214
rect 11244 14000 11296 14006
rect 11150 13968 11206 13977
rect 11244 13942 11296 13948
rect 11150 13903 11206 13912
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 10966 12744 11022 12753
rect 10876 12708 10928 12714
rect 10966 12679 11022 12688
rect 10876 12650 10928 12656
rect 10888 10606 10916 12650
rect 11256 12374 11284 13942
rect 11348 13802 11376 14418
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10416 10260 10468 10266
rect 10244 10220 10416 10248
rect 10796 10254 10916 10282
rect 10416 10202 10468 10208
rect 10428 10130 10456 10202
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 9968 9926 9996 10066
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9968 9178 9996 9522
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10060 9042 10088 9862
rect 10232 9648 10284 9654
rect 10230 9616 10232 9625
rect 10284 9616 10286 9625
rect 10230 9551 10286 9560
rect 10336 9518 10364 10066
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10428 9654 10456 9862
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10152 9178 10180 9454
rect 10232 9376 10284 9382
rect 10704 9364 10732 10066
rect 10796 9926 10824 10134
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10704 9336 10824 9364
rect 10232 9318 10284 9324
rect 10140 9172 10192 9178
rect 10244 9160 10272 9318
rect 10364 9276 10740 9285
rect 10420 9274 10444 9276
rect 10500 9274 10524 9276
rect 10580 9274 10604 9276
rect 10660 9274 10684 9276
rect 10420 9222 10430 9274
rect 10674 9222 10684 9274
rect 10420 9220 10444 9222
rect 10500 9220 10524 9222
rect 10580 9220 10604 9222
rect 10660 9220 10684 9222
rect 10364 9211 10740 9220
rect 10244 9132 10548 9160
rect 10140 9114 10192 9120
rect 10230 9072 10286 9081
rect 10048 9036 10100 9042
rect 10520 9042 10548 9132
rect 10796 9042 10824 9336
rect 10416 9036 10468 9042
rect 10230 9007 10286 9016
rect 10048 8978 10100 8984
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 10048 8424 10100 8430
rect 10244 8401 10272 9007
rect 10336 8996 10416 9024
rect 10336 8498 10364 8996
rect 10416 8978 10468 8984
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8945 10824 8978
rect 10782 8936 10838 8945
rect 10782 8871 10838 8880
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10048 8366 10100 8372
rect 10230 8392 10286 8401
rect 9968 6633 9996 8366
rect 10060 7750 10088 8366
rect 10230 8327 10232 8336
rect 10284 8327 10286 8336
rect 10232 8298 10284 8304
rect 10364 8188 10740 8197
rect 10420 8186 10444 8188
rect 10500 8186 10524 8188
rect 10580 8186 10604 8188
rect 10660 8186 10684 8188
rect 10420 8134 10430 8186
rect 10674 8134 10684 8186
rect 10420 8132 10444 8134
rect 10500 8132 10524 8134
rect 10580 8132 10604 8134
rect 10660 8132 10684 8134
rect 10364 8123 10740 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 6866 10088 7686
rect 10152 7546 10180 8026
rect 10796 7818 10824 8502
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10428 7546 10456 7686
rect 10704 7546 10732 7686
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10324 7472 10376 7478
rect 10376 7420 10548 7426
rect 10324 7414 10548 7420
rect 10336 7398 10548 7414
rect 10520 7342 10548 7398
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10152 6866 10180 7142
rect 10364 7100 10740 7109
rect 10420 7098 10444 7100
rect 10500 7098 10524 7100
rect 10580 7098 10604 7100
rect 10660 7098 10684 7100
rect 10420 7046 10430 7098
rect 10674 7046 10684 7098
rect 10420 7044 10444 7046
rect 10500 7044 10524 7046
rect 10580 7044 10604 7046
rect 10660 7044 10684 7046
rect 10364 7035 10740 7044
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10060 6746 10088 6802
rect 10324 6792 10376 6798
rect 10060 6718 10180 6746
rect 10416 6792 10468 6798
rect 10324 6734 10376 6740
rect 10414 6760 10416 6769
rect 10508 6792 10560 6798
rect 10468 6760 10470 6769
rect 9954 6624 10010 6633
rect 9954 6559 10010 6568
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9862 5264 9918 5273
rect 9862 5199 9918 5208
rect 9772 5160 9824 5166
rect 9588 5102 9640 5108
rect 9678 5128 9734 5137
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9600 4690 9628 5102
rect 9772 5102 9824 5108
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9678 5063 9734 5072
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4690 9720 4966
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9680 4684 9732 4690
rect 9732 4644 9812 4672
rect 9680 4626 9732 4632
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9416 3618 9444 4558
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9692 4010 9720 4490
rect 9784 4078 9812 4644
rect 9876 4554 9904 5102
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9416 3590 9628 3618
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9034 2479 9036 2488
rect 9088 2479 9090 2488
rect 9312 2508 9364 2514
rect 9036 2450 9088 2456
rect 9312 2450 9364 2456
rect 9126 2408 9182 2417
rect 9036 2372 9088 2378
rect 9126 2343 9182 2352
rect 9036 2314 9088 2320
rect 8944 1964 8996 1970
rect 8944 1906 8996 1912
rect 9048 1902 9076 2314
rect 9140 2038 9168 2343
rect 9128 2032 9180 2038
rect 9416 2020 9444 2790
rect 9128 1974 9180 1980
rect 9232 1992 9444 2020
rect 8852 1896 8904 1902
rect 8852 1838 8904 1844
rect 9036 1896 9088 1902
rect 9036 1838 9088 1844
rect 8484 1760 8536 1766
rect 8484 1702 8536 1708
rect 8576 1760 8628 1766
rect 8576 1702 8628 1708
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 8022 1527 8078 1536
rect 8116 1556 8168 1562
rect 7840 1498 7892 1504
rect 8036 1494 8064 1527
rect 8116 1498 8168 1504
rect 8496 1494 8524 1702
rect 8024 1488 8076 1494
rect 8024 1430 8076 1436
rect 8484 1488 8536 1494
rect 8484 1430 8536 1436
rect 8944 1488 8996 1494
rect 8944 1430 8996 1436
rect 7104 1420 7156 1426
rect 7104 1362 7156 1368
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 8484 1352 8536 1358
rect 8484 1294 8536 1300
rect 2780 1216 2832 1222
rect 2780 1158 2832 1164
rect 3608 1216 3660 1222
rect 3608 1158 3660 1164
rect 5356 1216 5408 1222
rect 5356 1158 5408 1164
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 6368 1216 6420 1222
rect 6368 1158 6420 1164
rect 6644 1216 6696 1222
rect 6644 1158 6696 1164
rect 6736 1216 6788 1222
rect 6736 1158 6788 1164
rect 6828 1216 6880 1222
rect 7760 1204 7788 1294
rect 8392 1216 8444 1222
rect 7760 1176 7880 1204
rect 6828 1158 6880 1164
rect 2504 1012 2556 1018
rect 2504 954 2556 960
rect 2412 876 2464 882
rect 2412 818 2464 824
rect 5368 814 5396 1158
rect 5828 1018 5856 1158
rect 5816 1012 5868 1018
rect 5816 954 5868 960
rect 2320 808 2372 814
rect 2320 750 2372 756
rect 4160 808 4212 814
rect 4160 750 4212 756
rect 5264 808 5316 814
rect 5264 750 5316 756
rect 5356 808 5408 814
rect 5356 750 5408 756
rect 6092 808 6144 814
rect 6092 750 6144 756
rect 2780 672 2832 678
rect 2780 614 2832 620
rect 3700 672 3752 678
rect 3700 614 3752 620
rect 2792 400 2820 614
rect 3712 456 3740 614
rect 3528 428 3740 456
rect 3528 400 3556 428
rect 570 0 626 400
rect 1306 0 1362 400
rect 2042 0 2098 400
rect 2778 0 2834 400
rect 3514 0 3570 400
rect 4172 202 4200 750
rect 4252 672 4304 678
rect 4252 614 4304 620
rect 5172 672 5224 678
rect 5172 614 5224 620
rect 4264 400 4292 614
rect 4364 572 4740 581
rect 4420 570 4444 572
rect 4500 570 4524 572
rect 4580 570 4604 572
rect 4660 570 4684 572
rect 4420 518 4430 570
rect 4674 518 4684 570
rect 4420 516 4444 518
rect 4500 516 4524 518
rect 4580 516 4604 518
rect 4660 516 4684 518
rect 4364 507 4740 516
rect 5184 456 5212 614
rect 5276 474 5304 750
rect 5908 672 5960 678
rect 5908 614 5960 620
rect 5000 428 5212 456
rect 5264 468 5316 474
rect 5000 400 5028 428
rect 5920 456 5948 614
rect 6104 474 6132 750
rect 5264 410 5316 416
rect 5736 428 5948 456
rect 6092 468 6144 474
rect 5736 400 5764 428
rect 6092 410 6144 416
rect 6380 406 6408 1158
rect 6656 814 6684 1158
rect 6748 814 6776 1158
rect 7364 1116 7740 1125
rect 7420 1114 7444 1116
rect 7500 1114 7524 1116
rect 7580 1114 7604 1116
rect 7660 1114 7684 1116
rect 7420 1062 7430 1114
rect 7674 1062 7684 1114
rect 7420 1060 7444 1062
rect 7500 1060 7524 1062
rect 7580 1060 7604 1062
rect 7660 1060 7684 1062
rect 7364 1051 7740 1060
rect 6644 808 6696 814
rect 6644 750 6696 756
rect 6736 808 6788 814
rect 6736 750 6788 756
rect 6644 672 6696 678
rect 6644 614 6696 620
rect 7196 672 7248 678
rect 7196 614 7248 620
rect 6656 456 6684 614
rect 6472 428 6684 456
rect 6368 400 6420 406
rect 6472 400 6500 428
rect 7208 400 7236 614
rect 4160 196 4212 202
rect 4160 138 4212 144
rect 4250 0 4306 400
rect 4986 0 5042 400
rect 5722 0 5778 400
rect 6368 342 6420 348
rect 6458 0 6514 400
rect 7194 0 7250 400
rect 7852 270 7880 1176
rect 8392 1158 8444 1164
rect 8116 876 8168 882
rect 8404 864 8432 1158
rect 8168 836 8432 864
rect 8116 818 8168 824
rect 8496 814 8524 1294
rect 8956 1290 8984 1430
rect 9232 1426 9260 1992
rect 9220 1420 9272 1426
rect 9600 1408 9628 3590
rect 9692 3584 9720 3946
rect 9784 3738 9812 4014
rect 9876 3738 9904 4014
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9864 3596 9916 3602
rect 9692 3556 9864 3584
rect 9864 3538 9916 3544
rect 9770 3360 9826 3369
rect 9770 3295 9826 3304
rect 9784 3058 9812 3295
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 1902 9812 2246
rect 9680 1896 9732 1902
rect 9680 1838 9732 1844
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 9692 1601 9720 1838
rect 9770 1728 9826 1737
rect 9770 1663 9826 1672
rect 9678 1592 9734 1601
rect 9784 1562 9812 1663
rect 9678 1527 9734 1536
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 9772 1420 9824 1426
rect 9600 1380 9772 1408
rect 9220 1362 9272 1368
rect 9772 1362 9824 1368
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 8852 1284 8904 1290
rect 8852 1226 8904 1232
rect 8944 1284 8996 1290
rect 8944 1226 8996 1232
rect 8864 1018 8892 1226
rect 9324 1018 9352 1294
rect 9678 1184 9734 1193
rect 9678 1119 9734 1128
rect 8852 1012 8904 1018
rect 8852 954 8904 960
rect 9312 1012 9364 1018
rect 9312 954 9364 960
rect 9404 944 9456 950
rect 9404 886 9456 892
rect 8484 808 8536 814
rect 8484 750 8536 756
rect 8116 740 8168 746
rect 8116 682 8168 688
rect 8128 456 8156 682
rect 8392 672 8444 678
rect 8392 614 8444 620
rect 7944 428 8156 456
rect 7944 400 7972 428
rect 7840 264 7892 270
rect 7840 206 7892 212
rect 7930 0 7986 400
rect 8404 354 8432 614
rect 8588 428 8708 456
rect 8588 354 8616 428
rect 8680 400 8708 428
rect 9416 400 9444 886
rect 9692 406 9720 1119
rect 9876 814 9904 1838
rect 9968 1018 9996 6190
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10060 5166 10088 5510
rect 10152 5166 10180 6718
rect 10336 6254 10364 6734
rect 10796 6780 10824 7754
rect 10560 6752 10824 6780
rect 10508 6734 10560 6740
rect 10414 6695 10470 6704
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10364 6012 10740 6021
rect 10420 6010 10444 6012
rect 10500 6010 10524 6012
rect 10580 6010 10604 6012
rect 10660 6010 10684 6012
rect 10420 5958 10430 6010
rect 10674 5958 10684 6010
rect 10420 5956 10444 5958
rect 10500 5956 10524 5958
rect 10580 5956 10604 5958
rect 10660 5956 10684 5958
rect 10364 5947 10740 5956
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10060 4078 10088 4966
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3738 10088 3878
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10060 3194 10088 3538
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10152 1850 10180 4966
rect 10244 3602 10272 5578
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5234 10824 5510
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10364 4924 10740 4933
rect 10420 4922 10444 4924
rect 10500 4922 10524 4924
rect 10580 4922 10604 4924
rect 10660 4922 10684 4924
rect 10420 4870 10430 4922
rect 10674 4870 10684 4922
rect 10420 4868 10444 4870
rect 10500 4868 10524 4870
rect 10580 4868 10604 4870
rect 10660 4868 10684 4870
rect 10364 4859 10740 4868
rect 10796 4622 10824 4966
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10364 3836 10740 3845
rect 10420 3834 10444 3836
rect 10500 3834 10524 3836
rect 10580 3834 10604 3836
rect 10660 3834 10684 3836
rect 10420 3782 10430 3834
rect 10674 3782 10684 3834
rect 10420 3780 10444 3782
rect 10500 3780 10524 3782
rect 10580 3780 10604 3782
rect 10660 3780 10684 3782
rect 10364 3771 10740 3780
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10428 3534 10456 3674
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10428 3398 10456 3470
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10364 2748 10740 2757
rect 10420 2746 10444 2748
rect 10500 2746 10524 2748
rect 10580 2746 10604 2748
rect 10660 2746 10684 2748
rect 10420 2694 10430 2746
rect 10674 2694 10684 2746
rect 10420 2692 10444 2694
rect 10500 2692 10524 2694
rect 10580 2692 10604 2694
rect 10660 2692 10684 2694
rect 10364 2683 10740 2692
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10612 2378 10640 2450
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 10888 2145 10916 10254
rect 10980 10130 11008 12242
rect 11348 12102 11376 13330
rect 11440 13326 11468 14758
rect 11532 14634 11560 15399
rect 11612 15370 11664 15376
rect 11716 14822 11744 15914
rect 11808 15094 11836 17546
rect 11992 17134 12020 17845
rect 12820 17678 12848 17845
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 13648 17542 13676 17845
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13004 17270 13032 17478
rect 13364 17436 13740 17445
rect 13420 17434 13444 17436
rect 13500 17434 13524 17436
rect 13580 17434 13604 17436
rect 13660 17434 13684 17436
rect 13420 17382 13430 17434
rect 13674 17382 13684 17434
rect 13420 17380 13444 17382
rect 13500 17380 13524 17382
rect 13580 17380 13604 17382
rect 13660 17380 13684 17382
rect 13364 17371 13740 17380
rect 12992 17264 13044 17270
rect 13820 17264 13872 17270
rect 12992 17206 13044 17212
rect 13740 17212 13820 17218
rect 13740 17206 13872 17212
rect 13740 17190 13860 17206
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11992 15450 12020 15574
rect 11900 15422 12020 15450
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11900 14958 11928 15422
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11532 14606 11836 14634
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11532 13394 11560 14214
rect 11624 13802 11652 14350
rect 11808 14278 11836 14606
rect 11900 14550 11928 14894
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11978 14512 12034 14521
rect 11978 14447 12034 14456
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11150 11100 11494
rect 11256 11354 11284 11630
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11348 11286 11376 12038
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9500 11008 10066
rect 11060 9512 11112 9518
rect 10980 9472 11060 9500
rect 11060 9454 11112 9460
rect 11164 9382 11192 10950
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11072 9178 11100 9318
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10980 7002 11008 8230
rect 11072 7410 11100 8230
rect 11256 7954 11284 10678
rect 11348 10266 11376 10678
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11348 9110 11376 10202
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11440 8566 11468 12786
rect 11716 12434 11744 14214
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11808 12918 11836 14010
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11900 13433 11928 13806
rect 11886 13424 11942 13433
rect 11886 13359 11942 13368
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11992 12850 12020 14447
rect 12084 14113 12112 16934
rect 12360 16510 12664 16538
rect 12360 16250 12388 16510
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15638 12204 15846
rect 12164 15632 12216 15638
rect 12164 15574 12216 15580
rect 12268 15337 12296 16050
rect 12348 15564 12400 15570
rect 12544 15552 12572 16390
rect 12636 16182 12664 16510
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12728 16046 12756 17002
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12820 15978 12848 16730
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13096 16182 13124 16390
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12400 15524 12572 15552
rect 12348 15506 12400 15512
rect 12254 15328 12310 15337
rect 12254 15263 12310 15272
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12176 14385 12204 14554
rect 12162 14376 12218 14385
rect 12162 14311 12218 14320
rect 12070 14104 12126 14113
rect 12070 14039 12126 14048
rect 12084 13938 12112 14039
rect 12176 14006 12204 14311
rect 12268 14006 12296 14894
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12360 14618 12388 14826
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12360 14482 12388 14554
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12452 14278 12480 15524
rect 12544 15348 12572 15524
rect 12716 15564 12768 15570
rect 12820 15552 12848 15914
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 12768 15524 12848 15552
rect 12716 15506 12768 15512
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12716 15360 12768 15366
rect 12544 15320 12716 15348
rect 12716 15302 12768 15308
rect 12820 15076 12848 15370
rect 12912 15337 12940 15846
rect 13096 15706 13124 15846
rect 13188 15706 13216 16594
rect 13372 16538 13400 16594
rect 13464 16590 13492 17070
rect 13740 16794 13768 17190
rect 14108 17134 14136 17614
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 14384 16726 14412 17070
rect 14476 16794 14504 17845
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 13280 16510 13400 16538
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13280 16250 13308 16510
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 13364 16348 13740 16357
rect 13420 16346 13444 16348
rect 13500 16346 13524 16348
rect 13580 16346 13604 16348
rect 13660 16346 13684 16348
rect 13420 16294 13430 16346
rect 13674 16294 13684 16346
rect 13420 16292 13444 16294
rect 13500 16292 13524 16294
rect 13580 16292 13604 16294
rect 13660 16292 13684 16294
rect 13364 16283 13740 16292
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12992 15496 13044 15502
rect 12990 15464 12992 15473
rect 13044 15464 13046 15473
rect 12990 15399 13046 15408
rect 13096 15416 13124 15506
rect 13096 15388 13130 15416
rect 12992 15360 13044 15366
rect 12898 15328 12954 15337
rect 12992 15302 13044 15308
rect 12898 15263 12954 15272
rect 12900 15088 12952 15094
rect 12820 15048 12900 15076
rect 12900 15030 12952 15036
rect 12900 14952 12952 14958
rect 12622 14920 12678 14929
rect 12900 14894 12952 14900
rect 12622 14855 12624 14864
rect 12676 14855 12678 14864
rect 12624 14826 12676 14832
rect 12912 14414 12940 14894
rect 12532 14408 12584 14414
rect 12900 14408 12952 14414
rect 12532 14350 12584 14356
rect 12820 14368 12900 14396
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12084 13530 12112 13874
rect 12544 13870 12572 14350
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12532 13864 12584 13870
rect 12530 13832 12532 13841
rect 12624 13864 12676 13870
rect 12584 13832 12586 13841
rect 12624 13806 12676 13812
rect 12530 13767 12586 13776
rect 12440 13728 12492 13734
rect 12636 13705 12664 13806
rect 12440 13670 12492 13676
rect 12622 13696 12678 13705
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 12850 12204 13330
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 11796 12640 11848 12646
rect 11848 12600 12112 12628
rect 11796 12582 11848 12588
rect 12084 12434 12112 12600
rect 11716 12406 11836 12434
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11716 11898 11744 12242
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11440 8362 11468 8502
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11072 6882 11100 7142
rect 10968 6860 11020 6866
rect 11072 6854 11192 6882
rect 10968 6802 11020 6808
rect 10980 6254 11008 6802
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6458 11100 6734
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11072 4214 11100 4762
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 3602 11008 4082
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10874 2136 10930 2145
rect 10692 2100 10744 2106
rect 10874 2071 10930 2080
rect 10692 2042 10744 2048
rect 10048 1828 10100 1834
rect 10152 1822 10272 1850
rect 10048 1770 10100 1776
rect 10060 1562 10088 1770
rect 10140 1760 10192 1766
rect 10140 1702 10192 1708
rect 10048 1556 10100 1562
rect 10048 1498 10100 1504
rect 10152 1442 10180 1702
rect 10060 1426 10180 1442
rect 10048 1420 10180 1426
rect 10100 1414 10180 1420
rect 10048 1362 10100 1368
rect 10244 1340 10272 1822
rect 10704 1766 10732 2042
rect 10980 2020 11008 3538
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 2990 11100 3334
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2446 11100 2926
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 10888 1992 11008 2020
rect 10888 1834 10916 1992
rect 11072 1970 11100 2382
rect 11060 1964 11112 1970
rect 11060 1906 11112 1912
rect 10876 1828 10928 1834
rect 10876 1770 10928 1776
rect 10692 1760 10744 1766
rect 10692 1702 10744 1708
rect 10968 1760 11020 1766
rect 10968 1702 11020 1708
rect 10364 1660 10740 1669
rect 10420 1658 10444 1660
rect 10500 1658 10524 1660
rect 10580 1658 10604 1660
rect 10660 1658 10684 1660
rect 10420 1606 10430 1658
rect 10674 1606 10684 1658
rect 10420 1604 10444 1606
rect 10500 1604 10524 1606
rect 10580 1604 10604 1606
rect 10660 1604 10684 1606
rect 10364 1595 10740 1604
rect 10692 1488 10744 1494
rect 10692 1430 10744 1436
rect 10508 1352 10560 1358
rect 10244 1312 10508 1340
rect 10704 1329 10732 1430
rect 10980 1358 11008 1702
rect 10968 1352 11020 1358
rect 10508 1294 10560 1300
rect 10690 1320 10746 1329
rect 10048 1284 10100 1290
rect 11060 1352 11112 1358
rect 10968 1294 11020 1300
rect 11058 1320 11060 1329
rect 11112 1320 11114 1329
rect 10690 1255 10746 1264
rect 10048 1226 10100 1232
rect 9956 1012 10008 1018
rect 9956 954 10008 960
rect 9864 808 9916 814
rect 9864 750 9916 756
rect 9680 400 9732 406
rect 8404 326 8616 354
rect 8666 0 8722 400
rect 9402 0 9458 400
rect 9680 342 9732 348
rect 10060 202 10088 1226
rect 10980 814 11008 1294
rect 11058 1255 11114 1264
rect 10968 808 11020 814
rect 10968 750 11020 756
rect 11072 746 11100 1255
rect 11164 1018 11192 6854
rect 11256 6458 11284 7890
rect 11532 7886 11560 11494
rect 11716 11354 11744 11630
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11624 10198 11652 11154
rect 11716 10606 11744 11290
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11624 9722 11652 10134
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11716 9110 11744 9454
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11716 8430 11744 9046
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11256 5574 11284 6394
rect 11348 6390 11376 6802
rect 11428 6792 11480 6798
rect 11532 6780 11560 7822
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11624 7546 11652 7686
rect 11716 7546 11744 7754
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11612 7336 11664 7342
rect 11808 7313 11836 12406
rect 11992 12406 12112 12434
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11612 7278 11664 7284
rect 11794 7304 11850 7313
rect 11480 6752 11560 6780
rect 11428 6734 11480 6740
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11440 6089 11468 6258
rect 11426 6080 11482 6089
rect 11426 6015 11482 6024
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11256 4282 11284 5102
rect 11348 4826 11376 5714
rect 11532 5234 11560 6752
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11532 4078 11560 4626
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11256 2650 11284 3674
rect 11532 3466 11560 4014
rect 11624 3738 11652 7278
rect 11794 7239 11850 7248
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11716 6118 11744 6666
rect 11808 6254 11836 7239
rect 11900 6934 11928 8298
rect 11992 7410 12020 12406
rect 12072 11620 12124 11626
rect 12072 11562 12124 11568
rect 12084 11014 12112 11562
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11354 12388 11494
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12256 11144 12308 11150
rect 12254 11112 12256 11121
rect 12308 11112 12310 11121
rect 12254 11047 12310 11056
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 9042 12112 10950
rect 12346 10568 12402 10577
rect 12346 10503 12402 10512
rect 12360 10266 12388 10503
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12452 10010 12480 13670
rect 12622 13631 12678 13640
rect 12636 13462 12664 13631
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12530 12880 12586 12889
rect 12530 12815 12532 12824
rect 12584 12815 12586 12824
rect 12532 12786 12584 12792
rect 12624 12776 12676 12782
rect 12544 12724 12624 12730
rect 12544 12718 12676 12724
rect 12544 12702 12664 12718
rect 12544 12442 12572 12702
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 10266 12572 12038
rect 12636 11801 12664 12582
rect 12622 11792 12678 11801
rect 12622 11727 12678 11736
rect 12728 11642 12756 14214
rect 12820 13530 12848 14368
rect 12900 14350 12952 14356
rect 13004 13716 13032 15302
rect 13102 15178 13130 15388
rect 13096 15150 13130 15178
rect 13096 14822 13124 15150
rect 13188 15042 13216 15642
rect 13280 15609 13308 15982
rect 13266 15600 13322 15609
rect 13322 15558 13492 15586
rect 13266 15535 13322 15544
rect 13464 15434 13492 15558
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13280 15144 13308 15370
rect 13364 15260 13740 15269
rect 13420 15258 13444 15260
rect 13500 15258 13524 15260
rect 13580 15258 13604 15260
rect 13660 15258 13684 15260
rect 13420 15206 13430 15258
rect 13674 15206 13684 15258
rect 13420 15204 13444 15206
rect 13500 15204 13524 15206
rect 13580 15204 13604 15206
rect 13660 15204 13684 15206
rect 13364 15195 13740 15204
rect 13452 15156 13504 15162
rect 13280 15116 13400 15144
rect 13188 15026 13308 15042
rect 13188 15020 13320 15026
rect 13188 15014 13268 15020
rect 13268 14962 13320 14968
rect 13372 14929 13400 15116
rect 13452 15098 13504 15104
rect 13358 14920 13414 14929
rect 13464 14890 13492 15098
rect 13358 14855 13414 14864
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 12988 13688 13032 13716
rect 12988 13546 13016 13688
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12900 13524 12952 13530
rect 12988 13518 13032 13546
rect 13096 13530 13124 14758
rect 13832 14634 13860 16050
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15570 13952 15846
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 14200 15434 14228 16390
rect 14384 16164 14412 16662
rect 14568 16658 14596 17478
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14844 16590 14872 17546
rect 15304 17338 15332 17845
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 16132 17202 16160 17845
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14464 16176 14516 16182
rect 14384 16136 14464 16164
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15570 14320 15846
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 14188 15428 14240 15434
rect 14188 15370 14240 15376
rect 13924 15162 13952 15370
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13910 15056 13966 15065
rect 13910 14991 13966 15000
rect 14188 15020 14240 15026
rect 13924 14890 13952 14991
rect 14188 14962 14240 14968
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13648 14606 13860 14634
rect 13648 14362 13676 14606
rect 14016 14482 14044 14894
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13188 14334 13676 14362
rect 12900 13466 12952 13472
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12646 12848 12786
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11762 12848 12038
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12728 11614 12848 11642
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12728 11218 12756 11494
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12820 10962 12848 11614
rect 12912 11354 12940 13466
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12820 10934 12940 10962
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12532 10260 12584 10266
rect 12584 10220 12664 10248
rect 12532 10202 12584 10208
rect 12348 9988 12400 9994
rect 12452 9982 12572 10010
rect 12348 9930 12400 9936
rect 12360 9722 12388 9930
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12256 9512 12308 9518
rect 12452 9500 12480 9862
rect 12308 9472 12480 9500
rect 12256 9454 12308 9460
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12268 8498 12296 8842
rect 12360 8634 12388 9318
rect 12452 9110 12480 9318
rect 12440 9104 12492 9110
rect 12438 9072 12440 9081
rect 12492 9072 12494 9081
rect 12438 9007 12494 9016
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12544 8514 12572 9982
rect 12636 9450 12664 10220
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12636 8838 12664 9386
rect 12728 9042 12756 10610
rect 12820 10266 12848 10746
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12806 9616 12862 9625
rect 12806 9551 12862 9560
rect 12820 9518 12848 9551
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 9066 12848 9318
rect 12808 9060 12860 9066
rect 12716 9036 12768 9042
rect 12808 9002 12860 9008
rect 12716 8978 12768 8984
rect 12808 8968 12860 8974
rect 12728 8916 12808 8922
rect 12728 8910 12860 8916
rect 12728 8894 12848 8910
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12728 8650 12756 8894
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12360 8486 12572 8514
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7954 12204 8230
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12360 7834 12388 8486
rect 12544 7954 12572 8486
rect 12636 8622 12756 8650
rect 12636 8401 12664 8622
rect 12622 8392 12678 8401
rect 12622 8327 12678 8336
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12084 7806 12388 7834
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11796 6248 11848 6254
rect 11848 6208 11928 6236
rect 11796 6190 11848 6196
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11716 4758 11744 5510
rect 11808 4758 11836 5578
rect 11900 5250 11928 6208
rect 11992 5574 12020 7346
rect 11980 5568 12032 5574
rect 11978 5536 11980 5545
rect 12032 5536 12034 5545
rect 11978 5471 12034 5480
rect 11900 5222 12020 5250
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11900 4826 11928 5102
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11992 3584 12020 5222
rect 12084 4826 12112 7806
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 7546 12388 7686
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12176 7449 12204 7482
rect 12162 7440 12218 7449
rect 12218 7398 12388 7426
rect 12162 7375 12218 7384
rect 12360 7342 12388 7398
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6186 12204 6598
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12268 6254 12296 6394
rect 12452 6304 12480 7482
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12360 6276 12480 6304
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12162 5808 12218 5817
rect 12268 5778 12296 6054
rect 12162 5743 12218 5752
rect 12256 5772 12308 5778
rect 12176 5234 12204 5743
rect 12256 5714 12308 5720
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12176 4826 12204 5034
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12268 4622 12296 5714
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12268 4146 12296 4558
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12254 3632 12310 3641
rect 12164 3596 12216 3602
rect 11992 3556 12164 3584
rect 12254 3567 12310 3576
rect 12164 3538 12216 3544
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11808 3194 11836 3402
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11256 1018 11284 2450
rect 11334 2000 11390 2009
rect 11390 1958 11468 1986
rect 11334 1935 11390 1944
rect 11440 1494 11468 1958
rect 11428 1488 11480 1494
rect 11428 1430 11480 1436
rect 11520 1216 11572 1222
rect 11520 1158 11572 1164
rect 11612 1216 11664 1222
rect 11612 1158 11664 1164
rect 11152 1012 11204 1018
rect 11152 954 11204 960
rect 11244 1012 11296 1018
rect 11244 954 11296 960
rect 11060 740 11112 746
rect 11060 682 11112 688
rect 11152 740 11204 746
rect 11152 682 11204 688
rect 10140 672 10192 678
rect 10140 614 10192 620
rect 10152 400 10180 614
rect 10364 572 10740 581
rect 10420 570 10444 572
rect 10500 570 10524 572
rect 10580 570 10604 572
rect 10660 570 10684 572
rect 10420 518 10430 570
rect 10674 518 10684 570
rect 10420 516 10444 518
rect 10500 516 10524 518
rect 10580 516 10604 518
rect 10660 516 10684 518
rect 10364 507 10740 516
rect 10888 428 11008 456
rect 10888 400 10916 428
rect 10048 196 10100 202
rect 10048 138 10100 144
rect 10138 0 10194 400
rect 10874 0 10930 400
rect 10980 354 11008 428
rect 11164 354 11192 682
rect 11428 672 11480 678
rect 11428 614 11480 620
rect 11440 406 11468 614
rect 10980 326 11192 354
rect 11428 400 11480 406
rect 11428 342 11480 348
rect 11532 202 11560 1158
rect 11624 400 11652 1158
rect 11808 814 11836 2926
rect 11900 1222 11928 3470
rect 12268 3398 12296 3567
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 2378 12112 2926
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 11980 1964 12032 1970
rect 11980 1906 12032 1912
rect 11888 1216 11940 1222
rect 11888 1158 11940 1164
rect 11796 808 11848 814
rect 11796 750 11848 756
rect 11520 196 11572 202
rect 11520 138 11572 144
rect 11610 0 11666 400
rect 11992 270 12020 1906
rect 12084 1358 12112 2042
rect 12164 1828 12216 1834
rect 12164 1770 12216 1776
rect 12176 1358 12204 1770
rect 12268 1748 12296 3334
rect 12360 2961 12388 6276
rect 12544 5658 12572 6598
rect 12636 5817 12664 8327
rect 12912 7546 12940 10934
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12806 6352 12862 6361
rect 12806 6287 12862 6296
rect 12820 6254 12848 6287
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12622 5808 12678 5817
rect 12678 5766 12756 5794
rect 12622 5743 12678 5752
rect 12452 5630 12572 5658
rect 12452 3738 12480 5630
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12544 3058 12572 5510
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12346 2952 12402 2961
rect 12346 2887 12402 2896
rect 12360 2582 12388 2887
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12544 2417 12572 2450
rect 12530 2408 12586 2417
rect 12440 2372 12492 2378
rect 12530 2343 12586 2352
rect 12440 2314 12492 2320
rect 12452 2038 12480 2314
rect 12440 2032 12492 2038
rect 12440 1974 12492 1980
rect 12636 1970 12664 5034
rect 12728 4842 12756 5766
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12820 5681 12848 5714
rect 12806 5672 12862 5681
rect 12912 5642 12940 7278
rect 13004 6236 13032 13518
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13188 13190 13216 14334
rect 13364 14172 13740 14181
rect 13420 14170 13444 14172
rect 13500 14170 13524 14172
rect 13580 14170 13604 14172
rect 13660 14170 13684 14172
rect 13420 14118 13430 14170
rect 13674 14118 13684 14170
rect 13420 14116 13444 14118
rect 13500 14116 13524 14118
rect 13580 14116 13604 14118
rect 13660 14116 13684 14118
rect 13364 14107 13740 14116
rect 13728 14068 13780 14074
rect 13832 14056 13860 14418
rect 13780 14028 13860 14056
rect 13728 14010 13780 14016
rect 13924 13938 13952 14418
rect 14016 14346 14044 14418
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 14006 14044 14282
rect 14108 14074 14136 14758
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 14002 13696 14058 13705
rect 13360 13456 13412 13462
rect 13280 13416 13360 13444
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13280 12986 13308 13416
rect 13360 13398 13412 13404
rect 13832 13394 13860 13670
rect 14108 13682 14136 13738
rect 14058 13654 14136 13682
rect 14002 13631 14058 13640
rect 14200 13546 14228 14962
rect 14108 13518 14228 13546
rect 14004 13456 14056 13462
rect 13924 13416 14004 13444
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13364 13084 13740 13093
rect 13420 13082 13444 13084
rect 13500 13082 13524 13084
rect 13580 13082 13604 13084
rect 13660 13082 13684 13084
rect 13420 13030 13430 13082
rect 13674 13030 13684 13082
rect 13420 13028 13444 13030
rect 13500 13028 13524 13030
rect 13580 13028 13604 13030
rect 13660 13028 13684 13030
rect 13364 13019 13740 13028
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 13096 11898 13124 12650
rect 13280 12442 13308 12922
rect 13728 12776 13780 12782
rect 13924 12764 13952 13416
rect 14004 13398 14056 13404
rect 13780 12736 13952 12764
rect 14004 12776 14056 12782
rect 13728 12718 13780 12724
rect 14108 12764 14136 13518
rect 14292 12866 14320 15302
rect 14384 15026 14412 16136
rect 14464 16118 14516 16124
rect 14844 15978 14872 16526
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15028 16114 15056 16458
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 15028 15706 15056 16050
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 15094 14596 15438
rect 15028 15162 15056 15642
rect 15120 15366 15148 17002
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 16046 15332 16390
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 15212 15570 15240 15914
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15396 15162 15424 17070
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 16590 15884 16934
rect 16224 16794 16252 17274
rect 16364 16892 16740 16901
rect 16420 16890 16444 16892
rect 16500 16890 16524 16892
rect 16580 16890 16604 16892
rect 16660 16890 16684 16892
rect 16420 16838 16430 16890
rect 16674 16838 16684 16890
rect 16420 16836 16444 16838
rect 16500 16836 16524 16838
rect 16580 16836 16604 16838
rect 16660 16836 16684 16838
rect 16364 16827 16740 16836
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15580 16046 15608 16390
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15488 15434 15516 15846
rect 15580 15706 15608 15846
rect 15764 15706 15792 15914
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14384 14482 14412 14962
rect 14556 14952 14608 14958
rect 14752 14940 14780 15030
rect 14608 14912 14780 14940
rect 15856 14906 15884 16526
rect 16040 15502 16068 16594
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 15706 16160 16390
rect 16364 15804 16740 15813
rect 16420 15802 16444 15804
rect 16500 15802 16524 15804
rect 16580 15802 16604 15804
rect 16660 15802 16684 15804
rect 16420 15750 16430 15802
rect 16674 15750 16684 15802
rect 16420 15748 16444 15750
rect 16500 15748 16524 15750
rect 16580 15748 16604 15750
rect 16660 15748 16684 15750
rect 16364 15739 16740 15748
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 14556 14894 14608 14900
rect 15672 14878 15884 14906
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14384 13870 14412 14418
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 12986 14596 13262
rect 14752 13258 14780 13738
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 14740 13252 14792 13258
rect 14660 13212 14740 13240
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14292 12838 14504 12866
rect 14056 12736 14136 12764
rect 14280 12776 14332 12782
rect 14004 12718 14056 12724
rect 14280 12718 14332 12724
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13096 11694 13124 11834
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13096 6662 13124 11290
rect 13188 10810 13216 11766
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13280 9586 13308 12378
rect 13648 12374 13676 12582
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13364 11996 13740 12005
rect 13420 11994 13444 11996
rect 13500 11994 13524 11996
rect 13580 11994 13604 11996
rect 13660 11994 13684 11996
rect 13420 11942 13430 11994
rect 13674 11942 13684 11994
rect 13420 11940 13444 11942
rect 13500 11940 13524 11942
rect 13580 11940 13604 11942
rect 13660 11940 13684 11942
rect 13364 11931 13740 11940
rect 13832 11880 13860 12242
rect 13740 11852 13860 11880
rect 13740 11558 13768 11852
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11132 13768 11494
rect 13832 11234 13860 11698
rect 13924 11354 13952 12242
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13832 11206 13952 11234
rect 13634 11112 13690 11121
rect 13740 11104 13860 11132
rect 13634 11047 13636 11056
rect 13688 11047 13690 11056
rect 13636 11018 13688 11024
rect 13364 10908 13740 10917
rect 13420 10906 13444 10908
rect 13500 10906 13524 10908
rect 13580 10906 13604 10908
rect 13660 10906 13684 10908
rect 13420 10854 13430 10906
rect 13674 10854 13684 10906
rect 13420 10852 13444 10854
rect 13500 10852 13524 10854
rect 13580 10852 13604 10854
rect 13660 10852 13684 10854
rect 13364 10843 13740 10852
rect 13358 10704 13414 10713
rect 13358 10639 13414 10648
rect 13372 10606 13400 10639
rect 13832 10606 13860 11104
rect 13924 10810 13952 11206
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14016 10674 14044 12718
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14108 10606 14136 11154
rect 13360 10600 13412 10606
rect 13820 10600 13872 10606
rect 13412 10560 13584 10588
rect 13360 10542 13412 10548
rect 13556 10470 13584 10560
rect 13820 10542 13872 10548
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10130 13584 10406
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13364 9820 13740 9829
rect 13420 9818 13444 9820
rect 13500 9818 13524 9820
rect 13580 9818 13604 9820
rect 13660 9818 13684 9820
rect 13420 9766 13430 9818
rect 13674 9766 13684 9818
rect 13420 9764 13444 9766
rect 13500 9764 13524 9766
rect 13580 9764 13604 9766
rect 13660 9764 13684 9766
rect 13364 9755 13740 9764
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13832 9178 13860 10202
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9722 13952 9998
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13188 8945 13216 9046
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13174 8936 13230 8945
rect 13174 8871 13230 8880
rect 13364 8732 13740 8741
rect 13420 8730 13444 8732
rect 13500 8730 13524 8732
rect 13580 8730 13604 8732
rect 13660 8730 13684 8732
rect 13420 8678 13430 8730
rect 13674 8678 13684 8730
rect 13420 8676 13444 8678
rect 13500 8676 13524 8678
rect 13580 8676 13604 8678
rect 13660 8676 13684 8678
rect 13364 8667 13740 8676
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13188 7954 13216 8570
rect 13832 8498 13860 8978
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13556 7954 13584 8230
rect 13648 7954 13676 8230
rect 13832 8090 13860 8230
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13832 7954 13860 8026
rect 13176 7948 13228 7954
rect 13544 7948 13596 7954
rect 13228 7908 13308 7936
rect 13176 7890 13228 7896
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13004 6208 13124 6236
rect 12990 5944 13046 5953
rect 12990 5879 13046 5888
rect 12806 5607 12862 5616
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12806 5536 12862 5545
rect 12806 5471 12862 5480
rect 12820 5370 12848 5471
rect 12898 5400 12954 5409
rect 12808 5364 12860 5370
rect 12898 5335 12954 5344
rect 12808 5306 12860 5312
rect 12912 5302 12940 5335
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12912 5166 12940 5238
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12728 4814 12848 4842
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12728 2582 12756 4558
rect 12820 4146 12848 4814
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12912 3126 12940 3470
rect 13004 3233 13032 5879
rect 12990 3224 13046 3233
rect 12990 3159 13046 3168
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12808 2372 12860 2378
rect 12728 2332 12808 2360
rect 12624 1964 12676 1970
rect 12624 1906 12676 1912
rect 12348 1896 12400 1902
rect 12346 1864 12348 1873
rect 12440 1896 12492 1902
rect 12400 1864 12402 1873
rect 12440 1838 12492 1844
rect 12346 1799 12402 1808
rect 12452 1748 12480 1838
rect 12268 1720 12480 1748
rect 12452 1562 12480 1720
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12440 1556 12492 1562
rect 12440 1498 12492 1504
rect 12532 1556 12584 1562
rect 12532 1498 12584 1504
rect 12544 1408 12572 1498
rect 12452 1380 12572 1408
rect 12072 1352 12124 1358
rect 12072 1294 12124 1300
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 12452 814 12480 1380
rect 12636 1306 12664 1702
rect 12728 1426 12756 2332
rect 12808 2314 12860 2320
rect 12806 2000 12862 2009
rect 12806 1935 12862 1944
rect 12716 1420 12768 1426
rect 12820 1408 12848 1935
rect 13004 1426 13032 2994
rect 13096 2145 13124 6208
rect 13188 4690 13216 7142
rect 13280 6934 13308 7908
rect 13544 7890 13596 7896
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13556 7818 13584 7890
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13832 7750 13860 7890
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13364 7644 13740 7653
rect 13420 7642 13444 7644
rect 13500 7642 13524 7644
rect 13580 7642 13604 7644
rect 13660 7642 13684 7644
rect 13420 7590 13430 7642
rect 13674 7590 13684 7642
rect 13420 7588 13444 7590
rect 13500 7588 13524 7590
rect 13580 7588 13604 7590
rect 13660 7588 13684 7590
rect 13364 7579 13740 7588
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13280 5778 13308 6870
rect 13364 6556 13740 6565
rect 13420 6554 13444 6556
rect 13500 6554 13524 6556
rect 13580 6554 13604 6556
rect 13660 6554 13684 6556
rect 13420 6502 13430 6554
rect 13674 6502 13684 6554
rect 13420 6500 13444 6502
rect 13500 6500 13524 6502
rect 13580 6500 13604 6502
rect 13660 6500 13684 6502
rect 13364 6491 13740 6500
rect 13832 6322 13860 7482
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13634 6216 13690 6225
rect 13634 6151 13690 6160
rect 13542 5808 13598 5817
rect 13268 5772 13320 5778
rect 13648 5778 13676 6151
rect 13542 5743 13598 5752
rect 13636 5772 13688 5778
rect 13268 5714 13320 5720
rect 13556 5642 13584 5743
rect 13636 5714 13688 5720
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13188 2854 13216 4014
rect 13280 3738 13308 5510
rect 13364 5468 13740 5477
rect 13420 5466 13444 5468
rect 13500 5466 13524 5468
rect 13580 5466 13604 5468
rect 13660 5466 13684 5468
rect 13420 5414 13430 5466
rect 13674 5414 13684 5466
rect 13420 5412 13444 5414
rect 13500 5412 13524 5414
rect 13580 5412 13604 5414
rect 13660 5412 13684 5414
rect 13364 5403 13740 5412
rect 13832 5352 13860 5714
rect 13740 5324 13860 5352
rect 13740 5166 13768 5324
rect 13924 5284 13952 9046
rect 13832 5256 13952 5284
rect 13360 5160 13412 5166
rect 13358 5128 13360 5137
rect 13728 5160 13780 5166
rect 13412 5128 13414 5137
rect 13728 5102 13780 5108
rect 13358 5063 13414 5072
rect 13364 4380 13740 4389
rect 13420 4378 13444 4380
rect 13500 4378 13524 4380
rect 13580 4378 13604 4380
rect 13660 4378 13684 4380
rect 13420 4326 13430 4378
rect 13674 4326 13684 4378
rect 13420 4324 13444 4326
rect 13500 4324 13524 4326
rect 13580 4324 13604 4326
rect 13660 4324 13684 4326
rect 13364 4315 13740 4324
rect 13832 4078 13860 5256
rect 14016 4622 14044 9318
rect 14108 7018 14136 10542
rect 14200 8430 14228 12650
rect 14292 12170 14320 12718
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14292 11257 14320 12106
rect 14370 11656 14426 11665
rect 14370 11591 14426 11600
rect 14384 11558 14412 11591
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14278 11248 14334 11257
rect 14278 11183 14334 11192
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14292 9654 14320 11018
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14384 9518 14412 10474
rect 14476 10130 14504 12838
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14568 11150 14596 12310
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14292 9178 14320 9454
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14384 8294 14412 9318
rect 14476 8906 14504 9454
rect 14568 9382 14596 10950
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14200 7954 14228 8230
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 7177 14228 7890
rect 14292 7342 14320 8230
rect 14370 7440 14426 7449
rect 14370 7375 14372 7384
rect 14424 7375 14426 7384
rect 14372 7346 14424 7352
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14186 7168 14242 7177
rect 14186 7103 14242 7112
rect 14108 6990 14320 7018
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 14108 5681 14136 6870
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14200 6089 14228 6190
rect 14186 6080 14242 6089
rect 14186 6015 14242 6024
rect 14094 5672 14150 5681
rect 14094 5607 14150 5616
rect 14108 5574 14136 5607
rect 14200 5574 14228 6015
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13372 3482 13400 3878
rect 13464 3738 13492 3946
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13556 3534 13584 3878
rect 13832 3738 13860 4014
rect 13924 3738 13952 4558
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 14016 3602 14044 4218
rect 14108 4078 14136 5170
rect 14292 5166 14320 6990
rect 14384 6934 14412 7346
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14200 4026 14228 4422
rect 14384 4282 14412 6666
rect 14476 4758 14504 8842
rect 14568 7954 14596 8978
rect 14660 8106 14688 13212
rect 14740 13194 14792 13200
rect 14936 12782 14964 13330
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 11830 14872 12582
rect 15212 12186 15240 12718
rect 15304 12714 15332 13194
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 14936 12158 15240 12186
rect 14936 12102 14964 12158
rect 14924 12096 14976 12102
rect 15200 12096 15252 12102
rect 14924 12038 14976 12044
rect 15120 12056 15200 12084
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14936 11694 14964 12038
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14752 11286 14780 11630
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14936 11218 14964 11630
rect 15120 11626 15148 12056
rect 15200 12038 15252 12044
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 15120 11218 15148 11562
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14752 8242 14780 9998
rect 14844 8537 14872 10746
rect 14936 9518 14964 11154
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14830 8528 14886 8537
rect 14936 8498 14964 9454
rect 14830 8463 14886 8472
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14752 8214 14964 8242
rect 14660 8078 14872 8106
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14568 6254 14596 7890
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 6934 14688 7754
rect 14752 7546 14780 7890
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14648 6928 14700 6934
rect 14700 6888 14780 6916
rect 14648 6870 14700 6876
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14568 5234 14596 5714
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14464 4752 14516 4758
rect 14516 4712 14596 4740
rect 14464 4694 14516 4700
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14200 3998 14412 4026
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 14200 3534 14228 3674
rect 13280 3454 13400 3482
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13082 2136 13138 2145
rect 13082 2071 13138 2080
rect 13084 2032 13136 2038
rect 13084 1974 13136 1980
rect 12900 1420 12952 1426
rect 12820 1380 12900 1408
rect 12716 1362 12768 1368
rect 12900 1362 12952 1368
rect 12992 1420 13044 1426
rect 12992 1362 13044 1368
rect 12544 1278 12664 1306
rect 12440 808 12492 814
rect 12440 750 12492 756
rect 12348 740 12400 746
rect 12348 682 12400 688
rect 12360 400 12388 682
rect 11980 264 12032 270
rect 11980 206 12032 212
rect 12346 0 12402 400
rect 12544 338 12572 1278
rect 12728 882 12756 1362
rect 12808 1012 12860 1018
rect 12808 954 12860 960
rect 12716 876 12768 882
rect 12716 818 12768 824
rect 12820 474 12848 954
rect 12912 678 12940 1362
rect 13096 898 13124 1974
rect 13188 1834 13216 2790
rect 13176 1828 13228 1834
rect 13176 1770 13228 1776
rect 13280 1494 13308 3454
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 14004 3392 14056 3398
rect 14292 3346 14320 3878
rect 14004 3334 14056 3340
rect 13364 3292 13740 3301
rect 13420 3290 13444 3292
rect 13500 3290 13524 3292
rect 13580 3290 13604 3292
rect 13660 3290 13684 3292
rect 13420 3238 13430 3290
rect 13674 3238 13684 3290
rect 13420 3236 13444 3238
rect 13500 3236 13524 3238
rect 13580 3236 13604 3238
rect 13660 3236 13684 3238
rect 13364 3227 13740 3236
rect 13924 3126 13952 3334
rect 13728 3120 13780 3126
rect 13912 3120 13964 3126
rect 13728 3062 13780 3068
rect 13818 3088 13874 3097
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13372 2854 13400 2926
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13740 2394 13768 3062
rect 13912 3062 13964 3068
rect 13818 3023 13820 3032
rect 13872 3023 13874 3032
rect 13820 2994 13872 3000
rect 14016 2582 14044 3334
rect 14108 3318 14320 3346
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 13740 2366 13860 2394
rect 13364 2204 13740 2213
rect 13420 2202 13444 2204
rect 13500 2202 13524 2204
rect 13580 2202 13604 2204
rect 13660 2202 13684 2204
rect 13420 2150 13430 2202
rect 13674 2150 13684 2202
rect 13420 2148 13444 2150
rect 13500 2148 13524 2150
rect 13580 2148 13604 2150
rect 13660 2148 13684 2150
rect 13364 2139 13740 2148
rect 13358 2000 13414 2009
rect 13832 1986 13860 2366
rect 14004 2304 14056 2310
rect 13910 2272 13966 2281
rect 14004 2246 14056 2252
rect 13910 2207 13966 2216
rect 13648 1970 13860 1986
rect 13924 1970 13952 2207
rect 13358 1935 13360 1944
rect 13412 1935 13414 1944
rect 13636 1964 13860 1970
rect 13360 1906 13412 1912
rect 13688 1958 13860 1964
rect 13912 1964 13964 1970
rect 13636 1906 13688 1912
rect 13912 1906 13964 1912
rect 13372 1850 13400 1906
rect 13820 1896 13872 1902
rect 13372 1822 13492 1850
rect 13820 1838 13872 1844
rect 13464 1562 13492 1822
rect 13832 1737 13860 1838
rect 13818 1728 13874 1737
rect 13818 1663 13874 1672
rect 13910 1592 13966 1601
rect 13452 1556 13504 1562
rect 13910 1527 13966 1536
rect 13452 1498 13504 1504
rect 13176 1488 13228 1494
rect 13176 1430 13228 1436
rect 13268 1488 13320 1494
rect 13268 1430 13320 1436
rect 13188 1018 13216 1430
rect 13360 1420 13412 1426
rect 13464 1408 13492 1498
rect 13924 1426 13952 1527
rect 13412 1380 13492 1408
rect 13912 1420 13964 1426
rect 13360 1362 13412 1368
rect 13912 1362 13964 1368
rect 13364 1116 13740 1125
rect 13420 1114 13444 1116
rect 13500 1114 13524 1116
rect 13580 1114 13604 1116
rect 13660 1114 13684 1116
rect 13420 1062 13430 1114
rect 13674 1062 13684 1114
rect 13420 1060 13444 1062
rect 13500 1060 13524 1062
rect 13580 1060 13604 1062
rect 13660 1060 13684 1062
rect 13364 1051 13740 1060
rect 13176 1012 13228 1018
rect 13176 954 13228 960
rect 13096 870 13308 898
rect 13280 814 13308 870
rect 13360 876 13412 882
rect 13360 818 13412 824
rect 13268 808 13320 814
rect 13268 750 13320 756
rect 12900 672 12952 678
rect 12900 614 12952 620
rect 12912 474 12940 614
rect 13372 490 13400 818
rect 13924 814 13952 1362
rect 14016 1193 14044 2246
rect 14108 1426 14136 3318
rect 14186 3088 14242 3097
rect 14186 3023 14242 3032
rect 14200 2938 14228 3023
rect 14200 2910 14320 2938
rect 14292 2854 14320 2910
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14200 2666 14228 2790
rect 14200 2638 14320 2666
rect 14292 2514 14320 2638
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14188 2100 14240 2106
rect 14188 2042 14240 2048
rect 14096 1420 14148 1426
rect 14096 1362 14148 1368
rect 14096 1284 14148 1290
rect 14096 1226 14148 1232
rect 14002 1184 14058 1193
rect 14002 1119 14058 1128
rect 14004 944 14056 950
rect 14004 886 14056 892
rect 13912 808 13964 814
rect 13912 750 13964 756
rect 14016 490 14044 886
rect 14108 814 14136 1226
rect 14200 1018 14228 2042
rect 14292 1018 14320 2246
rect 14384 1426 14412 3998
rect 14476 3602 14504 4422
rect 14568 4282 14596 4712
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3641 14596 3878
rect 14554 3632 14610 3641
rect 14464 3596 14516 3602
rect 14554 3567 14610 3576
rect 14464 3538 14516 3544
rect 14660 3534 14688 4422
rect 14752 3602 14780 6888
rect 14844 6730 14872 8078
rect 14936 7954 14964 8214
rect 14924 7948 14976 7954
rect 15028 7936 15056 11086
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15120 10062 15148 10474
rect 15212 10266 15240 10678
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15304 10266 15332 10610
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15212 8090 15240 8774
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15200 7948 15252 7954
rect 15028 7908 15148 7936
rect 14924 7890 14976 7896
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14936 7410 14964 7686
rect 15028 7410 15056 7686
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14936 7041 14964 7142
rect 14922 7032 14978 7041
rect 14922 6967 14978 6976
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14830 6352 14886 6361
rect 14936 6338 14964 6734
rect 14886 6310 14964 6338
rect 14830 6287 14832 6296
rect 14884 6287 14886 6296
rect 14832 6258 14884 6264
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14844 4146 14872 6054
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14568 3194 14596 3402
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14554 2680 14610 2689
rect 14554 2615 14610 2624
rect 14568 2514 14596 2615
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14568 1902 14596 2246
rect 14556 1896 14608 1902
rect 14556 1838 14608 1844
rect 14372 1420 14424 1426
rect 14372 1362 14424 1368
rect 14660 1018 14688 3334
rect 14752 2990 14780 3538
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14752 2310 14780 2586
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14844 2106 14872 3878
rect 15028 3738 15056 7142
rect 15120 4690 15148 7908
rect 15200 7890 15252 7896
rect 15212 7002 15240 7890
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15212 5846 15240 6122
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15120 4282 15148 4626
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15212 4146 15240 5510
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15198 4040 15254 4049
rect 15304 4026 15332 10066
rect 15396 7342 15424 13126
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15488 12442 15516 12650
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15580 12322 15608 13330
rect 15488 12294 15608 12322
rect 15488 10554 15516 12294
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15580 10674 15608 11834
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15488 10526 15608 10554
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15254 3998 15332 4026
rect 15198 3975 15254 3984
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 15396 3534 15424 6938
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15028 3126 15056 3470
rect 15488 3380 15516 9862
rect 15580 7478 15608 10526
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15672 7342 15700 14878
rect 15948 14770 15976 15302
rect 15856 14742 15976 14770
rect 15750 14376 15806 14385
rect 15750 14311 15752 14320
rect 15804 14311 15806 14320
rect 15752 14282 15804 14288
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15764 13530 15792 13806
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 10130 15792 13126
rect 15856 11098 15884 14742
rect 16364 14716 16740 14725
rect 16420 14714 16444 14716
rect 16500 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16420 14662 16430 14714
rect 16674 14662 16684 14714
rect 16420 14660 16444 14662
rect 16500 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16364 14651 16740 14660
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15948 14006 15976 14418
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 15936 14000 15988 14006
rect 15936 13942 15988 13948
rect 16040 13394 16068 14282
rect 16868 13954 16896 15302
rect 16960 14521 16988 17845
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15706 17080 15846
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 16946 14512 17002 14521
rect 16946 14447 17002 14456
rect 16212 13932 16264 13938
rect 16132 13892 16212 13920
rect 16132 13705 16160 13892
rect 16212 13874 16264 13880
rect 16396 13932 16448 13938
rect 16868 13926 16988 13954
rect 16396 13874 16448 13880
rect 16408 13818 16436 13874
rect 16224 13790 16436 13818
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16118 13696 16174 13705
rect 16118 13631 16174 13640
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15948 12646 15976 13330
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16224 12434 16252 13790
rect 16364 13628 16740 13637
rect 16420 13626 16444 13628
rect 16500 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16420 13574 16430 13626
rect 16674 13574 16684 13626
rect 16420 13572 16444 13574
rect 16500 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16364 13563 16740 13572
rect 16776 13394 16804 13806
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16408 12714 16436 13330
rect 16868 12986 16896 13806
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16364 12540 16740 12549
rect 16420 12538 16444 12540
rect 16500 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16420 12486 16430 12538
rect 16674 12486 16684 12538
rect 16420 12484 16444 12486
rect 16500 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16364 12475 16740 12484
rect 16960 12442 16988 13926
rect 17052 13802 17080 14758
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17040 13796 17092 13802
rect 17040 13738 17092 13744
rect 16040 12406 16252 12434
rect 16948 12436 17000 12442
rect 15856 11070 15976 11098
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15856 10742 15884 10950
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15750 9072 15806 9081
rect 15750 9007 15752 9016
rect 15804 9007 15806 9016
rect 15752 8978 15804 8984
rect 15750 8528 15806 8537
rect 15750 8463 15806 8472
rect 15764 8022 15792 8463
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15580 6458 15608 7278
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15580 6254 15608 6394
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5914 15608 6054
rect 15568 5908 15620 5914
rect 15764 5896 15792 7414
rect 15856 6458 15884 10542
rect 15948 6866 15976 11070
rect 16040 10062 16068 12406
rect 16948 12378 17000 12384
rect 17052 12238 17080 13738
rect 17144 13530 17172 13942
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17144 12782 17172 13126
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17236 12866 17264 12922
rect 17236 12838 17356 12866
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16132 11354 16160 11562
rect 16224 11354 16252 12038
rect 16364 11452 16740 11461
rect 16420 11450 16444 11452
rect 16500 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16420 11398 16430 11450
rect 16674 11398 16684 11450
rect 16420 11396 16444 11398
rect 16500 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16364 11387 16740 11396
rect 16960 11354 16988 12038
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16224 10674 16252 11290
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16316 10810 16344 11154
rect 16592 11121 16620 11154
rect 16578 11112 16634 11121
rect 16634 11070 16804 11098
rect 16578 11047 16634 11056
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16224 9625 16252 10406
rect 16364 10364 16740 10373
rect 16420 10362 16444 10364
rect 16500 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16420 10310 16430 10362
rect 16674 10310 16684 10362
rect 16420 10308 16444 10310
rect 16500 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16364 10299 16740 10308
rect 16776 10130 16804 11070
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16210 9616 16266 9625
rect 16210 9551 16266 9560
rect 16224 9518 16252 9551
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16364 9276 16740 9285
rect 16420 9274 16444 9276
rect 16500 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16420 9222 16430 9274
rect 16674 9222 16684 9274
rect 16420 9220 16444 9222
rect 16500 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16364 9211 16740 9220
rect 16776 9178 16804 10066
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16868 9042 16896 9318
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 16040 5914 16068 8910
rect 16868 8634 16896 8978
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16364 8188 16740 8197
rect 16420 8186 16444 8188
rect 16500 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16420 8134 16430 8186
rect 16674 8134 16684 8186
rect 16420 8132 16444 8134
rect 16500 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16364 8123 16740 8132
rect 16776 8090 16804 8298
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16224 6934 16252 7278
rect 16364 7100 16740 7109
rect 16420 7098 16444 7100
rect 16500 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16420 7046 16430 7098
rect 16674 7046 16684 7098
rect 16420 7044 16444 7046
rect 16500 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16364 7035 16740 7044
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16132 6254 16160 6802
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16132 5914 16160 6054
rect 16224 5914 16252 6394
rect 16500 6236 16528 6870
rect 16580 6248 16632 6254
rect 16500 6208 16580 6236
rect 16580 6190 16632 6196
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16364 6012 16740 6021
rect 16420 6010 16444 6012
rect 16500 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16420 5958 16430 6010
rect 16674 5958 16684 6010
rect 16420 5956 16444 5958
rect 16500 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16364 5947 16740 5956
rect 15568 5850 15620 5856
rect 15672 5868 15792 5896
rect 16028 5908 16080 5914
rect 15672 4758 15700 5868
rect 16028 5850 16080 5856
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16040 5794 16068 5850
rect 16868 5817 16896 6054
rect 16854 5808 16910 5817
rect 15752 5772 15804 5778
rect 16040 5766 16252 5794
rect 16224 5760 16252 5766
rect 16396 5772 16448 5778
rect 16224 5732 16396 5760
rect 15752 5714 15804 5720
rect 16854 5743 16910 5752
rect 16396 5714 16448 5720
rect 15764 5302 15792 5714
rect 16960 5658 16988 10406
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17052 9654 17080 10066
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17052 9178 17080 9590
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17144 8974 17172 9862
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17144 5778 17172 8774
rect 17236 7342 17264 12378
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17236 6254 17264 7278
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16868 5630 16988 5658
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 16364 4924 16740 4933
rect 16420 4922 16444 4924
rect 16500 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16420 4870 16430 4922
rect 16674 4870 16684 4922
rect 16420 4868 16444 4870
rect 16500 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16364 4859 16740 4868
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15672 4282 15700 4694
rect 16776 4690 16804 5578
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 15566 3904 15622 3913
rect 15566 3839 15622 3848
rect 15396 3352 15516 3380
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2514 14964 2790
rect 15028 2582 15056 3062
rect 15292 2984 15344 2990
rect 15290 2952 15292 2961
rect 15344 2952 15346 2961
rect 15290 2887 15346 2896
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 14924 2508 14976 2514
rect 14924 2450 14976 2456
rect 14832 2100 14884 2106
rect 14832 2042 14884 2048
rect 15120 1970 15148 2790
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 15108 1964 15160 1970
rect 15108 1906 15160 1912
rect 14924 1896 14976 1902
rect 14922 1864 14924 1873
rect 15016 1896 15068 1902
rect 14976 1864 14978 1873
rect 15016 1838 15068 1844
rect 14922 1799 14978 1808
rect 14740 1420 14792 1426
rect 14740 1362 14792 1368
rect 14188 1012 14240 1018
rect 14188 954 14240 960
rect 14280 1012 14332 1018
rect 14280 954 14332 960
rect 14648 1012 14700 1018
rect 14648 954 14700 960
rect 14096 808 14148 814
rect 14096 750 14148 756
rect 14372 808 14424 814
rect 14372 750 14424 756
rect 12808 468 12860 474
rect 12808 410 12860 416
rect 12900 468 12952 474
rect 12900 410 12952 416
rect 13096 462 13400 490
rect 13832 462 14044 490
rect 13096 400 13124 462
rect 13832 400 13860 462
rect 12532 332 12584 338
rect 12532 274 12584 280
rect 13082 0 13138 400
rect 13818 0 13874 400
rect 14108 270 14136 750
rect 14384 474 14412 750
rect 14372 468 14424 474
rect 14372 410 14424 416
rect 14568 462 14688 490
rect 14752 474 14780 1362
rect 14924 1216 14976 1222
rect 14924 1158 14976 1164
rect 14936 1034 14964 1158
rect 14844 1006 14964 1034
rect 15028 1018 15056 1838
rect 15120 1426 15148 1906
rect 15108 1420 15160 1426
rect 15108 1362 15160 1368
rect 15106 1320 15162 1329
rect 15212 1290 15240 2518
rect 15396 2514 15424 3352
rect 15580 2854 15608 3839
rect 16132 3194 16160 4014
rect 16224 3534 16252 4422
rect 16776 4214 16804 4626
rect 16868 4622 16896 5630
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16776 4078 16804 4150
rect 16960 4078 16988 5510
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16364 3836 16740 3845
rect 16420 3834 16444 3836
rect 16500 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16420 3782 16430 3834
rect 16674 3782 16684 3834
rect 16420 3780 16444 3782
rect 16500 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16364 3771 16740 3780
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16224 3194 16252 3470
rect 16776 3398 16804 4014
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16868 3602 16896 3946
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16868 3058 16896 3538
rect 17052 3534 17080 4558
rect 17328 4078 17356 12838
rect 17420 12238 17448 13670
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17420 8838 17448 9522
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17144 3046 17448 3074
rect 17144 2990 17172 3046
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15580 2514 15608 2790
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 2145 15332 2246
rect 15290 2136 15346 2145
rect 15290 2071 15346 2080
rect 15396 1902 15424 2450
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15488 2106 15516 2246
rect 15476 2100 15528 2106
rect 15476 2042 15528 2048
rect 15384 1896 15436 1902
rect 15384 1838 15436 1844
rect 15474 1864 15530 1873
rect 15292 1556 15344 1562
rect 15292 1498 15344 1504
rect 15106 1255 15162 1264
rect 15200 1284 15252 1290
rect 15016 1012 15068 1018
rect 14568 400 14596 462
rect 14096 264 14148 270
rect 14096 206 14148 212
rect 14554 0 14610 400
rect 14660 354 14688 462
rect 14740 468 14792 474
rect 14740 410 14792 416
rect 14844 354 14872 1006
rect 15016 954 15068 960
rect 15120 814 15148 1255
rect 15200 1226 15252 1232
rect 15198 1184 15254 1193
rect 15198 1119 15254 1128
rect 15212 814 15240 1119
rect 15108 808 15160 814
rect 15108 750 15160 756
rect 15200 808 15252 814
rect 15200 750 15252 756
rect 15304 400 15332 1498
rect 15396 1290 15424 1838
rect 15474 1799 15530 1808
rect 15488 1562 15516 1799
rect 15580 1766 15608 2314
rect 15844 2304 15896 2310
rect 16028 2304 16080 2310
rect 15844 2246 15896 2252
rect 16026 2272 16028 2281
rect 16080 2272 16082 2281
rect 15658 2136 15714 2145
rect 15658 2071 15714 2080
rect 15672 1970 15700 2071
rect 15660 1964 15712 1970
rect 15660 1906 15712 1912
rect 15568 1760 15620 1766
rect 15568 1702 15620 1708
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15750 1728 15806 1737
rect 15476 1556 15528 1562
rect 15476 1498 15528 1504
rect 15672 1465 15700 1702
rect 15750 1663 15806 1672
rect 15658 1456 15714 1465
rect 15764 1426 15792 1663
rect 15658 1391 15714 1400
rect 15752 1420 15804 1426
rect 15752 1362 15804 1368
rect 15384 1284 15436 1290
rect 15384 1226 15436 1232
rect 15856 1170 15884 2246
rect 16026 2207 16082 2216
rect 15936 1828 15988 1834
rect 15936 1770 15988 1776
rect 16028 1828 16080 1834
rect 16028 1770 16080 1776
rect 15948 1426 15976 1770
rect 16040 1562 16068 1770
rect 16028 1556 16080 1562
rect 16028 1498 16080 1504
rect 15936 1420 15988 1426
rect 15936 1362 15988 1368
rect 15856 1142 16068 1170
rect 16040 400 16068 1142
rect 16132 678 16160 2926
rect 16948 2916 17000 2922
rect 17224 2916 17276 2922
rect 17000 2876 17080 2904
rect 16948 2858 17000 2864
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16364 2748 16740 2757
rect 16420 2746 16444 2748
rect 16500 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16420 2694 16430 2746
rect 16674 2694 16684 2746
rect 16420 2692 16444 2694
rect 16500 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16364 2683 16740 2692
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16224 1873 16252 2586
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16408 1986 16436 2246
rect 16500 2106 16528 2246
rect 16488 2100 16540 2106
rect 16488 2042 16540 2048
rect 16580 2032 16632 2038
rect 16408 1980 16580 1986
rect 16408 1974 16632 1980
rect 16408 1958 16620 1974
rect 16210 1864 16266 1873
rect 16266 1822 16528 1850
rect 16210 1799 16266 1808
rect 16500 1766 16528 1822
rect 16488 1760 16540 1766
rect 16488 1702 16540 1708
rect 16364 1660 16740 1669
rect 16420 1658 16444 1660
rect 16500 1658 16524 1660
rect 16580 1658 16604 1660
rect 16660 1658 16684 1660
rect 16420 1606 16430 1658
rect 16674 1606 16684 1658
rect 16420 1604 16444 1606
rect 16500 1604 16524 1606
rect 16580 1604 16604 1606
rect 16660 1604 16684 1606
rect 16364 1595 16740 1604
rect 16212 740 16264 746
rect 16212 682 16264 688
rect 16120 672 16172 678
rect 16120 614 16172 620
rect 16224 474 16252 682
rect 16364 572 16740 581
rect 16420 570 16444 572
rect 16500 570 16524 572
rect 16580 570 16604 572
rect 16660 570 16684 572
rect 16420 518 16430 570
rect 16674 518 16684 570
rect 16420 516 16444 518
rect 16500 516 16524 518
rect 16580 516 16604 518
rect 16660 516 16684 518
rect 16364 507 16740 516
rect 16212 468 16264 474
rect 16212 410 16264 416
rect 16776 400 16804 2790
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 814 16896 2246
rect 17052 1902 17080 2876
rect 17224 2858 17276 2864
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17040 1896 17092 1902
rect 17040 1838 17092 1844
rect 17040 1420 17092 1426
rect 17040 1362 17092 1368
rect 17052 1018 17080 1362
rect 17040 1012 17092 1018
rect 17040 954 17092 960
rect 17144 882 17172 2586
rect 17236 1494 17264 2858
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17328 1902 17356 2790
rect 17316 1896 17368 1902
rect 17316 1838 17368 1844
rect 17420 1494 17448 3046
rect 17512 2582 17540 11018
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17604 2582 17632 10202
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 17224 1488 17276 1494
rect 17224 1430 17276 1436
rect 17408 1488 17460 1494
rect 17408 1430 17460 1436
rect 17132 876 17184 882
rect 17132 818 17184 824
rect 16856 808 16908 814
rect 16856 750 16908 756
rect 17512 400 17540 2314
rect 14660 326 14872 354
rect 15290 0 15346 400
rect 16026 0 16082 400
rect 16762 0 16818 400
rect 17498 0 17554 400
<< via2 >>
rect 1364 17434 1420 17436
rect 1444 17434 1500 17436
rect 1524 17434 1580 17436
rect 1604 17434 1660 17436
rect 1684 17434 1740 17436
rect 1364 17382 1366 17434
rect 1366 17382 1418 17434
rect 1418 17382 1420 17434
rect 1444 17382 1482 17434
rect 1482 17382 1494 17434
rect 1494 17382 1500 17434
rect 1524 17382 1546 17434
rect 1546 17382 1558 17434
rect 1558 17382 1580 17434
rect 1604 17382 1610 17434
rect 1610 17382 1622 17434
rect 1622 17382 1660 17434
rect 1684 17382 1686 17434
rect 1686 17382 1738 17434
rect 1738 17382 1740 17434
rect 1364 17380 1420 17382
rect 1444 17380 1500 17382
rect 1524 17380 1580 17382
rect 1604 17380 1660 17382
rect 1684 17380 1740 17382
rect 4364 16890 4420 16892
rect 4444 16890 4500 16892
rect 4524 16890 4580 16892
rect 4604 16890 4660 16892
rect 4684 16890 4740 16892
rect 4364 16838 4366 16890
rect 4366 16838 4418 16890
rect 4418 16838 4420 16890
rect 4444 16838 4482 16890
rect 4482 16838 4494 16890
rect 4494 16838 4500 16890
rect 4524 16838 4546 16890
rect 4546 16838 4558 16890
rect 4558 16838 4580 16890
rect 4604 16838 4610 16890
rect 4610 16838 4622 16890
rect 4622 16838 4660 16890
rect 4684 16838 4686 16890
rect 4686 16838 4738 16890
rect 4738 16838 4740 16890
rect 4364 16836 4420 16838
rect 4444 16836 4500 16838
rect 4524 16836 4580 16838
rect 4604 16836 4660 16838
rect 4684 16836 4740 16838
rect 4894 16632 4950 16688
rect 1364 16346 1420 16348
rect 1444 16346 1500 16348
rect 1524 16346 1580 16348
rect 1604 16346 1660 16348
rect 1684 16346 1740 16348
rect 1364 16294 1366 16346
rect 1366 16294 1418 16346
rect 1418 16294 1420 16346
rect 1444 16294 1482 16346
rect 1482 16294 1494 16346
rect 1494 16294 1500 16346
rect 1524 16294 1546 16346
rect 1546 16294 1558 16346
rect 1558 16294 1580 16346
rect 1604 16294 1610 16346
rect 1610 16294 1622 16346
rect 1622 16294 1660 16346
rect 1684 16294 1686 16346
rect 1686 16294 1738 16346
rect 1738 16294 1740 16346
rect 1364 16292 1420 16294
rect 1444 16292 1500 16294
rect 1524 16292 1580 16294
rect 1604 16292 1660 16294
rect 1684 16292 1740 16294
rect 2042 15700 2098 15736
rect 2042 15680 2044 15700
rect 2044 15680 2096 15700
rect 2096 15680 2098 15700
rect 1364 15258 1420 15260
rect 1444 15258 1500 15260
rect 1524 15258 1580 15260
rect 1604 15258 1660 15260
rect 1684 15258 1740 15260
rect 1364 15206 1366 15258
rect 1366 15206 1418 15258
rect 1418 15206 1420 15258
rect 1444 15206 1482 15258
rect 1482 15206 1494 15258
rect 1494 15206 1500 15258
rect 1524 15206 1546 15258
rect 1546 15206 1558 15258
rect 1558 15206 1580 15258
rect 1604 15206 1610 15258
rect 1610 15206 1622 15258
rect 1622 15206 1660 15258
rect 1684 15206 1686 15258
rect 1686 15206 1738 15258
rect 1738 15206 1740 15258
rect 1364 15204 1420 15206
rect 1444 15204 1500 15206
rect 1524 15204 1580 15206
rect 1604 15204 1660 15206
rect 1684 15204 1740 15206
rect 2686 14864 2742 14920
rect 1364 14170 1420 14172
rect 1444 14170 1500 14172
rect 1524 14170 1580 14172
rect 1604 14170 1660 14172
rect 1684 14170 1740 14172
rect 1364 14118 1366 14170
rect 1366 14118 1418 14170
rect 1418 14118 1420 14170
rect 1444 14118 1482 14170
rect 1482 14118 1494 14170
rect 1494 14118 1500 14170
rect 1524 14118 1546 14170
rect 1546 14118 1558 14170
rect 1558 14118 1580 14170
rect 1604 14118 1610 14170
rect 1610 14118 1622 14170
rect 1622 14118 1660 14170
rect 1684 14118 1686 14170
rect 1686 14118 1738 14170
rect 1738 14118 1740 14170
rect 1364 14116 1420 14118
rect 1444 14116 1500 14118
rect 1524 14116 1580 14118
rect 1604 14116 1660 14118
rect 1684 14116 1740 14118
rect 1364 13082 1420 13084
rect 1444 13082 1500 13084
rect 1524 13082 1580 13084
rect 1604 13082 1660 13084
rect 1684 13082 1740 13084
rect 1364 13030 1366 13082
rect 1366 13030 1418 13082
rect 1418 13030 1420 13082
rect 1444 13030 1482 13082
rect 1482 13030 1494 13082
rect 1494 13030 1500 13082
rect 1524 13030 1546 13082
rect 1546 13030 1558 13082
rect 1558 13030 1580 13082
rect 1604 13030 1610 13082
rect 1610 13030 1622 13082
rect 1622 13030 1660 13082
rect 1684 13030 1686 13082
rect 1686 13030 1738 13082
rect 1738 13030 1740 13082
rect 1364 13028 1420 13030
rect 1444 13028 1500 13030
rect 1524 13028 1580 13030
rect 1604 13028 1660 13030
rect 1684 13028 1740 13030
rect 1364 11994 1420 11996
rect 1444 11994 1500 11996
rect 1524 11994 1580 11996
rect 1604 11994 1660 11996
rect 1684 11994 1740 11996
rect 1364 11942 1366 11994
rect 1366 11942 1418 11994
rect 1418 11942 1420 11994
rect 1444 11942 1482 11994
rect 1482 11942 1494 11994
rect 1494 11942 1500 11994
rect 1524 11942 1546 11994
rect 1546 11942 1558 11994
rect 1558 11942 1580 11994
rect 1604 11942 1610 11994
rect 1610 11942 1622 11994
rect 1622 11942 1660 11994
rect 1684 11942 1686 11994
rect 1686 11942 1738 11994
rect 1738 11942 1740 11994
rect 1364 11940 1420 11942
rect 1444 11940 1500 11942
rect 1524 11940 1580 11942
rect 1604 11940 1660 11942
rect 1684 11940 1740 11942
rect 2686 14320 2742 14376
rect 1364 10906 1420 10908
rect 1444 10906 1500 10908
rect 1524 10906 1580 10908
rect 1604 10906 1660 10908
rect 1684 10906 1740 10908
rect 1364 10854 1366 10906
rect 1366 10854 1418 10906
rect 1418 10854 1420 10906
rect 1444 10854 1482 10906
rect 1482 10854 1494 10906
rect 1494 10854 1500 10906
rect 1524 10854 1546 10906
rect 1546 10854 1558 10906
rect 1558 10854 1580 10906
rect 1604 10854 1610 10906
rect 1610 10854 1622 10906
rect 1622 10854 1660 10906
rect 1684 10854 1686 10906
rect 1686 10854 1738 10906
rect 1738 10854 1740 10906
rect 1364 10852 1420 10854
rect 1444 10852 1500 10854
rect 1524 10852 1580 10854
rect 1604 10852 1660 10854
rect 1684 10852 1740 10854
rect 1364 9818 1420 9820
rect 1444 9818 1500 9820
rect 1524 9818 1580 9820
rect 1604 9818 1660 9820
rect 1684 9818 1740 9820
rect 1364 9766 1366 9818
rect 1366 9766 1418 9818
rect 1418 9766 1420 9818
rect 1444 9766 1482 9818
rect 1482 9766 1494 9818
rect 1494 9766 1500 9818
rect 1524 9766 1546 9818
rect 1546 9766 1558 9818
rect 1558 9766 1580 9818
rect 1604 9766 1610 9818
rect 1610 9766 1622 9818
rect 1622 9766 1660 9818
rect 1684 9766 1686 9818
rect 1686 9766 1738 9818
rect 1738 9766 1740 9818
rect 1364 9764 1420 9766
rect 1444 9764 1500 9766
rect 1524 9764 1580 9766
rect 1604 9764 1660 9766
rect 1684 9764 1740 9766
rect 1858 8880 1914 8936
rect 1364 8730 1420 8732
rect 1444 8730 1500 8732
rect 1524 8730 1580 8732
rect 1604 8730 1660 8732
rect 1684 8730 1740 8732
rect 1364 8678 1366 8730
rect 1366 8678 1418 8730
rect 1418 8678 1420 8730
rect 1444 8678 1482 8730
rect 1482 8678 1494 8730
rect 1494 8678 1500 8730
rect 1524 8678 1546 8730
rect 1546 8678 1558 8730
rect 1558 8678 1580 8730
rect 1604 8678 1610 8730
rect 1610 8678 1622 8730
rect 1622 8678 1660 8730
rect 1684 8678 1686 8730
rect 1686 8678 1738 8730
rect 1738 8678 1740 8730
rect 1364 8676 1420 8678
rect 1444 8676 1500 8678
rect 1524 8676 1580 8678
rect 1604 8676 1660 8678
rect 1684 8676 1740 8678
rect 1364 7642 1420 7644
rect 1444 7642 1500 7644
rect 1524 7642 1580 7644
rect 1604 7642 1660 7644
rect 1684 7642 1740 7644
rect 1364 7590 1366 7642
rect 1366 7590 1418 7642
rect 1418 7590 1420 7642
rect 1444 7590 1482 7642
rect 1482 7590 1494 7642
rect 1494 7590 1500 7642
rect 1524 7590 1546 7642
rect 1546 7590 1558 7642
rect 1558 7590 1580 7642
rect 1604 7590 1610 7642
rect 1610 7590 1622 7642
rect 1622 7590 1660 7642
rect 1684 7590 1686 7642
rect 1686 7590 1738 7642
rect 1738 7590 1740 7642
rect 1364 7588 1420 7590
rect 1444 7588 1500 7590
rect 1524 7588 1580 7590
rect 1604 7588 1660 7590
rect 1684 7588 1740 7590
rect 1364 6554 1420 6556
rect 1444 6554 1500 6556
rect 1524 6554 1580 6556
rect 1604 6554 1660 6556
rect 1684 6554 1740 6556
rect 1364 6502 1366 6554
rect 1366 6502 1418 6554
rect 1418 6502 1420 6554
rect 1444 6502 1482 6554
rect 1482 6502 1494 6554
rect 1494 6502 1500 6554
rect 1524 6502 1546 6554
rect 1546 6502 1558 6554
rect 1558 6502 1580 6554
rect 1604 6502 1610 6554
rect 1610 6502 1622 6554
rect 1622 6502 1660 6554
rect 1684 6502 1686 6554
rect 1686 6502 1738 6554
rect 1738 6502 1740 6554
rect 1364 6500 1420 6502
rect 1444 6500 1500 6502
rect 1524 6500 1580 6502
rect 1604 6500 1660 6502
rect 1684 6500 1740 6502
rect 1364 5466 1420 5468
rect 1444 5466 1500 5468
rect 1524 5466 1580 5468
rect 1604 5466 1660 5468
rect 1684 5466 1740 5468
rect 1364 5414 1366 5466
rect 1366 5414 1418 5466
rect 1418 5414 1420 5466
rect 1444 5414 1482 5466
rect 1482 5414 1494 5466
rect 1494 5414 1500 5466
rect 1524 5414 1546 5466
rect 1546 5414 1558 5466
rect 1558 5414 1580 5466
rect 1604 5414 1610 5466
rect 1610 5414 1622 5466
rect 1622 5414 1660 5466
rect 1684 5414 1686 5466
rect 1686 5414 1738 5466
rect 1738 5414 1740 5466
rect 1364 5412 1420 5414
rect 1444 5412 1500 5414
rect 1524 5412 1580 5414
rect 1604 5412 1660 5414
rect 1684 5412 1740 5414
rect 1364 4378 1420 4380
rect 1444 4378 1500 4380
rect 1524 4378 1580 4380
rect 1604 4378 1660 4380
rect 1684 4378 1740 4380
rect 1364 4326 1366 4378
rect 1366 4326 1418 4378
rect 1418 4326 1420 4378
rect 1444 4326 1482 4378
rect 1482 4326 1494 4378
rect 1494 4326 1500 4378
rect 1524 4326 1546 4378
rect 1546 4326 1558 4378
rect 1558 4326 1580 4378
rect 1604 4326 1610 4378
rect 1610 4326 1622 4378
rect 1622 4326 1660 4378
rect 1684 4326 1686 4378
rect 1686 4326 1738 4378
rect 1738 4326 1740 4378
rect 1364 4324 1420 4326
rect 1444 4324 1500 4326
rect 1524 4324 1580 4326
rect 1604 4324 1660 4326
rect 1684 4324 1740 4326
rect 1364 3290 1420 3292
rect 1444 3290 1500 3292
rect 1524 3290 1580 3292
rect 1604 3290 1660 3292
rect 1684 3290 1740 3292
rect 1364 3238 1366 3290
rect 1366 3238 1418 3290
rect 1418 3238 1420 3290
rect 1444 3238 1482 3290
rect 1482 3238 1494 3290
rect 1494 3238 1500 3290
rect 1524 3238 1546 3290
rect 1546 3238 1558 3290
rect 1558 3238 1580 3290
rect 1604 3238 1610 3290
rect 1610 3238 1622 3290
rect 1622 3238 1660 3290
rect 1684 3238 1686 3290
rect 1686 3238 1738 3290
rect 1738 3238 1740 3290
rect 1364 3236 1420 3238
rect 1444 3236 1500 3238
rect 1524 3236 1580 3238
rect 1604 3236 1660 3238
rect 1684 3236 1740 3238
rect 1306 2488 1362 2544
rect 1364 2202 1420 2204
rect 1444 2202 1500 2204
rect 1524 2202 1580 2204
rect 1604 2202 1660 2204
rect 1684 2202 1740 2204
rect 1364 2150 1366 2202
rect 1366 2150 1418 2202
rect 1418 2150 1420 2202
rect 1444 2150 1482 2202
rect 1482 2150 1494 2202
rect 1494 2150 1500 2202
rect 1524 2150 1546 2202
rect 1546 2150 1558 2202
rect 1558 2150 1580 2202
rect 1604 2150 1610 2202
rect 1610 2150 1622 2202
rect 1622 2150 1660 2202
rect 1684 2150 1686 2202
rect 1686 2150 1738 2202
rect 1738 2150 1740 2202
rect 1364 2148 1420 2150
rect 1444 2148 1500 2150
rect 1524 2148 1580 2150
rect 1604 2148 1660 2150
rect 1684 2148 1740 2150
rect 2686 12688 2742 12744
rect 3238 15700 3294 15736
rect 3238 15680 3240 15700
rect 3240 15680 3292 15700
rect 3292 15680 3294 15700
rect 2870 12824 2926 12880
rect 2134 7792 2190 7848
rect 2594 9036 2650 9072
rect 2594 9016 2596 9036
rect 2596 9016 2648 9036
rect 2648 9016 2650 9036
rect 3514 13912 3570 13968
rect 4364 15802 4420 15804
rect 4444 15802 4500 15804
rect 4524 15802 4580 15804
rect 4604 15802 4660 15804
rect 4684 15802 4740 15804
rect 4364 15750 4366 15802
rect 4366 15750 4418 15802
rect 4418 15750 4420 15802
rect 4444 15750 4482 15802
rect 4482 15750 4494 15802
rect 4494 15750 4500 15802
rect 4524 15750 4546 15802
rect 4546 15750 4558 15802
rect 4558 15750 4580 15802
rect 4604 15750 4610 15802
rect 4610 15750 4622 15802
rect 4622 15750 4660 15802
rect 4684 15750 4686 15802
rect 4686 15750 4738 15802
rect 4738 15750 4740 15802
rect 4364 15748 4420 15750
rect 4444 15748 4500 15750
rect 4524 15748 4580 15750
rect 4604 15748 4660 15750
rect 4684 15748 4740 15750
rect 4066 14456 4122 14512
rect 4364 14714 4420 14716
rect 4444 14714 4500 14716
rect 4524 14714 4580 14716
rect 4604 14714 4660 14716
rect 4684 14714 4740 14716
rect 4364 14662 4366 14714
rect 4366 14662 4418 14714
rect 4418 14662 4420 14714
rect 4444 14662 4482 14714
rect 4482 14662 4494 14714
rect 4494 14662 4500 14714
rect 4524 14662 4546 14714
rect 4546 14662 4558 14714
rect 4558 14662 4580 14714
rect 4604 14662 4610 14714
rect 4610 14662 4622 14714
rect 4622 14662 4660 14714
rect 4684 14662 4686 14714
rect 4686 14662 4738 14714
rect 4738 14662 4740 14714
rect 4364 14660 4420 14662
rect 4444 14660 4500 14662
rect 4524 14660 4580 14662
rect 4604 14660 4660 14662
rect 4684 14660 4740 14662
rect 4526 14492 4528 14512
rect 4528 14492 4580 14512
rect 4580 14492 4582 14512
rect 4526 14456 4582 14492
rect 4618 14048 4674 14104
rect 4342 13932 4398 13968
rect 4342 13912 4344 13932
rect 4344 13912 4396 13932
rect 4396 13912 4398 13932
rect 4894 14864 4950 14920
rect 5078 15000 5134 15056
rect 4066 13368 4122 13424
rect 4364 13626 4420 13628
rect 4444 13626 4500 13628
rect 4524 13626 4580 13628
rect 4604 13626 4660 13628
rect 4684 13626 4740 13628
rect 4364 13574 4366 13626
rect 4366 13574 4418 13626
rect 4418 13574 4420 13626
rect 4444 13574 4482 13626
rect 4482 13574 4494 13626
rect 4494 13574 4500 13626
rect 4524 13574 4546 13626
rect 4546 13574 4558 13626
rect 4558 13574 4580 13626
rect 4604 13574 4610 13626
rect 4610 13574 4622 13626
rect 4622 13574 4660 13626
rect 4684 13574 4686 13626
rect 4686 13574 4738 13626
rect 4738 13574 4740 13626
rect 4364 13572 4420 13574
rect 4444 13572 4500 13574
rect 4524 13572 4580 13574
rect 4604 13572 4660 13574
rect 4684 13572 4740 13574
rect 2870 7248 2926 7304
rect 2594 4972 2596 4992
rect 2596 4972 2648 4992
rect 2648 4972 2650 4992
rect 2594 4936 2650 4972
rect 5262 13812 5264 13832
rect 5264 13812 5316 13832
rect 5316 13812 5318 13832
rect 5262 13776 5318 13812
rect 4364 12538 4420 12540
rect 4444 12538 4500 12540
rect 4524 12538 4580 12540
rect 4604 12538 4660 12540
rect 4684 12538 4740 12540
rect 4364 12486 4366 12538
rect 4366 12486 4418 12538
rect 4418 12486 4420 12538
rect 4444 12486 4482 12538
rect 4482 12486 4494 12538
rect 4494 12486 4500 12538
rect 4524 12486 4546 12538
rect 4546 12486 4558 12538
rect 4558 12486 4580 12538
rect 4604 12486 4610 12538
rect 4610 12486 4622 12538
rect 4622 12486 4660 12538
rect 4684 12486 4686 12538
rect 4686 12486 4738 12538
rect 4738 12486 4740 12538
rect 4364 12484 4420 12486
rect 4444 12484 4500 12486
rect 4524 12484 4580 12486
rect 4604 12484 4660 12486
rect 4684 12484 4740 12486
rect 3882 10920 3938 10976
rect 4066 10784 4122 10840
rect 4364 11450 4420 11452
rect 4444 11450 4500 11452
rect 4524 11450 4580 11452
rect 4604 11450 4660 11452
rect 4684 11450 4740 11452
rect 4364 11398 4366 11450
rect 4366 11398 4418 11450
rect 4418 11398 4420 11450
rect 4444 11398 4482 11450
rect 4482 11398 4494 11450
rect 4494 11398 4500 11450
rect 4524 11398 4546 11450
rect 4546 11398 4558 11450
rect 4558 11398 4580 11450
rect 4604 11398 4610 11450
rect 4610 11398 4622 11450
rect 4622 11398 4660 11450
rect 4684 11398 4686 11450
rect 4686 11398 4738 11450
rect 4738 11398 4740 11450
rect 4364 11396 4420 11398
rect 4444 11396 4500 11398
rect 4524 11396 4580 11398
rect 4604 11396 4660 11398
rect 4684 11396 4740 11398
rect 4618 10548 4620 10568
rect 4620 10548 4672 10568
rect 4672 10548 4674 10568
rect 4618 10512 4674 10548
rect 3790 9968 3846 10024
rect 4364 10362 4420 10364
rect 4444 10362 4500 10364
rect 4524 10362 4580 10364
rect 4604 10362 4660 10364
rect 4684 10362 4740 10364
rect 4364 10310 4366 10362
rect 4366 10310 4418 10362
rect 4418 10310 4420 10362
rect 4444 10310 4482 10362
rect 4482 10310 4494 10362
rect 4494 10310 4500 10362
rect 4524 10310 4546 10362
rect 4546 10310 4558 10362
rect 4558 10310 4580 10362
rect 4604 10310 4610 10362
rect 4610 10310 4622 10362
rect 4622 10310 4660 10362
rect 4684 10310 4686 10362
rect 4686 10310 4738 10362
rect 4738 10310 4740 10362
rect 4364 10308 4420 10310
rect 4444 10308 4500 10310
rect 4524 10308 4580 10310
rect 4604 10308 4660 10310
rect 4684 10308 4740 10310
rect 4342 10104 4398 10160
rect 3698 9832 3754 9888
rect 3514 9580 3570 9616
rect 4618 9968 4674 10024
rect 5078 11056 5134 11112
rect 6458 16496 6514 16552
rect 6274 15000 6330 15056
rect 6366 14884 6422 14920
rect 6366 14864 6368 14884
rect 6368 14864 6420 14884
rect 6420 14864 6422 14884
rect 6182 13912 6238 13968
rect 5998 13676 6000 13696
rect 6000 13676 6052 13696
rect 6052 13676 6054 13696
rect 5998 13640 6054 13676
rect 6550 15408 6606 15464
rect 6366 13504 6422 13560
rect 6090 13388 6146 13424
rect 6090 13368 6092 13388
rect 6092 13368 6144 13388
rect 6144 13368 6146 13388
rect 6366 12688 6422 12744
rect 6274 12416 6330 12472
rect 6918 13232 6974 13288
rect 7364 17434 7420 17436
rect 7444 17434 7500 17436
rect 7524 17434 7580 17436
rect 7604 17434 7660 17436
rect 7684 17434 7740 17436
rect 7364 17382 7366 17434
rect 7366 17382 7418 17434
rect 7418 17382 7420 17434
rect 7444 17382 7482 17434
rect 7482 17382 7494 17434
rect 7494 17382 7500 17434
rect 7524 17382 7546 17434
rect 7546 17382 7558 17434
rect 7558 17382 7580 17434
rect 7604 17382 7610 17434
rect 7610 17382 7622 17434
rect 7622 17382 7660 17434
rect 7684 17382 7686 17434
rect 7686 17382 7738 17434
rect 7738 17382 7740 17434
rect 7364 17380 7420 17382
rect 7444 17380 7500 17382
rect 7524 17380 7580 17382
rect 7604 17380 7660 17382
rect 7684 17380 7740 17382
rect 7378 16516 7434 16552
rect 7378 16496 7380 16516
rect 7380 16496 7432 16516
rect 7432 16496 7434 16516
rect 7364 16346 7420 16348
rect 7444 16346 7500 16348
rect 7524 16346 7580 16348
rect 7604 16346 7660 16348
rect 7684 16346 7740 16348
rect 7364 16294 7366 16346
rect 7366 16294 7418 16346
rect 7418 16294 7420 16346
rect 7444 16294 7482 16346
rect 7482 16294 7494 16346
rect 7494 16294 7500 16346
rect 7524 16294 7546 16346
rect 7546 16294 7558 16346
rect 7558 16294 7580 16346
rect 7604 16294 7610 16346
rect 7610 16294 7622 16346
rect 7622 16294 7660 16346
rect 7684 16294 7686 16346
rect 7686 16294 7738 16346
rect 7738 16294 7740 16346
rect 7364 16292 7420 16294
rect 7444 16292 7500 16294
rect 7524 16292 7580 16294
rect 7604 16292 7660 16294
rect 7684 16292 7740 16294
rect 9034 16632 9090 16688
rect 10364 16890 10420 16892
rect 10444 16890 10500 16892
rect 10524 16890 10580 16892
rect 10604 16890 10660 16892
rect 10684 16890 10740 16892
rect 10364 16838 10366 16890
rect 10366 16838 10418 16890
rect 10418 16838 10420 16890
rect 10444 16838 10482 16890
rect 10482 16838 10494 16890
rect 10494 16838 10500 16890
rect 10524 16838 10546 16890
rect 10546 16838 10558 16890
rect 10558 16838 10580 16890
rect 10604 16838 10610 16890
rect 10610 16838 10622 16890
rect 10622 16838 10660 16890
rect 10684 16838 10686 16890
rect 10686 16838 10738 16890
rect 10738 16838 10740 16890
rect 10364 16836 10420 16838
rect 10444 16836 10500 16838
rect 10524 16836 10580 16838
rect 10604 16836 10660 16838
rect 10684 16836 10740 16838
rect 7102 15272 7158 15328
rect 7102 15000 7158 15056
rect 5814 11212 5870 11248
rect 5814 11192 5816 11212
rect 5816 11192 5868 11212
rect 5868 11192 5870 11212
rect 4526 9832 4582 9888
rect 3514 9560 3516 9580
rect 3516 9560 3568 9580
rect 3568 9560 3570 9580
rect 4364 9274 4420 9276
rect 4444 9274 4500 9276
rect 4524 9274 4580 9276
rect 4604 9274 4660 9276
rect 4684 9274 4740 9276
rect 4364 9222 4366 9274
rect 4366 9222 4418 9274
rect 4418 9222 4420 9274
rect 4444 9222 4482 9274
rect 4482 9222 4494 9274
rect 4494 9222 4500 9274
rect 4524 9222 4546 9274
rect 4546 9222 4558 9274
rect 4558 9222 4580 9274
rect 4604 9222 4610 9274
rect 4610 9222 4622 9274
rect 4622 9222 4660 9274
rect 4684 9222 4686 9274
rect 4686 9222 4738 9274
rect 4738 9222 4740 9274
rect 4364 9220 4420 9222
rect 4444 9220 4500 9222
rect 4524 9220 4580 9222
rect 4604 9220 4660 9222
rect 4684 9220 4740 9222
rect 5262 10668 5318 10704
rect 5262 10648 5264 10668
rect 5264 10648 5316 10668
rect 5316 10648 5318 10668
rect 5538 10956 5540 10976
rect 5540 10956 5592 10976
rect 5592 10956 5594 10976
rect 5538 10920 5594 10956
rect 4364 8186 4420 8188
rect 4444 8186 4500 8188
rect 4524 8186 4580 8188
rect 4604 8186 4660 8188
rect 4684 8186 4740 8188
rect 4364 8134 4366 8186
rect 4366 8134 4418 8186
rect 4418 8134 4420 8186
rect 4444 8134 4482 8186
rect 4482 8134 4494 8186
rect 4494 8134 4500 8186
rect 4524 8134 4546 8186
rect 4546 8134 4558 8186
rect 4558 8134 4580 8186
rect 4604 8134 4610 8186
rect 4610 8134 4622 8186
rect 4622 8134 4660 8186
rect 4684 8134 4686 8186
rect 4686 8134 4738 8186
rect 4738 8134 4740 8186
rect 4364 8132 4420 8134
rect 4444 8132 4500 8134
rect 4524 8132 4580 8134
rect 4604 8132 4660 8134
rect 4684 8132 4740 8134
rect 1766 1808 1822 1864
rect 1364 1114 1420 1116
rect 1444 1114 1500 1116
rect 1524 1114 1580 1116
rect 1604 1114 1660 1116
rect 1684 1114 1740 1116
rect 1364 1062 1366 1114
rect 1366 1062 1418 1114
rect 1418 1062 1420 1114
rect 1444 1062 1482 1114
rect 1482 1062 1494 1114
rect 1494 1062 1500 1114
rect 1524 1062 1546 1114
rect 1546 1062 1558 1114
rect 1558 1062 1580 1114
rect 1604 1062 1610 1114
rect 1610 1062 1622 1114
rect 1622 1062 1660 1114
rect 1684 1062 1686 1114
rect 1686 1062 1738 1114
rect 1738 1062 1740 1114
rect 1364 1060 1420 1062
rect 1444 1060 1500 1062
rect 1524 1060 1580 1062
rect 1604 1060 1660 1062
rect 1684 1060 1740 1062
rect 4364 7098 4420 7100
rect 4444 7098 4500 7100
rect 4524 7098 4580 7100
rect 4604 7098 4660 7100
rect 4684 7098 4740 7100
rect 4364 7046 4366 7098
rect 4366 7046 4418 7098
rect 4418 7046 4420 7098
rect 4444 7046 4482 7098
rect 4482 7046 4494 7098
rect 4494 7046 4500 7098
rect 4524 7046 4546 7098
rect 4546 7046 4558 7098
rect 4558 7046 4580 7098
rect 4604 7046 4610 7098
rect 4610 7046 4622 7098
rect 4622 7046 4660 7098
rect 4684 7046 4686 7098
rect 4686 7046 4738 7098
rect 4738 7046 4740 7098
rect 4364 7044 4420 7046
rect 4444 7044 4500 7046
rect 4524 7044 4580 7046
rect 4604 7044 4660 7046
rect 4684 7044 4740 7046
rect 4158 4972 4160 4992
rect 4160 4972 4212 4992
rect 4212 4972 4214 4992
rect 4158 4936 4214 4972
rect 4364 6010 4420 6012
rect 4444 6010 4500 6012
rect 4524 6010 4580 6012
rect 4604 6010 4660 6012
rect 4684 6010 4740 6012
rect 4364 5958 4366 6010
rect 4366 5958 4418 6010
rect 4418 5958 4420 6010
rect 4444 5958 4482 6010
rect 4482 5958 4494 6010
rect 4494 5958 4500 6010
rect 4524 5958 4546 6010
rect 4546 5958 4558 6010
rect 4558 5958 4580 6010
rect 4604 5958 4610 6010
rect 4610 5958 4622 6010
rect 4622 5958 4660 6010
rect 4684 5958 4686 6010
rect 4686 5958 4738 6010
rect 4738 5958 4740 6010
rect 4364 5956 4420 5958
rect 4444 5956 4500 5958
rect 4524 5956 4580 5958
rect 4604 5956 4660 5958
rect 4684 5956 4740 5958
rect 4364 4922 4420 4924
rect 4444 4922 4500 4924
rect 4524 4922 4580 4924
rect 4604 4922 4660 4924
rect 4684 4922 4740 4924
rect 4364 4870 4366 4922
rect 4366 4870 4418 4922
rect 4418 4870 4420 4922
rect 4444 4870 4482 4922
rect 4482 4870 4494 4922
rect 4494 4870 4500 4922
rect 4524 4870 4546 4922
rect 4546 4870 4558 4922
rect 4558 4870 4580 4922
rect 4604 4870 4610 4922
rect 4610 4870 4622 4922
rect 4622 4870 4660 4922
rect 4684 4870 4686 4922
rect 4686 4870 4738 4922
rect 4738 4870 4740 4922
rect 4364 4868 4420 4870
rect 4444 4868 4500 4870
rect 4524 4868 4580 4870
rect 4604 4868 4660 4870
rect 4684 4868 4740 4870
rect 4364 3834 4420 3836
rect 4444 3834 4500 3836
rect 4524 3834 4580 3836
rect 4604 3834 4660 3836
rect 4684 3834 4740 3836
rect 4364 3782 4366 3834
rect 4366 3782 4418 3834
rect 4418 3782 4420 3834
rect 4444 3782 4482 3834
rect 4482 3782 4494 3834
rect 4494 3782 4500 3834
rect 4524 3782 4546 3834
rect 4546 3782 4558 3834
rect 4558 3782 4580 3834
rect 4604 3782 4610 3834
rect 4610 3782 4622 3834
rect 4622 3782 4660 3834
rect 4684 3782 4686 3834
rect 4686 3782 4738 3834
rect 4738 3782 4740 3834
rect 4364 3780 4420 3782
rect 4444 3780 4500 3782
rect 4524 3780 4580 3782
rect 4604 3780 4660 3782
rect 4684 3780 4740 3782
rect 4434 3304 4490 3360
rect 4986 5072 5042 5128
rect 4894 4528 4950 4584
rect 4894 3984 4950 4040
rect 3514 2488 3570 2544
rect 4364 2746 4420 2748
rect 4444 2746 4500 2748
rect 4524 2746 4580 2748
rect 4604 2746 4660 2748
rect 4684 2746 4740 2748
rect 4364 2694 4366 2746
rect 4366 2694 4418 2746
rect 4418 2694 4420 2746
rect 4444 2694 4482 2746
rect 4482 2694 4494 2746
rect 4494 2694 4500 2746
rect 4524 2694 4546 2746
rect 4546 2694 4558 2746
rect 4558 2694 4580 2746
rect 4604 2694 4610 2746
rect 4610 2694 4622 2746
rect 4622 2694 4660 2746
rect 4684 2694 4686 2746
rect 4686 2694 4738 2746
rect 4738 2694 4740 2746
rect 4364 2692 4420 2694
rect 4444 2692 4500 2694
rect 4524 2692 4580 2694
rect 4604 2692 4660 2694
rect 4684 2692 4740 2694
rect 4066 1420 4122 1456
rect 4364 1658 4420 1660
rect 4444 1658 4500 1660
rect 4524 1658 4580 1660
rect 4604 1658 4660 1660
rect 4684 1658 4740 1660
rect 4364 1606 4366 1658
rect 4366 1606 4418 1658
rect 4418 1606 4420 1658
rect 4444 1606 4482 1658
rect 4482 1606 4494 1658
rect 4494 1606 4500 1658
rect 4524 1606 4546 1658
rect 4546 1606 4558 1658
rect 4558 1606 4580 1658
rect 4604 1606 4610 1658
rect 4610 1606 4622 1658
rect 4622 1606 4660 1658
rect 4684 1606 4686 1658
rect 4686 1606 4738 1658
rect 4738 1606 4740 1658
rect 4364 1604 4420 1606
rect 4444 1604 4500 1606
rect 4524 1604 4580 1606
rect 4604 1604 4660 1606
rect 4684 1604 4740 1606
rect 5906 8372 5908 8392
rect 5908 8372 5960 8392
rect 5960 8372 5962 8392
rect 5906 8336 5962 8372
rect 6090 11464 6146 11520
rect 7364 15258 7420 15260
rect 7444 15258 7500 15260
rect 7524 15258 7580 15260
rect 7604 15258 7660 15260
rect 7684 15258 7740 15260
rect 7364 15206 7366 15258
rect 7366 15206 7418 15258
rect 7418 15206 7420 15258
rect 7444 15206 7482 15258
rect 7482 15206 7494 15258
rect 7494 15206 7500 15258
rect 7524 15206 7546 15258
rect 7546 15206 7558 15258
rect 7558 15206 7580 15258
rect 7604 15206 7610 15258
rect 7610 15206 7622 15258
rect 7622 15206 7660 15258
rect 7684 15206 7686 15258
rect 7686 15206 7738 15258
rect 7738 15206 7740 15258
rect 7364 15204 7420 15206
rect 7444 15204 7500 15206
rect 7524 15204 7580 15206
rect 7604 15204 7660 15206
rect 7684 15204 7740 15206
rect 7746 14900 7748 14920
rect 7748 14900 7800 14920
rect 7800 14900 7802 14920
rect 7746 14864 7802 14900
rect 7286 14320 7342 14376
rect 7364 14170 7420 14172
rect 7444 14170 7500 14172
rect 7524 14170 7580 14172
rect 7604 14170 7660 14172
rect 7684 14170 7740 14172
rect 7364 14118 7366 14170
rect 7366 14118 7418 14170
rect 7418 14118 7420 14170
rect 7444 14118 7482 14170
rect 7482 14118 7494 14170
rect 7494 14118 7500 14170
rect 7524 14118 7546 14170
rect 7546 14118 7558 14170
rect 7558 14118 7580 14170
rect 7604 14118 7610 14170
rect 7610 14118 7622 14170
rect 7622 14118 7660 14170
rect 7684 14118 7686 14170
rect 7686 14118 7738 14170
rect 7738 14118 7740 14170
rect 7364 14116 7420 14118
rect 7444 14116 7500 14118
rect 7524 14116 7580 14118
rect 7604 14116 7660 14118
rect 7684 14116 7740 14118
rect 7838 14048 7894 14104
rect 7470 13912 7526 13968
rect 7654 13912 7710 13968
rect 7364 13082 7420 13084
rect 7444 13082 7500 13084
rect 7524 13082 7580 13084
rect 7604 13082 7660 13084
rect 7684 13082 7740 13084
rect 7364 13030 7366 13082
rect 7366 13030 7418 13082
rect 7418 13030 7420 13082
rect 7444 13030 7482 13082
rect 7482 13030 7494 13082
rect 7494 13030 7500 13082
rect 7524 13030 7546 13082
rect 7546 13030 7558 13082
rect 7558 13030 7580 13082
rect 7604 13030 7610 13082
rect 7610 13030 7622 13082
rect 7622 13030 7660 13082
rect 7684 13030 7686 13082
rect 7686 13030 7738 13082
rect 7738 13030 7740 13082
rect 7364 13028 7420 13030
rect 7444 13028 7500 13030
rect 7524 13028 7580 13030
rect 7604 13028 7660 13030
rect 7684 13028 7740 13030
rect 8390 14864 8446 14920
rect 8390 14184 8446 14240
rect 6918 11736 6974 11792
rect 7930 12552 7986 12608
rect 7930 12436 7986 12472
rect 7930 12416 7932 12436
rect 7932 12416 7984 12436
rect 7984 12416 7986 12436
rect 6366 10668 6422 10704
rect 6366 10648 6368 10668
rect 6368 10648 6420 10668
rect 6420 10648 6422 10668
rect 6182 10376 6238 10432
rect 6734 11056 6790 11112
rect 7010 10804 7066 10840
rect 7010 10784 7012 10804
rect 7012 10784 7064 10804
rect 7064 10784 7066 10804
rect 6826 9968 6882 10024
rect 5170 3032 5226 3088
rect 5814 4564 5816 4584
rect 5816 4564 5868 4584
rect 5868 4564 5870 4584
rect 5814 4528 5870 4564
rect 5630 3848 5686 3904
rect 6458 8880 6514 8936
rect 7364 11994 7420 11996
rect 7444 11994 7500 11996
rect 7524 11994 7580 11996
rect 7604 11994 7660 11996
rect 7684 11994 7740 11996
rect 7364 11942 7366 11994
rect 7366 11942 7418 11994
rect 7418 11942 7420 11994
rect 7444 11942 7482 11994
rect 7482 11942 7494 11994
rect 7494 11942 7500 11994
rect 7524 11942 7546 11994
rect 7546 11942 7558 11994
rect 7558 11942 7580 11994
rect 7604 11942 7610 11994
rect 7610 11942 7622 11994
rect 7622 11942 7660 11994
rect 7684 11942 7686 11994
rect 7686 11942 7738 11994
rect 7738 11942 7740 11994
rect 7364 11940 7420 11942
rect 7444 11940 7500 11942
rect 7524 11940 7580 11942
rect 7604 11940 7660 11942
rect 7684 11940 7740 11942
rect 7286 11736 7342 11792
rect 7654 11736 7710 11792
rect 8022 11212 8078 11248
rect 8022 11192 8024 11212
rect 8024 11192 8076 11212
rect 8076 11192 8078 11212
rect 7364 10906 7420 10908
rect 7444 10906 7500 10908
rect 7524 10906 7580 10908
rect 7604 10906 7660 10908
rect 7684 10906 7740 10908
rect 7364 10854 7366 10906
rect 7366 10854 7418 10906
rect 7418 10854 7420 10906
rect 7444 10854 7482 10906
rect 7482 10854 7494 10906
rect 7494 10854 7500 10906
rect 7524 10854 7546 10906
rect 7546 10854 7558 10906
rect 7558 10854 7580 10906
rect 7604 10854 7610 10906
rect 7610 10854 7622 10906
rect 7622 10854 7660 10906
rect 7684 10854 7686 10906
rect 7686 10854 7738 10906
rect 7738 10854 7740 10906
rect 7364 10852 7420 10854
rect 7444 10852 7500 10854
rect 7524 10852 7580 10854
rect 7604 10852 7660 10854
rect 7684 10852 7740 10854
rect 8114 10920 8170 10976
rect 6734 8492 6790 8528
rect 7654 9968 7710 10024
rect 6734 8472 6736 8492
rect 6736 8472 6788 8492
rect 6788 8472 6790 8492
rect 7364 9818 7420 9820
rect 7444 9818 7500 9820
rect 7524 9818 7580 9820
rect 7604 9818 7660 9820
rect 7684 9818 7740 9820
rect 7364 9766 7366 9818
rect 7366 9766 7418 9818
rect 7418 9766 7420 9818
rect 7444 9766 7482 9818
rect 7482 9766 7494 9818
rect 7494 9766 7500 9818
rect 7524 9766 7546 9818
rect 7546 9766 7558 9818
rect 7558 9766 7580 9818
rect 7604 9766 7610 9818
rect 7610 9766 7622 9818
rect 7622 9766 7660 9818
rect 7684 9766 7686 9818
rect 7686 9766 7738 9818
rect 7738 9766 7740 9818
rect 7364 9764 7420 9766
rect 7444 9764 7500 9766
rect 7524 9764 7580 9766
rect 7604 9764 7660 9766
rect 7684 9764 7740 9766
rect 7364 8730 7420 8732
rect 7444 8730 7500 8732
rect 7524 8730 7580 8732
rect 7604 8730 7660 8732
rect 7684 8730 7740 8732
rect 7364 8678 7366 8730
rect 7366 8678 7418 8730
rect 7418 8678 7420 8730
rect 7444 8678 7482 8730
rect 7482 8678 7494 8730
rect 7494 8678 7500 8730
rect 7524 8678 7546 8730
rect 7546 8678 7558 8730
rect 7558 8678 7580 8730
rect 7604 8678 7610 8730
rect 7610 8678 7622 8730
rect 7622 8678 7660 8730
rect 7684 8678 7686 8730
rect 7686 8678 7738 8730
rect 7738 8678 7740 8730
rect 7364 8676 7420 8678
rect 7444 8676 7500 8678
rect 7524 8676 7580 8678
rect 7604 8676 7660 8678
rect 7684 8676 7740 8678
rect 7378 8492 7434 8528
rect 7378 8472 7380 8492
rect 7380 8472 7432 8492
rect 7432 8472 7434 8492
rect 7470 8372 7472 8392
rect 7472 8372 7524 8392
rect 7524 8372 7526 8392
rect 7470 8336 7526 8372
rect 7364 7642 7420 7644
rect 7444 7642 7500 7644
rect 7524 7642 7580 7644
rect 7604 7642 7660 7644
rect 7684 7642 7740 7644
rect 7364 7590 7366 7642
rect 7366 7590 7418 7642
rect 7418 7590 7420 7642
rect 7444 7590 7482 7642
rect 7482 7590 7494 7642
rect 7494 7590 7500 7642
rect 7524 7590 7546 7642
rect 7546 7590 7558 7642
rect 7558 7590 7580 7642
rect 7604 7590 7610 7642
rect 7610 7590 7622 7642
rect 7622 7590 7660 7642
rect 7684 7590 7686 7642
rect 7686 7590 7738 7642
rect 7738 7590 7740 7642
rect 7364 7588 7420 7590
rect 7444 7588 7500 7590
rect 7524 7588 7580 7590
rect 7604 7588 7660 7590
rect 7684 7588 7740 7590
rect 7470 7248 7526 7304
rect 5814 2644 5870 2680
rect 5814 2624 5816 2644
rect 5816 2624 5868 2644
rect 5868 2624 5870 2644
rect 4986 1844 4988 1864
rect 4988 1844 5040 1864
rect 5040 1844 5042 1864
rect 4986 1808 5042 1844
rect 4066 1400 4068 1420
rect 4068 1400 4120 1420
rect 4120 1400 4122 1420
rect 4802 1420 4858 1456
rect 6090 2352 6146 2408
rect 6550 4156 6552 4176
rect 6552 4156 6604 4176
rect 6604 4156 6606 4176
rect 6550 4120 6606 4156
rect 6366 1536 6422 1592
rect 4802 1400 4804 1420
rect 4804 1400 4856 1420
rect 4856 1400 4858 1420
rect 7010 4664 7066 4720
rect 7746 6740 7748 6760
rect 7748 6740 7800 6760
rect 7800 6740 7802 6760
rect 7746 6704 7802 6740
rect 7364 6554 7420 6556
rect 7444 6554 7500 6556
rect 7524 6554 7580 6556
rect 7604 6554 7660 6556
rect 7684 6554 7740 6556
rect 7364 6502 7366 6554
rect 7366 6502 7418 6554
rect 7418 6502 7420 6554
rect 7444 6502 7482 6554
rect 7482 6502 7494 6554
rect 7494 6502 7500 6554
rect 7524 6502 7546 6554
rect 7546 6502 7558 6554
rect 7558 6502 7580 6554
rect 7604 6502 7610 6554
rect 7610 6502 7622 6554
rect 7622 6502 7660 6554
rect 7684 6502 7686 6554
rect 7686 6502 7738 6554
rect 7738 6502 7740 6554
rect 7364 6500 7420 6502
rect 7444 6500 7500 6502
rect 7524 6500 7580 6502
rect 7604 6500 7660 6502
rect 7684 6500 7740 6502
rect 7364 5466 7420 5468
rect 7444 5466 7500 5468
rect 7524 5466 7580 5468
rect 7604 5466 7660 5468
rect 7684 5466 7740 5468
rect 7364 5414 7366 5466
rect 7366 5414 7418 5466
rect 7418 5414 7420 5466
rect 7444 5414 7482 5466
rect 7482 5414 7494 5466
rect 7494 5414 7500 5466
rect 7524 5414 7546 5466
rect 7546 5414 7558 5466
rect 7558 5414 7580 5466
rect 7604 5414 7610 5466
rect 7610 5414 7622 5466
rect 7622 5414 7660 5466
rect 7684 5414 7686 5466
rect 7686 5414 7738 5466
rect 7738 5414 7740 5466
rect 7364 5412 7420 5414
rect 7444 5412 7500 5414
rect 7524 5412 7580 5414
rect 7604 5412 7660 5414
rect 7684 5412 7740 5414
rect 7562 5108 7564 5128
rect 7564 5108 7616 5128
rect 7616 5108 7618 5128
rect 7562 5072 7618 5108
rect 8114 9560 8170 9616
rect 7930 5072 7986 5128
rect 7930 4800 7986 4856
rect 7364 4378 7420 4380
rect 7444 4378 7500 4380
rect 7524 4378 7580 4380
rect 7604 4378 7660 4380
rect 7684 4378 7740 4380
rect 7364 4326 7366 4378
rect 7366 4326 7418 4378
rect 7418 4326 7420 4378
rect 7444 4326 7482 4378
rect 7482 4326 7494 4378
rect 7494 4326 7500 4378
rect 7524 4326 7546 4378
rect 7546 4326 7558 4378
rect 7558 4326 7580 4378
rect 7604 4326 7610 4378
rect 7610 4326 7622 4378
rect 7622 4326 7660 4378
rect 7684 4326 7686 4378
rect 7686 4326 7738 4378
rect 7738 4326 7740 4378
rect 7364 4324 7420 4326
rect 7444 4324 7500 4326
rect 7524 4324 7580 4326
rect 7604 4324 7660 4326
rect 7684 4324 7740 4326
rect 7746 4020 7748 4040
rect 7748 4020 7800 4040
rect 7800 4020 7802 4040
rect 7746 3984 7802 4020
rect 7364 3290 7420 3292
rect 7444 3290 7500 3292
rect 7524 3290 7580 3292
rect 7604 3290 7660 3292
rect 7684 3290 7740 3292
rect 7364 3238 7366 3290
rect 7366 3238 7418 3290
rect 7418 3238 7420 3290
rect 7444 3238 7482 3290
rect 7482 3238 7494 3290
rect 7494 3238 7500 3290
rect 7524 3238 7546 3290
rect 7546 3238 7558 3290
rect 7558 3238 7580 3290
rect 7604 3238 7610 3290
rect 7610 3238 7622 3290
rect 7622 3238 7660 3290
rect 7684 3238 7686 3290
rect 7686 3238 7738 3290
rect 7738 3238 7740 3290
rect 7364 3236 7420 3238
rect 7444 3236 7500 3238
rect 7524 3236 7580 3238
rect 7604 3236 7660 3238
rect 7684 3236 7740 3238
rect 7838 3032 7894 3088
rect 7654 2896 7710 2952
rect 7364 2202 7420 2204
rect 7444 2202 7500 2204
rect 7524 2202 7580 2204
rect 7604 2202 7660 2204
rect 7684 2202 7740 2204
rect 7364 2150 7366 2202
rect 7366 2150 7418 2202
rect 7418 2150 7420 2202
rect 7444 2150 7482 2202
rect 7482 2150 7494 2202
rect 7494 2150 7500 2202
rect 7524 2150 7546 2202
rect 7546 2150 7558 2202
rect 7558 2150 7580 2202
rect 7604 2150 7610 2202
rect 7610 2150 7622 2202
rect 7622 2150 7660 2202
rect 7684 2150 7686 2202
rect 7686 2150 7738 2202
rect 7738 2150 7740 2202
rect 7364 2148 7420 2150
rect 7444 2148 7500 2150
rect 7524 2148 7580 2150
rect 7604 2148 7660 2150
rect 7684 2148 7740 2150
rect 8666 14184 8722 14240
rect 8666 13388 8722 13424
rect 8666 13368 8668 13388
rect 8668 13368 8720 13388
rect 8720 13368 8722 13388
rect 8666 13096 8722 13152
rect 8666 12688 8722 12744
rect 8298 12008 8354 12064
rect 8482 10412 8484 10432
rect 8484 10412 8536 10432
rect 8536 10412 8538 10432
rect 8482 10376 8538 10412
rect 8482 8472 8538 8528
rect 8482 7792 8538 7848
rect 8206 4936 8262 4992
rect 8022 1536 8078 1592
rect 8390 6160 8446 6216
rect 8390 5480 8446 5536
rect 8574 5364 8630 5400
rect 8574 5344 8576 5364
rect 8576 5344 8628 5364
rect 8628 5344 8630 5364
rect 10364 15802 10420 15804
rect 10444 15802 10500 15804
rect 10524 15802 10580 15804
rect 10604 15802 10660 15804
rect 10684 15802 10740 15804
rect 10364 15750 10366 15802
rect 10366 15750 10418 15802
rect 10418 15750 10420 15802
rect 10444 15750 10482 15802
rect 10482 15750 10494 15802
rect 10494 15750 10500 15802
rect 10524 15750 10546 15802
rect 10546 15750 10558 15802
rect 10558 15750 10580 15802
rect 10604 15750 10610 15802
rect 10610 15750 10622 15802
rect 10622 15750 10660 15802
rect 10684 15750 10686 15802
rect 10686 15750 10738 15802
rect 10738 15750 10740 15802
rect 10364 15748 10420 15750
rect 10444 15748 10500 15750
rect 10524 15748 10580 15750
rect 10604 15748 10660 15750
rect 10684 15748 10740 15750
rect 9310 15000 9366 15056
rect 9126 13096 9182 13152
rect 8666 5208 8722 5264
rect 8482 5108 8484 5128
rect 8484 5108 8536 5128
rect 8536 5108 8538 5128
rect 8482 5072 8538 5108
rect 8482 4684 8538 4720
rect 8482 4664 8484 4684
rect 8484 4664 8536 4684
rect 8536 4664 8538 4684
rect 8482 4528 8538 4584
rect 9678 13640 9734 13696
rect 9586 13504 9642 13560
rect 10046 13368 10102 13424
rect 10364 14714 10420 14716
rect 10444 14714 10500 14716
rect 10524 14714 10580 14716
rect 10604 14714 10660 14716
rect 10684 14714 10740 14716
rect 10364 14662 10366 14714
rect 10366 14662 10418 14714
rect 10418 14662 10420 14714
rect 10444 14662 10482 14714
rect 10482 14662 10494 14714
rect 10494 14662 10500 14714
rect 10524 14662 10546 14714
rect 10546 14662 10558 14714
rect 10558 14662 10580 14714
rect 10604 14662 10610 14714
rect 10610 14662 10622 14714
rect 10622 14662 10660 14714
rect 10684 14662 10686 14714
rect 10686 14662 10738 14714
rect 10738 14662 10740 14714
rect 10364 14660 10420 14662
rect 10444 14660 10500 14662
rect 10524 14660 10580 14662
rect 10604 14660 10660 14662
rect 10684 14660 10740 14662
rect 10506 14456 10562 14512
rect 10598 14320 10654 14376
rect 10364 13626 10420 13628
rect 10444 13626 10500 13628
rect 10524 13626 10580 13628
rect 10604 13626 10660 13628
rect 10684 13626 10740 13628
rect 10364 13574 10366 13626
rect 10366 13574 10418 13626
rect 10418 13574 10420 13626
rect 10444 13574 10482 13626
rect 10482 13574 10494 13626
rect 10494 13574 10500 13626
rect 10524 13574 10546 13626
rect 10546 13574 10558 13626
rect 10558 13574 10580 13626
rect 10604 13574 10610 13626
rect 10610 13574 10622 13626
rect 10622 13574 10660 13626
rect 10684 13574 10686 13626
rect 10686 13574 10738 13626
rect 10738 13574 10740 13626
rect 10364 13572 10420 13574
rect 10444 13572 10500 13574
rect 10524 13572 10580 13574
rect 10604 13572 10660 13574
rect 10684 13572 10740 13574
rect 10322 13252 10378 13288
rect 10322 13232 10324 13252
rect 10324 13232 10376 13252
rect 10376 13232 10378 13252
rect 9310 12008 9366 12064
rect 9402 11736 9458 11792
rect 9034 10920 9090 10976
rect 9770 11192 9826 11248
rect 9678 10376 9734 10432
rect 8942 9052 8944 9072
rect 8944 9052 8996 9072
rect 8996 9052 8998 9072
rect 8942 9016 8998 9052
rect 9678 10104 9734 10160
rect 9770 9016 9826 9072
rect 9586 7384 9642 7440
rect 9126 7284 9128 7304
rect 9128 7284 9180 7304
rect 9180 7284 9182 7304
rect 9126 7248 9182 7284
rect 8942 6432 8998 6488
rect 9126 6296 9182 6352
rect 9034 6160 9090 6216
rect 8942 5480 8998 5536
rect 9034 4120 9090 4176
rect 9126 3848 9182 3904
rect 8574 1808 8630 1864
rect 9034 2508 9090 2544
rect 9770 7420 9772 7440
rect 9772 7420 9824 7440
rect 9824 7420 9826 7440
rect 9770 7384 9826 7420
rect 10364 12538 10420 12540
rect 10444 12538 10500 12540
rect 10524 12538 10580 12540
rect 10604 12538 10660 12540
rect 10684 12538 10740 12540
rect 10364 12486 10366 12538
rect 10366 12486 10418 12538
rect 10418 12486 10420 12538
rect 10444 12486 10482 12538
rect 10482 12486 10494 12538
rect 10494 12486 10500 12538
rect 10524 12486 10546 12538
rect 10546 12486 10558 12538
rect 10558 12486 10580 12538
rect 10604 12486 10610 12538
rect 10610 12486 10622 12538
rect 10622 12486 10660 12538
rect 10684 12486 10686 12538
rect 10686 12486 10738 12538
rect 10738 12486 10740 12538
rect 10364 12484 10420 12486
rect 10444 12484 10500 12486
rect 10524 12484 10580 12486
rect 10604 12484 10660 12486
rect 10684 12484 10740 12486
rect 10364 11450 10420 11452
rect 10444 11450 10500 11452
rect 10524 11450 10580 11452
rect 10604 11450 10660 11452
rect 10684 11450 10740 11452
rect 10364 11398 10366 11450
rect 10366 11398 10418 11450
rect 10418 11398 10420 11450
rect 10444 11398 10482 11450
rect 10482 11398 10494 11450
rect 10494 11398 10500 11450
rect 10524 11398 10546 11450
rect 10546 11398 10558 11450
rect 10558 11398 10580 11450
rect 10604 11398 10610 11450
rect 10610 11398 10622 11450
rect 10622 11398 10660 11450
rect 10684 11398 10686 11450
rect 10686 11398 10738 11450
rect 10738 11398 10740 11450
rect 10364 11396 10420 11398
rect 10444 11396 10500 11398
rect 10524 11396 10580 11398
rect 10604 11396 10660 11398
rect 10684 11396 10740 11398
rect 10364 10362 10420 10364
rect 10444 10362 10500 10364
rect 10524 10362 10580 10364
rect 10604 10362 10660 10364
rect 10684 10362 10740 10364
rect 10364 10310 10366 10362
rect 10366 10310 10418 10362
rect 10418 10310 10420 10362
rect 10444 10310 10482 10362
rect 10482 10310 10494 10362
rect 10494 10310 10500 10362
rect 10524 10310 10546 10362
rect 10546 10310 10558 10362
rect 10558 10310 10580 10362
rect 10604 10310 10610 10362
rect 10610 10310 10622 10362
rect 10622 10310 10660 10362
rect 10684 10310 10686 10362
rect 10686 10310 10738 10362
rect 10738 10310 10740 10362
rect 10364 10308 10420 10310
rect 10444 10308 10500 10310
rect 10524 10308 10580 10310
rect 10604 10308 10660 10310
rect 10684 10308 10740 10310
rect 11334 15544 11390 15600
rect 11518 15408 11574 15464
rect 11150 13912 11206 13968
rect 10966 12688 11022 12744
rect 10230 9596 10232 9616
rect 10232 9596 10284 9616
rect 10284 9596 10286 9616
rect 10230 9560 10286 9596
rect 10364 9274 10420 9276
rect 10444 9274 10500 9276
rect 10524 9274 10580 9276
rect 10604 9274 10660 9276
rect 10684 9274 10740 9276
rect 10364 9222 10366 9274
rect 10366 9222 10418 9274
rect 10418 9222 10420 9274
rect 10444 9222 10482 9274
rect 10482 9222 10494 9274
rect 10494 9222 10500 9274
rect 10524 9222 10546 9274
rect 10546 9222 10558 9274
rect 10558 9222 10580 9274
rect 10604 9222 10610 9274
rect 10610 9222 10622 9274
rect 10622 9222 10660 9274
rect 10684 9222 10686 9274
rect 10686 9222 10738 9274
rect 10738 9222 10740 9274
rect 10364 9220 10420 9222
rect 10444 9220 10500 9222
rect 10524 9220 10580 9222
rect 10604 9220 10660 9222
rect 10684 9220 10740 9222
rect 10230 9016 10286 9072
rect 10782 8880 10838 8936
rect 10230 8356 10286 8392
rect 10230 8336 10232 8356
rect 10232 8336 10284 8356
rect 10284 8336 10286 8356
rect 10364 8186 10420 8188
rect 10444 8186 10500 8188
rect 10524 8186 10580 8188
rect 10604 8186 10660 8188
rect 10684 8186 10740 8188
rect 10364 8134 10366 8186
rect 10366 8134 10418 8186
rect 10418 8134 10420 8186
rect 10444 8134 10482 8186
rect 10482 8134 10494 8186
rect 10494 8134 10500 8186
rect 10524 8134 10546 8186
rect 10546 8134 10558 8186
rect 10558 8134 10580 8186
rect 10604 8134 10610 8186
rect 10610 8134 10622 8186
rect 10622 8134 10660 8186
rect 10684 8134 10686 8186
rect 10686 8134 10738 8186
rect 10738 8134 10740 8186
rect 10364 8132 10420 8134
rect 10444 8132 10500 8134
rect 10524 8132 10580 8134
rect 10604 8132 10660 8134
rect 10684 8132 10740 8134
rect 10364 7098 10420 7100
rect 10444 7098 10500 7100
rect 10524 7098 10580 7100
rect 10604 7098 10660 7100
rect 10684 7098 10740 7100
rect 10364 7046 10366 7098
rect 10366 7046 10418 7098
rect 10418 7046 10420 7098
rect 10444 7046 10482 7098
rect 10482 7046 10494 7098
rect 10494 7046 10500 7098
rect 10524 7046 10546 7098
rect 10546 7046 10558 7098
rect 10558 7046 10580 7098
rect 10604 7046 10610 7098
rect 10610 7046 10622 7098
rect 10622 7046 10660 7098
rect 10684 7046 10686 7098
rect 10686 7046 10738 7098
rect 10738 7046 10740 7098
rect 10364 7044 10420 7046
rect 10444 7044 10500 7046
rect 10524 7044 10580 7046
rect 10604 7044 10660 7046
rect 10684 7044 10740 7046
rect 10414 6740 10416 6760
rect 10416 6740 10468 6760
rect 10468 6740 10470 6760
rect 9954 6568 10010 6624
rect 9862 5208 9918 5264
rect 9678 5072 9734 5128
rect 9034 2488 9036 2508
rect 9036 2488 9088 2508
rect 9088 2488 9090 2508
rect 9126 2352 9182 2408
rect 4364 570 4420 572
rect 4444 570 4500 572
rect 4524 570 4580 572
rect 4604 570 4660 572
rect 4684 570 4740 572
rect 4364 518 4366 570
rect 4366 518 4418 570
rect 4418 518 4420 570
rect 4444 518 4482 570
rect 4482 518 4494 570
rect 4494 518 4500 570
rect 4524 518 4546 570
rect 4546 518 4558 570
rect 4558 518 4580 570
rect 4604 518 4610 570
rect 4610 518 4622 570
rect 4622 518 4660 570
rect 4684 518 4686 570
rect 4686 518 4738 570
rect 4738 518 4740 570
rect 4364 516 4420 518
rect 4444 516 4500 518
rect 4524 516 4580 518
rect 4604 516 4660 518
rect 4684 516 4740 518
rect 7364 1114 7420 1116
rect 7444 1114 7500 1116
rect 7524 1114 7580 1116
rect 7604 1114 7660 1116
rect 7684 1114 7740 1116
rect 7364 1062 7366 1114
rect 7366 1062 7418 1114
rect 7418 1062 7420 1114
rect 7444 1062 7482 1114
rect 7482 1062 7494 1114
rect 7494 1062 7500 1114
rect 7524 1062 7546 1114
rect 7546 1062 7558 1114
rect 7558 1062 7580 1114
rect 7604 1062 7610 1114
rect 7610 1062 7622 1114
rect 7622 1062 7660 1114
rect 7684 1062 7686 1114
rect 7686 1062 7738 1114
rect 7738 1062 7740 1114
rect 7364 1060 7420 1062
rect 7444 1060 7500 1062
rect 7524 1060 7580 1062
rect 7604 1060 7660 1062
rect 7684 1060 7740 1062
rect 9770 3304 9826 3360
rect 9770 1672 9826 1728
rect 9678 1536 9734 1592
rect 9678 1128 9734 1184
rect 10414 6704 10470 6740
rect 10364 6010 10420 6012
rect 10444 6010 10500 6012
rect 10524 6010 10580 6012
rect 10604 6010 10660 6012
rect 10684 6010 10740 6012
rect 10364 5958 10366 6010
rect 10366 5958 10418 6010
rect 10418 5958 10420 6010
rect 10444 5958 10482 6010
rect 10482 5958 10494 6010
rect 10494 5958 10500 6010
rect 10524 5958 10546 6010
rect 10546 5958 10558 6010
rect 10558 5958 10580 6010
rect 10604 5958 10610 6010
rect 10610 5958 10622 6010
rect 10622 5958 10660 6010
rect 10684 5958 10686 6010
rect 10686 5958 10738 6010
rect 10738 5958 10740 6010
rect 10364 5956 10420 5958
rect 10444 5956 10500 5958
rect 10524 5956 10580 5958
rect 10604 5956 10660 5958
rect 10684 5956 10740 5958
rect 10364 4922 10420 4924
rect 10444 4922 10500 4924
rect 10524 4922 10580 4924
rect 10604 4922 10660 4924
rect 10684 4922 10740 4924
rect 10364 4870 10366 4922
rect 10366 4870 10418 4922
rect 10418 4870 10420 4922
rect 10444 4870 10482 4922
rect 10482 4870 10494 4922
rect 10494 4870 10500 4922
rect 10524 4870 10546 4922
rect 10546 4870 10558 4922
rect 10558 4870 10580 4922
rect 10604 4870 10610 4922
rect 10610 4870 10622 4922
rect 10622 4870 10660 4922
rect 10684 4870 10686 4922
rect 10686 4870 10738 4922
rect 10738 4870 10740 4922
rect 10364 4868 10420 4870
rect 10444 4868 10500 4870
rect 10524 4868 10580 4870
rect 10604 4868 10660 4870
rect 10684 4868 10740 4870
rect 10364 3834 10420 3836
rect 10444 3834 10500 3836
rect 10524 3834 10580 3836
rect 10604 3834 10660 3836
rect 10684 3834 10740 3836
rect 10364 3782 10366 3834
rect 10366 3782 10418 3834
rect 10418 3782 10420 3834
rect 10444 3782 10482 3834
rect 10482 3782 10494 3834
rect 10494 3782 10500 3834
rect 10524 3782 10546 3834
rect 10546 3782 10558 3834
rect 10558 3782 10580 3834
rect 10604 3782 10610 3834
rect 10610 3782 10622 3834
rect 10622 3782 10660 3834
rect 10684 3782 10686 3834
rect 10686 3782 10738 3834
rect 10738 3782 10740 3834
rect 10364 3780 10420 3782
rect 10444 3780 10500 3782
rect 10524 3780 10580 3782
rect 10604 3780 10660 3782
rect 10684 3780 10740 3782
rect 10364 2746 10420 2748
rect 10444 2746 10500 2748
rect 10524 2746 10580 2748
rect 10604 2746 10660 2748
rect 10684 2746 10740 2748
rect 10364 2694 10366 2746
rect 10366 2694 10418 2746
rect 10418 2694 10420 2746
rect 10444 2694 10482 2746
rect 10482 2694 10494 2746
rect 10494 2694 10500 2746
rect 10524 2694 10546 2746
rect 10546 2694 10558 2746
rect 10558 2694 10580 2746
rect 10604 2694 10610 2746
rect 10610 2694 10622 2746
rect 10622 2694 10660 2746
rect 10684 2694 10686 2746
rect 10686 2694 10738 2746
rect 10738 2694 10740 2746
rect 10364 2692 10420 2694
rect 10444 2692 10500 2694
rect 10524 2692 10580 2694
rect 10604 2692 10660 2694
rect 10684 2692 10740 2694
rect 13364 17434 13420 17436
rect 13444 17434 13500 17436
rect 13524 17434 13580 17436
rect 13604 17434 13660 17436
rect 13684 17434 13740 17436
rect 13364 17382 13366 17434
rect 13366 17382 13418 17434
rect 13418 17382 13420 17434
rect 13444 17382 13482 17434
rect 13482 17382 13494 17434
rect 13494 17382 13500 17434
rect 13524 17382 13546 17434
rect 13546 17382 13558 17434
rect 13558 17382 13580 17434
rect 13604 17382 13610 17434
rect 13610 17382 13622 17434
rect 13622 17382 13660 17434
rect 13684 17382 13686 17434
rect 13686 17382 13738 17434
rect 13738 17382 13740 17434
rect 13364 17380 13420 17382
rect 13444 17380 13500 17382
rect 13524 17380 13580 17382
rect 13604 17380 13660 17382
rect 13684 17380 13740 17382
rect 11978 14456 12034 14512
rect 11886 13368 11942 13424
rect 12254 15272 12310 15328
rect 12162 14320 12218 14376
rect 12070 14048 12126 14104
rect 13364 16346 13420 16348
rect 13444 16346 13500 16348
rect 13524 16346 13580 16348
rect 13604 16346 13660 16348
rect 13684 16346 13740 16348
rect 13364 16294 13366 16346
rect 13366 16294 13418 16346
rect 13418 16294 13420 16346
rect 13444 16294 13482 16346
rect 13482 16294 13494 16346
rect 13494 16294 13500 16346
rect 13524 16294 13546 16346
rect 13546 16294 13558 16346
rect 13558 16294 13580 16346
rect 13604 16294 13610 16346
rect 13610 16294 13622 16346
rect 13622 16294 13660 16346
rect 13684 16294 13686 16346
rect 13686 16294 13738 16346
rect 13738 16294 13740 16346
rect 13364 16292 13420 16294
rect 13444 16292 13500 16294
rect 13524 16292 13580 16294
rect 13604 16292 13660 16294
rect 13684 16292 13740 16294
rect 12990 15444 12992 15464
rect 12992 15444 13044 15464
rect 13044 15444 13046 15464
rect 12990 15408 13046 15444
rect 12898 15272 12954 15328
rect 12622 14884 12678 14920
rect 12622 14864 12624 14884
rect 12624 14864 12676 14884
rect 12676 14864 12678 14884
rect 12530 13812 12532 13832
rect 12532 13812 12584 13832
rect 12584 13812 12586 13832
rect 12530 13776 12586 13812
rect 10874 2080 10930 2136
rect 10364 1658 10420 1660
rect 10444 1658 10500 1660
rect 10524 1658 10580 1660
rect 10604 1658 10660 1660
rect 10684 1658 10740 1660
rect 10364 1606 10366 1658
rect 10366 1606 10418 1658
rect 10418 1606 10420 1658
rect 10444 1606 10482 1658
rect 10482 1606 10494 1658
rect 10494 1606 10500 1658
rect 10524 1606 10546 1658
rect 10546 1606 10558 1658
rect 10558 1606 10580 1658
rect 10604 1606 10610 1658
rect 10610 1606 10622 1658
rect 10622 1606 10660 1658
rect 10684 1606 10686 1658
rect 10686 1606 10738 1658
rect 10738 1606 10740 1658
rect 10364 1604 10420 1606
rect 10444 1604 10500 1606
rect 10524 1604 10580 1606
rect 10604 1604 10660 1606
rect 10684 1604 10740 1606
rect 10690 1264 10746 1320
rect 11058 1300 11060 1320
rect 11060 1300 11112 1320
rect 11112 1300 11114 1320
rect 11058 1264 11114 1300
rect 11426 6024 11482 6080
rect 11794 7248 11850 7304
rect 12254 11092 12256 11112
rect 12256 11092 12308 11112
rect 12308 11092 12310 11112
rect 12254 11056 12310 11092
rect 12346 10512 12402 10568
rect 12622 13640 12678 13696
rect 12530 12844 12586 12880
rect 12530 12824 12532 12844
rect 12532 12824 12584 12844
rect 12584 12824 12586 12844
rect 12622 11736 12678 11792
rect 13266 15544 13322 15600
rect 13364 15258 13420 15260
rect 13444 15258 13500 15260
rect 13524 15258 13580 15260
rect 13604 15258 13660 15260
rect 13684 15258 13740 15260
rect 13364 15206 13366 15258
rect 13366 15206 13418 15258
rect 13418 15206 13420 15258
rect 13444 15206 13482 15258
rect 13482 15206 13494 15258
rect 13494 15206 13500 15258
rect 13524 15206 13546 15258
rect 13546 15206 13558 15258
rect 13558 15206 13580 15258
rect 13604 15206 13610 15258
rect 13610 15206 13622 15258
rect 13622 15206 13660 15258
rect 13684 15206 13686 15258
rect 13686 15206 13738 15258
rect 13738 15206 13740 15258
rect 13364 15204 13420 15206
rect 13444 15204 13500 15206
rect 13524 15204 13580 15206
rect 13604 15204 13660 15206
rect 13684 15204 13740 15206
rect 13358 14864 13414 14920
rect 13910 15000 13966 15056
rect 12438 9052 12440 9072
rect 12440 9052 12492 9072
rect 12492 9052 12494 9072
rect 12438 9016 12494 9052
rect 12806 9560 12862 9616
rect 12622 8336 12678 8392
rect 11978 5516 11980 5536
rect 11980 5516 12032 5536
rect 12032 5516 12034 5536
rect 11978 5480 12034 5516
rect 12162 7384 12218 7440
rect 12162 5752 12218 5808
rect 12254 3576 12310 3632
rect 11334 1944 11390 2000
rect 10364 570 10420 572
rect 10444 570 10500 572
rect 10524 570 10580 572
rect 10604 570 10660 572
rect 10684 570 10740 572
rect 10364 518 10366 570
rect 10366 518 10418 570
rect 10418 518 10420 570
rect 10444 518 10482 570
rect 10482 518 10494 570
rect 10494 518 10500 570
rect 10524 518 10546 570
rect 10546 518 10558 570
rect 10558 518 10580 570
rect 10604 518 10610 570
rect 10610 518 10622 570
rect 10622 518 10660 570
rect 10684 518 10686 570
rect 10686 518 10738 570
rect 10738 518 10740 570
rect 10364 516 10420 518
rect 10444 516 10500 518
rect 10524 516 10580 518
rect 10604 516 10660 518
rect 10684 516 10740 518
rect 12806 6296 12862 6352
rect 12622 5752 12678 5808
rect 12346 2896 12402 2952
rect 12530 2352 12586 2408
rect 12806 5616 12862 5672
rect 13364 14170 13420 14172
rect 13444 14170 13500 14172
rect 13524 14170 13580 14172
rect 13604 14170 13660 14172
rect 13684 14170 13740 14172
rect 13364 14118 13366 14170
rect 13366 14118 13418 14170
rect 13418 14118 13420 14170
rect 13444 14118 13482 14170
rect 13482 14118 13494 14170
rect 13494 14118 13500 14170
rect 13524 14118 13546 14170
rect 13546 14118 13558 14170
rect 13558 14118 13580 14170
rect 13604 14118 13610 14170
rect 13610 14118 13622 14170
rect 13622 14118 13660 14170
rect 13684 14118 13686 14170
rect 13686 14118 13738 14170
rect 13738 14118 13740 14170
rect 13364 14116 13420 14118
rect 13444 14116 13500 14118
rect 13524 14116 13580 14118
rect 13604 14116 13660 14118
rect 13684 14116 13740 14118
rect 14002 13640 14058 13696
rect 13364 13082 13420 13084
rect 13444 13082 13500 13084
rect 13524 13082 13580 13084
rect 13604 13082 13660 13084
rect 13684 13082 13740 13084
rect 13364 13030 13366 13082
rect 13366 13030 13418 13082
rect 13418 13030 13420 13082
rect 13444 13030 13482 13082
rect 13482 13030 13494 13082
rect 13494 13030 13500 13082
rect 13524 13030 13546 13082
rect 13546 13030 13558 13082
rect 13558 13030 13580 13082
rect 13604 13030 13610 13082
rect 13610 13030 13622 13082
rect 13622 13030 13660 13082
rect 13684 13030 13686 13082
rect 13686 13030 13738 13082
rect 13738 13030 13740 13082
rect 13364 13028 13420 13030
rect 13444 13028 13500 13030
rect 13524 13028 13580 13030
rect 13604 13028 13660 13030
rect 13684 13028 13740 13030
rect 16364 16890 16420 16892
rect 16444 16890 16500 16892
rect 16524 16890 16580 16892
rect 16604 16890 16660 16892
rect 16684 16890 16740 16892
rect 16364 16838 16366 16890
rect 16366 16838 16418 16890
rect 16418 16838 16420 16890
rect 16444 16838 16482 16890
rect 16482 16838 16494 16890
rect 16494 16838 16500 16890
rect 16524 16838 16546 16890
rect 16546 16838 16558 16890
rect 16558 16838 16580 16890
rect 16604 16838 16610 16890
rect 16610 16838 16622 16890
rect 16622 16838 16660 16890
rect 16684 16838 16686 16890
rect 16686 16838 16738 16890
rect 16738 16838 16740 16890
rect 16364 16836 16420 16838
rect 16444 16836 16500 16838
rect 16524 16836 16580 16838
rect 16604 16836 16660 16838
rect 16684 16836 16740 16838
rect 16364 15802 16420 15804
rect 16444 15802 16500 15804
rect 16524 15802 16580 15804
rect 16604 15802 16660 15804
rect 16684 15802 16740 15804
rect 16364 15750 16366 15802
rect 16366 15750 16418 15802
rect 16418 15750 16420 15802
rect 16444 15750 16482 15802
rect 16482 15750 16494 15802
rect 16494 15750 16500 15802
rect 16524 15750 16546 15802
rect 16546 15750 16558 15802
rect 16558 15750 16580 15802
rect 16604 15750 16610 15802
rect 16610 15750 16622 15802
rect 16622 15750 16660 15802
rect 16684 15750 16686 15802
rect 16686 15750 16738 15802
rect 16738 15750 16740 15802
rect 16364 15748 16420 15750
rect 16444 15748 16500 15750
rect 16524 15748 16580 15750
rect 16604 15748 16660 15750
rect 16684 15748 16740 15750
rect 13364 11994 13420 11996
rect 13444 11994 13500 11996
rect 13524 11994 13580 11996
rect 13604 11994 13660 11996
rect 13684 11994 13740 11996
rect 13364 11942 13366 11994
rect 13366 11942 13418 11994
rect 13418 11942 13420 11994
rect 13444 11942 13482 11994
rect 13482 11942 13494 11994
rect 13494 11942 13500 11994
rect 13524 11942 13546 11994
rect 13546 11942 13558 11994
rect 13558 11942 13580 11994
rect 13604 11942 13610 11994
rect 13610 11942 13622 11994
rect 13622 11942 13660 11994
rect 13684 11942 13686 11994
rect 13686 11942 13738 11994
rect 13738 11942 13740 11994
rect 13364 11940 13420 11942
rect 13444 11940 13500 11942
rect 13524 11940 13580 11942
rect 13604 11940 13660 11942
rect 13684 11940 13740 11942
rect 13634 11076 13690 11112
rect 13634 11056 13636 11076
rect 13636 11056 13688 11076
rect 13688 11056 13690 11076
rect 13364 10906 13420 10908
rect 13444 10906 13500 10908
rect 13524 10906 13580 10908
rect 13604 10906 13660 10908
rect 13684 10906 13740 10908
rect 13364 10854 13366 10906
rect 13366 10854 13418 10906
rect 13418 10854 13420 10906
rect 13444 10854 13482 10906
rect 13482 10854 13494 10906
rect 13494 10854 13500 10906
rect 13524 10854 13546 10906
rect 13546 10854 13558 10906
rect 13558 10854 13580 10906
rect 13604 10854 13610 10906
rect 13610 10854 13622 10906
rect 13622 10854 13660 10906
rect 13684 10854 13686 10906
rect 13686 10854 13738 10906
rect 13738 10854 13740 10906
rect 13364 10852 13420 10854
rect 13444 10852 13500 10854
rect 13524 10852 13580 10854
rect 13604 10852 13660 10854
rect 13684 10852 13740 10854
rect 13358 10648 13414 10704
rect 13364 9818 13420 9820
rect 13444 9818 13500 9820
rect 13524 9818 13580 9820
rect 13604 9818 13660 9820
rect 13684 9818 13740 9820
rect 13364 9766 13366 9818
rect 13366 9766 13418 9818
rect 13418 9766 13420 9818
rect 13444 9766 13482 9818
rect 13482 9766 13494 9818
rect 13494 9766 13500 9818
rect 13524 9766 13546 9818
rect 13546 9766 13558 9818
rect 13558 9766 13580 9818
rect 13604 9766 13610 9818
rect 13610 9766 13622 9818
rect 13622 9766 13660 9818
rect 13684 9766 13686 9818
rect 13686 9766 13738 9818
rect 13738 9766 13740 9818
rect 13364 9764 13420 9766
rect 13444 9764 13500 9766
rect 13524 9764 13580 9766
rect 13604 9764 13660 9766
rect 13684 9764 13740 9766
rect 13174 8880 13230 8936
rect 13364 8730 13420 8732
rect 13444 8730 13500 8732
rect 13524 8730 13580 8732
rect 13604 8730 13660 8732
rect 13684 8730 13740 8732
rect 13364 8678 13366 8730
rect 13366 8678 13418 8730
rect 13418 8678 13420 8730
rect 13444 8678 13482 8730
rect 13482 8678 13494 8730
rect 13494 8678 13500 8730
rect 13524 8678 13546 8730
rect 13546 8678 13558 8730
rect 13558 8678 13580 8730
rect 13604 8678 13610 8730
rect 13610 8678 13622 8730
rect 13622 8678 13660 8730
rect 13684 8678 13686 8730
rect 13686 8678 13738 8730
rect 13738 8678 13740 8730
rect 13364 8676 13420 8678
rect 13444 8676 13500 8678
rect 13524 8676 13580 8678
rect 13604 8676 13660 8678
rect 13684 8676 13740 8678
rect 12990 5888 13046 5944
rect 12806 5480 12862 5536
rect 12898 5344 12954 5400
rect 12990 3168 13046 3224
rect 12346 1844 12348 1864
rect 12348 1844 12400 1864
rect 12400 1844 12402 1864
rect 12346 1808 12402 1844
rect 12806 1944 12862 2000
rect 13364 7642 13420 7644
rect 13444 7642 13500 7644
rect 13524 7642 13580 7644
rect 13604 7642 13660 7644
rect 13684 7642 13740 7644
rect 13364 7590 13366 7642
rect 13366 7590 13418 7642
rect 13418 7590 13420 7642
rect 13444 7590 13482 7642
rect 13482 7590 13494 7642
rect 13494 7590 13500 7642
rect 13524 7590 13546 7642
rect 13546 7590 13558 7642
rect 13558 7590 13580 7642
rect 13604 7590 13610 7642
rect 13610 7590 13622 7642
rect 13622 7590 13660 7642
rect 13684 7590 13686 7642
rect 13686 7590 13738 7642
rect 13738 7590 13740 7642
rect 13364 7588 13420 7590
rect 13444 7588 13500 7590
rect 13524 7588 13580 7590
rect 13604 7588 13660 7590
rect 13684 7588 13740 7590
rect 13364 6554 13420 6556
rect 13444 6554 13500 6556
rect 13524 6554 13580 6556
rect 13604 6554 13660 6556
rect 13684 6554 13740 6556
rect 13364 6502 13366 6554
rect 13366 6502 13418 6554
rect 13418 6502 13420 6554
rect 13444 6502 13482 6554
rect 13482 6502 13494 6554
rect 13494 6502 13500 6554
rect 13524 6502 13546 6554
rect 13546 6502 13558 6554
rect 13558 6502 13580 6554
rect 13604 6502 13610 6554
rect 13610 6502 13622 6554
rect 13622 6502 13660 6554
rect 13684 6502 13686 6554
rect 13686 6502 13738 6554
rect 13738 6502 13740 6554
rect 13364 6500 13420 6502
rect 13444 6500 13500 6502
rect 13524 6500 13580 6502
rect 13604 6500 13660 6502
rect 13684 6500 13740 6502
rect 13634 6160 13690 6216
rect 13542 5752 13598 5808
rect 13364 5466 13420 5468
rect 13444 5466 13500 5468
rect 13524 5466 13580 5468
rect 13604 5466 13660 5468
rect 13684 5466 13740 5468
rect 13364 5414 13366 5466
rect 13366 5414 13418 5466
rect 13418 5414 13420 5466
rect 13444 5414 13482 5466
rect 13482 5414 13494 5466
rect 13494 5414 13500 5466
rect 13524 5414 13546 5466
rect 13546 5414 13558 5466
rect 13558 5414 13580 5466
rect 13604 5414 13610 5466
rect 13610 5414 13622 5466
rect 13622 5414 13660 5466
rect 13684 5414 13686 5466
rect 13686 5414 13738 5466
rect 13738 5414 13740 5466
rect 13364 5412 13420 5414
rect 13444 5412 13500 5414
rect 13524 5412 13580 5414
rect 13604 5412 13660 5414
rect 13684 5412 13740 5414
rect 13358 5108 13360 5128
rect 13360 5108 13412 5128
rect 13412 5108 13414 5128
rect 13358 5072 13414 5108
rect 13364 4378 13420 4380
rect 13444 4378 13500 4380
rect 13524 4378 13580 4380
rect 13604 4378 13660 4380
rect 13684 4378 13740 4380
rect 13364 4326 13366 4378
rect 13366 4326 13418 4378
rect 13418 4326 13420 4378
rect 13444 4326 13482 4378
rect 13482 4326 13494 4378
rect 13494 4326 13500 4378
rect 13524 4326 13546 4378
rect 13546 4326 13558 4378
rect 13558 4326 13580 4378
rect 13604 4326 13610 4378
rect 13610 4326 13622 4378
rect 13622 4326 13660 4378
rect 13684 4326 13686 4378
rect 13686 4326 13738 4378
rect 13738 4326 13740 4378
rect 13364 4324 13420 4326
rect 13444 4324 13500 4326
rect 13524 4324 13580 4326
rect 13604 4324 13660 4326
rect 13684 4324 13740 4326
rect 14370 11600 14426 11656
rect 14278 11192 14334 11248
rect 14370 7404 14426 7440
rect 14370 7384 14372 7404
rect 14372 7384 14424 7404
rect 14424 7384 14426 7404
rect 14186 7112 14242 7168
rect 14186 6024 14242 6080
rect 14094 5616 14150 5672
rect 14830 8472 14886 8528
rect 13082 2080 13138 2136
rect 13364 3290 13420 3292
rect 13444 3290 13500 3292
rect 13524 3290 13580 3292
rect 13604 3290 13660 3292
rect 13684 3290 13740 3292
rect 13364 3238 13366 3290
rect 13366 3238 13418 3290
rect 13418 3238 13420 3290
rect 13444 3238 13482 3290
rect 13482 3238 13494 3290
rect 13494 3238 13500 3290
rect 13524 3238 13546 3290
rect 13546 3238 13558 3290
rect 13558 3238 13580 3290
rect 13604 3238 13610 3290
rect 13610 3238 13622 3290
rect 13622 3238 13660 3290
rect 13684 3238 13686 3290
rect 13686 3238 13738 3290
rect 13738 3238 13740 3290
rect 13364 3236 13420 3238
rect 13444 3236 13500 3238
rect 13524 3236 13580 3238
rect 13604 3236 13660 3238
rect 13684 3236 13740 3238
rect 13818 3052 13874 3088
rect 13818 3032 13820 3052
rect 13820 3032 13872 3052
rect 13872 3032 13874 3052
rect 13364 2202 13420 2204
rect 13444 2202 13500 2204
rect 13524 2202 13580 2204
rect 13604 2202 13660 2204
rect 13684 2202 13740 2204
rect 13364 2150 13366 2202
rect 13366 2150 13418 2202
rect 13418 2150 13420 2202
rect 13444 2150 13482 2202
rect 13482 2150 13494 2202
rect 13494 2150 13500 2202
rect 13524 2150 13546 2202
rect 13546 2150 13558 2202
rect 13558 2150 13580 2202
rect 13604 2150 13610 2202
rect 13610 2150 13622 2202
rect 13622 2150 13660 2202
rect 13684 2150 13686 2202
rect 13686 2150 13738 2202
rect 13738 2150 13740 2202
rect 13364 2148 13420 2150
rect 13444 2148 13500 2150
rect 13524 2148 13580 2150
rect 13604 2148 13660 2150
rect 13684 2148 13740 2150
rect 13358 1964 13414 2000
rect 13910 2216 13966 2272
rect 13358 1944 13360 1964
rect 13360 1944 13412 1964
rect 13412 1944 13414 1964
rect 13818 1672 13874 1728
rect 13910 1536 13966 1592
rect 13364 1114 13420 1116
rect 13444 1114 13500 1116
rect 13524 1114 13580 1116
rect 13604 1114 13660 1116
rect 13684 1114 13740 1116
rect 13364 1062 13366 1114
rect 13366 1062 13418 1114
rect 13418 1062 13420 1114
rect 13444 1062 13482 1114
rect 13482 1062 13494 1114
rect 13494 1062 13500 1114
rect 13524 1062 13546 1114
rect 13546 1062 13558 1114
rect 13558 1062 13580 1114
rect 13604 1062 13610 1114
rect 13610 1062 13622 1114
rect 13622 1062 13660 1114
rect 13684 1062 13686 1114
rect 13686 1062 13738 1114
rect 13738 1062 13740 1114
rect 13364 1060 13420 1062
rect 13444 1060 13500 1062
rect 13524 1060 13580 1062
rect 13604 1060 13660 1062
rect 13684 1060 13740 1062
rect 14186 3032 14242 3088
rect 14002 1128 14058 1184
rect 14554 3576 14610 3632
rect 14922 6976 14978 7032
rect 14830 6316 14886 6352
rect 14830 6296 14832 6316
rect 14832 6296 14884 6316
rect 14884 6296 14886 6316
rect 14554 2624 14610 2680
rect 15198 3984 15254 4040
rect 15750 14340 15806 14376
rect 15750 14320 15752 14340
rect 15752 14320 15804 14340
rect 15804 14320 15806 14340
rect 16364 14714 16420 14716
rect 16444 14714 16500 14716
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16364 14662 16366 14714
rect 16366 14662 16418 14714
rect 16418 14662 16420 14714
rect 16444 14662 16482 14714
rect 16482 14662 16494 14714
rect 16494 14662 16500 14714
rect 16524 14662 16546 14714
rect 16546 14662 16558 14714
rect 16558 14662 16580 14714
rect 16604 14662 16610 14714
rect 16610 14662 16622 14714
rect 16622 14662 16660 14714
rect 16684 14662 16686 14714
rect 16686 14662 16738 14714
rect 16738 14662 16740 14714
rect 16364 14660 16420 14662
rect 16444 14660 16500 14662
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16946 14456 17002 14512
rect 16118 13640 16174 13696
rect 16364 13626 16420 13628
rect 16444 13626 16500 13628
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16364 13574 16366 13626
rect 16366 13574 16418 13626
rect 16418 13574 16420 13626
rect 16444 13574 16482 13626
rect 16482 13574 16494 13626
rect 16494 13574 16500 13626
rect 16524 13574 16546 13626
rect 16546 13574 16558 13626
rect 16558 13574 16580 13626
rect 16604 13574 16610 13626
rect 16610 13574 16622 13626
rect 16622 13574 16660 13626
rect 16684 13574 16686 13626
rect 16686 13574 16738 13626
rect 16738 13574 16740 13626
rect 16364 13572 16420 13574
rect 16444 13572 16500 13574
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16364 12538 16420 12540
rect 16444 12538 16500 12540
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16364 12486 16366 12538
rect 16366 12486 16418 12538
rect 16418 12486 16420 12538
rect 16444 12486 16482 12538
rect 16482 12486 16494 12538
rect 16494 12486 16500 12538
rect 16524 12486 16546 12538
rect 16546 12486 16558 12538
rect 16558 12486 16580 12538
rect 16604 12486 16610 12538
rect 16610 12486 16622 12538
rect 16622 12486 16660 12538
rect 16684 12486 16686 12538
rect 16686 12486 16738 12538
rect 16738 12486 16740 12538
rect 16364 12484 16420 12486
rect 16444 12484 16500 12486
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 15750 9036 15806 9072
rect 15750 9016 15752 9036
rect 15752 9016 15804 9036
rect 15804 9016 15806 9036
rect 15750 8472 15806 8528
rect 16364 11450 16420 11452
rect 16444 11450 16500 11452
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16364 11398 16366 11450
rect 16366 11398 16418 11450
rect 16418 11398 16420 11450
rect 16444 11398 16482 11450
rect 16482 11398 16494 11450
rect 16494 11398 16500 11450
rect 16524 11398 16546 11450
rect 16546 11398 16558 11450
rect 16558 11398 16580 11450
rect 16604 11398 16610 11450
rect 16610 11398 16622 11450
rect 16622 11398 16660 11450
rect 16684 11398 16686 11450
rect 16686 11398 16738 11450
rect 16738 11398 16740 11450
rect 16364 11396 16420 11398
rect 16444 11396 16500 11398
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16578 11056 16634 11112
rect 16364 10362 16420 10364
rect 16444 10362 16500 10364
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16364 10310 16366 10362
rect 16366 10310 16418 10362
rect 16418 10310 16420 10362
rect 16444 10310 16482 10362
rect 16482 10310 16494 10362
rect 16494 10310 16500 10362
rect 16524 10310 16546 10362
rect 16546 10310 16558 10362
rect 16558 10310 16580 10362
rect 16604 10310 16610 10362
rect 16610 10310 16622 10362
rect 16622 10310 16660 10362
rect 16684 10310 16686 10362
rect 16686 10310 16738 10362
rect 16738 10310 16740 10362
rect 16364 10308 16420 10310
rect 16444 10308 16500 10310
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16210 9560 16266 9616
rect 16364 9274 16420 9276
rect 16444 9274 16500 9276
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16364 9222 16366 9274
rect 16366 9222 16418 9274
rect 16418 9222 16420 9274
rect 16444 9222 16482 9274
rect 16482 9222 16494 9274
rect 16494 9222 16500 9274
rect 16524 9222 16546 9274
rect 16546 9222 16558 9274
rect 16558 9222 16580 9274
rect 16604 9222 16610 9274
rect 16610 9222 16622 9274
rect 16622 9222 16660 9274
rect 16684 9222 16686 9274
rect 16686 9222 16738 9274
rect 16738 9222 16740 9274
rect 16364 9220 16420 9222
rect 16444 9220 16500 9222
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16364 8186 16420 8188
rect 16444 8186 16500 8188
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16364 8134 16366 8186
rect 16366 8134 16418 8186
rect 16418 8134 16420 8186
rect 16444 8134 16482 8186
rect 16482 8134 16494 8186
rect 16494 8134 16500 8186
rect 16524 8134 16546 8186
rect 16546 8134 16558 8186
rect 16558 8134 16580 8186
rect 16604 8134 16610 8186
rect 16610 8134 16622 8186
rect 16622 8134 16660 8186
rect 16684 8134 16686 8186
rect 16686 8134 16738 8186
rect 16738 8134 16740 8186
rect 16364 8132 16420 8134
rect 16444 8132 16500 8134
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16364 7098 16420 7100
rect 16444 7098 16500 7100
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16364 7046 16366 7098
rect 16366 7046 16418 7098
rect 16418 7046 16420 7098
rect 16444 7046 16482 7098
rect 16482 7046 16494 7098
rect 16494 7046 16500 7098
rect 16524 7046 16546 7098
rect 16546 7046 16558 7098
rect 16558 7046 16580 7098
rect 16604 7046 16610 7098
rect 16610 7046 16622 7098
rect 16622 7046 16660 7098
rect 16684 7046 16686 7098
rect 16686 7046 16738 7098
rect 16738 7046 16740 7098
rect 16364 7044 16420 7046
rect 16444 7044 16500 7046
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16364 6010 16420 6012
rect 16444 6010 16500 6012
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16364 5958 16366 6010
rect 16366 5958 16418 6010
rect 16418 5958 16420 6010
rect 16444 5958 16482 6010
rect 16482 5958 16494 6010
rect 16494 5958 16500 6010
rect 16524 5958 16546 6010
rect 16546 5958 16558 6010
rect 16558 5958 16580 6010
rect 16604 5958 16610 6010
rect 16610 5958 16622 6010
rect 16622 5958 16660 6010
rect 16684 5958 16686 6010
rect 16686 5958 16738 6010
rect 16738 5958 16740 6010
rect 16364 5956 16420 5958
rect 16444 5956 16500 5958
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16854 5752 16910 5808
rect 16364 4922 16420 4924
rect 16444 4922 16500 4924
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16364 4870 16366 4922
rect 16366 4870 16418 4922
rect 16418 4870 16420 4922
rect 16444 4870 16482 4922
rect 16482 4870 16494 4922
rect 16494 4870 16500 4922
rect 16524 4870 16546 4922
rect 16546 4870 16558 4922
rect 16558 4870 16580 4922
rect 16604 4870 16610 4922
rect 16610 4870 16622 4922
rect 16622 4870 16660 4922
rect 16684 4870 16686 4922
rect 16686 4870 16738 4922
rect 16738 4870 16740 4922
rect 16364 4868 16420 4870
rect 16444 4868 16500 4870
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 15566 3848 15622 3904
rect 15290 2932 15292 2952
rect 15292 2932 15344 2952
rect 15344 2932 15346 2952
rect 15290 2896 15346 2932
rect 14922 1844 14924 1864
rect 14924 1844 14976 1864
rect 14976 1844 14978 1864
rect 14922 1808 14978 1844
rect 15106 1264 15162 1320
rect 16364 3834 16420 3836
rect 16444 3834 16500 3836
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16364 3782 16366 3834
rect 16366 3782 16418 3834
rect 16418 3782 16420 3834
rect 16444 3782 16482 3834
rect 16482 3782 16494 3834
rect 16494 3782 16500 3834
rect 16524 3782 16546 3834
rect 16546 3782 16558 3834
rect 16558 3782 16580 3834
rect 16604 3782 16610 3834
rect 16610 3782 16622 3834
rect 16622 3782 16660 3834
rect 16684 3782 16686 3834
rect 16686 3782 16738 3834
rect 16738 3782 16740 3834
rect 16364 3780 16420 3782
rect 16444 3780 16500 3782
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 15290 2080 15346 2136
rect 15198 1128 15254 1184
rect 15474 1808 15530 1864
rect 16026 2252 16028 2272
rect 16028 2252 16080 2272
rect 16080 2252 16082 2272
rect 15658 2080 15714 2136
rect 15750 1672 15806 1728
rect 15658 1400 15714 1456
rect 16026 2216 16082 2252
rect 16364 2746 16420 2748
rect 16444 2746 16500 2748
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16364 2694 16366 2746
rect 16366 2694 16418 2746
rect 16418 2694 16420 2746
rect 16444 2694 16482 2746
rect 16482 2694 16494 2746
rect 16494 2694 16500 2746
rect 16524 2694 16546 2746
rect 16546 2694 16558 2746
rect 16558 2694 16580 2746
rect 16604 2694 16610 2746
rect 16610 2694 16622 2746
rect 16622 2694 16660 2746
rect 16684 2694 16686 2746
rect 16686 2694 16738 2746
rect 16738 2694 16740 2746
rect 16364 2692 16420 2694
rect 16444 2692 16500 2694
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16210 1808 16266 1864
rect 16364 1658 16420 1660
rect 16444 1658 16500 1660
rect 16524 1658 16580 1660
rect 16604 1658 16660 1660
rect 16684 1658 16740 1660
rect 16364 1606 16366 1658
rect 16366 1606 16418 1658
rect 16418 1606 16420 1658
rect 16444 1606 16482 1658
rect 16482 1606 16494 1658
rect 16494 1606 16500 1658
rect 16524 1606 16546 1658
rect 16546 1606 16558 1658
rect 16558 1606 16580 1658
rect 16604 1606 16610 1658
rect 16610 1606 16622 1658
rect 16622 1606 16660 1658
rect 16684 1606 16686 1658
rect 16686 1606 16738 1658
rect 16738 1606 16740 1658
rect 16364 1604 16420 1606
rect 16444 1604 16500 1606
rect 16524 1604 16580 1606
rect 16604 1604 16660 1606
rect 16684 1604 16740 1606
rect 16364 570 16420 572
rect 16444 570 16500 572
rect 16524 570 16580 572
rect 16604 570 16660 572
rect 16684 570 16740 572
rect 16364 518 16366 570
rect 16366 518 16418 570
rect 16418 518 16420 570
rect 16444 518 16482 570
rect 16482 518 16494 570
rect 16494 518 16500 570
rect 16524 518 16546 570
rect 16546 518 16558 570
rect 16558 518 16580 570
rect 16604 518 16610 570
rect 16610 518 16622 570
rect 16622 518 16660 570
rect 16684 518 16686 570
rect 16686 518 16738 570
rect 16738 518 16740 570
rect 16364 516 16420 518
rect 16444 516 16500 518
rect 16524 516 16580 518
rect 16604 516 16660 518
rect 16684 516 16740 518
<< metal3 >>
rect 1354 17440 1750 17441
rect 1354 17376 1360 17440
rect 1424 17376 1440 17440
rect 1504 17376 1520 17440
rect 1584 17376 1600 17440
rect 1664 17376 1680 17440
rect 1744 17376 1750 17440
rect 1354 17375 1750 17376
rect 7354 17440 7750 17441
rect 7354 17376 7360 17440
rect 7424 17376 7440 17440
rect 7504 17376 7520 17440
rect 7584 17376 7600 17440
rect 7664 17376 7680 17440
rect 7744 17376 7750 17440
rect 7354 17375 7750 17376
rect 13354 17440 13750 17441
rect 13354 17376 13360 17440
rect 13424 17376 13440 17440
rect 13504 17376 13520 17440
rect 13584 17376 13600 17440
rect 13664 17376 13680 17440
rect 13744 17376 13750 17440
rect 13354 17375 13750 17376
rect 4354 16896 4750 16897
rect 4354 16832 4360 16896
rect 4424 16832 4440 16896
rect 4504 16832 4520 16896
rect 4584 16832 4600 16896
rect 4664 16832 4680 16896
rect 4744 16832 4750 16896
rect 4354 16831 4750 16832
rect 10354 16896 10750 16897
rect 10354 16832 10360 16896
rect 10424 16832 10440 16896
rect 10504 16832 10520 16896
rect 10584 16832 10600 16896
rect 10664 16832 10680 16896
rect 10744 16832 10750 16896
rect 10354 16831 10750 16832
rect 16354 16896 16750 16897
rect 16354 16832 16360 16896
rect 16424 16832 16440 16896
rect 16504 16832 16520 16896
rect 16584 16832 16600 16896
rect 16664 16832 16680 16896
rect 16744 16832 16750 16896
rect 16354 16831 16750 16832
rect 4889 16690 4955 16693
rect 6494 16690 6500 16692
rect 4889 16688 6500 16690
rect 4889 16632 4894 16688
rect 4950 16632 6500 16688
rect 4889 16630 6500 16632
rect 4889 16627 4955 16630
rect 6494 16628 6500 16630
rect 6564 16628 6570 16692
rect 8702 16628 8708 16692
rect 8772 16690 8778 16692
rect 9029 16690 9095 16693
rect 8772 16688 9095 16690
rect 8772 16632 9034 16688
rect 9090 16632 9095 16688
rect 8772 16630 9095 16632
rect 8772 16628 8778 16630
rect 9029 16627 9095 16630
rect 6453 16554 6519 16557
rect 7373 16554 7439 16557
rect 6453 16552 7439 16554
rect 6453 16496 6458 16552
rect 6514 16496 7378 16552
rect 7434 16496 7439 16552
rect 6453 16494 7439 16496
rect 6453 16491 6519 16494
rect 7373 16491 7439 16494
rect 1354 16352 1750 16353
rect 1354 16288 1360 16352
rect 1424 16288 1440 16352
rect 1504 16288 1520 16352
rect 1584 16288 1600 16352
rect 1664 16288 1680 16352
rect 1744 16288 1750 16352
rect 1354 16287 1750 16288
rect 7354 16352 7750 16353
rect 7354 16288 7360 16352
rect 7424 16288 7440 16352
rect 7504 16288 7520 16352
rect 7584 16288 7600 16352
rect 7664 16288 7680 16352
rect 7744 16288 7750 16352
rect 7354 16287 7750 16288
rect 13354 16352 13750 16353
rect 13354 16288 13360 16352
rect 13424 16288 13440 16352
rect 13504 16288 13520 16352
rect 13584 16288 13600 16352
rect 13664 16288 13680 16352
rect 13744 16288 13750 16352
rect 13354 16287 13750 16288
rect 4354 15808 4750 15809
rect 4354 15744 4360 15808
rect 4424 15744 4440 15808
rect 4504 15744 4520 15808
rect 4584 15744 4600 15808
rect 4664 15744 4680 15808
rect 4744 15744 4750 15808
rect 4354 15743 4750 15744
rect 10354 15808 10750 15809
rect 10354 15744 10360 15808
rect 10424 15744 10440 15808
rect 10504 15744 10520 15808
rect 10584 15744 10600 15808
rect 10664 15744 10680 15808
rect 10744 15744 10750 15808
rect 10354 15743 10750 15744
rect 16354 15808 16750 15809
rect 16354 15744 16360 15808
rect 16424 15744 16440 15808
rect 16504 15744 16520 15808
rect 16584 15744 16600 15808
rect 16664 15744 16680 15808
rect 16744 15744 16750 15808
rect 16354 15743 16750 15744
rect 2037 15738 2103 15741
rect 3233 15738 3299 15741
rect 2037 15736 3299 15738
rect 2037 15680 2042 15736
rect 2098 15680 3238 15736
rect 3294 15680 3299 15736
rect 2037 15678 3299 15680
rect 2037 15675 2103 15678
rect 3233 15675 3299 15678
rect 11329 15602 11395 15605
rect 13261 15602 13327 15605
rect 11329 15600 13327 15602
rect 11329 15544 11334 15600
rect 11390 15544 13266 15600
rect 13322 15544 13327 15600
rect 11329 15542 13327 15544
rect 11329 15539 11395 15542
rect 13261 15539 13327 15542
rect 6545 15466 6611 15469
rect 9254 15466 9260 15468
rect 6545 15464 9260 15466
rect 6545 15408 6550 15464
rect 6606 15408 9260 15464
rect 6545 15406 9260 15408
rect 6545 15403 6611 15406
rect 9254 15404 9260 15406
rect 9324 15404 9330 15468
rect 11513 15466 11579 15469
rect 12985 15466 13051 15469
rect 11513 15464 13051 15466
rect 11513 15408 11518 15464
rect 11574 15408 12990 15464
rect 13046 15408 13051 15464
rect 11513 15406 13051 15408
rect 11513 15403 11579 15406
rect 12985 15403 13051 15406
rect 6126 15268 6132 15332
rect 6196 15330 6202 15332
rect 7097 15330 7163 15333
rect 6196 15328 7163 15330
rect 6196 15272 7102 15328
rect 7158 15272 7163 15328
rect 6196 15270 7163 15272
rect 6196 15268 6202 15270
rect 7097 15267 7163 15270
rect 11278 15268 11284 15332
rect 11348 15330 11354 15332
rect 12249 15330 12315 15333
rect 11348 15328 12315 15330
rect 11348 15272 12254 15328
rect 12310 15272 12315 15328
rect 11348 15270 12315 15272
rect 11348 15268 11354 15270
rect 12249 15267 12315 15270
rect 12893 15330 12959 15333
rect 13118 15330 13124 15332
rect 12893 15328 13124 15330
rect 12893 15272 12898 15328
rect 12954 15272 13124 15328
rect 12893 15270 13124 15272
rect 12893 15267 12959 15270
rect 13118 15268 13124 15270
rect 13188 15268 13194 15332
rect 1354 15264 1750 15265
rect 1354 15200 1360 15264
rect 1424 15200 1440 15264
rect 1504 15200 1520 15264
rect 1584 15200 1600 15264
rect 1664 15200 1680 15264
rect 1744 15200 1750 15264
rect 1354 15199 1750 15200
rect 7354 15264 7750 15265
rect 7354 15200 7360 15264
rect 7424 15200 7440 15264
rect 7504 15200 7520 15264
rect 7584 15200 7600 15264
rect 7664 15200 7680 15264
rect 7744 15200 7750 15264
rect 7354 15199 7750 15200
rect 13354 15264 13750 15265
rect 13354 15200 13360 15264
rect 13424 15200 13440 15264
rect 13504 15200 13520 15264
rect 13584 15200 13600 15264
rect 13664 15200 13680 15264
rect 13744 15200 13750 15264
rect 13354 15199 13750 15200
rect 5073 15058 5139 15061
rect 6269 15058 6335 15061
rect 5073 15056 6335 15058
rect 5073 15000 5078 15056
rect 5134 15000 6274 15056
rect 6330 15000 6335 15056
rect 5073 14998 6335 15000
rect 5073 14995 5139 14998
rect 6269 14995 6335 14998
rect 7097 15058 7163 15061
rect 9305 15058 9371 15061
rect 13905 15058 13971 15061
rect 7097 15056 13971 15058
rect 7097 15000 7102 15056
rect 7158 15000 9310 15056
rect 9366 15000 13910 15056
rect 13966 15000 13971 15056
rect 7097 14998 13971 15000
rect 7097 14995 7163 14998
rect 9305 14995 9371 14998
rect 13905 14995 13971 14998
rect 2681 14922 2747 14925
rect 4889 14922 4955 14925
rect 2681 14920 4955 14922
rect 2681 14864 2686 14920
rect 2742 14864 4894 14920
rect 4950 14864 4955 14920
rect 2681 14862 4955 14864
rect 2681 14859 2747 14862
rect 4889 14859 4955 14862
rect 6361 14922 6427 14925
rect 7741 14922 7807 14925
rect 8385 14922 8451 14925
rect 6361 14920 8451 14922
rect 6361 14864 6366 14920
rect 6422 14864 7746 14920
rect 7802 14864 8390 14920
rect 8446 14864 8451 14920
rect 6361 14862 8451 14864
rect 6361 14859 6427 14862
rect 7741 14859 7807 14862
rect 8385 14859 8451 14862
rect 12617 14922 12683 14925
rect 13353 14922 13419 14925
rect 12617 14920 13419 14922
rect 12617 14864 12622 14920
rect 12678 14864 13358 14920
rect 13414 14864 13419 14920
rect 12617 14862 13419 14864
rect 12617 14859 12683 14862
rect 13353 14859 13419 14862
rect 4354 14720 4750 14721
rect 4354 14656 4360 14720
rect 4424 14656 4440 14720
rect 4504 14656 4520 14720
rect 4584 14656 4600 14720
rect 4664 14656 4680 14720
rect 4744 14656 4750 14720
rect 4354 14655 4750 14656
rect 10354 14720 10750 14721
rect 10354 14656 10360 14720
rect 10424 14656 10440 14720
rect 10504 14656 10520 14720
rect 10584 14656 10600 14720
rect 10664 14656 10680 14720
rect 10744 14656 10750 14720
rect 10354 14655 10750 14656
rect 16354 14720 16750 14721
rect 16354 14656 16360 14720
rect 16424 14656 16440 14720
rect 16504 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16750 14720
rect 16354 14655 16750 14656
rect 4061 14514 4127 14517
rect 4521 14514 4587 14517
rect 10501 14514 10567 14517
rect 4061 14512 4587 14514
rect 4061 14456 4066 14512
rect 4122 14456 4526 14512
rect 4582 14456 4587 14512
rect 4061 14454 4587 14456
rect 4061 14451 4127 14454
rect 4521 14451 4587 14454
rect 7054 14512 10567 14514
rect 7054 14456 10506 14512
rect 10562 14456 10567 14512
rect 7054 14454 10567 14456
rect 2681 14378 2747 14381
rect 7054 14378 7114 14454
rect 10501 14451 10567 14454
rect 11973 14514 12039 14517
rect 16941 14514 17007 14517
rect 11973 14512 17007 14514
rect 11973 14456 11978 14512
rect 12034 14456 16946 14512
rect 17002 14456 17007 14512
rect 11973 14454 17007 14456
rect 11973 14451 12039 14454
rect 16941 14451 17007 14454
rect 2681 14376 7114 14378
rect 2681 14320 2686 14376
rect 2742 14320 7114 14376
rect 2681 14318 7114 14320
rect 7281 14378 7347 14381
rect 10593 14378 10659 14381
rect 7281 14376 10659 14378
rect 7281 14320 7286 14376
rect 7342 14320 10598 14376
rect 10654 14320 10659 14376
rect 7281 14318 10659 14320
rect 2681 14315 2747 14318
rect 7281 14315 7347 14318
rect 10593 14315 10659 14318
rect 12157 14378 12223 14381
rect 15745 14378 15811 14381
rect 12157 14376 15811 14378
rect 12157 14320 12162 14376
rect 12218 14320 15750 14376
rect 15806 14320 15811 14376
rect 12157 14318 15811 14320
rect 12157 14315 12223 14318
rect 15745 14315 15811 14318
rect 8385 14242 8451 14245
rect 8661 14242 8727 14245
rect 8385 14240 8727 14242
rect 8385 14184 8390 14240
rect 8446 14184 8666 14240
rect 8722 14184 8727 14240
rect 8385 14182 8727 14184
rect 8385 14179 8451 14182
rect 8661 14179 8727 14182
rect 1354 14176 1750 14177
rect 1354 14112 1360 14176
rect 1424 14112 1440 14176
rect 1504 14112 1520 14176
rect 1584 14112 1600 14176
rect 1664 14112 1680 14176
rect 1744 14112 1750 14176
rect 1354 14111 1750 14112
rect 7354 14176 7750 14177
rect 7354 14112 7360 14176
rect 7424 14112 7440 14176
rect 7504 14112 7520 14176
rect 7584 14112 7600 14176
rect 7664 14112 7680 14176
rect 7744 14112 7750 14176
rect 7354 14111 7750 14112
rect 13354 14176 13750 14177
rect 13354 14112 13360 14176
rect 13424 14112 13440 14176
rect 13504 14112 13520 14176
rect 13584 14112 13600 14176
rect 13664 14112 13680 14176
rect 13744 14112 13750 14176
rect 13354 14111 13750 14112
rect 4613 14106 4679 14109
rect 7833 14106 7899 14109
rect 12065 14106 12131 14109
rect 4613 14104 6378 14106
rect 4613 14048 4618 14104
rect 4674 14048 6378 14104
rect 4613 14046 6378 14048
rect 4613 14043 4679 14046
rect 3509 13970 3575 13973
rect 4337 13970 4403 13973
rect 6177 13970 6243 13973
rect 3509 13968 6243 13970
rect 3509 13912 3514 13968
rect 3570 13912 4342 13968
rect 4398 13912 6182 13968
rect 6238 13912 6243 13968
rect 3509 13910 6243 13912
rect 6318 13970 6378 14046
rect 7833 14104 12131 14106
rect 7833 14048 7838 14104
rect 7894 14048 12070 14104
rect 12126 14048 12131 14104
rect 7833 14046 12131 14048
rect 7833 14043 7899 14046
rect 12065 14043 12131 14046
rect 7465 13970 7531 13973
rect 6318 13968 7531 13970
rect 6318 13912 7470 13968
rect 7526 13912 7531 13968
rect 6318 13910 7531 13912
rect 3509 13907 3575 13910
rect 4337 13907 4403 13910
rect 6177 13907 6243 13910
rect 7465 13907 7531 13910
rect 7649 13970 7715 13973
rect 11145 13970 11211 13973
rect 7649 13968 11211 13970
rect 7649 13912 7654 13968
rect 7710 13912 11150 13968
rect 11206 13912 11211 13968
rect 7649 13910 11211 13912
rect 7649 13907 7715 13910
rect 11145 13907 11211 13910
rect 5257 13834 5323 13837
rect 12525 13834 12591 13837
rect 5257 13832 12591 13834
rect 5257 13776 5262 13832
rect 5318 13776 12530 13832
rect 12586 13776 12591 13832
rect 5257 13774 12591 13776
rect 5257 13771 5323 13774
rect 12525 13771 12591 13774
rect 5993 13698 6059 13701
rect 9673 13698 9739 13701
rect 5993 13696 9739 13698
rect 5993 13640 5998 13696
rect 6054 13640 9678 13696
rect 9734 13640 9739 13696
rect 5993 13638 9739 13640
rect 5993 13635 6059 13638
rect 9673 13635 9739 13638
rect 12617 13698 12683 13701
rect 13997 13698 14063 13701
rect 16113 13698 16179 13701
rect 12617 13696 16179 13698
rect 12617 13640 12622 13696
rect 12678 13640 14002 13696
rect 14058 13640 16118 13696
rect 16174 13640 16179 13696
rect 12617 13638 16179 13640
rect 12617 13635 12683 13638
rect 13997 13635 14063 13638
rect 16113 13635 16179 13638
rect 4354 13632 4750 13633
rect 4354 13568 4360 13632
rect 4424 13568 4440 13632
rect 4504 13568 4520 13632
rect 4584 13568 4600 13632
rect 4664 13568 4680 13632
rect 4744 13568 4750 13632
rect 4354 13567 4750 13568
rect 10354 13632 10750 13633
rect 10354 13568 10360 13632
rect 10424 13568 10440 13632
rect 10504 13568 10520 13632
rect 10584 13568 10600 13632
rect 10664 13568 10680 13632
rect 10744 13568 10750 13632
rect 10354 13567 10750 13568
rect 16354 13632 16750 13633
rect 16354 13568 16360 13632
rect 16424 13568 16440 13632
rect 16504 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16750 13632
rect 16354 13567 16750 13568
rect 6361 13562 6427 13565
rect 9581 13562 9647 13565
rect 6361 13560 9647 13562
rect 6361 13504 6366 13560
rect 6422 13504 9586 13560
rect 9642 13504 9647 13560
rect 6361 13502 9647 13504
rect 6361 13499 6427 13502
rect 9581 13499 9647 13502
rect 4061 13426 4127 13429
rect 6085 13426 6151 13429
rect 8661 13426 8727 13429
rect 4061 13424 8727 13426
rect 4061 13368 4066 13424
rect 4122 13368 6090 13424
rect 6146 13368 8666 13424
rect 8722 13368 8727 13424
rect 4061 13366 8727 13368
rect 4061 13363 4127 13366
rect 6085 13363 6151 13366
rect 8661 13363 8727 13366
rect 10041 13426 10107 13429
rect 11881 13426 11947 13429
rect 10041 13424 11947 13426
rect 10041 13368 10046 13424
rect 10102 13368 11886 13424
rect 11942 13368 11947 13424
rect 10041 13366 11947 13368
rect 10041 13363 10107 13366
rect 11881 13363 11947 13366
rect 6913 13290 6979 13293
rect 10317 13290 10383 13293
rect 6913 13288 10383 13290
rect 6913 13232 6918 13288
rect 6974 13232 10322 13288
rect 10378 13232 10383 13288
rect 6913 13230 10383 13232
rect 6913 13227 6979 13230
rect 10317 13227 10383 13230
rect 8661 13154 8727 13157
rect 9121 13154 9187 13157
rect 8661 13152 9187 13154
rect 8661 13096 8666 13152
rect 8722 13096 9126 13152
rect 9182 13096 9187 13152
rect 8661 13094 9187 13096
rect 8661 13091 8727 13094
rect 9121 13091 9187 13094
rect 1354 13088 1750 13089
rect 1354 13024 1360 13088
rect 1424 13024 1440 13088
rect 1504 13024 1520 13088
rect 1584 13024 1600 13088
rect 1664 13024 1680 13088
rect 1744 13024 1750 13088
rect 1354 13023 1750 13024
rect 7354 13088 7750 13089
rect 7354 13024 7360 13088
rect 7424 13024 7440 13088
rect 7504 13024 7520 13088
rect 7584 13024 7600 13088
rect 7664 13024 7680 13088
rect 7744 13024 7750 13088
rect 7354 13023 7750 13024
rect 13354 13088 13750 13089
rect 13354 13024 13360 13088
rect 13424 13024 13440 13088
rect 13504 13024 13520 13088
rect 13584 13024 13600 13088
rect 13664 13024 13680 13088
rect 13744 13024 13750 13088
rect 13354 13023 13750 13024
rect 2865 12882 2931 12885
rect 12525 12882 12591 12885
rect 2865 12880 12591 12882
rect 2865 12824 2870 12880
rect 2926 12824 12530 12880
rect 12586 12824 12591 12880
rect 2865 12822 12591 12824
rect 2865 12819 2931 12822
rect 12525 12819 12591 12822
rect 2681 12746 2747 12749
rect 6361 12746 6427 12749
rect 8661 12746 8727 12749
rect 2681 12744 8727 12746
rect 2681 12688 2686 12744
rect 2742 12688 6366 12744
rect 6422 12688 8666 12744
rect 8722 12688 8727 12744
rect 2681 12686 8727 12688
rect 2681 12683 2747 12686
rect 6361 12683 6427 12686
rect 8661 12683 8727 12686
rect 10961 12746 11027 12749
rect 14038 12746 14044 12748
rect 10961 12744 14044 12746
rect 10961 12688 10966 12744
rect 11022 12688 14044 12744
rect 10961 12686 14044 12688
rect 10961 12683 11027 12686
rect 14038 12684 14044 12686
rect 14108 12684 14114 12748
rect 7925 12610 7991 12613
rect 8886 12610 8892 12612
rect 7925 12608 8892 12610
rect 7925 12552 7930 12608
rect 7986 12552 8892 12608
rect 7925 12550 8892 12552
rect 7925 12547 7991 12550
rect 8886 12548 8892 12550
rect 8956 12548 8962 12612
rect 4354 12544 4750 12545
rect 4354 12480 4360 12544
rect 4424 12480 4440 12544
rect 4504 12480 4520 12544
rect 4584 12480 4600 12544
rect 4664 12480 4680 12544
rect 4744 12480 4750 12544
rect 4354 12479 4750 12480
rect 10354 12544 10750 12545
rect 10354 12480 10360 12544
rect 10424 12480 10440 12544
rect 10504 12480 10520 12544
rect 10584 12480 10600 12544
rect 10664 12480 10680 12544
rect 10744 12480 10750 12544
rect 10354 12479 10750 12480
rect 16354 12544 16750 12545
rect 16354 12480 16360 12544
rect 16424 12480 16440 12544
rect 16504 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16750 12544
rect 16354 12479 16750 12480
rect 6269 12474 6335 12477
rect 7925 12474 7991 12477
rect 6269 12472 7991 12474
rect 6269 12416 6274 12472
rect 6330 12416 7930 12472
rect 7986 12416 7991 12472
rect 6269 12414 7991 12416
rect 6269 12411 6335 12414
rect 7925 12411 7991 12414
rect 8293 12066 8359 12069
rect 9305 12066 9371 12069
rect 8293 12064 9371 12066
rect 8293 12008 8298 12064
rect 8354 12008 9310 12064
rect 9366 12008 9371 12064
rect 8293 12006 9371 12008
rect 8293 12003 8359 12006
rect 9305 12003 9371 12006
rect 1354 12000 1750 12001
rect 1354 11936 1360 12000
rect 1424 11936 1440 12000
rect 1504 11936 1520 12000
rect 1584 11936 1600 12000
rect 1664 11936 1680 12000
rect 1744 11936 1750 12000
rect 1354 11935 1750 11936
rect 7354 12000 7750 12001
rect 7354 11936 7360 12000
rect 7424 11936 7440 12000
rect 7504 11936 7520 12000
rect 7584 11936 7600 12000
rect 7664 11936 7680 12000
rect 7744 11936 7750 12000
rect 7354 11935 7750 11936
rect 13354 12000 13750 12001
rect 13354 11936 13360 12000
rect 13424 11936 13440 12000
rect 13504 11936 13520 12000
rect 13584 11936 13600 12000
rect 13664 11936 13680 12000
rect 13744 11936 13750 12000
rect 13354 11935 13750 11936
rect 6913 11794 6979 11797
rect 7281 11794 7347 11797
rect 6913 11792 7347 11794
rect 6913 11736 6918 11792
rect 6974 11736 7286 11792
rect 7342 11736 7347 11792
rect 6913 11734 7347 11736
rect 6913 11731 6979 11734
rect 7281 11731 7347 11734
rect 7649 11794 7715 11797
rect 9397 11794 9463 11797
rect 7649 11792 9463 11794
rect 7649 11736 7654 11792
rect 7710 11736 9402 11792
rect 9458 11736 9463 11792
rect 7649 11734 9463 11736
rect 7649 11731 7715 11734
rect 9397 11731 9463 11734
rect 12617 11794 12683 11797
rect 12750 11794 12756 11796
rect 12617 11792 12756 11794
rect 12617 11736 12622 11792
rect 12678 11736 12756 11792
rect 12617 11734 12756 11736
rect 12617 11731 12683 11734
rect 12750 11732 12756 11734
rect 12820 11732 12826 11796
rect 14365 11658 14431 11661
rect 8526 11656 14431 11658
rect 8526 11600 14370 11656
rect 14426 11600 14431 11656
rect 8526 11598 14431 11600
rect 6085 11522 6151 11525
rect 8526 11522 8586 11598
rect 14365 11595 14431 11598
rect 6085 11520 8586 11522
rect 6085 11464 6090 11520
rect 6146 11464 8586 11520
rect 6085 11462 8586 11464
rect 6085 11459 6151 11462
rect 4354 11456 4750 11457
rect 4354 11392 4360 11456
rect 4424 11392 4440 11456
rect 4504 11392 4520 11456
rect 4584 11392 4600 11456
rect 4664 11392 4680 11456
rect 4744 11392 4750 11456
rect 4354 11391 4750 11392
rect 10354 11456 10750 11457
rect 10354 11392 10360 11456
rect 10424 11392 10440 11456
rect 10504 11392 10520 11456
rect 10584 11392 10600 11456
rect 10664 11392 10680 11456
rect 10744 11392 10750 11456
rect 10354 11391 10750 11392
rect 16354 11456 16750 11457
rect 16354 11392 16360 11456
rect 16424 11392 16440 11456
rect 16504 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16750 11456
rect 16354 11391 16750 11392
rect 5809 11250 5875 11253
rect 8017 11250 8083 11253
rect 5809 11248 8083 11250
rect 5809 11192 5814 11248
rect 5870 11192 8022 11248
rect 8078 11192 8083 11248
rect 5809 11190 8083 11192
rect 5809 11187 5875 11190
rect 8017 11187 8083 11190
rect 9765 11250 9831 11253
rect 14273 11250 14339 11253
rect 9765 11248 14339 11250
rect 9765 11192 9770 11248
rect 9826 11192 14278 11248
rect 14334 11192 14339 11248
rect 9765 11190 14339 11192
rect 9765 11187 9831 11190
rect 14273 11187 14339 11190
rect 5073 11114 5139 11117
rect 6729 11114 6795 11117
rect 12249 11116 12315 11117
rect 12198 11114 12204 11116
rect 5073 11112 8172 11114
rect 5073 11056 5078 11112
rect 5134 11056 6734 11112
rect 6790 11056 8172 11112
rect 5073 11054 8172 11056
rect 12158 11054 12204 11114
rect 12268 11112 12315 11116
rect 12310 11056 12315 11112
rect 5073 11051 5139 11054
rect 6729 11051 6795 11054
rect 8112 10981 8172 11054
rect 12198 11052 12204 11054
rect 12268 11052 12315 11056
rect 12249 11051 12315 11052
rect 13629 11114 13695 11117
rect 16573 11114 16639 11117
rect 13629 11112 16639 11114
rect 13629 11056 13634 11112
rect 13690 11056 16578 11112
rect 16634 11056 16639 11112
rect 13629 11054 16639 11056
rect 13629 11051 13695 11054
rect 16573 11051 16639 11054
rect 3877 10978 3943 10981
rect 5533 10978 5599 10981
rect 3877 10976 5599 10978
rect 3877 10920 3882 10976
rect 3938 10920 5538 10976
rect 5594 10920 5599 10976
rect 3877 10918 5599 10920
rect 3877 10915 3943 10918
rect 5533 10915 5599 10918
rect 8109 10976 8175 10981
rect 8109 10920 8114 10976
rect 8170 10920 8175 10976
rect 8109 10915 8175 10920
rect 8886 10916 8892 10980
rect 8956 10978 8962 10980
rect 9029 10978 9095 10981
rect 8956 10976 9095 10978
rect 8956 10920 9034 10976
rect 9090 10920 9095 10976
rect 8956 10918 9095 10920
rect 8956 10916 8962 10918
rect 9029 10915 9095 10918
rect 1354 10912 1750 10913
rect 1354 10848 1360 10912
rect 1424 10848 1440 10912
rect 1504 10848 1520 10912
rect 1584 10848 1600 10912
rect 1664 10848 1680 10912
rect 1744 10848 1750 10912
rect 1354 10847 1750 10848
rect 7354 10912 7750 10913
rect 7354 10848 7360 10912
rect 7424 10848 7440 10912
rect 7504 10848 7520 10912
rect 7584 10848 7600 10912
rect 7664 10848 7680 10912
rect 7744 10848 7750 10912
rect 7354 10847 7750 10848
rect 13354 10912 13750 10913
rect 13354 10848 13360 10912
rect 13424 10848 13440 10912
rect 13504 10848 13520 10912
rect 13584 10848 13600 10912
rect 13664 10848 13680 10912
rect 13744 10848 13750 10912
rect 13354 10847 13750 10848
rect 4061 10842 4127 10845
rect 7005 10842 7071 10845
rect 4061 10840 7071 10842
rect 4061 10784 4066 10840
rect 4122 10784 7010 10840
rect 7066 10784 7071 10840
rect 4061 10782 7071 10784
rect 4061 10779 4127 10782
rect 7005 10779 7071 10782
rect 5257 10706 5323 10709
rect 6361 10706 6427 10709
rect 13353 10706 13419 10709
rect 5257 10704 5872 10706
rect 5257 10648 5262 10704
rect 5318 10648 5872 10704
rect 5257 10646 5872 10648
rect 5257 10643 5323 10646
rect 4613 10570 4679 10573
rect 5812 10570 5872 10646
rect 6361 10704 13419 10706
rect 6361 10648 6366 10704
rect 6422 10648 13358 10704
rect 13414 10648 13419 10704
rect 6361 10646 13419 10648
rect 6361 10643 6427 10646
rect 13353 10643 13419 10646
rect 12341 10570 12407 10573
rect 4613 10568 4906 10570
rect 4613 10512 4618 10568
rect 4674 10512 4906 10568
rect 4613 10510 4906 10512
rect 5812 10568 12407 10570
rect 5812 10512 12346 10568
rect 12402 10512 12407 10568
rect 5812 10510 12407 10512
rect 4613 10507 4679 10510
rect 4354 10368 4750 10369
rect 4354 10304 4360 10368
rect 4424 10304 4440 10368
rect 4504 10304 4520 10368
rect 4584 10304 4600 10368
rect 4664 10304 4680 10368
rect 4744 10304 4750 10368
rect 4354 10303 4750 10304
rect 4337 10162 4403 10165
rect 4846 10162 4906 10510
rect 12341 10507 12407 10510
rect 6177 10434 6243 10437
rect 8477 10434 8543 10437
rect 6177 10432 8543 10434
rect 6177 10376 6182 10432
rect 6238 10376 8482 10432
rect 8538 10376 8543 10432
rect 6177 10374 8543 10376
rect 6177 10371 6243 10374
rect 8477 10371 8543 10374
rect 9673 10432 9739 10437
rect 9673 10376 9678 10432
rect 9734 10376 9739 10432
rect 9673 10371 9739 10376
rect 9676 10165 9736 10371
rect 10354 10368 10750 10369
rect 10354 10304 10360 10368
rect 10424 10304 10440 10368
rect 10504 10304 10520 10368
rect 10584 10304 10600 10368
rect 10664 10304 10680 10368
rect 10744 10304 10750 10368
rect 10354 10303 10750 10304
rect 16354 10368 16750 10369
rect 16354 10304 16360 10368
rect 16424 10304 16440 10368
rect 16504 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16750 10368
rect 16354 10303 16750 10304
rect 4337 10160 4906 10162
rect 4337 10104 4342 10160
rect 4398 10104 4906 10160
rect 4337 10102 4906 10104
rect 9673 10160 9739 10165
rect 9673 10104 9678 10160
rect 9734 10104 9739 10160
rect 4337 10099 4403 10102
rect 9673 10099 9739 10104
rect 3785 10026 3851 10029
rect 4613 10026 4679 10029
rect 3785 10024 4679 10026
rect 3785 9968 3790 10024
rect 3846 9968 4618 10024
rect 4674 9968 4679 10024
rect 3785 9966 4679 9968
rect 3785 9963 3851 9966
rect 4613 9963 4679 9966
rect 6821 10026 6887 10029
rect 7649 10026 7715 10029
rect 6821 10024 7715 10026
rect 6821 9968 6826 10024
rect 6882 9968 7654 10024
rect 7710 9968 7715 10024
rect 6821 9966 7715 9968
rect 6821 9963 6887 9966
rect 7649 9963 7715 9966
rect 3693 9890 3759 9893
rect 4521 9890 4587 9893
rect 3693 9888 4587 9890
rect 3693 9832 3698 9888
rect 3754 9832 4526 9888
rect 4582 9832 4587 9888
rect 3693 9830 4587 9832
rect 3693 9827 3759 9830
rect 4521 9827 4587 9830
rect 1354 9824 1750 9825
rect 1354 9760 1360 9824
rect 1424 9760 1440 9824
rect 1504 9760 1520 9824
rect 1584 9760 1600 9824
rect 1664 9760 1680 9824
rect 1744 9760 1750 9824
rect 1354 9759 1750 9760
rect 7354 9824 7750 9825
rect 7354 9760 7360 9824
rect 7424 9760 7440 9824
rect 7504 9760 7520 9824
rect 7584 9760 7600 9824
rect 7664 9760 7680 9824
rect 7744 9760 7750 9824
rect 7354 9759 7750 9760
rect 13354 9824 13750 9825
rect 13354 9760 13360 9824
rect 13424 9760 13440 9824
rect 13504 9760 13520 9824
rect 13584 9760 13600 9824
rect 13664 9760 13680 9824
rect 13744 9760 13750 9824
rect 13354 9759 13750 9760
rect 3509 9618 3575 9621
rect 8109 9618 8175 9621
rect 3509 9616 8175 9618
rect 3509 9560 3514 9616
rect 3570 9560 8114 9616
rect 8170 9560 8175 9616
rect 3509 9558 8175 9560
rect 3509 9555 3575 9558
rect 8109 9555 8175 9558
rect 10225 9618 10291 9621
rect 12801 9618 12867 9621
rect 16205 9618 16271 9621
rect 10225 9616 16271 9618
rect 10225 9560 10230 9616
rect 10286 9560 12806 9616
rect 12862 9560 16210 9616
rect 16266 9560 16271 9616
rect 10225 9558 16271 9560
rect 10225 9555 10291 9558
rect 12801 9555 12867 9558
rect 16205 9555 16271 9558
rect 4354 9280 4750 9281
rect 4354 9216 4360 9280
rect 4424 9216 4440 9280
rect 4504 9216 4520 9280
rect 4584 9216 4600 9280
rect 4664 9216 4680 9280
rect 4744 9216 4750 9280
rect 4354 9215 4750 9216
rect 10354 9280 10750 9281
rect 10354 9216 10360 9280
rect 10424 9216 10440 9280
rect 10504 9216 10520 9280
rect 10584 9216 10600 9280
rect 10664 9216 10680 9280
rect 10744 9216 10750 9280
rect 10354 9215 10750 9216
rect 16354 9280 16750 9281
rect 16354 9216 16360 9280
rect 16424 9216 16440 9280
rect 16504 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16750 9280
rect 16354 9215 16750 9216
rect 2589 9074 2655 9077
rect 8937 9074 9003 9077
rect 2589 9072 9003 9074
rect 2589 9016 2594 9072
rect 2650 9016 8942 9072
rect 8998 9016 9003 9072
rect 2589 9014 9003 9016
rect 2589 9011 2655 9014
rect 8937 9011 9003 9014
rect 9765 9074 9831 9077
rect 10225 9074 10291 9077
rect 9765 9072 10291 9074
rect 9765 9016 9770 9072
rect 9826 9016 10230 9072
rect 10286 9016 10291 9072
rect 9765 9014 10291 9016
rect 9765 9011 9831 9014
rect 10225 9011 10291 9014
rect 12433 9074 12499 9077
rect 15745 9074 15811 9077
rect 12433 9072 15811 9074
rect 12433 9016 12438 9072
rect 12494 9016 15750 9072
rect 15806 9016 15811 9072
rect 12433 9014 15811 9016
rect 12433 9011 12499 9014
rect 15745 9011 15811 9014
rect 1853 8938 1919 8941
rect 6453 8938 6519 8941
rect 1853 8936 6519 8938
rect 1853 8880 1858 8936
rect 1914 8880 6458 8936
rect 6514 8880 6519 8936
rect 1853 8878 6519 8880
rect 1853 8875 1919 8878
rect 6453 8875 6519 8878
rect 10777 8938 10843 8941
rect 13169 8938 13235 8941
rect 10777 8936 13235 8938
rect 10777 8880 10782 8936
rect 10838 8880 13174 8936
rect 13230 8880 13235 8936
rect 10777 8878 13235 8880
rect 10777 8875 10843 8878
rect 13169 8875 13235 8878
rect 1354 8736 1750 8737
rect 1354 8672 1360 8736
rect 1424 8672 1440 8736
rect 1504 8672 1520 8736
rect 1584 8672 1600 8736
rect 1664 8672 1680 8736
rect 1744 8672 1750 8736
rect 1354 8671 1750 8672
rect 7354 8736 7750 8737
rect 7354 8672 7360 8736
rect 7424 8672 7440 8736
rect 7504 8672 7520 8736
rect 7584 8672 7600 8736
rect 7664 8672 7680 8736
rect 7744 8672 7750 8736
rect 7354 8671 7750 8672
rect 13354 8736 13750 8737
rect 13354 8672 13360 8736
rect 13424 8672 13440 8736
rect 13504 8672 13520 8736
rect 13584 8672 13600 8736
rect 13664 8672 13680 8736
rect 13744 8672 13750 8736
rect 13354 8671 13750 8672
rect 6729 8530 6795 8533
rect 7373 8530 7439 8533
rect 6729 8528 7439 8530
rect 6729 8472 6734 8528
rect 6790 8472 7378 8528
rect 7434 8472 7439 8528
rect 6729 8470 7439 8472
rect 6729 8467 6795 8470
rect 7373 8467 7439 8470
rect 8477 8530 8543 8533
rect 14825 8530 14891 8533
rect 15745 8530 15811 8533
rect 8477 8528 15811 8530
rect 8477 8472 8482 8528
rect 8538 8472 14830 8528
rect 14886 8472 15750 8528
rect 15806 8472 15811 8528
rect 8477 8470 15811 8472
rect 8477 8467 8543 8470
rect 14825 8467 14891 8470
rect 15745 8467 15811 8470
rect 5901 8394 5967 8397
rect 7465 8394 7531 8397
rect 5901 8392 7531 8394
rect 5901 8336 5906 8392
rect 5962 8336 7470 8392
rect 7526 8336 7531 8392
rect 5901 8334 7531 8336
rect 5901 8331 5967 8334
rect 7465 8331 7531 8334
rect 10225 8394 10291 8397
rect 12617 8394 12683 8397
rect 10225 8392 12683 8394
rect 10225 8336 10230 8392
rect 10286 8336 12622 8392
rect 12678 8336 12683 8392
rect 10225 8334 12683 8336
rect 10225 8331 10291 8334
rect 12617 8331 12683 8334
rect 4354 8192 4750 8193
rect 4354 8128 4360 8192
rect 4424 8128 4440 8192
rect 4504 8128 4520 8192
rect 4584 8128 4600 8192
rect 4664 8128 4680 8192
rect 4744 8128 4750 8192
rect 4354 8127 4750 8128
rect 10354 8192 10750 8193
rect 10354 8128 10360 8192
rect 10424 8128 10440 8192
rect 10504 8128 10520 8192
rect 10584 8128 10600 8192
rect 10664 8128 10680 8192
rect 10744 8128 10750 8192
rect 10354 8127 10750 8128
rect 16354 8192 16750 8193
rect 16354 8128 16360 8192
rect 16424 8128 16440 8192
rect 16504 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16750 8192
rect 16354 8127 16750 8128
rect 2129 7850 2195 7853
rect 8477 7850 8543 7853
rect 2129 7848 8543 7850
rect 2129 7792 2134 7848
rect 2190 7792 8482 7848
rect 8538 7792 8543 7848
rect 2129 7790 8543 7792
rect 2129 7787 2195 7790
rect 8477 7787 8543 7790
rect 1354 7648 1750 7649
rect 1354 7584 1360 7648
rect 1424 7584 1440 7648
rect 1504 7584 1520 7648
rect 1584 7584 1600 7648
rect 1664 7584 1680 7648
rect 1744 7584 1750 7648
rect 1354 7583 1750 7584
rect 7354 7648 7750 7649
rect 7354 7584 7360 7648
rect 7424 7584 7440 7648
rect 7504 7584 7520 7648
rect 7584 7584 7600 7648
rect 7664 7584 7680 7648
rect 7744 7584 7750 7648
rect 7354 7583 7750 7584
rect 13354 7648 13750 7649
rect 13354 7584 13360 7648
rect 13424 7584 13440 7648
rect 13504 7584 13520 7648
rect 13584 7584 13600 7648
rect 13664 7584 13680 7648
rect 13744 7584 13750 7648
rect 13354 7583 13750 7584
rect 5942 7380 5948 7444
rect 6012 7442 6018 7444
rect 9581 7442 9647 7445
rect 6012 7440 9647 7442
rect 6012 7384 9586 7440
rect 9642 7384 9647 7440
rect 6012 7382 9647 7384
rect 6012 7380 6018 7382
rect 9581 7379 9647 7382
rect 9765 7442 9831 7445
rect 12157 7442 12223 7445
rect 9765 7440 12223 7442
rect 9765 7384 9770 7440
rect 9826 7384 12162 7440
rect 12218 7384 12223 7440
rect 9765 7382 12223 7384
rect 9765 7379 9831 7382
rect 12157 7379 12223 7382
rect 14038 7380 14044 7444
rect 14108 7442 14114 7444
rect 14365 7442 14431 7445
rect 14108 7440 14431 7442
rect 14108 7384 14370 7440
rect 14426 7384 14431 7440
rect 14108 7382 14431 7384
rect 14108 7380 14114 7382
rect 14365 7379 14431 7382
rect 2865 7306 2931 7309
rect 7465 7306 7531 7309
rect 2865 7304 7531 7306
rect 2865 7248 2870 7304
rect 2926 7248 7470 7304
rect 7526 7248 7531 7304
rect 2865 7246 7531 7248
rect 2865 7243 2931 7246
rect 7465 7243 7531 7246
rect 9121 7306 9187 7309
rect 11789 7306 11855 7309
rect 9121 7304 11855 7306
rect 9121 7248 9126 7304
rect 9182 7248 11794 7304
rect 11850 7248 11855 7304
rect 9121 7246 11855 7248
rect 9121 7243 9187 7246
rect 11789 7243 11855 7246
rect 13854 7108 13860 7172
rect 13924 7170 13930 7172
rect 14181 7170 14247 7173
rect 13924 7168 14247 7170
rect 13924 7112 14186 7168
rect 14242 7112 14247 7168
rect 13924 7110 14247 7112
rect 13924 7108 13930 7110
rect 14181 7107 14247 7110
rect 4354 7104 4750 7105
rect 4354 7040 4360 7104
rect 4424 7040 4440 7104
rect 4504 7040 4520 7104
rect 4584 7040 4600 7104
rect 4664 7040 4680 7104
rect 4744 7040 4750 7104
rect 4354 7039 4750 7040
rect 10354 7104 10750 7105
rect 10354 7040 10360 7104
rect 10424 7040 10440 7104
rect 10504 7040 10520 7104
rect 10584 7040 10600 7104
rect 10664 7040 10680 7104
rect 10744 7040 10750 7104
rect 10354 7039 10750 7040
rect 16354 7104 16750 7105
rect 16354 7040 16360 7104
rect 16424 7040 16440 7104
rect 16504 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16750 7104
rect 16354 7039 16750 7040
rect 14774 6972 14780 7036
rect 14844 7034 14850 7036
rect 14917 7034 14983 7037
rect 14844 7032 14983 7034
rect 14844 6976 14922 7032
rect 14978 6976 14983 7032
rect 14844 6974 14983 6976
rect 14844 6972 14850 6974
rect 14917 6971 14983 6974
rect 7741 6762 7807 6765
rect 10409 6762 10475 6765
rect 7741 6760 10475 6762
rect 7741 6704 7746 6760
rect 7802 6704 10414 6760
rect 10470 6704 10475 6760
rect 7741 6702 10475 6704
rect 7741 6699 7807 6702
rect 10409 6699 10475 6702
rect 9806 6564 9812 6628
rect 9876 6626 9882 6628
rect 9949 6626 10015 6629
rect 9876 6624 10015 6626
rect 9876 6568 9954 6624
rect 10010 6568 10015 6624
rect 9876 6566 10015 6568
rect 9876 6564 9882 6566
rect 9949 6563 10015 6566
rect 1354 6560 1750 6561
rect 1354 6496 1360 6560
rect 1424 6496 1440 6560
rect 1504 6496 1520 6560
rect 1584 6496 1600 6560
rect 1664 6496 1680 6560
rect 1744 6496 1750 6560
rect 1354 6495 1750 6496
rect 7354 6560 7750 6561
rect 7354 6496 7360 6560
rect 7424 6496 7440 6560
rect 7504 6496 7520 6560
rect 7584 6496 7600 6560
rect 7664 6496 7680 6560
rect 7744 6496 7750 6560
rect 7354 6495 7750 6496
rect 13354 6560 13750 6561
rect 13354 6496 13360 6560
rect 13424 6496 13440 6560
rect 13504 6496 13520 6560
rect 13584 6496 13600 6560
rect 13664 6496 13680 6560
rect 13744 6496 13750 6560
rect 13354 6495 13750 6496
rect 8937 6488 9003 6493
rect 8937 6432 8942 6488
rect 8998 6432 9003 6488
rect 8937 6427 9003 6432
rect 8940 6354 9000 6427
rect 9121 6354 9187 6357
rect 8940 6352 9187 6354
rect 8940 6296 9126 6352
rect 9182 6296 9187 6352
rect 8940 6294 9187 6296
rect 9121 6291 9187 6294
rect 12801 6354 12867 6357
rect 14825 6354 14891 6357
rect 12801 6352 14891 6354
rect 12801 6296 12806 6352
rect 12862 6296 14830 6352
rect 14886 6296 14891 6352
rect 12801 6294 14891 6296
rect 12801 6291 12867 6294
rect 14825 6291 14891 6294
rect 8385 6218 8451 6221
rect 9029 6218 9095 6221
rect 8385 6216 9095 6218
rect 8385 6160 8390 6216
rect 8446 6160 9034 6216
rect 9090 6160 9095 6216
rect 8385 6158 9095 6160
rect 8385 6155 8451 6158
rect 9029 6155 9095 6158
rect 13629 6218 13695 6221
rect 13854 6218 13860 6220
rect 13629 6216 13860 6218
rect 13629 6160 13634 6216
rect 13690 6160 13860 6216
rect 13629 6158 13860 6160
rect 13629 6155 13695 6158
rect 13854 6156 13860 6158
rect 13924 6156 13930 6220
rect 11421 6082 11487 6085
rect 14181 6082 14247 6085
rect 11421 6080 14247 6082
rect 11421 6024 11426 6080
rect 11482 6024 14186 6080
rect 14242 6024 14247 6080
rect 11421 6022 14247 6024
rect 11421 6019 11487 6022
rect 14181 6019 14247 6022
rect 4354 6016 4750 6017
rect 4354 5952 4360 6016
rect 4424 5952 4440 6016
rect 4504 5952 4520 6016
rect 4584 5952 4600 6016
rect 4664 5952 4680 6016
rect 4744 5952 4750 6016
rect 4354 5951 4750 5952
rect 10354 6016 10750 6017
rect 10354 5952 10360 6016
rect 10424 5952 10440 6016
rect 10504 5952 10520 6016
rect 10584 5952 10600 6016
rect 10664 5952 10680 6016
rect 10744 5952 10750 6016
rect 10354 5951 10750 5952
rect 16354 6016 16750 6017
rect 16354 5952 16360 6016
rect 16424 5952 16440 6016
rect 16504 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16750 6016
rect 16354 5951 16750 5952
rect 12750 5884 12756 5948
rect 12820 5946 12826 5948
rect 12985 5946 13051 5949
rect 12820 5944 13051 5946
rect 12820 5888 12990 5944
rect 13046 5888 13051 5944
rect 12820 5886 13051 5888
rect 12820 5884 12826 5886
rect 12985 5883 13051 5886
rect 12157 5810 12223 5813
rect 12617 5810 12683 5813
rect 12157 5808 12683 5810
rect 12157 5752 12162 5808
rect 12218 5752 12622 5808
rect 12678 5752 12683 5808
rect 12157 5750 12683 5752
rect 12157 5747 12223 5750
rect 12617 5747 12683 5750
rect 13537 5810 13603 5813
rect 16849 5810 16915 5813
rect 13537 5808 16915 5810
rect 13537 5752 13542 5808
rect 13598 5752 16854 5808
rect 16910 5752 16915 5808
rect 13537 5750 16915 5752
rect 13537 5747 13603 5750
rect 16849 5747 16915 5750
rect 12801 5674 12867 5677
rect 14089 5674 14155 5677
rect 12801 5672 14155 5674
rect 12801 5616 12806 5672
rect 12862 5616 14094 5672
rect 14150 5616 14155 5672
rect 12801 5614 14155 5616
rect 12801 5611 12867 5614
rect 14089 5611 14155 5614
rect 8385 5538 8451 5541
rect 8937 5538 9003 5541
rect 8385 5536 9003 5538
rect 8385 5480 8390 5536
rect 8446 5480 8942 5536
rect 8998 5480 9003 5536
rect 8385 5478 9003 5480
rect 8385 5475 8451 5478
rect 8937 5475 9003 5478
rect 11973 5538 12039 5541
rect 12801 5538 12867 5541
rect 11973 5536 12867 5538
rect 11973 5480 11978 5536
rect 12034 5480 12806 5536
rect 12862 5480 12867 5536
rect 11973 5478 12867 5480
rect 11973 5475 12039 5478
rect 12801 5475 12867 5478
rect 1354 5472 1750 5473
rect 1354 5408 1360 5472
rect 1424 5408 1440 5472
rect 1504 5408 1520 5472
rect 1584 5408 1600 5472
rect 1664 5408 1680 5472
rect 1744 5408 1750 5472
rect 1354 5407 1750 5408
rect 7354 5472 7750 5473
rect 7354 5408 7360 5472
rect 7424 5408 7440 5472
rect 7504 5408 7520 5472
rect 7584 5408 7600 5472
rect 7664 5408 7680 5472
rect 7744 5408 7750 5472
rect 7354 5407 7750 5408
rect 13354 5472 13750 5473
rect 13354 5408 13360 5472
rect 13424 5408 13440 5472
rect 13504 5408 13520 5472
rect 13584 5408 13600 5472
rect 13664 5408 13680 5472
rect 13744 5408 13750 5472
rect 13354 5407 13750 5408
rect 8569 5402 8635 5405
rect 12893 5402 12959 5405
rect 8569 5400 12959 5402
rect 8569 5344 8574 5400
rect 8630 5344 12898 5400
rect 12954 5344 12959 5400
rect 8569 5342 12959 5344
rect 8569 5339 8635 5342
rect 12893 5339 12959 5342
rect 8661 5266 8727 5269
rect 8526 5264 8727 5266
rect 8526 5208 8666 5264
rect 8722 5208 8727 5264
rect 8526 5206 8727 5208
rect 8526 5133 8586 5206
rect 8661 5203 8727 5206
rect 9857 5266 9923 5269
rect 9990 5266 9996 5268
rect 9857 5264 9996 5266
rect 9857 5208 9862 5264
rect 9918 5208 9996 5264
rect 9857 5206 9996 5208
rect 9857 5203 9923 5206
rect 9990 5204 9996 5206
rect 10060 5204 10066 5268
rect 4981 5130 5047 5133
rect 7557 5130 7623 5133
rect 7925 5130 7991 5133
rect 4981 5128 7623 5130
rect 4981 5072 4986 5128
rect 5042 5072 7562 5128
rect 7618 5072 7623 5128
rect 4981 5070 7623 5072
rect 4981 5067 5047 5070
rect 7557 5067 7623 5070
rect 7790 5128 7991 5130
rect 7790 5072 7930 5128
rect 7986 5072 7991 5128
rect 7790 5070 7991 5072
rect 2589 4994 2655 4997
rect 4153 4994 4219 4997
rect 2589 4992 4219 4994
rect 2589 4936 2594 4992
rect 2650 4936 4158 4992
rect 4214 4936 4219 4992
rect 2589 4934 4219 4936
rect 2589 4931 2655 4934
rect 4153 4931 4219 4934
rect 4354 4928 4750 4929
rect 4354 4864 4360 4928
rect 4424 4864 4440 4928
rect 4504 4864 4520 4928
rect 4584 4864 4600 4928
rect 4664 4864 4680 4928
rect 4744 4864 4750 4928
rect 4354 4863 4750 4864
rect 7790 4858 7850 5070
rect 7925 5067 7991 5070
rect 8477 5128 8586 5133
rect 8477 5072 8482 5128
rect 8538 5072 8586 5128
rect 8477 5070 8586 5072
rect 9673 5130 9739 5133
rect 13353 5130 13419 5133
rect 9673 5128 13419 5130
rect 9673 5072 9678 5128
rect 9734 5072 13358 5128
rect 13414 5072 13419 5128
rect 9673 5070 13419 5072
rect 8477 5067 8543 5070
rect 9673 5067 9739 5070
rect 13353 5067 13419 5070
rect 7966 4932 7972 4996
rect 8036 4994 8042 4996
rect 8201 4994 8267 4997
rect 8036 4992 8267 4994
rect 8036 4936 8206 4992
rect 8262 4936 8267 4992
rect 8036 4934 8267 4936
rect 8036 4932 8042 4934
rect 8201 4931 8267 4934
rect 10354 4928 10750 4929
rect 10354 4864 10360 4928
rect 10424 4864 10440 4928
rect 10504 4864 10520 4928
rect 10584 4864 10600 4928
rect 10664 4864 10680 4928
rect 10744 4864 10750 4928
rect 10354 4863 10750 4864
rect 16354 4928 16750 4929
rect 16354 4864 16360 4928
rect 16424 4864 16440 4928
rect 16504 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16750 4928
rect 16354 4863 16750 4864
rect 7925 4858 7991 4861
rect 7790 4856 7991 4858
rect 7790 4800 7930 4856
rect 7986 4800 7991 4856
rect 7790 4798 7991 4800
rect 7925 4795 7991 4798
rect 7005 4722 7071 4725
rect 8477 4722 8543 4725
rect 7005 4720 8543 4722
rect 7005 4664 7010 4720
rect 7066 4664 8482 4720
rect 8538 4664 8543 4720
rect 7005 4662 8543 4664
rect 7005 4659 7071 4662
rect 8477 4659 8543 4662
rect 4889 4586 4955 4589
rect 5809 4586 5875 4589
rect 8477 4586 8543 4589
rect 4889 4584 8543 4586
rect 4889 4528 4894 4584
rect 4950 4528 5814 4584
rect 5870 4528 8482 4584
rect 8538 4528 8543 4584
rect 4889 4526 8543 4528
rect 4889 4523 4955 4526
rect 5809 4523 5875 4526
rect 8477 4523 8543 4526
rect 1354 4384 1750 4385
rect 1354 4320 1360 4384
rect 1424 4320 1440 4384
rect 1504 4320 1520 4384
rect 1584 4320 1600 4384
rect 1664 4320 1680 4384
rect 1744 4320 1750 4384
rect 1354 4319 1750 4320
rect 7354 4384 7750 4385
rect 7354 4320 7360 4384
rect 7424 4320 7440 4384
rect 7504 4320 7520 4384
rect 7584 4320 7600 4384
rect 7664 4320 7680 4384
rect 7744 4320 7750 4384
rect 7354 4319 7750 4320
rect 13354 4384 13750 4385
rect 13354 4320 13360 4384
rect 13424 4320 13440 4384
rect 13504 4320 13520 4384
rect 13584 4320 13600 4384
rect 13664 4320 13680 4384
rect 13744 4320 13750 4384
rect 13354 4319 13750 4320
rect 6545 4178 6611 4181
rect 9029 4178 9095 4181
rect 6545 4176 9095 4178
rect 6545 4120 6550 4176
rect 6606 4120 9034 4176
rect 9090 4120 9095 4176
rect 6545 4118 9095 4120
rect 6545 4115 6611 4118
rect 9029 4115 9095 4118
rect 4889 4042 4955 4045
rect 7741 4042 7807 4045
rect 15193 4044 15259 4045
rect 4889 4040 7807 4042
rect 4889 3984 4894 4040
rect 4950 3984 7746 4040
rect 7802 3984 7807 4040
rect 4889 3982 7807 3984
rect 4889 3979 4955 3982
rect 7741 3979 7807 3982
rect 15142 3980 15148 4044
rect 15212 4042 15259 4044
rect 15212 4040 15304 4042
rect 15254 3984 15304 4040
rect 15212 3982 15304 3984
rect 15212 3980 15259 3982
rect 15193 3979 15259 3980
rect 5625 3906 5691 3909
rect 9121 3906 9187 3909
rect 5625 3904 9187 3906
rect 5625 3848 5630 3904
rect 5686 3848 9126 3904
rect 9182 3848 9187 3904
rect 5625 3846 9187 3848
rect 5625 3843 5691 3846
rect 9121 3843 9187 3846
rect 12198 3844 12204 3908
rect 12268 3906 12274 3908
rect 15561 3906 15627 3909
rect 12268 3904 15627 3906
rect 12268 3848 15566 3904
rect 15622 3848 15627 3904
rect 12268 3846 15627 3848
rect 12268 3844 12274 3846
rect 15561 3843 15627 3846
rect 4354 3840 4750 3841
rect 4354 3776 4360 3840
rect 4424 3776 4440 3840
rect 4504 3776 4520 3840
rect 4584 3776 4600 3840
rect 4664 3776 4680 3840
rect 4744 3776 4750 3840
rect 4354 3775 4750 3776
rect 10354 3840 10750 3841
rect 10354 3776 10360 3840
rect 10424 3776 10440 3840
rect 10504 3776 10520 3840
rect 10584 3776 10600 3840
rect 10664 3776 10680 3840
rect 10744 3776 10750 3840
rect 10354 3775 10750 3776
rect 16354 3840 16750 3841
rect 16354 3776 16360 3840
rect 16424 3776 16440 3840
rect 16504 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16750 3840
rect 16354 3775 16750 3776
rect 12249 3634 12315 3637
rect 14549 3634 14615 3637
rect 12249 3632 14615 3634
rect 12249 3576 12254 3632
rect 12310 3576 14554 3632
rect 14610 3576 14615 3632
rect 12249 3574 14615 3576
rect 12249 3571 12315 3574
rect 14549 3571 14615 3574
rect 4429 3362 4495 3365
rect 9765 3364 9831 3365
rect 5942 3362 5948 3364
rect 4429 3360 5948 3362
rect 4429 3304 4434 3360
rect 4490 3304 5948 3360
rect 4429 3302 5948 3304
rect 4429 3299 4495 3302
rect 5942 3300 5948 3302
rect 6012 3300 6018 3364
rect 9765 3360 9812 3364
rect 9876 3362 9882 3364
rect 9765 3304 9770 3360
rect 9765 3300 9812 3304
rect 9876 3302 9922 3362
rect 9876 3300 9882 3302
rect 9765 3299 9831 3300
rect 1354 3296 1750 3297
rect 1354 3232 1360 3296
rect 1424 3232 1440 3296
rect 1504 3232 1520 3296
rect 1584 3232 1600 3296
rect 1664 3232 1680 3296
rect 1744 3232 1750 3296
rect 1354 3231 1750 3232
rect 7354 3296 7750 3297
rect 7354 3232 7360 3296
rect 7424 3232 7440 3296
rect 7504 3232 7520 3296
rect 7584 3232 7600 3296
rect 7664 3232 7680 3296
rect 7744 3232 7750 3296
rect 7354 3231 7750 3232
rect 13354 3296 13750 3297
rect 13354 3232 13360 3296
rect 13424 3232 13440 3296
rect 13504 3232 13520 3296
rect 13584 3232 13600 3296
rect 13664 3232 13680 3296
rect 13744 3232 13750 3296
rect 13354 3231 13750 3232
rect 12985 3226 13051 3229
rect 12985 3224 13186 3226
rect 12985 3168 12990 3224
rect 13046 3168 13186 3224
rect 12985 3166 13186 3168
rect 12985 3163 13051 3166
rect 5165 3090 5231 3093
rect 7833 3090 7899 3093
rect 5165 3088 7899 3090
rect 5165 3032 5170 3088
rect 5226 3032 7838 3088
rect 7894 3032 7899 3088
rect 5165 3030 7899 3032
rect 13126 3090 13186 3166
rect 13813 3090 13879 3093
rect 14181 3090 14247 3093
rect 13126 3088 14247 3090
rect 13126 3032 13818 3088
rect 13874 3032 14186 3088
rect 14242 3032 14247 3088
rect 13126 3030 14247 3032
rect 5165 3027 5231 3030
rect 7833 3027 7899 3030
rect 13813 3027 13879 3030
rect 14181 3027 14247 3030
rect 7649 2954 7715 2957
rect 7966 2954 7972 2956
rect 7649 2952 7972 2954
rect 7649 2896 7654 2952
rect 7710 2896 7972 2952
rect 7649 2894 7972 2896
rect 7649 2891 7715 2894
rect 7966 2892 7972 2894
rect 8036 2892 8042 2956
rect 12341 2954 12407 2957
rect 15285 2954 15351 2957
rect 12341 2952 15351 2954
rect 12341 2896 12346 2952
rect 12402 2896 15290 2952
rect 15346 2896 15351 2952
rect 12341 2894 15351 2896
rect 12341 2891 12407 2894
rect 15285 2891 15351 2894
rect 4354 2752 4750 2753
rect 4354 2688 4360 2752
rect 4424 2688 4440 2752
rect 4504 2688 4520 2752
rect 4584 2688 4600 2752
rect 4664 2688 4680 2752
rect 4744 2688 4750 2752
rect 4354 2687 4750 2688
rect 10354 2752 10750 2753
rect 10354 2688 10360 2752
rect 10424 2688 10440 2752
rect 10504 2688 10520 2752
rect 10584 2688 10600 2752
rect 10664 2688 10680 2752
rect 10744 2688 10750 2752
rect 10354 2687 10750 2688
rect 16354 2752 16750 2753
rect 16354 2688 16360 2752
rect 16424 2688 16440 2752
rect 16504 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16750 2752
rect 16354 2687 16750 2688
rect 5809 2682 5875 2685
rect 6494 2682 6500 2684
rect 5809 2680 6500 2682
rect 5809 2624 5814 2680
rect 5870 2624 6500 2680
rect 5809 2622 6500 2624
rect 5809 2619 5875 2622
rect 6494 2620 6500 2622
rect 6564 2620 6570 2684
rect 14549 2682 14615 2685
rect 14774 2682 14780 2684
rect 14549 2680 14780 2682
rect 14549 2624 14554 2680
rect 14610 2624 14780 2680
rect 14549 2622 14780 2624
rect 14549 2619 14615 2622
rect 14774 2620 14780 2622
rect 14844 2620 14850 2684
rect 1301 2546 1367 2549
rect 3509 2546 3575 2549
rect 9029 2546 9095 2549
rect 1301 2544 2790 2546
rect 1301 2488 1306 2544
rect 1362 2488 2790 2544
rect 1301 2486 2790 2488
rect 1301 2483 1367 2486
rect 2730 2410 2790 2486
rect 3509 2544 9095 2546
rect 3509 2488 3514 2544
rect 3570 2488 9034 2544
rect 9090 2488 9095 2544
rect 3509 2486 9095 2488
rect 3509 2483 3575 2486
rect 9029 2483 9095 2486
rect 6085 2412 6151 2413
rect 6085 2410 6132 2412
rect 2730 2408 6132 2410
rect 6196 2410 6202 2412
rect 9121 2410 9187 2413
rect 9254 2410 9260 2412
rect 2730 2352 6090 2408
rect 2730 2350 6132 2352
rect 6085 2348 6132 2350
rect 6196 2350 6242 2410
rect 9121 2408 9260 2410
rect 9121 2352 9126 2408
rect 9182 2352 9260 2408
rect 9121 2350 9260 2352
rect 6196 2348 6202 2350
rect 6085 2347 6151 2348
rect 9121 2347 9187 2350
rect 9254 2348 9260 2350
rect 9324 2410 9330 2412
rect 12525 2410 12591 2413
rect 9324 2408 12591 2410
rect 9324 2352 12530 2408
rect 12586 2352 12591 2408
rect 9324 2350 12591 2352
rect 9324 2348 9330 2350
rect 12525 2347 12591 2350
rect 13905 2274 13971 2277
rect 16021 2274 16087 2277
rect 13905 2272 16087 2274
rect 13905 2216 13910 2272
rect 13966 2216 16026 2272
rect 16082 2216 16087 2272
rect 13905 2214 16087 2216
rect 13905 2211 13971 2214
rect 16021 2211 16087 2214
rect 1354 2208 1750 2209
rect 1354 2144 1360 2208
rect 1424 2144 1440 2208
rect 1504 2144 1520 2208
rect 1584 2144 1600 2208
rect 1664 2144 1680 2208
rect 1744 2144 1750 2208
rect 1354 2143 1750 2144
rect 7354 2208 7750 2209
rect 7354 2144 7360 2208
rect 7424 2144 7440 2208
rect 7504 2144 7520 2208
rect 7584 2144 7600 2208
rect 7664 2144 7680 2208
rect 7744 2144 7750 2208
rect 7354 2143 7750 2144
rect 13354 2208 13750 2209
rect 13354 2144 13360 2208
rect 13424 2144 13440 2208
rect 13504 2144 13520 2208
rect 13584 2144 13600 2208
rect 13664 2144 13680 2208
rect 13744 2144 13750 2208
rect 13354 2143 13750 2144
rect 10869 2138 10935 2141
rect 13077 2138 13143 2141
rect 10869 2136 10978 2138
rect 10869 2080 10874 2136
rect 10930 2080 10978 2136
rect 10869 2075 10978 2080
rect 10918 2002 10978 2075
rect 12942 2136 13143 2138
rect 12942 2080 13082 2136
rect 13138 2080 13143 2136
rect 12942 2078 13143 2080
rect 11329 2002 11395 2005
rect 8342 2000 11395 2002
rect 8342 1944 11334 2000
rect 11390 1944 11395 2000
rect 8342 1942 11395 1944
rect 1761 1866 1827 1869
rect 4981 1866 5047 1869
rect 1761 1864 5047 1866
rect 1761 1808 1766 1864
rect 1822 1808 4986 1864
rect 5042 1808 5047 1864
rect 1761 1806 5047 1808
rect 1761 1803 1827 1806
rect 4981 1803 5047 1806
rect 4354 1664 4750 1665
rect 4354 1600 4360 1664
rect 4424 1600 4440 1664
rect 4504 1600 4520 1664
rect 4584 1600 4600 1664
rect 4664 1600 4680 1664
rect 4744 1600 4750 1664
rect 4354 1599 4750 1600
rect 6361 1594 6427 1597
rect 8017 1594 8083 1597
rect 8342 1594 8402 1942
rect 11329 1939 11395 1942
rect 12801 2002 12867 2005
rect 12942 2002 13002 2078
rect 13077 2075 13143 2078
rect 15285 2138 15351 2141
rect 15653 2138 15719 2141
rect 15285 2136 15719 2138
rect 15285 2080 15290 2136
rect 15346 2080 15658 2136
rect 15714 2080 15719 2136
rect 15285 2078 15719 2080
rect 15285 2075 15351 2078
rect 15653 2075 15719 2078
rect 12801 2000 13002 2002
rect 12801 1944 12806 2000
rect 12862 1944 13002 2000
rect 12801 1942 13002 1944
rect 12801 1939 12867 1942
rect 13118 1940 13124 2004
rect 13188 2002 13194 2004
rect 13353 2002 13419 2005
rect 13188 2000 13419 2002
rect 13188 1944 13358 2000
rect 13414 1944 13419 2000
rect 13188 1942 13419 1944
rect 13188 1940 13194 1942
rect 13353 1939 13419 1942
rect 8569 1866 8635 1869
rect 8702 1866 8708 1868
rect 8569 1864 8708 1866
rect 8569 1808 8574 1864
rect 8630 1808 8708 1864
rect 8569 1806 8708 1808
rect 8569 1803 8635 1806
rect 8702 1804 8708 1806
rect 8772 1866 8778 1868
rect 12341 1866 12407 1869
rect 8772 1864 12407 1866
rect 8772 1808 12346 1864
rect 12402 1808 12407 1864
rect 8772 1806 12407 1808
rect 8772 1804 8778 1806
rect 12341 1803 12407 1806
rect 14917 1866 14983 1869
rect 15469 1866 15535 1869
rect 16205 1866 16271 1869
rect 14917 1864 16271 1866
rect 14917 1808 14922 1864
rect 14978 1808 15474 1864
rect 15530 1808 16210 1864
rect 16266 1808 16271 1864
rect 14917 1806 16271 1808
rect 14917 1803 14983 1806
rect 15469 1803 15535 1806
rect 16205 1803 16271 1806
rect 9765 1730 9831 1733
rect 9990 1730 9996 1732
rect 9765 1728 9996 1730
rect 9765 1672 9770 1728
rect 9826 1672 9996 1728
rect 9765 1670 9996 1672
rect 9765 1667 9831 1670
rect 9990 1668 9996 1670
rect 10060 1668 10066 1732
rect 13813 1730 13879 1733
rect 15745 1730 15811 1733
rect 13813 1728 15811 1730
rect 13813 1672 13818 1728
rect 13874 1672 15750 1728
rect 15806 1672 15811 1728
rect 13813 1670 15811 1672
rect 13813 1667 13879 1670
rect 15745 1667 15811 1670
rect 10354 1664 10750 1665
rect 10354 1600 10360 1664
rect 10424 1600 10440 1664
rect 10504 1600 10520 1664
rect 10584 1600 10600 1664
rect 10664 1600 10680 1664
rect 10744 1600 10750 1664
rect 10354 1599 10750 1600
rect 16354 1664 16750 1665
rect 16354 1600 16360 1664
rect 16424 1600 16440 1664
rect 16504 1600 16520 1664
rect 16584 1600 16600 1664
rect 16664 1600 16680 1664
rect 16744 1600 16750 1664
rect 16354 1599 16750 1600
rect 6361 1592 8402 1594
rect 6361 1536 6366 1592
rect 6422 1536 8022 1592
rect 8078 1536 8402 1592
rect 6361 1534 8402 1536
rect 9673 1594 9739 1597
rect 9806 1594 9812 1596
rect 9673 1592 9812 1594
rect 9673 1536 9678 1592
rect 9734 1536 9812 1592
rect 9673 1534 9812 1536
rect 6361 1531 6427 1534
rect 8017 1531 8083 1534
rect 9673 1531 9739 1534
rect 9806 1532 9812 1534
rect 9876 1532 9882 1596
rect 13905 1594 13971 1597
rect 15142 1594 15148 1596
rect 13905 1592 15148 1594
rect 13905 1536 13910 1592
rect 13966 1536 15148 1592
rect 13905 1534 15148 1536
rect 13905 1531 13971 1534
rect 15142 1532 15148 1534
rect 15212 1532 15218 1596
rect 4061 1458 4127 1461
rect 4797 1458 4863 1461
rect 15653 1458 15719 1461
rect 4061 1456 15719 1458
rect 4061 1400 4066 1456
rect 4122 1400 4802 1456
rect 4858 1400 15658 1456
rect 15714 1400 15719 1456
rect 4061 1398 15719 1400
rect 4061 1395 4127 1398
rect 4797 1395 4863 1398
rect 15653 1395 15719 1398
rect 9990 1260 9996 1324
rect 10060 1322 10066 1324
rect 10685 1322 10751 1325
rect 10060 1320 10751 1322
rect 10060 1264 10690 1320
rect 10746 1264 10751 1320
rect 10060 1262 10751 1264
rect 10060 1260 10066 1262
rect 10685 1259 10751 1262
rect 11053 1322 11119 1325
rect 15101 1324 15167 1325
rect 11278 1322 11284 1324
rect 11053 1320 11284 1322
rect 11053 1264 11058 1320
rect 11114 1264 11284 1320
rect 11053 1262 11284 1264
rect 11053 1259 11119 1262
rect 11278 1260 11284 1262
rect 11348 1260 11354 1324
rect 15101 1322 15148 1324
rect 15056 1320 15148 1322
rect 15056 1264 15106 1320
rect 15056 1262 15148 1264
rect 15101 1260 15148 1262
rect 15212 1260 15218 1324
rect 15101 1259 15167 1260
rect 9673 1186 9739 1189
rect 9806 1186 9812 1188
rect 9673 1184 9812 1186
rect 9673 1128 9678 1184
rect 9734 1128 9812 1184
rect 9673 1126 9812 1128
rect 9673 1123 9739 1126
rect 9806 1124 9812 1126
rect 9876 1124 9882 1188
rect 13997 1186 14063 1189
rect 15193 1186 15259 1189
rect 13997 1184 15259 1186
rect 13997 1128 14002 1184
rect 14058 1128 15198 1184
rect 15254 1128 15259 1184
rect 13997 1126 15259 1128
rect 13997 1123 14063 1126
rect 15193 1123 15259 1126
rect 1354 1120 1750 1121
rect 1354 1056 1360 1120
rect 1424 1056 1440 1120
rect 1504 1056 1520 1120
rect 1584 1056 1600 1120
rect 1664 1056 1680 1120
rect 1744 1056 1750 1120
rect 1354 1055 1750 1056
rect 7354 1120 7750 1121
rect 7354 1056 7360 1120
rect 7424 1056 7440 1120
rect 7504 1056 7520 1120
rect 7584 1056 7600 1120
rect 7664 1056 7680 1120
rect 7744 1056 7750 1120
rect 7354 1055 7750 1056
rect 13354 1120 13750 1121
rect 13354 1056 13360 1120
rect 13424 1056 13440 1120
rect 13504 1056 13520 1120
rect 13584 1056 13600 1120
rect 13664 1056 13680 1120
rect 13744 1056 13750 1120
rect 13354 1055 13750 1056
rect 4354 576 4750 577
rect 4354 512 4360 576
rect 4424 512 4440 576
rect 4504 512 4520 576
rect 4584 512 4600 576
rect 4664 512 4680 576
rect 4744 512 4750 576
rect 4354 511 4750 512
rect 10354 576 10750 577
rect 10354 512 10360 576
rect 10424 512 10440 576
rect 10504 512 10520 576
rect 10584 512 10600 576
rect 10664 512 10680 576
rect 10744 512 10750 576
rect 10354 511 10750 512
rect 16354 576 16750 577
rect 16354 512 16360 576
rect 16424 512 16440 576
rect 16504 512 16520 576
rect 16584 512 16600 576
rect 16664 512 16680 576
rect 16744 512 16750 576
rect 16354 511 16750 512
<< via3 >>
rect 1360 17436 1424 17440
rect 1360 17380 1364 17436
rect 1364 17380 1420 17436
rect 1420 17380 1424 17436
rect 1360 17376 1424 17380
rect 1440 17436 1504 17440
rect 1440 17380 1444 17436
rect 1444 17380 1500 17436
rect 1500 17380 1504 17436
rect 1440 17376 1504 17380
rect 1520 17436 1584 17440
rect 1520 17380 1524 17436
rect 1524 17380 1580 17436
rect 1580 17380 1584 17436
rect 1520 17376 1584 17380
rect 1600 17436 1664 17440
rect 1600 17380 1604 17436
rect 1604 17380 1660 17436
rect 1660 17380 1664 17436
rect 1600 17376 1664 17380
rect 1680 17436 1744 17440
rect 1680 17380 1684 17436
rect 1684 17380 1740 17436
rect 1740 17380 1744 17436
rect 1680 17376 1744 17380
rect 7360 17436 7424 17440
rect 7360 17380 7364 17436
rect 7364 17380 7420 17436
rect 7420 17380 7424 17436
rect 7360 17376 7424 17380
rect 7440 17436 7504 17440
rect 7440 17380 7444 17436
rect 7444 17380 7500 17436
rect 7500 17380 7504 17436
rect 7440 17376 7504 17380
rect 7520 17436 7584 17440
rect 7520 17380 7524 17436
rect 7524 17380 7580 17436
rect 7580 17380 7584 17436
rect 7520 17376 7584 17380
rect 7600 17436 7664 17440
rect 7600 17380 7604 17436
rect 7604 17380 7660 17436
rect 7660 17380 7664 17436
rect 7600 17376 7664 17380
rect 7680 17436 7744 17440
rect 7680 17380 7684 17436
rect 7684 17380 7740 17436
rect 7740 17380 7744 17436
rect 7680 17376 7744 17380
rect 13360 17436 13424 17440
rect 13360 17380 13364 17436
rect 13364 17380 13420 17436
rect 13420 17380 13424 17436
rect 13360 17376 13424 17380
rect 13440 17436 13504 17440
rect 13440 17380 13444 17436
rect 13444 17380 13500 17436
rect 13500 17380 13504 17436
rect 13440 17376 13504 17380
rect 13520 17436 13584 17440
rect 13520 17380 13524 17436
rect 13524 17380 13580 17436
rect 13580 17380 13584 17436
rect 13520 17376 13584 17380
rect 13600 17436 13664 17440
rect 13600 17380 13604 17436
rect 13604 17380 13660 17436
rect 13660 17380 13664 17436
rect 13600 17376 13664 17380
rect 13680 17436 13744 17440
rect 13680 17380 13684 17436
rect 13684 17380 13740 17436
rect 13740 17380 13744 17436
rect 13680 17376 13744 17380
rect 4360 16892 4424 16896
rect 4360 16836 4364 16892
rect 4364 16836 4420 16892
rect 4420 16836 4424 16892
rect 4360 16832 4424 16836
rect 4440 16892 4504 16896
rect 4440 16836 4444 16892
rect 4444 16836 4500 16892
rect 4500 16836 4504 16892
rect 4440 16832 4504 16836
rect 4520 16892 4584 16896
rect 4520 16836 4524 16892
rect 4524 16836 4580 16892
rect 4580 16836 4584 16892
rect 4520 16832 4584 16836
rect 4600 16892 4664 16896
rect 4600 16836 4604 16892
rect 4604 16836 4660 16892
rect 4660 16836 4664 16892
rect 4600 16832 4664 16836
rect 4680 16892 4744 16896
rect 4680 16836 4684 16892
rect 4684 16836 4740 16892
rect 4740 16836 4744 16892
rect 4680 16832 4744 16836
rect 10360 16892 10424 16896
rect 10360 16836 10364 16892
rect 10364 16836 10420 16892
rect 10420 16836 10424 16892
rect 10360 16832 10424 16836
rect 10440 16892 10504 16896
rect 10440 16836 10444 16892
rect 10444 16836 10500 16892
rect 10500 16836 10504 16892
rect 10440 16832 10504 16836
rect 10520 16892 10584 16896
rect 10520 16836 10524 16892
rect 10524 16836 10580 16892
rect 10580 16836 10584 16892
rect 10520 16832 10584 16836
rect 10600 16892 10664 16896
rect 10600 16836 10604 16892
rect 10604 16836 10660 16892
rect 10660 16836 10664 16892
rect 10600 16832 10664 16836
rect 10680 16892 10744 16896
rect 10680 16836 10684 16892
rect 10684 16836 10740 16892
rect 10740 16836 10744 16892
rect 10680 16832 10744 16836
rect 16360 16892 16424 16896
rect 16360 16836 16364 16892
rect 16364 16836 16420 16892
rect 16420 16836 16424 16892
rect 16360 16832 16424 16836
rect 16440 16892 16504 16896
rect 16440 16836 16444 16892
rect 16444 16836 16500 16892
rect 16500 16836 16504 16892
rect 16440 16832 16504 16836
rect 16520 16892 16584 16896
rect 16520 16836 16524 16892
rect 16524 16836 16580 16892
rect 16580 16836 16584 16892
rect 16520 16832 16584 16836
rect 16600 16892 16664 16896
rect 16600 16836 16604 16892
rect 16604 16836 16660 16892
rect 16660 16836 16664 16892
rect 16600 16832 16664 16836
rect 16680 16892 16744 16896
rect 16680 16836 16684 16892
rect 16684 16836 16740 16892
rect 16740 16836 16744 16892
rect 16680 16832 16744 16836
rect 6500 16628 6564 16692
rect 8708 16628 8772 16692
rect 1360 16348 1424 16352
rect 1360 16292 1364 16348
rect 1364 16292 1420 16348
rect 1420 16292 1424 16348
rect 1360 16288 1424 16292
rect 1440 16348 1504 16352
rect 1440 16292 1444 16348
rect 1444 16292 1500 16348
rect 1500 16292 1504 16348
rect 1440 16288 1504 16292
rect 1520 16348 1584 16352
rect 1520 16292 1524 16348
rect 1524 16292 1580 16348
rect 1580 16292 1584 16348
rect 1520 16288 1584 16292
rect 1600 16348 1664 16352
rect 1600 16292 1604 16348
rect 1604 16292 1660 16348
rect 1660 16292 1664 16348
rect 1600 16288 1664 16292
rect 1680 16348 1744 16352
rect 1680 16292 1684 16348
rect 1684 16292 1740 16348
rect 1740 16292 1744 16348
rect 1680 16288 1744 16292
rect 7360 16348 7424 16352
rect 7360 16292 7364 16348
rect 7364 16292 7420 16348
rect 7420 16292 7424 16348
rect 7360 16288 7424 16292
rect 7440 16348 7504 16352
rect 7440 16292 7444 16348
rect 7444 16292 7500 16348
rect 7500 16292 7504 16348
rect 7440 16288 7504 16292
rect 7520 16348 7584 16352
rect 7520 16292 7524 16348
rect 7524 16292 7580 16348
rect 7580 16292 7584 16348
rect 7520 16288 7584 16292
rect 7600 16348 7664 16352
rect 7600 16292 7604 16348
rect 7604 16292 7660 16348
rect 7660 16292 7664 16348
rect 7600 16288 7664 16292
rect 7680 16348 7744 16352
rect 7680 16292 7684 16348
rect 7684 16292 7740 16348
rect 7740 16292 7744 16348
rect 7680 16288 7744 16292
rect 13360 16348 13424 16352
rect 13360 16292 13364 16348
rect 13364 16292 13420 16348
rect 13420 16292 13424 16348
rect 13360 16288 13424 16292
rect 13440 16348 13504 16352
rect 13440 16292 13444 16348
rect 13444 16292 13500 16348
rect 13500 16292 13504 16348
rect 13440 16288 13504 16292
rect 13520 16348 13584 16352
rect 13520 16292 13524 16348
rect 13524 16292 13580 16348
rect 13580 16292 13584 16348
rect 13520 16288 13584 16292
rect 13600 16348 13664 16352
rect 13600 16292 13604 16348
rect 13604 16292 13660 16348
rect 13660 16292 13664 16348
rect 13600 16288 13664 16292
rect 13680 16348 13744 16352
rect 13680 16292 13684 16348
rect 13684 16292 13740 16348
rect 13740 16292 13744 16348
rect 13680 16288 13744 16292
rect 4360 15804 4424 15808
rect 4360 15748 4364 15804
rect 4364 15748 4420 15804
rect 4420 15748 4424 15804
rect 4360 15744 4424 15748
rect 4440 15804 4504 15808
rect 4440 15748 4444 15804
rect 4444 15748 4500 15804
rect 4500 15748 4504 15804
rect 4440 15744 4504 15748
rect 4520 15804 4584 15808
rect 4520 15748 4524 15804
rect 4524 15748 4580 15804
rect 4580 15748 4584 15804
rect 4520 15744 4584 15748
rect 4600 15804 4664 15808
rect 4600 15748 4604 15804
rect 4604 15748 4660 15804
rect 4660 15748 4664 15804
rect 4600 15744 4664 15748
rect 4680 15804 4744 15808
rect 4680 15748 4684 15804
rect 4684 15748 4740 15804
rect 4740 15748 4744 15804
rect 4680 15744 4744 15748
rect 10360 15804 10424 15808
rect 10360 15748 10364 15804
rect 10364 15748 10420 15804
rect 10420 15748 10424 15804
rect 10360 15744 10424 15748
rect 10440 15804 10504 15808
rect 10440 15748 10444 15804
rect 10444 15748 10500 15804
rect 10500 15748 10504 15804
rect 10440 15744 10504 15748
rect 10520 15804 10584 15808
rect 10520 15748 10524 15804
rect 10524 15748 10580 15804
rect 10580 15748 10584 15804
rect 10520 15744 10584 15748
rect 10600 15804 10664 15808
rect 10600 15748 10604 15804
rect 10604 15748 10660 15804
rect 10660 15748 10664 15804
rect 10600 15744 10664 15748
rect 10680 15804 10744 15808
rect 10680 15748 10684 15804
rect 10684 15748 10740 15804
rect 10740 15748 10744 15804
rect 10680 15744 10744 15748
rect 16360 15804 16424 15808
rect 16360 15748 16364 15804
rect 16364 15748 16420 15804
rect 16420 15748 16424 15804
rect 16360 15744 16424 15748
rect 16440 15804 16504 15808
rect 16440 15748 16444 15804
rect 16444 15748 16500 15804
rect 16500 15748 16504 15804
rect 16440 15744 16504 15748
rect 16520 15804 16584 15808
rect 16520 15748 16524 15804
rect 16524 15748 16580 15804
rect 16580 15748 16584 15804
rect 16520 15744 16584 15748
rect 16600 15804 16664 15808
rect 16600 15748 16604 15804
rect 16604 15748 16660 15804
rect 16660 15748 16664 15804
rect 16600 15744 16664 15748
rect 16680 15804 16744 15808
rect 16680 15748 16684 15804
rect 16684 15748 16740 15804
rect 16740 15748 16744 15804
rect 16680 15744 16744 15748
rect 9260 15404 9324 15468
rect 6132 15268 6196 15332
rect 11284 15268 11348 15332
rect 13124 15268 13188 15332
rect 1360 15260 1424 15264
rect 1360 15204 1364 15260
rect 1364 15204 1420 15260
rect 1420 15204 1424 15260
rect 1360 15200 1424 15204
rect 1440 15260 1504 15264
rect 1440 15204 1444 15260
rect 1444 15204 1500 15260
rect 1500 15204 1504 15260
rect 1440 15200 1504 15204
rect 1520 15260 1584 15264
rect 1520 15204 1524 15260
rect 1524 15204 1580 15260
rect 1580 15204 1584 15260
rect 1520 15200 1584 15204
rect 1600 15260 1664 15264
rect 1600 15204 1604 15260
rect 1604 15204 1660 15260
rect 1660 15204 1664 15260
rect 1600 15200 1664 15204
rect 1680 15260 1744 15264
rect 1680 15204 1684 15260
rect 1684 15204 1740 15260
rect 1740 15204 1744 15260
rect 1680 15200 1744 15204
rect 7360 15260 7424 15264
rect 7360 15204 7364 15260
rect 7364 15204 7420 15260
rect 7420 15204 7424 15260
rect 7360 15200 7424 15204
rect 7440 15260 7504 15264
rect 7440 15204 7444 15260
rect 7444 15204 7500 15260
rect 7500 15204 7504 15260
rect 7440 15200 7504 15204
rect 7520 15260 7584 15264
rect 7520 15204 7524 15260
rect 7524 15204 7580 15260
rect 7580 15204 7584 15260
rect 7520 15200 7584 15204
rect 7600 15260 7664 15264
rect 7600 15204 7604 15260
rect 7604 15204 7660 15260
rect 7660 15204 7664 15260
rect 7600 15200 7664 15204
rect 7680 15260 7744 15264
rect 7680 15204 7684 15260
rect 7684 15204 7740 15260
rect 7740 15204 7744 15260
rect 7680 15200 7744 15204
rect 13360 15260 13424 15264
rect 13360 15204 13364 15260
rect 13364 15204 13420 15260
rect 13420 15204 13424 15260
rect 13360 15200 13424 15204
rect 13440 15260 13504 15264
rect 13440 15204 13444 15260
rect 13444 15204 13500 15260
rect 13500 15204 13504 15260
rect 13440 15200 13504 15204
rect 13520 15260 13584 15264
rect 13520 15204 13524 15260
rect 13524 15204 13580 15260
rect 13580 15204 13584 15260
rect 13520 15200 13584 15204
rect 13600 15260 13664 15264
rect 13600 15204 13604 15260
rect 13604 15204 13660 15260
rect 13660 15204 13664 15260
rect 13600 15200 13664 15204
rect 13680 15260 13744 15264
rect 13680 15204 13684 15260
rect 13684 15204 13740 15260
rect 13740 15204 13744 15260
rect 13680 15200 13744 15204
rect 4360 14716 4424 14720
rect 4360 14660 4364 14716
rect 4364 14660 4420 14716
rect 4420 14660 4424 14716
rect 4360 14656 4424 14660
rect 4440 14716 4504 14720
rect 4440 14660 4444 14716
rect 4444 14660 4500 14716
rect 4500 14660 4504 14716
rect 4440 14656 4504 14660
rect 4520 14716 4584 14720
rect 4520 14660 4524 14716
rect 4524 14660 4580 14716
rect 4580 14660 4584 14716
rect 4520 14656 4584 14660
rect 4600 14716 4664 14720
rect 4600 14660 4604 14716
rect 4604 14660 4660 14716
rect 4660 14660 4664 14716
rect 4600 14656 4664 14660
rect 4680 14716 4744 14720
rect 4680 14660 4684 14716
rect 4684 14660 4740 14716
rect 4740 14660 4744 14716
rect 4680 14656 4744 14660
rect 10360 14716 10424 14720
rect 10360 14660 10364 14716
rect 10364 14660 10420 14716
rect 10420 14660 10424 14716
rect 10360 14656 10424 14660
rect 10440 14716 10504 14720
rect 10440 14660 10444 14716
rect 10444 14660 10500 14716
rect 10500 14660 10504 14716
rect 10440 14656 10504 14660
rect 10520 14716 10584 14720
rect 10520 14660 10524 14716
rect 10524 14660 10580 14716
rect 10580 14660 10584 14716
rect 10520 14656 10584 14660
rect 10600 14716 10664 14720
rect 10600 14660 10604 14716
rect 10604 14660 10660 14716
rect 10660 14660 10664 14716
rect 10600 14656 10664 14660
rect 10680 14716 10744 14720
rect 10680 14660 10684 14716
rect 10684 14660 10740 14716
rect 10740 14660 10744 14716
rect 10680 14656 10744 14660
rect 16360 14716 16424 14720
rect 16360 14660 16364 14716
rect 16364 14660 16420 14716
rect 16420 14660 16424 14716
rect 16360 14656 16424 14660
rect 16440 14716 16504 14720
rect 16440 14660 16444 14716
rect 16444 14660 16500 14716
rect 16500 14660 16504 14716
rect 16440 14656 16504 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 1360 14172 1424 14176
rect 1360 14116 1364 14172
rect 1364 14116 1420 14172
rect 1420 14116 1424 14172
rect 1360 14112 1424 14116
rect 1440 14172 1504 14176
rect 1440 14116 1444 14172
rect 1444 14116 1500 14172
rect 1500 14116 1504 14172
rect 1440 14112 1504 14116
rect 1520 14172 1584 14176
rect 1520 14116 1524 14172
rect 1524 14116 1580 14172
rect 1580 14116 1584 14172
rect 1520 14112 1584 14116
rect 1600 14172 1664 14176
rect 1600 14116 1604 14172
rect 1604 14116 1660 14172
rect 1660 14116 1664 14172
rect 1600 14112 1664 14116
rect 1680 14172 1744 14176
rect 1680 14116 1684 14172
rect 1684 14116 1740 14172
rect 1740 14116 1744 14172
rect 1680 14112 1744 14116
rect 7360 14172 7424 14176
rect 7360 14116 7364 14172
rect 7364 14116 7420 14172
rect 7420 14116 7424 14172
rect 7360 14112 7424 14116
rect 7440 14172 7504 14176
rect 7440 14116 7444 14172
rect 7444 14116 7500 14172
rect 7500 14116 7504 14172
rect 7440 14112 7504 14116
rect 7520 14172 7584 14176
rect 7520 14116 7524 14172
rect 7524 14116 7580 14172
rect 7580 14116 7584 14172
rect 7520 14112 7584 14116
rect 7600 14172 7664 14176
rect 7600 14116 7604 14172
rect 7604 14116 7660 14172
rect 7660 14116 7664 14172
rect 7600 14112 7664 14116
rect 7680 14172 7744 14176
rect 7680 14116 7684 14172
rect 7684 14116 7740 14172
rect 7740 14116 7744 14172
rect 7680 14112 7744 14116
rect 13360 14172 13424 14176
rect 13360 14116 13364 14172
rect 13364 14116 13420 14172
rect 13420 14116 13424 14172
rect 13360 14112 13424 14116
rect 13440 14172 13504 14176
rect 13440 14116 13444 14172
rect 13444 14116 13500 14172
rect 13500 14116 13504 14172
rect 13440 14112 13504 14116
rect 13520 14172 13584 14176
rect 13520 14116 13524 14172
rect 13524 14116 13580 14172
rect 13580 14116 13584 14172
rect 13520 14112 13584 14116
rect 13600 14172 13664 14176
rect 13600 14116 13604 14172
rect 13604 14116 13660 14172
rect 13660 14116 13664 14172
rect 13600 14112 13664 14116
rect 13680 14172 13744 14176
rect 13680 14116 13684 14172
rect 13684 14116 13740 14172
rect 13740 14116 13744 14172
rect 13680 14112 13744 14116
rect 4360 13628 4424 13632
rect 4360 13572 4364 13628
rect 4364 13572 4420 13628
rect 4420 13572 4424 13628
rect 4360 13568 4424 13572
rect 4440 13628 4504 13632
rect 4440 13572 4444 13628
rect 4444 13572 4500 13628
rect 4500 13572 4504 13628
rect 4440 13568 4504 13572
rect 4520 13628 4584 13632
rect 4520 13572 4524 13628
rect 4524 13572 4580 13628
rect 4580 13572 4584 13628
rect 4520 13568 4584 13572
rect 4600 13628 4664 13632
rect 4600 13572 4604 13628
rect 4604 13572 4660 13628
rect 4660 13572 4664 13628
rect 4600 13568 4664 13572
rect 4680 13628 4744 13632
rect 4680 13572 4684 13628
rect 4684 13572 4740 13628
rect 4740 13572 4744 13628
rect 4680 13568 4744 13572
rect 10360 13628 10424 13632
rect 10360 13572 10364 13628
rect 10364 13572 10420 13628
rect 10420 13572 10424 13628
rect 10360 13568 10424 13572
rect 10440 13628 10504 13632
rect 10440 13572 10444 13628
rect 10444 13572 10500 13628
rect 10500 13572 10504 13628
rect 10440 13568 10504 13572
rect 10520 13628 10584 13632
rect 10520 13572 10524 13628
rect 10524 13572 10580 13628
rect 10580 13572 10584 13628
rect 10520 13568 10584 13572
rect 10600 13628 10664 13632
rect 10600 13572 10604 13628
rect 10604 13572 10660 13628
rect 10660 13572 10664 13628
rect 10600 13568 10664 13572
rect 10680 13628 10744 13632
rect 10680 13572 10684 13628
rect 10684 13572 10740 13628
rect 10740 13572 10744 13628
rect 10680 13568 10744 13572
rect 16360 13628 16424 13632
rect 16360 13572 16364 13628
rect 16364 13572 16420 13628
rect 16420 13572 16424 13628
rect 16360 13568 16424 13572
rect 16440 13628 16504 13632
rect 16440 13572 16444 13628
rect 16444 13572 16500 13628
rect 16500 13572 16504 13628
rect 16440 13568 16504 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 1360 13084 1424 13088
rect 1360 13028 1364 13084
rect 1364 13028 1420 13084
rect 1420 13028 1424 13084
rect 1360 13024 1424 13028
rect 1440 13084 1504 13088
rect 1440 13028 1444 13084
rect 1444 13028 1500 13084
rect 1500 13028 1504 13084
rect 1440 13024 1504 13028
rect 1520 13084 1584 13088
rect 1520 13028 1524 13084
rect 1524 13028 1580 13084
rect 1580 13028 1584 13084
rect 1520 13024 1584 13028
rect 1600 13084 1664 13088
rect 1600 13028 1604 13084
rect 1604 13028 1660 13084
rect 1660 13028 1664 13084
rect 1600 13024 1664 13028
rect 1680 13084 1744 13088
rect 1680 13028 1684 13084
rect 1684 13028 1740 13084
rect 1740 13028 1744 13084
rect 1680 13024 1744 13028
rect 7360 13084 7424 13088
rect 7360 13028 7364 13084
rect 7364 13028 7420 13084
rect 7420 13028 7424 13084
rect 7360 13024 7424 13028
rect 7440 13084 7504 13088
rect 7440 13028 7444 13084
rect 7444 13028 7500 13084
rect 7500 13028 7504 13084
rect 7440 13024 7504 13028
rect 7520 13084 7584 13088
rect 7520 13028 7524 13084
rect 7524 13028 7580 13084
rect 7580 13028 7584 13084
rect 7520 13024 7584 13028
rect 7600 13084 7664 13088
rect 7600 13028 7604 13084
rect 7604 13028 7660 13084
rect 7660 13028 7664 13084
rect 7600 13024 7664 13028
rect 7680 13084 7744 13088
rect 7680 13028 7684 13084
rect 7684 13028 7740 13084
rect 7740 13028 7744 13084
rect 7680 13024 7744 13028
rect 13360 13084 13424 13088
rect 13360 13028 13364 13084
rect 13364 13028 13420 13084
rect 13420 13028 13424 13084
rect 13360 13024 13424 13028
rect 13440 13084 13504 13088
rect 13440 13028 13444 13084
rect 13444 13028 13500 13084
rect 13500 13028 13504 13084
rect 13440 13024 13504 13028
rect 13520 13084 13584 13088
rect 13520 13028 13524 13084
rect 13524 13028 13580 13084
rect 13580 13028 13584 13084
rect 13520 13024 13584 13028
rect 13600 13084 13664 13088
rect 13600 13028 13604 13084
rect 13604 13028 13660 13084
rect 13660 13028 13664 13084
rect 13600 13024 13664 13028
rect 13680 13084 13744 13088
rect 13680 13028 13684 13084
rect 13684 13028 13740 13084
rect 13740 13028 13744 13084
rect 13680 13024 13744 13028
rect 14044 12684 14108 12748
rect 8892 12548 8956 12612
rect 4360 12540 4424 12544
rect 4360 12484 4364 12540
rect 4364 12484 4420 12540
rect 4420 12484 4424 12540
rect 4360 12480 4424 12484
rect 4440 12540 4504 12544
rect 4440 12484 4444 12540
rect 4444 12484 4500 12540
rect 4500 12484 4504 12540
rect 4440 12480 4504 12484
rect 4520 12540 4584 12544
rect 4520 12484 4524 12540
rect 4524 12484 4580 12540
rect 4580 12484 4584 12540
rect 4520 12480 4584 12484
rect 4600 12540 4664 12544
rect 4600 12484 4604 12540
rect 4604 12484 4660 12540
rect 4660 12484 4664 12540
rect 4600 12480 4664 12484
rect 4680 12540 4744 12544
rect 4680 12484 4684 12540
rect 4684 12484 4740 12540
rect 4740 12484 4744 12540
rect 4680 12480 4744 12484
rect 10360 12540 10424 12544
rect 10360 12484 10364 12540
rect 10364 12484 10420 12540
rect 10420 12484 10424 12540
rect 10360 12480 10424 12484
rect 10440 12540 10504 12544
rect 10440 12484 10444 12540
rect 10444 12484 10500 12540
rect 10500 12484 10504 12540
rect 10440 12480 10504 12484
rect 10520 12540 10584 12544
rect 10520 12484 10524 12540
rect 10524 12484 10580 12540
rect 10580 12484 10584 12540
rect 10520 12480 10584 12484
rect 10600 12540 10664 12544
rect 10600 12484 10604 12540
rect 10604 12484 10660 12540
rect 10660 12484 10664 12540
rect 10600 12480 10664 12484
rect 10680 12540 10744 12544
rect 10680 12484 10684 12540
rect 10684 12484 10740 12540
rect 10740 12484 10744 12540
rect 10680 12480 10744 12484
rect 16360 12540 16424 12544
rect 16360 12484 16364 12540
rect 16364 12484 16420 12540
rect 16420 12484 16424 12540
rect 16360 12480 16424 12484
rect 16440 12540 16504 12544
rect 16440 12484 16444 12540
rect 16444 12484 16500 12540
rect 16500 12484 16504 12540
rect 16440 12480 16504 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 1360 11996 1424 12000
rect 1360 11940 1364 11996
rect 1364 11940 1420 11996
rect 1420 11940 1424 11996
rect 1360 11936 1424 11940
rect 1440 11996 1504 12000
rect 1440 11940 1444 11996
rect 1444 11940 1500 11996
rect 1500 11940 1504 11996
rect 1440 11936 1504 11940
rect 1520 11996 1584 12000
rect 1520 11940 1524 11996
rect 1524 11940 1580 11996
rect 1580 11940 1584 11996
rect 1520 11936 1584 11940
rect 1600 11996 1664 12000
rect 1600 11940 1604 11996
rect 1604 11940 1660 11996
rect 1660 11940 1664 11996
rect 1600 11936 1664 11940
rect 1680 11996 1744 12000
rect 1680 11940 1684 11996
rect 1684 11940 1740 11996
rect 1740 11940 1744 11996
rect 1680 11936 1744 11940
rect 7360 11996 7424 12000
rect 7360 11940 7364 11996
rect 7364 11940 7420 11996
rect 7420 11940 7424 11996
rect 7360 11936 7424 11940
rect 7440 11996 7504 12000
rect 7440 11940 7444 11996
rect 7444 11940 7500 11996
rect 7500 11940 7504 11996
rect 7440 11936 7504 11940
rect 7520 11996 7584 12000
rect 7520 11940 7524 11996
rect 7524 11940 7580 11996
rect 7580 11940 7584 11996
rect 7520 11936 7584 11940
rect 7600 11996 7664 12000
rect 7600 11940 7604 11996
rect 7604 11940 7660 11996
rect 7660 11940 7664 11996
rect 7600 11936 7664 11940
rect 7680 11996 7744 12000
rect 7680 11940 7684 11996
rect 7684 11940 7740 11996
rect 7740 11940 7744 11996
rect 7680 11936 7744 11940
rect 13360 11996 13424 12000
rect 13360 11940 13364 11996
rect 13364 11940 13420 11996
rect 13420 11940 13424 11996
rect 13360 11936 13424 11940
rect 13440 11996 13504 12000
rect 13440 11940 13444 11996
rect 13444 11940 13500 11996
rect 13500 11940 13504 11996
rect 13440 11936 13504 11940
rect 13520 11996 13584 12000
rect 13520 11940 13524 11996
rect 13524 11940 13580 11996
rect 13580 11940 13584 11996
rect 13520 11936 13584 11940
rect 13600 11996 13664 12000
rect 13600 11940 13604 11996
rect 13604 11940 13660 11996
rect 13660 11940 13664 11996
rect 13600 11936 13664 11940
rect 13680 11996 13744 12000
rect 13680 11940 13684 11996
rect 13684 11940 13740 11996
rect 13740 11940 13744 11996
rect 13680 11936 13744 11940
rect 12756 11732 12820 11796
rect 4360 11452 4424 11456
rect 4360 11396 4364 11452
rect 4364 11396 4420 11452
rect 4420 11396 4424 11452
rect 4360 11392 4424 11396
rect 4440 11452 4504 11456
rect 4440 11396 4444 11452
rect 4444 11396 4500 11452
rect 4500 11396 4504 11452
rect 4440 11392 4504 11396
rect 4520 11452 4584 11456
rect 4520 11396 4524 11452
rect 4524 11396 4580 11452
rect 4580 11396 4584 11452
rect 4520 11392 4584 11396
rect 4600 11452 4664 11456
rect 4600 11396 4604 11452
rect 4604 11396 4660 11452
rect 4660 11396 4664 11452
rect 4600 11392 4664 11396
rect 4680 11452 4744 11456
rect 4680 11396 4684 11452
rect 4684 11396 4740 11452
rect 4740 11396 4744 11452
rect 4680 11392 4744 11396
rect 10360 11452 10424 11456
rect 10360 11396 10364 11452
rect 10364 11396 10420 11452
rect 10420 11396 10424 11452
rect 10360 11392 10424 11396
rect 10440 11452 10504 11456
rect 10440 11396 10444 11452
rect 10444 11396 10500 11452
rect 10500 11396 10504 11452
rect 10440 11392 10504 11396
rect 10520 11452 10584 11456
rect 10520 11396 10524 11452
rect 10524 11396 10580 11452
rect 10580 11396 10584 11452
rect 10520 11392 10584 11396
rect 10600 11452 10664 11456
rect 10600 11396 10604 11452
rect 10604 11396 10660 11452
rect 10660 11396 10664 11452
rect 10600 11392 10664 11396
rect 10680 11452 10744 11456
rect 10680 11396 10684 11452
rect 10684 11396 10740 11452
rect 10740 11396 10744 11452
rect 10680 11392 10744 11396
rect 16360 11452 16424 11456
rect 16360 11396 16364 11452
rect 16364 11396 16420 11452
rect 16420 11396 16424 11452
rect 16360 11392 16424 11396
rect 16440 11452 16504 11456
rect 16440 11396 16444 11452
rect 16444 11396 16500 11452
rect 16500 11396 16504 11452
rect 16440 11392 16504 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 12204 11112 12268 11116
rect 12204 11056 12254 11112
rect 12254 11056 12268 11112
rect 12204 11052 12268 11056
rect 8892 10916 8956 10980
rect 1360 10908 1424 10912
rect 1360 10852 1364 10908
rect 1364 10852 1420 10908
rect 1420 10852 1424 10908
rect 1360 10848 1424 10852
rect 1440 10908 1504 10912
rect 1440 10852 1444 10908
rect 1444 10852 1500 10908
rect 1500 10852 1504 10908
rect 1440 10848 1504 10852
rect 1520 10908 1584 10912
rect 1520 10852 1524 10908
rect 1524 10852 1580 10908
rect 1580 10852 1584 10908
rect 1520 10848 1584 10852
rect 1600 10908 1664 10912
rect 1600 10852 1604 10908
rect 1604 10852 1660 10908
rect 1660 10852 1664 10908
rect 1600 10848 1664 10852
rect 1680 10908 1744 10912
rect 1680 10852 1684 10908
rect 1684 10852 1740 10908
rect 1740 10852 1744 10908
rect 1680 10848 1744 10852
rect 7360 10908 7424 10912
rect 7360 10852 7364 10908
rect 7364 10852 7420 10908
rect 7420 10852 7424 10908
rect 7360 10848 7424 10852
rect 7440 10908 7504 10912
rect 7440 10852 7444 10908
rect 7444 10852 7500 10908
rect 7500 10852 7504 10908
rect 7440 10848 7504 10852
rect 7520 10908 7584 10912
rect 7520 10852 7524 10908
rect 7524 10852 7580 10908
rect 7580 10852 7584 10908
rect 7520 10848 7584 10852
rect 7600 10908 7664 10912
rect 7600 10852 7604 10908
rect 7604 10852 7660 10908
rect 7660 10852 7664 10908
rect 7600 10848 7664 10852
rect 7680 10908 7744 10912
rect 7680 10852 7684 10908
rect 7684 10852 7740 10908
rect 7740 10852 7744 10908
rect 7680 10848 7744 10852
rect 13360 10908 13424 10912
rect 13360 10852 13364 10908
rect 13364 10852 13420 10908
rect 13420 10852 13424 10908
rect 13360 10848 13424 10852
rect 13440 10908 13504 10912
rect 13440 10852 13444 10908
rect 13444 10852 13500 10908
rect 13500 10852 13504 10908
rect 13440 10848 13504 10852
rect 13520 10908 13584 10912
rect 13520 10852 13524 10908
rect 13524 10852 13580 10908
rect 13580 10852 13584 10908
rect 13520 10848 13584 10852
rect 13600 10908 13664 10912
rect 13600 10852 13604 10908
rect 13604 10852 13660 10908
rect 13660 10852 13664 10908
rect 13600 10848 13664 10852
rect 13680 10908 13744 10912
rect 13680 10852 13684 10908
rect 13684 10852 13740 10908
rect 13740 10852 13744 10908
rect 13680 10848 13744 10852
rect 4360 10364 4424 10368
rect 4360 10308 4364 10364
rect 4364 10308 4420 10364
rect 4420 10308 4424 10364
rect 4360 10304 4424 10308
rect 4440 10364 4504 10368
rect 4440 10308 4444 10364
rect 4444 10308 4500 10364
rect 4500 10308 4504 10364
rect 4440 10304 4504 10308
rect 4520 10364 4584 10368
rect 4520 10308 4524 10364
rect 4524 10308 4580 10364
rect 4580 10308 4584 10364
rect 4520 10304 4584 10308
rect 4600 10364 4664 10368
rect 4600 10308 4604 10364
rect 4604 10308 4660 10364
rect 4660 10308 4664 10364
rect 4600 10304 4664 10308
rect 4680 10364 4744 10368
rect 4680 10308 4684 10364
rect 4684 10308 4740 10364
rect 4740 10308 4744 10364
rect 4680 10304 4744 10308
rect 10360 10364 10424 10368
rect 10360 10308 10364 10364
rect 10364 10308 10420 10364
rect 10420 10308 10424 10364
rect 10360 10304 10424 10308
rect 10440 10364 10504 10368
rect 10440 10308 10444 10364
rect 10444 10308 10500 10364
rect 10500 10308 10504 10364
rect 10440 10304 10504 10308
rect 10520 10364 10584 10368
rect 10520 10308 10524 10364
rect 10524 10308 10580 10364
rect 10580 10308 10584 10364
rect 10520 10304 10584 10308
rect 10600 10364 10664 10368
rect 10600 10308 10604 10364
rect 10604 10308 10660 10364
rect 10660 10308 10664 10364
rect 10600 10304 10664 10308
rect 10680 10364 10744 10368
rect 10680 10308 10684 10364
rect 10684 10308 10740 10364
rect 10740 10308 10744 10364
rect 10680 10304 10744 10308
rect 16360 10364 16424 10368
rect 16360 10308 16364 10364
rect 16364 10308 16420 10364
rect 16420 10308 16424 10364
rect 16360 10304 16424 10308
rect 16440 10364 16504 10368
rect 16440 10308 16444 10364
rect 16444 10308 16500 10364
rect 16500 10308 16504 10364
rect 16440 10304 16504 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 1360 9820 1424 9824
rect 1360 9764 1364 9820
rect 1364 9764 1420 9820
rect 1420 9764 1424 9820
rect 1360 9760 1424 9764
rect 1440 9820 1504 9824
rect 1440 9764 1444 9820
rect 1444 9764 1500 9820
rect 1500 9764 1504 9820
rect 1440 9760 1504 9764
rect 1520 9820 1584 9824
rect 1520 9764 1524 9820
rect 1524 9764 1580 9820
rect 1580 9764 1584 9820
rect 1520 9760 1584 9764
rect 1600 9820 1664 9824
rect 1600 9764 1604 9820
rect 1604 9764 1660 9820
rect 1660 9764 1664 9820
rect 1600 9760 1664 9764
rect 1680 9820 1744 9824
rect 1680 9764 1684 9820
rect 1684 9764 1740 9820
rect 1740 9764 1744 9820
rect 1680 9760 1744 9764
rect 7360 9820 7424 9824
rect 7360 9764 7364 9820
rect 7364 9764 7420 9820
rect 7420 9764 7424 9820
rect 7360 9760 7424 9764
rect 7440 9820 7504 9824
rect 7440 9764 7444 9820
rect 7444 9764 7500 9820
rect 7500 9764 7504 9820
rect 7440 9760 7504 9764
rect 7520 9820 7584 9824
rect 7520 9764 7524 9820
rect 7524 9764 7580 9820
rect 7580 9764 7584 9820
rect 7520 9760 7584 9764
rect 7600 9820 7664 9824
rect 7600 9764 7604 9820
rect 7604 9764 7660 9820
rect 7660 9764 7664 9820
rect 7600 9760 7664 9764
rect 7680 9820 7744 9824
rect 7680 9764 7684 9820
rect 7684 9764 7740 9820
rect 7740 9764 7744 9820
rect 7680 9760 7744 9764
rect 13360 9820 13424 9824
rect 13360 9764 13364 9820
rect 13364 9764 13420 9820
rect 13420 9764 13424 9820
rect 13360 9760 13424 9764
rect 13440 9820 13504 9824
rect 13440 9764 13444 9820
rect 13444 9764 13500 9820
rect 13500 9764 13504 9820
rect 13440 9760 13504 9764
rect 13520 9820 13584 9824
rect 13520 9764 13524 9820
rect 13524 9764 13580 9820
rect 13580 9764 13584 9820
rect 13520 9760 13584 9764
rect 13600 9820 13664 9824
rect 13600 9764 13604 9820
rect 13604 9764 13660 9820
rect 13660 9764 13664 9820
rect 13600 9760 13664 9764
rect 13680 9820 13744 9824
rect 13680 9764 13684 9820
rect 13684 9764 13740 9820
rect 13740 9764 13744 9820
rect 13680 9760 13744 9764
rect 4360 9276 4424 9280
rect 4360 9220 4364 9276
rect 4364 9220 4420 9276
rect 4420 9220 4424 9276
rect 4360 9216 4424 9220
rect 4440 9276 4504 9280
rect 4440 9220 4444 9276
rect 4444 9220 4500 9276
rect 4500 9220 4504 9276
rect 4440 9216 4504 9220
rect 4520 9276 4584 9280
rect 4520 9220 4524 9276
rect 4524 9220 4580 9276
rect 4580 9220 4584 9276
rect 4520 9216 4584 9220
rect 4600 9276 4664 9280
rect 4600 9220 4604 9276
rect 4604 9220 4660 9276
rect 4660 9220 4664 9276
rect 4600 9216 4664 9220
rect 4680 9276 4744 9280
rect 4680 9220 4684 9276
rect 4684 9220 4740 9276
rect 4740 9220 4744 9276
rect 4680 9216 4744 9220
rect 10360 9276 10424 9280
rect 10360 9220 10364 9276
rect 10364 9220 10420 9276
rect 10420 9220 10424 9276
rect 10360 9216 10424 9220
rect 10440 9276 10504 9280
rect 10440 9220 10444 9276
rect 10444 9220 10500 9276
rect 10500 9220 10504 9276
rect 10440 9216 10504 9220
rect 10520 9276 10584 9280
rect 10520 9220 10524 9276
rect 10524 9220 10580 9276
rect 10580 9220 10584 9276
rect 10520 9216 10584 9220
rect 10600 9276 10664 9280
rect 10600 9220 10604 9276
rect 10604 9220 10660 9276
rect 10660 9220 10664 9276
rect 10600 9216 10664 9220
rect 10680 9276 10744 9280
rect 10680 9220 10684 9276
rect 10684 9220 10740 9276
rect 10740 9220 10744 9276
rect 10680 9216 10744 9220
rect 16360 9276 16424 9280
rect 16360 9220 16364 9276
rect 16364 9220 16420 9276
rect 16420 9220 16424 9276
rect 16360 9216 16424 9220
rect 16440 9276 16504 9280
rect 16440 9220 16444 9276
rect 16444 9220 16500 9276
rect 16500 9220 16504 9276
rect 16440 9216 16504 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 1360 8732 1424 8736
rect 1360 8676 1364 8732
rect 1364 8676 1420 8732
rect 1420 8676 1424 8732
rect 1360 8672 1424 8676
rect 1440 8732 1504 8736
rect 1440 8676 1444 8732
rect 1444 8676 1500 8732
rect 1500 8676 1504 8732
rect 1440 8672 1504 8676
rect 1520 8732 1584 8736
rect 1520 8676 1524 8732
rect 1524 8676 1580 8732
rect 1580 8676 1584 8732
rect 1520 8672 1584 8676
rect 1600 8732 1664 8736
rect 1600 8676 1604 8732
rect 1604 8676 1660 8732
rect 1660 8676 1664 8732
rect 1600 8672 1664 8676
rect 1680 8732 1744 8736
rect 1680 8676 1684 8732
rect 1684 8676 1740 8732
rect 1740 8676 1744 8732
rect 1680 8672 1744 8676
rect 7360 8732 7424 8736
rect 7360 8676 7364 8732
rect 7364 8676 7420 8732
rect 7420 8676 7424 8732
rect 7360 8672 7424 8676
rect 7440 8732 7504 8736
rect 7440 8676 7444 8732
rect 7444 8676 7500 8732
rect 7500 8676 7504 8732
rect 7440 8672 7504 8676
rect 7520 8732 7584 8736
rect 7520 8676 7524 8732
rect 7524 8676 7580 8732
rect 7580 8676 7584 8732
rect 7520 8672 7584 8676
rect 7600 8732 7664 8736
rect 7600 8676 7604 8732
rect 7604 8676 7660 8732
rect 7660 8676 7664 8732
rect 7600 8672 7664 8676
rect 7680 8732 7744 8736
rect 7680 8676 7684 8732
rect 7684 8676 7740 8732
rect 7740 8676 7744 8732
rect 7680 8672 7744 8676
rect 13360 8732 13424 8736
rect 13360 8676 13364 8732
rect 13364 8676 13420 8732
rect 13420 8676 13424 8732
rect 13360 8672 13424 8676
rect 13440 8732 13504 8736
rect 13440 8676 13444 8732
rect 13444 8676 13500 8732
rect 13500 8676 13504 8732
rect 13440 8672 13504 8676
rect 13520 8732 13584 8736
rect 13520 8676 13524 8732
rect 13524 8676 13580 8732
rect 13580 8676 13584 8732
rect 13520 8672 13584 8676
rect 13600 8732 13664 8736
rect 13600 8676 13604 8732
rect 13604 8676 13660 8732
rect 13660 8676 13664 8732
rect 13600 8672 13664 8676
rect 13680 8732 13744 8736
rect 13680 8676 13684 8732
rect 13684 8676 13740 8732
rect 13740 8676 13744 8732
rect 13680 8672 13744 8676
rect 4360 8188 4424 8192
rect 4360 8132 4364 8188
rect 4364 8132 4420 8188
rect 4420 8132 4424 8188
rect 4360 8128 4424 8132
rect 4440 8188 4504 8192
rect 4440 8132 4444 8188
rect 4444 8132 4500 8188
rect 4500 8132 4504 8188
rect 4440 8128 4504 8132
rect 4520 8188 4584 8192
rect 4520 8132 4524 8188
rect 4524 8132 4580 8188
rect 4580 8132 4584 8188
rect 4520 8128 4584 8132
rect 4600 8188 4664 8192
rect 4600 8132 4604 8188
rect 4604 8132 4660 8188
rect 4660 8132 4664 8188
rect 4600 8128 4664 8132
rect 4680 8188 4744 8192
rect 4680 8132 4684 8188
rect 4684 8132 4740 8188
rect 4740 8132 4744 8188
rect 4680 8128 4744 8132
rect 10360 8188 10424 8192
rect 10360 8132 10364 8188
rect 10364 8132 10420 8188
rect 10420 8132 10424 8188
rect 10360 8128 10424 8132
rect 10440 8188 10504 8192
rect 10440 8132 10444 8188
rect 10444 8132 10500 8188
rect 10500 8132 10504 8188
rect 10440 8128 10504 8132
rect 10520 8188 10584 8192
rect 10520 8132 10524 8188
rect 10524 8132 10580 8188
rect 10580 8132 10584 8188
rect 10520 8128 10584 8132
rect 10600 8188 10664 8192
rect 10600 8132 10604 8188
rect 10604 8132 10660 8188
rect 10660 8132 10664 8188
rect 10600 8128 10664 8132
rect 10680 8188 10744 8192
rect 10680 8132 10684 8188
rect 10684 8132 10740 8188
rect 10740 8132 10744 8188
rect 10680 8128 10744 8132
rect 16360 8188 16424 8192
rect 16360 8132 16364 8188
rect 16364 8132 16420 8188
rect 16420 8132 16424 8188
rect 16360 8128 16424 8132
rect 16440 8188 16504 8192
rect 16440 8132 16444 8188
rect 16444 8132 16500 8188
rect 16500 8132 16504 8188
rect 16440 8128 16504 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 1360 7644 1424 7648
rect 1360 7588 1364 7644
rect 1364 7588 1420 7644
rect 1420 7588 1424 7644
rect 1360 7584 1424 7588
rect 1440 7644 1504 7648
rect 1440 7588 1444 7644
rect 1444 7588 1500 7644
rect 1500 7588 1504 7644
rect 1440 7584 1504 7588
rect 1520 7644 1584 7648
rect 1520 7588 1524 7644
rect 1524 7588 1580 7644
rect 1580 7588 1584 7644
rect 1520 7584 1584 7588
rect 1600 7644 1664 7648
rect 1600 7588 1604 7644
rect 1604 7588 1660 7644
rect 1660 7588 1664 7644
rect 1600 7584 1664 7588
rect 1680 7644 1744 7648
rect 1680 7588 1684 7644
rect 1684 7588 1740 7644
rect 1740 7588 1744 7644
rect 1680 7584 1744 7588
rect 7360 7644 7424 7648
rect 7360 7588 7364 7644
rect 7364 7588 7420 7644
rect 7420 7588 7424 7644
rect 7360 7584 7424 7588
rect 7440 7644 7504 7648
rect 7440 7588 7444 7644
rect 7444 7588 7500 7644
rect 7500 7588 7504 7644
rect 7440 7584 7504 7588
rect 7520 7644 7584 7648
rect 7520 7588 7524 7644
rect 7524 7588 7580 7644
rect 7580 7588 7584 7644
rect 7520 7584 7584 7588
rect 7600 7644 7664 7648
rect 7600 7588 7604 7644
rect 7604 7588 7660 7644
rect 7660 7588 7664 7644
rect 7600 7584 7664 7588
rect 7680 7644 7744 7648
rect 7680 7588 7684 7644
rect 7684 7588 7740 7644
rect 7740 7588 7744 7644
rect 7680 7584 7744 7588
rect 13360 7644 13424 7648
rect 13360 7588 13364 7644
rect 13364 7588 13420 7644
rect 13420 7588 13424 7644
rect 13360 7584 13424 7588
rect 13440 7644 13504 7648
rect 13440 7588 13444 7644
rect 13444 7588 13500 7644
rect 13500 7588 13504 7644
rect 13440 7584 13504 7588
rect 13520 7644 13584 7648
rect 13520 7588 13524 7644
rect 13524 7588 13580 7644
rect 13580 7588 13584 7644
rect 13520 7584 13584 7588
rect 13600 7644 13664 7648
rect 13600 7588 13604 7644
rect 13604 7588 13660 7644
rect 13660 7588 13664 7644
rect 13600 7584 13664 7588
rect 13680 7644 13744 7648
rect 13680 7588 13684 7644
rect 13684 7588 13740 7644
rect 13740 7588 13744 7644
rect 13680 7584 13744 7588
rect 5948 7380 6012 7444
rect 14044 7380 14108 7444
rect 13860 7108 13924 7172
rect 4360 7100 4424 7104
rect 4360 7044 4364 7100
rect 4364 7044 4420 7100
rect 4420 7044 4424 7100
rect 4360 7040 4424 7044
rect 4440 7100 4504 7104
rect 4440 7044 4444 7100
rect 4444 7044 4500 7100
rect 4500 7044 4504 7100
rect 4440 7040 4504 7044
rect 4520 7100 4584 7104
rect 4520 7044 4524 7100
rect 4524 7044 4580 7100
rect 4580 7044 4584 7100
rect 4520 7040 4584 7044
rect 4600 7100 4664 7104
rect 4600 7044 4604 7100
rect 4604 7044 4660 7100
rect 4660 7044 4664 7100
rect 4600 7040 4664 7044
rect 4680 7100 4744 7104
rect 4680 7044 4684 7100
rect 4684 7044 4740 7100
rect 4740 7044 4744 7100
rect 4680 7040 4744 7044
rect 10360 7100 10424 7104
rect 10360 7044 10364 7100
rect 10364 7044 10420 7100
rect 10420 7044 10424 7100
rect 10360 7040 10424 7044
rect 10440 7100 10504 7104
rect 10440 7044 10444 7100
rect 10444 7044 10500 7100
rect 10500 7044 10504 7100
rect 10440 7040 10504 7044
rect 10520 7100 10584 7104
rect 10520 7044 10524 7100
rect 10524 7044 10580 7100
rect 10580 7044 10584 7100
rect 10520 7040 10584 7044
rect 10600 7100 10664 7104
rect 10600 7044 10604 7100
rect 10604 7044 10660 7100
rect 10660 7044 10664 7100
rect 10600 7040 10664 7044
rect 10680 7100 10744 7104
rect 10680 7044 10684 7100
rect 10684 7044 10740 7100
rect 10740 7044 10744 7100
rect 10680 7040 10744 7044
rect 16360 7100 16424 7104
rect 16360 7044 16364 7100
rect 16364 7044 16420 7100
rect 16420 7044 16424 7100
rect 16360 7040 16424 7044
rect 16440 7100 16504 7104
rect 16440 7044 16444 7100
rect 16444 7044 16500 7100
rect 16500 7044 16504 7100
rect 16440 7040 16504 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 14780 6972 14844 7036
rect 9812 6564 9876 6628
rect 1360 6556 1424 6560
rect 1360 6500 1364 6556
rect 1364 6500 1420 6556
rect 1420 6500 1424 6556
rect 1360 6496 1424 6500
rect 1440 6556 1504 6560
rect 1440 6500 1444 6556
rect 1444 6500 1500 6556
rect 1500 6500 1504 6556
rect 1440 6496 1504 6500
rect 1520 6556 1584 6560
rect 1520 6500 1524 6556
rect 1524 6500 1580 6556
rect 1580 6500 1584 6556
rect 1520 6496 1584 6500
rect 1600 6556 1664 6560
rect 1600 6500 1604 6556
rect 1604 6500 1660 6556
rect 1660 6500 1664 6556
rect 1600 6496 1664 6500
rect 1680 6556 1744 6560
rect 1680 6500 1684 6556
rect 1684 6500 1740 6556
rect 1740 6500 1744 6556
rect 1680 6496 1744 6500
rect 7360 6556 7424 6560
rect 7360 6500 7364 6556
rect 7364 6500 7420 6556
rect 7420 6500 7424 6556
rect 7360 6496 7424 6500
rect 7440 6556 7504 6560
rect 7440 6500 7444 6556
rect 7444 6500 7500 6556
rect 7500 6500 7504 6556
rect 7440 6496 7504 6500
rect 7520 6556 7584 6560
rect 7520 6500 7524 6556
rect 7524 6500 7580 6556
rect 7580 6500 7584 6556
rect 7520 6496 7584 6500
rect 7600 6556 7664 6560
rect 7600 6500 7604 6556
rect 7604 6500 7660 6556
rect 7660 6500 7664 6556
rect 7600 6496 7664 6500
rect 7680 6556 7744 6560
rect 7680 6500 7684 6556
rect 7684 6500 7740 6556
rect 7740 6500 7744 6556
rect 7680 6496 7744 6500
rect 13360 6556 13424 6560
rect 13360 6500 13364 6556
rect 13364 6500 13420 6556
rect 13420 6500 13424 6556
rect 13360 6496 13424 6500
rect 13440 6556 13504 6560
rect 13440 6500 13444 6556
rect 13444 6500 13500 6556
rect 13500 6500 13504 6556
rect 13440 6496 13504 6500
rect 13520 6556 13584 6560
rect 13520 6500 13524 6556
rect 13524 6500 13580 6556
rect 13580 6500 13584 6556
rect 13520 6496 13584 6500
rect 13600 6556 13664 6560
rect 13600 6500 13604 6556
rect 13604 6500 13660 6556
rect 13660 6500 13664 6556
rect 13600 6496 13664 6500
rect 13680 6556 13744 6560
rect 13680 6500 13684 6556
rect 13684 6500 13740 6556
rect 13740 6500 13744 6556
rect 13680 6496 13744 6500
rect 13860 6156 13924 6220
rect 4360 6012 4424 6016
rect 4360 5956 4364 6012
rect 4364 5956 4420 6012
rect 4420 5956 4424 6012
rect 4360 5952 4424 5956
rect 4440 6012 4504 6016
rect 4440 5956 4444 6012
rect 4444 5956 4500 6012
rect 4500 5956 4504 6012
rect 4440 5952 4504 5956
rect 4520 6012 4584 6016
rect 4520 5956 4524 6012
rect 4524 5956 4580 6012
rect 4580 5956 4584 6012
rect 4520 5952 4584 5956
rect 4600 6012 4664 6016
rect 4600 5956 4604 6012
rect 4604 5956 4660 6012
rect 4660 5956 4664 6012
rect 4600 5952 4664 5956
rect 4680 6012 4744 6016
rect 4680 5956 4684 6012
rect 4684 5956 4740 6012
rect 4740 5956 4744 6012
rect 4680 5952 4744 5956
rect 10360 6012 10424 6016
rect 10360 5956 10364 6012
rect 10364 5956 10420 6012
rect 10420 5956 10424 6012
rect 10360 5952 10424 5956
rect 10440 6012 10504 6016
rect 10440 5956 10444 6012
rect 10444 5956 10500 6012
rect 10500 5956 10504 6012
rect 10440 5952 10504 5956
rect 10520 6012 10584 6016
rect 10520 5956 10524 6012
rect 10524 5956 10580 6012
rect 10580 5956 10584 6012
rect 10520 5952 10584 5956
rect 10600 6012 10664 6016
rect 10600 5956 10604 6012
rect 10604 5956 10660 6012
rect 10660 5956 10664 6012
rect 10600 5952 10664 5956
rect 10680 6012 10744 6016
rect 10680 5956 10684 6012
rect 10684 5956 10740 6012
rect 10740 5956 10744 6012
rect 10680 5952 10744 5956
rect 16360 6012 16424 6016
rect 16360 5956 16364 6012
rect 16364 5956 16420 6012
rect 16420 5956 16424 6012
rect 16360 5952 16424 5956
rect 16440 6012 16504 6016
rect 16440 5956 16444 6012
rect 16444 5956 16500 6012
rect 16500 5956 16504 6012
rect 16440 5952 16504 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 12756 5884 12820 5948
rect 1360 5468 1424 5472
rect 1360 5412 1364 5468
rect 1364 5412 1420 5468
rect 1420 5412 1424 5468
rect 1360 5408 1424 5412
rect 1440 5468 1504 5472
rect 1440 5412 1444 5468
rect 1444 5412 1500 5468
rect 1500 5412 1504 5468
rect 1440 5408 1504 5412
rect 1520 5468 1584 5472
rect 1520 5412 1524 5468
rect 1524 5412 1580 5468
rect 1580 5412 1584 5468
rect 1520 5408 1584 5412
rect 1600 5468 1664 5472
rect 1600 5412 1604 5468
rect 1604 5412 1660 5468
rect 1660 5412 1664 5468
rect 1600 5408 1664 5412
rect 1680 5468 1744 5472
rect 1680 5412 1684 5468
rect 1684 5412 1740 5468
rect 1740 5412 1744 5468
rect 1680 5408 1744 5412
rect 7360 5468 7424 5472
rect 7360 5412 7364 5468
rect 7364 5412 7420 5468
rect 7420 5412 7424 5468
rect 7360 5408 7424 5412
rect 7440 5468 7504 5472
rect 7440 5412 7444 5468
rect 7444 5412 7500 5468
rect 7500 5412 7504 5468
rect 7440 5408 7504 5412
rect 7520 5468 7584 5472
rect 7520 5412 7524 5468
rect 7524 5412 7580 5468
rect 7580 5412 7584 5468
rect 7520 5408 7584 5412
rect 7600 5468 7664 5472
rect 7600 5412 7604 5468
rect 7604 5412 7660 5468
rect 7660 5412 7664 5468
rect 7600 5408 7664 5412
rect 7680 5468 7744 5472
rect 7680 5412 7684 5468
rect 7684 5412 7740 5468
rect 7740 5412 7744 5468
rect 7680 5408 7744 5412
rect 13360 5468 13424 5472
rect 13360 5412 13364 5468
rect 13364 5412 13420 5468
rect 13420 5412 13424 5468
rect 13360 5408 13424 5412
rect 13440 5468 13504 5472
rect 13440 5412 13444 5468
rect 13444 5412 13500 5468
rect 13500 5412 13504 5468
rect 13440 5408 13504 5412
rect 13520 5468 13584 5472
rect 13520 5412 13524 5468
rect 13524 5412 13580 5468
rect 13580 5412 13584 5468
rect 13520 5408 13584 5412
rect 13600 5468 13664 5472
rect 13600 5412 13604 5468
rect 13604 5412 13660 5468
rect 13660 5412 13664 5468
rect 13600 5408 13664 5412
rect 13680 5468 13744 5472
rect 13680 5412 13684 5468
rect 13684 5412 13740 5468
rect 13740 5412 13744 5468
rect 13680 5408 13744 5412
rect 9996 5204 10060 5268
rect 4360 4924 4424 4928
rect 4360 4868 4364 4924
rect 4364 4868 4420 4924
rect 4420 4868 4424 4924
rect 4360 4864 4424 4868
rect 4440 4924 4504 4928
rect 4440 4868 4444 4924
rect 4444 4868 4500 4924
rect 4500 4868 4504 4924
rect 4440 4864 4504 4868
rect 4520 4924 4584 4928
rect 4520 4868 4524 4924
rect 4524 4868 4580 4924
rect 4580 4868 4584 4924
rect 4520 4864 4584 4868
rect 4600 4924 4664 4928
rect 4600 4868 4604 4924
rect 4604 4868 4660 4924
rect 4660 4868 4664 4924
rect 4600 4864 4664 4868
rect 4680 4924 4744 4928
rect 4680 4868 4684 4924
rect 4684 4868 4740 4924
rect 4740 4868 4744 4924
rect 4680 4864 4744 4868
rect 7972 4932 8036 4996
rect 10360 4924 10424 4928
rect 10360 4868 10364 4924
rect 10364 4868 10420 4924
rect 10420 4868 10424 4924
rect 10360 4864 10424 4868
rect 10440 4924 10504 4928
rect 10440 4868 10444 4924
rect 10444 4868 10500 4924
rect 10500 4868 10504 4924
rect 10440 4864 10504 4868
rect 10520 4924 10584 4928
rect 10520 4868 10524 4924
rect 10524 4868 10580 4924
rect 10580 4868 10584 4924
rect 10520 4864 10584 4868
rect 10600 4924 10664 4928
rect 10600 4868 10604 4924
rect 10604 4868 10660 4924
rect 10660 4868 10664 4924
rect 10600 4864 10664 4868
rect 10680 4924 10744 4928
rect 10680 4868 10684 4924
rect 10684 4868 10740 4924
rect 10740 4868 10744 4924
rect 10680 4864 10744 4868
rect 16360 4924 16424 4928
rect 16360 4868 16364 4924
rect 16364 4868 16420 4924
rect 16420 4868 16424 4924
rect 16360 4864 16424 4868
rect 16440 4924 16504 4928
rect 16440 4868 16444 4924
rect 16444 4868 16500 4924
rect 16500 4868 16504 4924
rect 16440 4864 16504 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 1360 4380 1424 4384
rect 1360 4324 1364 4380
rect 1364 4324 1420 4380
rect 1420 4324 1424 4380
rect 1360 4320 1424 4324
rect 1440 4380 1504 4384
rect 1440 4324 1444 4380
rect 1444 4324 1500 4380
rect 1500 4324 1504 4380
rect 1440 4320 1504 4324
rect 1520 4380 1584 4384
rect 1520 4324 1524 4380
rect 1524 4324 1580 4380
rect 1580 4324 1584 4380
rect 1520 4320 1584 4324
rect 1600 4380 1664 4384
rect 1600 4324 1604 4380
rect 1604 4324 1660 4380
rect 1660 4324 1664 4380
rect 1600 4320 1664 4324
rect 1680 4380 1744 4384
rect 1680 4324 1684 4380
rect 1684 4324 1740 4380
rect 1740 4324 1744 4380
rect 1680 4320 1744 4324
rect 7360 4380 7424 4384
rect 7360 4324 7364 4380
rect 7364 4324 7420 4380
rect 7420 4324 7424 4380
rect 7360 4320 7424 4324
rect 7440 4380 7504 4384
rect 7440 4324 7444 4380
rect 7444 4324 7500 4380
rect 7500 4324 7504 4380
rect 7440 4320 7504 4324
rect 7520 4380 7584 4384
rect 7520 4324 7524 4380
rect 7524 4324 7580 4380
rect 7580 4324 7584 4380
rect 7520 4320 7584 4324
rect 7600 4380 7664 4384
rect 7600 4324 7604 4380
rect 7604 4324 7660 4380
rect 7660 4324 7664 4380
rect 7600 4320 7664 4324
rect 7680 4380 7744 4384
rect 7680 4324 7684 4380
rect 7684 4324 7740 4380
rect 7740 4324 7744 4380
rect 7680 4320 7744 4324
rect 13360 4380 13424 4384
rect 13360 4324 13364 4380
rect 13364 4324 13420 4380
rect 13420 4324 13424 4380
rect 13360 4320 13424 4324
rect 13440 4380 13504 4384
rect 13440 4324 13444 4380
rect 13444 4324 13500 4380
rect 13500 4324 13504 4380
rect 13440 4320 13504 4324
rect 13520 4380 13584 4384
rect 13520 4324 13524 4380
rect 13524 4324 13580 4380
rect 13580 4324 13584 4380
rect 13520 4320 13584 4324
rect 13600 4380 13664 4384
rect 13600 4324 13604 4380
rect 13604 4324 13660 4380
rect 13660 4324 13664 4380
rect 13600 4320 13664 4324
rect 13680 4380 13744 4384
rect 13680 4324 13684 4380
rect 13684 4324 13740 4380
rect 13740 4324 13744 4380
rect 13680 4320 13744 4324
rect 15148 4040 15212 4044
rect 15148 3984 15198 4040
rect 15198 3984 15212 4040
rect 15148 3980 15212 3984
rect 12204 3844 12268 3908
rect 4360 3836 4424 3840
rect 4360 3780 4364 3836
rect 4364 3780 4420 3836
rect 4420 3780 4424 3836
rect 4360 3776 4424 3780
rect 4440 3836 4504 3840
rect 4440 3780 4444 3836
rect 4444 3780 4500 3836
rect 4500 3780 4504 3836
rect 4440 3776 4504 3780
rect 4520 3836 4584 3840
rect 4520 3780 4524 3836
rect 4524 3780 4580 3836
rect 4580 3780 4584 3836
rect 4520 3776 4584 3780
rect 4600 3836 4664 3840
rect 4600 3780 4604 3836
rect 4604 3780 4660 3836
rect 4660 3780 4664 3836
rect 4600 3776 4664 3780
rect 4680 3836 4744 3840
rect 4680 3780 4684 3836
rect 4684 3780 4740 3836
rect 4740 3780 4744 3836
rect 4680 3776 4744 3780
rect 10360 3836 10424 3840
rect 10360 3780 10364 3836
rect 10364 3780 10420 3836
rect 10420 3780 10424 3836
rect 10360 3776 10424 3780
rect 10440 3836 10504 3840
rect 10440 3780 10444 3836
rect 10444 3780 10500 3836
rect 10500 3780 10504 3836
rect 10440 3776 10504 3780
rect 10520 3836 10584 3840
rect 10520 3780 10524 3836
rect 10524 3780 10580 3836
rect 10580 3780 10584 3836
rect 10520 3776 10584 3780
rect 10600 3836 10664 3840
rect 10600 3780 10604 3836
rect 10604 3780 10660 3836
rect 10660 3780 10664 3836
rect 10600 3776 10664 3780
rect 10680 3836 10744 3840
rect 10680 3780 10684 3836
rect 10684 3780 10740 3836
rect 10740 3780 10744 3836
rect 10680 3776 10744 3780
rect 16360 3836 16424 3840
rect 16360 3780 16364 3836
rect 16364 3780 16420 3836
rect 16420 3780 16424 3836
rect 16360 3776 16424 3780
rect 16440 3836 16504 3840
rect 16440 3780 16444 3836
rect 16444 3780 16500 3836
rect 16500 3780 16504 3836
rect 16440 3776 16504 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 5948 3300 6012 3364
rect 9812 3360 9876 3364
rect 9812 3304 9826 3360
rect 9826 3304 9876 3360
rect 9812 3300 9876 3304
rect 1360 3292 1424 3296
rect 1360 3236 1364 3292
rect 1364 3236 1420 3292
rect 1420 3236 1424 3292
rect 1360 3232 1424 3236
rect 1440 3292 1504 3296
rect 1440 3236 1444 3292
rect 1444 3236 1500 3292
rect 1500 3236 1504 3292
rect 1440 3232 1504 3236
rect 1520 3292 1584 3296
rect 1520 3236 1524 3292
rect 1524 3236 1580 3292
rect 1580 3236 1584 3292
rect 1520 3232 1584 3236
rect 1600 3292 1664 3296
rect 1600 3236 1604 3292
rect 1604 3236 1660 3292
rect 1660 3236 1664 3292
rect 1600 3232 1664 3236
rect 1680 3292 1744 3296
rect 1680 3236 1684 3292
rect 1684 3236 1740 3292
rect 1740 3236 1744 3292
rect 1680 3232 1744 3236
rect 7360 3292 7424 3296
rect 7360 3236 7364 3292
rect 7364 3236 7420 3292
rect 7420 3236 7424 3292
rect 7360 3232 7424 3236
rect 7440 3292 7504 3296
rect 7440 3236 7444 3292
rect 7444 3236 7500 3292
rect 7500 3236 7504 3292
rect 7440 3232 7504 3236
rect 7520 3292 7584 3296
rect 7520 3236 7524 3292
rect 7524 3236 7580 3292
rect 7580 3236 7584 3292
rect 7520 3232 7584 3236
rect 7600 3292 7664 3296
rect 7600 3236 7604 3292
rect 7604 3236 7660 3292
rect 7660 3236 7664 3292
rect 7600 3232 7664 3236
rect 7680 3292 7744 3296
rect 7680 3236 7684 3292
rect 7684 3236 7740 3292
rect 7740 3236 7744 3292
rect 7680 3232 7744 3236
rect 13360 3292 13424 3296
rect 13360 3236 13364 3292
rect 13364 3236 13420 3292
rect 13420 3236 13424 3292
rect 13360 3232 13424 3236
rect 13440 3292 13504 3296
rect 13440 3236 13444 3292
rect 13444 3236 13500 3292
rect 13500 3236 13504 3292
rect 13440 3232 13504 3236
rect 13520 3292 13584 3296
rect 13520 3236 13524 3292
rect 13524 3236 13580 3292
rect 13580 3236 13584 3292
rect 13520 3232 13584 3236
rect 13600 3292 13664 3296
rect 13600 3236 13604 3292
rect 13604 3236 13660 3292
rect 13660 3236 13664 3292
rect 13600 3232 13664 3236
rect 13680 3292 13744 3296
rect 13680 3236 13684 3292
rect 13684 3236 13740 3292
rect 13740 3236 13744 3292
rect 13680 3232 13744 3236
rect 7972 2892 8036 2956
rect 4360 2748 4424 2752
rect 4360 2692 4364 2748
rect 4364 2692 4420 2748
rect 4420 2692 4424 2748
rect 4360 2688 4424 2692
rect 4440 2748 4504 2752
rect 4440 2692 4444 2748
rect 4444 2692 4500 2748
rect 4500 2692 4504 2748
rect 4440 2688 4504 2692
rect 4520 2748 4584 2752
rect 4520 2692 4524 2748
rect 4524 2692 4580 2748
rect 4580 2692 4584 2748
rect 4520 2688 4584 2692
rect 4600 2748 4664 2752
rect 4600 2692 4604 2748
rect 4604 2692 4660 2748
rect 4660 2692 4664 2748
rect 4600 2688 4664 2692
rect 4680 2748 4744 2752
rect 4680 2692 4684 2748
rect 4684 2692 4740 2748
rect 4740 2692 4744 2748
rect 4680 2688 4744 2692
rect 10360 2748 10424 2752
rect 10360 2692 10364 2748
rect 10364 2692 10420 2748
rect 10420 2692 10424 2748
rect 10360 2688 10424 2692
rect 10440 2748 10504 2752
rect 10440 2692 10444 2748
rect 10444 2692 10500 2748
rect 10500 2692 10504 2748
rect 10440 2688 10504 2692
rect 10520 2748 10584 2752
rect 10520 2692 10524 2748
rect 10524 2692 10580 2748
rect 10580 2692 10584 2748
rect 10520 2688 10584 2692
rect 10600 2748 10664 2752
rect 10600 2692 10604 2748
rect 10604 2692 10660 2748
rect 10660 2692 10664 2748
rect 10600 2688 10664 2692
rect 10680 2748 10744 2752
rect 10680 2692 10684 2748
rect 10684 2692 10740 2748
rect 10740 2692 10744 2748
rect 10680 2688 10744 2692
rect 16360 2748 16424 2752
rect 16360 2692 16364 2748
rect 16364 2692 16420 2748
rect 16420 2692 16424 2748
rect 16360 2688 16424 2692
rect 16440 2748 16504 2752
rect 16440 2692 16444 2748
rect 16444 2692 16500 2748
rect 16500 2692 16504 2748
rect 16440 2688 16504 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 6500 2620 6564 2684
rect 14780 2620 14844 2684
rect 6132 2408 6196 2412
rect 6132 2352 6146 2408
rect 6146 2352 6196 2408
rect 6132 2348 6196 2352
rect 9260 2348 9324 2412
rect 1360 2204 1424 2208
rect 1360 2148 1364 2204
rect 1364 2148 1420 2204
rect 1420 2148 1424 2204
rect 1360 2144 1424 2148
rect 1440 2204 1504 2208
rect 1440 2148 1444 2204
rect 1444 2148 1500 2204
rect 1500 2148 1504 2204
rect 1440 2144 1504 2148
rect 1520 2204 1584 2208
rect 1520 2148 1524 2204
rect 1524 2148 1580 2204
rect 1580 2148 1584 2204
rect 1520 2144 1584 2148
rect 1600 2204 1664 2208
rect 1600 2148 1604 2204
rect 1604 2148 1660 2204
rect 1660 2148 1664 2204
rect 1600 2144 1664 2148
rect 1680 2204 1744 2208
rect 1680 2148 1684 2204
rect 1684 2148 1740 2204
rect 1740 2148 1744 2204
rect 1680 2144 1744 2148
rect 7360 2204 7424 2208
rect 7360 2148 7364 2204
rect 7364 2148 7420 2204
rect 7420 2148 7424 2204
rect 7360 2144 7424 2148
rect 7440 2204 7504 2208
rect 7440 2148 7444 2204
rect 7444 2148 7500 2204
rect 7500 2148 7504 2204
rect 7440 2144 7504 2148
rect 7520 2204 7584 2208
rect 7520 2148 7524 2204
rect 7524 2148 7580 2204
rect 7580 2148 7584 2204
rect 7520 2144 7584 2148
rect 7600 2204 7664 2208
rect 7600 2148 7604 2204
rect 7604 2148 7660 2204
rect 7660 2148 7664 2204
rect 7600 2144 7664 2148
rect 7680 2204 7744 2208
rect 7680 2148 7684 2204
rect 7684 2148 7740 2204
rect 7740 2148 7744 2204
rect 7680 2144 7744 2148
rect 13360 2204 13424 2208
rect 13360 2148 13364 2204
rect 13364 2148 13420 2204
rect 13420 2148 13424 2204
rect 13360 2144 13424 2148
rect 13440 2204 13504 2208
rect 13440 2148 13444 2204
rect 13444 2148 13500 2204
rect 13500 2148 13504 2204
rect 13440 2144 13504 2148
rect 13520 2204 13584 2208
rect 13520 2148 13524 2204
rect 13524 2148 13580 2204
rect 13580 2148 13584 2204
rect 13520 2144 13584 2148
rect 13600 2204 13664 2208
rect 13600 2148 13604 2204
rect 13604 2148 13660 2204
rect 13660 2148 13664 2204
rect 13600 2144 13664 2148
rect 13680 2204 13744 2208
rect 13680 2148 13684 2204
rect 13684 2148 13740 2204
rect 13740 2148 13744 2204
rect 13680 2144 13744 2148
rect 4360 1660 4424 1664
rect 4360 1604 4364 1660
rect 4364 1604 4420 1660
rect 4420 1604 4424 1660
rect 4360 1600 4424 1604
rect 4440 1660 4504 1664
rect 4440 1604 4444 1660
rect 4444 1604 4500 1660
rect 4500 1604 4504 1660
rect 4440 1600 4504 1604
rect 4520 1660 4584 1664
rect 4520 1604 4524 1660
rect 4524 1604 4580 1660
rect 4580 1604 4584 1660
rect 4520 1600 4584 1604
rect 4600 1660 4664 1664
rect 4600 1604 4604 1660
rect 4604 1604 4660 1660
rect 4660 1604 4664 1660
rect 4600 1600 4664 1604
rect 4680 1660 4744 1664
rect 4680 1604 4684 1660
rect 4684 1604 4740 1660
rect 4740 1604 4744 1660
rect 4680 1600 4744 1604
rect 13124 1940 13188 2004
rect 8708 1804 8772 1868
rect 9996 1668 10060 1732
rect 10360 1660 10424 1664
rect 10360 1604 10364 1660
rect 10364 1604 10420 1660
rect 10420 1604 10424 1660
rect 10360 1600 10424 1604
rect 10440 1660 10504 1664
rect 10440 1604 10444 1660
rect 10444 1604 10500 1660
rect 10500 1604 10504 1660
rect 10440 1600 10504 1604
rect 10520 1660 10584 1664
rect 10520 1604 10524 1660
rect 10524 1604 10580 1660
rect 10580 1604 10584 1660
rect 10520 1600 10584 1604
rect 10600 1660 10664 1664
rect 10600 1604 10604 1660
rect 10604 1604 10660 1660
rect 10660 1604 10664 1660
rect 10600 1600 10664 1604
rect 10680 1660 10744 1664
rect 10680 1604 10684 1660
rect 10684 1604 10740 1660
rect 10740 1604 10744 1660
rect 10680 1600 10744 1604
rect 16360 1660 16424 1664
rect 16360 1604 16364 1660
rect 16364 1604 16420 1660
rect 16420 1604 16424 1660
rect 16360 1600 16424 1604
rect 16440 1660 16504 1664
rect 16440 1604 16444 1660
rect 16444 1604 16500 1660
rect 16500 1604 16504 1660
rect 16440 1600 16504 1604
rect 16520 1660 16584 1664
rect 16520 1604 16524 1660
rect 16524 1604 16580 1660
rect 16580 1604 16584 1660
rect 16520 1600 16584 1604
rect 16600 1660 16664 1664
rect 16600 1604 16604 1660
rect 16604 1604 16660 1660
rect 16660 1604 16664 1660
rect 16600 1600 16664 1604
rect 16680 1660 16744 1664
rect 16680 1604 16684 1660
rect 16684 1604 16740 1660
rect 16740 1604 16744 1660
rect 16680 1600 16744 1604
rect 9812 1532 9876 1596
rect 15148 1532 15212 1596
rect 9996 1260 10060 1324
rect 11284 1260 11348 1324
rect 15148 1320 15212 1324
rect 15148 1264 15162 1320
rect 15162 1264 15212 1320
rect 15148 1260 15212 1264
rect 9812 1124 9876 1188
rect 1360 1116 1424 1120
rect 1360 1060 1364 1116
rect 1364 1060 1420 1116
rect 1420 1060 1424 1116
rect 1360 1056 1424 1060
rect 1440 1116 1504 1120
rect 1440 1060 1444 1116
rect 1444 1060 1500 1116
rect 1500 1060 1504 1116
rect 1440 1056 1504 1060
rect 1520 1116 1584 1120
rect 1520 1060 1524 1116
rect 1524 1060 1580 1116
rect 1580 1060 1584 1116
rect 1520 1056 1584 1060
rect 1600 1116 1664 1120
rect 1600 1060 1604 1116
rect 1604 1060 1660 1116
rect 1660 1060 1664 1116
rect 1600 1056 1664 1060
rect 1680 1116 1744 1120
rect 1680 1060 1684 1116
rect 1684 1060 1740 1116
rect 1740 1060 1744 1116
rect 1680 1056 1744 1060
rect 7360 1116 7424 1120
rect 7360 1060 7364 1116
rect 7364 1060 7420 1116
rect 7420 1060 7424 1116
rect 7360 1056 7424 1060
rect 7440 1116 7504 1120
rect 7440 1060 7444 1116
rect 7444 1060 7500 1116
rect 7500 1060 7504 1116
rect 7440 1056 7504 1060
rect 7520 1116 7584 1120
rect 7520 1060 7524 1116
rect 7524 1060 7580 1116
rect 7580 1060 7584 1116
rect 7520 1056 7584 1060
rect 7600 1116 7664 1120
rect 7600 1060 7604 1116
rect 7604 1060 7660 1116
rect 7660 1060 7664 1116
rect 7600 1056 7664 1060
rect 7680 1116 7744 1120
rect 7680 1060 7684 1116
rect 7684 1060 7740 1116
rect 7740 1060 7744 1116
rect 7680 1056 7744 1060
rect 13360 1116 13424 1120
rect 13360 1060 13364 1116
rect 13364 1060 13420 1116
rect 13420 1060 13424 1116
rect 13360 1056 13424 1060
rect 13440 1116 13504 1120
rect 13440 1060 13444 1116
rect 13444 1060 13500 1116
rect 13500 1060 13504 1116
rect 13440 1056 13504 1060
rect 13520 1116 13584 1120
rect 13520 1060 13524 1116
rect 13524 1060 13580 1116
rect 13580 1060 13584 1116
rect 13520 1056 13584 1060
rect 13600 1116 13664 1120
rect 13600 1060 13604 1116
rect 13604 1060 13660 1116
rect 13660 1060 13664 1116
rect 13600 1056 13664 1060
rect 13680 1116 13744 1120
rect 13680 1060 13684 1116
rect 13684 1060 13740 1116
rect 13740 1060 13744 1116
rect 13680 1056 13744 1060
rect 4360 572 4424 576
rect 4360 516 4364 572
rect 4364 516 4420 572
rect 4420 516 4424 572
rect 4360 512 4424 516
rect 4440 572 4504 576
rect 4440 516 4444 572
rect 4444 516 4500 572
rect 4500 516 4504 572
rect 4440 512 4504 516
rect 4520 572 4584 576
rect 4520 516 4524 572
rect 4524 516 4580 572
rect 4580 516 4584 572
rect 4520 512 4584 516
rect 4600 572 4664 576
rect 4600 516 4604 572
rect 4604 516 4660 572
rect 4660 516 4664 572
rect 4600 512 4664 516
rect 4680 572 4744 576
rect 4680 516 4684 572
rect 4684 516 4740 572
rect 4740 516 4744 572
rect 4680 512 4744 516
rect 10360 572 10424 576
rect 10360 516 10364 572
rect 10364 516 10420 572
rect 10420 516 10424 572
rect 10360 512 10424 516
rect 10440 572 10504 576
rect 10440 516 10444 572
rect 10444 516 10500 572
rect 10500 516 10504 572
rect 10440 512 10504 516
rect 10520 572 10584 576
rect 10520 516 10524 572
rect 10524 516 10580 572
rect 10580 516 10584 572
rect 10520 512 10584 516
rect 10600 572 10664 576
rect 10600 516 10604 572
rect 10604 516 10660 572
rect 10660 516 10664 572
rect 10600 512 10664 516
rect 10680 572 10744 576
rect 10680 516 10684 572
rect 10684 516 10740 572
rect 10740 516 10744 572
rect 10680 512 10744 516
rect 16360 572 16424 576
rect 16360 516 16364 572
rect 16364 516 16420 572
rect 16420 516 16424 572
rect 16360 512 16424 516
rect 16440 572 16504 576
rect 16440 516 16444 572
rect 16444 516 16500 572
rect 16500 516 16504 572
rect 16440 512 16504 516
rect 16520 572 16584 576
rect 16520 516 16524 572
rect 16524 516 16580 572
rect 16580 516 16584 572
rect 16520 512 16584 516
rect 16600 572 16664 576
rect 16600 516 16604 572
rect 16604 516 16660 572
rect 16660 516 16664 572
rect 16600 512 16664 516
rect 16680 572 16744 576
rect 16680 516 16684 572
rect 16684 516 16740 572
rect 16740 516 16744 572
rect 16680 512 16744 516
<< metal4 >>
rect 1352 17440 1752 17456
rect 1352 17376 1360 17440
rect 1424 17376 1440 17440
rect 1504 17376 1520 17440
rect 1584 17376 1600 17440
rect 1664 17376 1680 17440
rect 1744 17376 1752 17440
rect 1352 16352 1752 17376
rect 1352 16288 1360 16352
rect 1424 16288 1440 16352
rect 1504 16288 1520 16352
rect 1584 16288 1600 16352
rect 1664 16288 1680 16352
rect 1744 16288 1752 16352
rect 1352 15264 1752 16288
rect 1352 15200 1360 15264
rect 1424 15200 1440 15264
rect 1504 15200 1520 15264
rect 1584 15200 1600 15264
rect 1664 15200 1680 15264
rect 1744 15200 1752 15264
rect 1352 14176 1752 15200
rect 1352 14112 1360 14176
rect 1424 14112 1440 14176
rect 1504 14112 1520 14176
rect 1584 14112 1600 14176
rect 1664 14112 1680 14176
rect 1744 14112 1752 14176
rect 1352 13088 1752 14112
rect 1352 13024 1360 13088
rect 1424 13024 1440 13088
rect 1504 13024 1520 13088
rect 1584 13024 1600 13088
rect 1664 13024 1680 13088
rect 1744 13024 1752 13088
rect 1352 12000 1752 13024
rect 1352 11936 1360 12000
rect 1424 11936 1440 12000
rect 1504 11936 1520 12000
rect 1584 11936 1600 12000
rect 1664 11936 1680 12000
rect 1744 11936 1752 12000
rect 1352 10912 1752 11936
rect 1352 10848 1360 10912
rect 1424 10848 1440 10912
rect 1504 10848 1520 10912
rect 1584 10848 1600 10912
rect 1664 10848 1680 10912
rect 1744 10848 1752 10912
rect 1352 9824 1752 10848
rect 1352 9760 1360 9824
rect 1424 9760 1440 9824
rect 1504 9760 1520 9824
rect 1584 9760 1600 9824
rect 1664 9760 1680 9824
rect 1744 9760 1752 9824
rect 1352 8736 1752 9760
rect 1352 8672 1360 8736
rect 1424 8672 1440 8736
rect 1504 8672 1520 8736
rect 1584 8672 1600 8736
rect 1664 8672 1680 8736
rect 1744 8672 1752 8736
rect 1352 7648 1752 8672
rect 1352 7584 1360 7648
rect 1424 7584 1440 7648
rect 1504 7584 1520 7648
rect 1584 7584 1600 7648
rect 1664 7584 1680 7648
rect 1744 7584 1752 7648
rect 1352 6560 1752 7584
rect 1352 6496 1360 6560
rect 1424 6496 1440 6560
rect 1504 6496 1520 6560
rect 1584 6496 1600 6560
rect 1664 6496 1680 6560
rect 1744 6496 1752 6560
rect 1352 5472 1752 6496
rect 1352 5408 1360 5472
rect 1424 5408 1440 5472
rect 1504 5408 1520 5472
rect 1584 5408 1600 5472
rect 1664 5408 1680 5472
rect 1744 5408 1752 5472
rect 1352 4384 1752 5408
rect 1352 4320 1360 4384
rect 1424 4320 1440 4384
rect 1504 4320 1520 4384
rect 1584 4320 1600 4384
rect 1664 4320 1680 4384
rect 1744 4320 1752 4384
rect 1352 3296 1752 4320
rect 1352 3232 1360 3296
rect 1424 3232 1440 3296
rect 1504 3232 1520 3296
rect 1584 3232 1600 3296
rect 1664 3232 1680 3296
rect 1744 3232 1752 3296
rect 1352 2208 1752 3232
rect 1352 2144 1360 2208
rect 1424 2144 1440 2208
rect 1504 2144 1520 2208
rect 1584 2144 1600 2208
rect 1664 2144 1680 2208
rect 1744 2144 1752 2208
rect 1352 1120 1752 2144
rect 1352 1056 1360 1120
rect 1424 1056 1440 1120
rect 1504 1056 1520 1120
rect 1584 1056 1600 1120
rect 1664 1056 1680 1120
rect 1744 1056 1752 1120
rect 1352 496 1752 1056
rect 4352 16896 4752 17456
rect 4352 16832 4360 16896
rect 4424 16832 4440 16896
rect 4504 16832 4520 16896
rect 4584 16832 4600 16896
rect 4664 16832 4680 16896
rect 4744 16832 4752 16896
rect 4352 15808 4752 16832
rect 7352 17440 7752 17456
rect 7352 17376 7360 17440
rect 7424 17376 7440 17440
rect 7504 17376 7520 17440
rect 7584 17376 7600 17440
rect 7664 17376 7680 17440
rect 7744 17376 7752 17440
rect 6499 16692 6565 16693
rect 6499 16628 6500 16692
rect 6564 16628 6565 16692
rect 6499 16627 6565 16628
rect 4352 15744 4360 15808
rect 4424 15744 4440 15808
rect 4504 15744 4520 15808
rect 4584 15744 4600 15808
rect 4664 15744 4680 15808
rect 4744 15744 4752 15808
rect 4352 14720 4752 15744
rect 6131 15332 6197 15333
rect 6131 15268 6132 15332
rect 6196 15268 6197 15332
rect 6131 15267 6197 15268
rect 4352 14656 4360 14720
rect 4424 14656 4440 14720
rect 4504 14656 4520 14720
rect 4584 14656 4600 14720
rect 4664 14656 4680 14720
rect 4744 14656 4752 14720
rect 4352 13632 4752 14656
rect 4352 13568 4360 13632
rect 4424 13568 4440 13632
rect 4504 13568 4520 13632
rect 4584 13568 4600 13632
rect 4664 13568 4680 13632
rect 4744 13568 4752 13632
rect 4352 12544 4752 13568
rect 4352 12480 4360 12544
rect 4424 12480 4440 12544
rect 4504 12480 4520 12544
rect 4584 12480 4600 12544
rect 4664 12480 4680 12544
rect 4744 12480 4752 12544
rect 4352 11456 4752 12480
rect 4352 11392 4360 11456
rect 4424 11392 4440 11456
rect 4504 11392 4520 11456
rect 4584 11392 4600 11456
rect 4664 11392 4680 11456
rect 4744 11392 4752 11456
rect 4352 10368 4752 11392
rect 4352 10304 4360 10368
rect 4424 10304 4440 10368
rect 4504 10304 4520 10368
rect 4584 10304 4600 10368
rect 4664 10304 4680 10368
rect 4744 10304 4752 10368
rect 4352 9280 4752 10304
rect 4352 9216 4360 9280
rect 4424 9216 4440 9280
rect 4504 9216 4520 9280
rect 4584 9216 4600 9280
rect 4664 9216 4680 9280
rect 4744 9216 4752 9280
rect 4352 8192 4752 9216
rect 4352 8128 4360 8192
rect 4424 8128 4440 8192
rect 4504 8128 4520 8192
rect 4584 8128 4600 8192
rect 4664 8128 4680 8192
rect 4744 8128 4752 8192
rect 4352 7104 4752 8128
rect 5947 7444 6013 7445
rect 5947 7380 5948 7444
rect 6012 7380 6013 7444
rect 5947 7379 6013 7380
rect 4352 7040 4360 7104
rect 4424 7040 4440 7104
rect 4504 7040 4520 7104
rect 4584 7040 4600 7104
rect 4664 7040 4680 7104
rect 4744 7040 4752 7104
rect 4352 6016 4752 7040
rect 4352 5952 4360 6016
rect 4424 5952 4440 6016
rect 4504 5952 4520 6016
rect 4584 5952 4600 6016
rect 4664 5952 4680 6016
rect 4744 5952 4752 6016
rect 4352 4928 4752 5952
rect 4352 4864 4360 4928
rect 4424 4864 4440 4928
rect 4504 4864 4520 4928
rect 4584 4864 4600 4928
rect 4664 4864 4680 4928
rect 4744 4864 4752 4928
rect 4352 3840 4752 4864
rect 4352 3776 4360 3840
rect 4424 3776 4440 3840
rect 4504 3776 4520 3840
rect 4584 3776 4600 3840
rect 4664 3776 4680 3840
rect 4744 3776 4752 3840
rect 4352 2752 4752 3776
rect 5950 3365 6010 7379
rect 5947 3364 6013 3365
rect 5947 3300 5948 3364
rect 6012 3300 6013 3364
rect 5947 3299 6013 3300
rect 4352 2688 4360 2752
rect 4424 2688 4440 2752
rect 4504 2688 4520 2752
rect 4584 2688 4600 2752
rect 4664 2688 4680 2752
rect 4744 2688 4752 2752
rect 4352 1664 4752 2688
rect 6134 2413 6194 15267
rect 6502 2685 6562 16627
rect 7352 16352 7752 17376
rect 10352 16896 10752 17456
rect 10352 16832 10360 16896
rect 10424 16832 10440 16896
rect 10504 16832 10520 16896
rect 10584 16832 10600 16896
rect 10664 16832 10680 16896
rect 10744 16832 10752 16896
rect 8707 16692 8773 16693
rect 8707 16628 8708 16692
rect 8772 16628 8773 16692
rect 8707 16627 8773 16628
rect 7352 16288 7360 16352
rect 7424 16288 7440 16352
rect 7504 16288 7520 16352
rect 7584 16288 7600 16352
rect 7664 16288 7680 16352
rect 7744 16288 7752 16352
rect 7352 15264 7752 16288
rect 7352 15200 7360 15264
rect 7424 15200 7440 15264
rect 7504 15200 7520 15264
rect 7584 15200 7600 15264
rect 7664 15200 7680 15264
rect 7744 15200 7752 15264
rect 7352 14176 7752 15200
rect 7352 14112 7360 14176
rect 7424 14112 7440 14176
rect 7504 14112 7520 14176
rect 7584 14112 7600 14176
rect 7664 14112 7680 14176
rect 7744 14112 7752 14176
rect 7352 13088 7752 14112
rect 7352 13024 7360 13088
rect 7424 13024 7440 13088
rect 7504 13024 7520 13088
rect 7584 13024 7600 13088
rect 7664 13024 7680 13088
rect 7744 13024 7752 13088
rect 7352 12000 7752 13024
rect 7352 11936 7360 12000
rect 7424 11936 7440 12000
rect 7504 11936 7520 12000
rect 7584 11936 7600 12000
rect 7664 11936 7680 12000
rect 7744 11936 7752 12000
rect 7352 10912 7752 11936
rect 7352 10848 7360 10912
rect 7424 10848 7440 10912
rect 7504 10848 7520 10912
rect 7584 10848 7600 10912
rect 7664 10848 7680 10912
rect 7744 10848 7752 10912
rect 7352 9824 7752 10848
rect 7352 9760 7360 9824
rect 7424 9760 7440 9824
rect 7504 9760 7520 9824
rect 7584 9760 7600 9824
rect 7664 9760 7680 9824
rect 7744 9760 7752 9824
rect 7352 8736 7752 9760
rect 7352 8672 7360 8736
rect 7424 8672 7440 8736
rect 7504 8672 7520 8736
rect 7584 8672 7600 8736
rect 7664 8672 7680 8736
rect 7744 8672 7752 8736
rect 7352 7648 7752 8672
rect 7352 7584 7360 7648
rect 7424 7584 7440 7648
rect 7504 7584 7520 7648
rect 7584 7584 7600 7648
rect 7664 7584 7680 7648
rect 7744 7584 7752 7648
rect 7352 6560 7752 7584
rect 7352 6496 7360 6560
rect 7424 6496 7440 6560
rect 7504 6496 7520 6560
rect 7584 6496 7600 6560
rect 7664 6496 7680 6560
rect 7744 6496 7752 6560
rect 7352 5472 7752 6496
rect 7352 5408 7360 5472
rect 7424 5408 7440 5472
rect 7504 5408 7520 5472
rect 7584 5408 7600 5472
rect 7664 5408 7680 5472
rect 7744 5408 7752 5472
rect 7352 4384 7752 5408
rect 7971 4996 8037 4997
rect 7971 4932 7972 4996
rect 8036 4932 8037 4996
rect 7971 4931 8037 4932
rect 7352 4320 7360 4384
rect 7424 4320 7440 4384
rect 7504 4320 7520 4384
rect 7584 4320 7600 4384
rect 7664 4320 7680 4384
rect 7744 4320 7752 4384
rect 7352 3296 7752 4320
rect 7352 3232 7360 3296
rect 7424 3232 7440 3296
rect 7504 3232 7520 3296
rect 7584 3232 7600 3296
rect 7664 3232 7680 3296
rect 7744 3232 7752 3296
rect 6499 2684 6565 2685
rect 6499 2620 6500 2684
rect 6564 2620 6565 2684
rect 6499 2619 6565 2620
rect 6131 2412 6197 2413
rect 6131 2348 6132 2412
rect 6196 2348 6197 2412
rect 6131 2347 6197 2348
rect 4352 1600 4360 1664
rect 4424 1600 4440 1664
rect 4504 1600 4520 1664
rect 4584 1600 4600 1664
rect 4664 1600 4680 1664
rect 4744 1600 4752 1664
rect 4352 576 4752 1600
rect 4352 512 4360 576
rect 4424 512 4440 576
rect 4504 512 4520 576
rect 4584 512 4600 576
rect 4664 512 4680 576
rect 4744 512 4752 576
rect 4352 496 4752 512
rect 7352 2208 7752 3232
rect 7974 2957 8034 4931
rect 7971 2956 8037 2957
rect 7971 2892 7972 2956
rect 8036 2892 8037 2956
rect 7971 2891 8037 2892
rect 7352 2144 7360 2208
rect 7424 2144 7440 2208
rect 7504 2144 7520 2208
rect 7584 2144 7600 2208
rect 7664 2144 7680 2208
rect 7744 2144 7752 2208
rect 7352 1120 7752 2144
rect 8710 1869 8770 16627
rect 10352 15808 10752 16832
rect 10352 15744 10360 15808
rect 10424 15744 10440 15808
rect 10504 15744 10520 15808
rect 10584 15744 10600 15808
rect 10664 15744 10680 15808
rect 10744 15744 10752 15808
rect 9259 15468 9325 15469
rect 9259 15404 9260 15468
rect 9324 15404 9325 15468
rect 9259 15403 9325 15404
rect 8891 12612 8957 12613
rect 8891 12548 8892 12612
rect 8956 12548 8957 12612
rect 8891 12547 8957 12548
rect 8894 10981 8954 12547
rect 8891 10980 8957 10981
rect 8891 10916 8892 10980
rect 8956 10916 8957 10980
rect 8891 10915 8957 10916
rect 9262 2413 9322 15403
rect 10352 14720 10752 15744
rect 13352 17440 13752 17456
rect 13352 17376 13360 17440
rect 13424 17376 13440 17440
rect 13504 17376 13520 17440
rect 13584 17376 13600 17440
rect 13664 17376 13680 17440
rect 13744 17376 13752 17440
rect 13352 16352 13752 17376
rect 13352 16288 13360 16352
rect 13424 16288 13440 16352
rect 13504 16288 13520 16352
rect 13584 16288 13600 16352
rect 13664 16288 13680 16352
rect 13744 16288 13752 16352
rect 11283 15332 11349 15333
rect 11283 15268 11284 15332
rect 11348 15268 11349 15332
rect 11283 15267 11349 15268
rect 13123 15332 13189 15333
rect 13123 15268 13124 15332
rect 13188 15268 13189 15332
rect 13123 15267 13189 15268
rect 10352 14656 10360 14720
rect 10424 14656 10440 14720
rect 10504 14656 10520 14720
rect 10584 14656 10600 14720
rect 10664 14656 10680 14720
rect 10744 14656 10752 14720
rect 10352 13632 10752 14656
rect 10352 13568 10360 13632
rect 10424 13568 10440 13632
rect 10504 13568 10520 13632
rect 10584 13568 10600 13632
rect 10664 13568 10680 13632
rect 10744 13568 10752 13632
rect 10352 12544 10752 13568
rect 10352 12480 10360 12544
rect 10424 12480 10440 12544
rect 10504 12480 10520 12544
rect 10584 12480 10600 12544
rect 10664 12480 10680 12544
rect 10744 12480 10752 12544
rect 10352 11456 10752 12480
rect 10352 11392 10360 11456
rect 10424 11392 10440 11456
rect 10504 11392 10520 11456
rect 10584 11392 10600 11456
rect 10664 11392 10680 11456
rect 10744 11392 10752 11456
rect 10352 10368 10752 11392
rect 10352 10304 10360 10368
rect 10424 10304 10440 10368
rect 10504 10304 10520 10368
rect 10584 10304 10600 10368
rect 10664 10304 10680 10368
rect 10744 10304 10752 10368
rect 10352 9280 10752 10304
rect 10352 9216 10360 9280
rect 10424 9216 10440 9280
rect 10504 9216 10520 9280
rect 10584 9216 10600 9280
rect 10664 9216 10680 9280
rect 10744 9216 10752 9280
rect 10352 8192 10752 9216
rect 10352 8128 10360 8192
rect 10424 8128 10440 8192
rect 10504 8128 10520 8192
rect 10584 8128 10600 8192
rect 10664 8128 10680 8192
rect 10744 8128 10752 8192
rect 10352 7104 10752 8128
rect 10352 7040 10360 7104
rect 10424 7040 10440 7104
rect 10504 7040 10520 7104
rect 10584 7040 10600 7104
rect 10664 7040 10680 7104
rect 10744 7040 10752 7104
rect 9811 6628 9877 6629
rect 9811 6564 9812 6628
rect 9876 6564 9877 6628
rect 9811 6563 9877 6564
rect 9814 3365 9874 6563
rect 10352 6016 10752 7040
rect 10352 5952 10360 6016
rect 10424 5952 10440 6016
rect 10504 5952 10520 6016
rect 10584 5952 10600 6016
rect 10664 5952 10680 6016
rect 10744 5952 10752 6016
rect 9995 5268 10061 5269
rect 9995 5204 9996 5268
rect 10060 5204 10061 5268
rect 9995 5203 10061 5204
rect 9811 3364 9877 3365
rect 9811 3300 9812 3364
rect 9876 3300 9877 3364
rect 9811 3299 9877 3300
rect 9259 2412 9325 2413
rect 9259 2348 9260 2412
rect 9324 2348 9325 2412
rect 9259 2347 9325 2348
rect 8707 1868 8773 1869
rect 8707 1804 8708 1868
rect 8772 1804 8773 1868
rect 8707 1803 8773 1804
rect 9998 1733 10058 5203
rect 10352 4928 10752 5952
rect 10352 4864 10360 4928
rect 10424 4864 10440 4928
rect 10504 4864 10520 4928
rect 10584 4864 10600 4928
rect 10664 4864 10680 4928
rect 10744 4864 10752 4928
rect 10352 3840 10752 4864
rect 10352 3776 10360 3840
rect 10424 3776 10440 3840
rect 10504 3776 10520 3840
rect 10584 3776 10600 3840
rect 10664 3776 10680 3840
rect 10744 3776 10752 3840
rect 10352 2752 10752 3776
rect 10352 2688 10360 2752
rect 10424 2688 10440 2752
rect 10504 2688 10520 2752
rect 10584 2688 10600 2752
rect 10664 2688 10680 2752
rect 10744 2688 10752 2752
rect 9995 1732 10061 1733
rect 9995 1668 9996 1732
rect 10060 1668 10061 1732
rect 9995 1667 10061 1668
rect 9811 1596 9877 1597
rect 9811 1532 9812 1596
rect 9876 1532 9877 1596
rect 9811 1531 9877 1532
rect 9814 1189 9874 1531
rect 9998 1325 10058 1667
rect 10352 1664 10752 2688
rect 10352 1600 10360 1664
rect 10424 1600 10440 1664
rect 10504 1600 10520 1664
rect 10584 1600 10600 1664
rect 10664 1600 10680 1664
rect 10744 1600 10752 1664
rect 9995 1324 10061 1325
rect 9995 1260 9996 1324
rect 10060 1260 10061 1324
rect 9995 1259 10061 1260
rect 9811 1188 9877 1189
rect 9811 1124 9812 1188
rect 9876 1124 9877 1188
rect 9811 1123 9877 1124
rect 7352 1056 7360 1120
rect 7424 1056 7440 1120
rect 7504 1056 7520 1120
rect 7584 1056 7600 1120
rect 7664 1056 7680 1120
rect 7744 1056 7752 1120
rect 7352 496 7752 1056
rect 10352 576 10752 1600
rect 11286 1325 11346 15267
rect 12755 11796 12821 11797
rect 12755 11732 12756 11796
rect 12820 11732 12821 11796
rect 12755 11731 12821 11732
rect 12203 11116 12269 11117
rect 12203 11052 12204 11116
rect 12268 11052 12269 11116
rect 12203 11051 12269 11052
rect 12206 3909 12266 11051
rect 12758 5949 12818 11731
rect 12755 5948 12821 5949
rect 12755 5884 12756 5948
rect 12820 5884 12821 5948
rect 12755 5883 12821 5884
rect 12203 3908 12269 3909
rect 12203 3844 12204 3908
rect 12268 3844 12269 3908
rect 12203 3843 12269 3844
rect 13126 2005 13186 15267
rect 13352 15264 13752 16288
rect 13352 15200 13360 15264
rect 13424 15200 13440 15264
rect 13504 15200 13520 15264
rect 13584 15200 13600 15264
rect 13664 15200 13680 15264
rect 13744 15200 13752 15264
rect 13352 14176 13752 15200
rect 13352 14112 13360 14176
rect 13424 14112 13440 14176
rect 13504 14112 13520 14176
rect 13584 14112 13600 14176
rect 13664 14112 13680 14176
rect 13744 14112 13752 14176
rect 13352 13088 13752 14112
rect 13352 13024 13360 13088
rect 13424 13024 13440 13088
rect 13504 13024 13520 13088
rect 13584 13024 13600 13088
rect 13664 13024 13680 13088
rect 13744 13024 13752 13088
rect 13352 12000 13752 13024
rect 16352 16896 16752 17456
rect 16352 16832 16360 16896
rect 16424 16832 16440 16896
rect 16504 16832 16520 16896
rect 16584 16832 16600 16896
rect 16664 16832 16680 16896
rect 16744 16832 16752 16896
rect 16352 15808 16752 16832
rect 16352 15744 16360 15808
rect 16424 15744 16440 15808
rect 16504 15744 16520 15808
rect 16584 15744 16600 15808
rect 16664 15744 16680 15808
rect 16744 15744 16752 15808
rect 16352 14720 16752 15744
rect 16352 14656 16360 14720
rect 16424 14656 16440 14720
rect 16504 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16752 14720
rect 16352 13632 16752 14656
rect 16352 13568 16360 13632
rect 16424 13568 16440 13632
rect 16504 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16752 13632
rect 14043 12748 14109 12749
rect 14043 12684 14044 12748
rect 14108 12684 14109 12748
rect 14043 12683 14109 12684
rect 13352 11936 13360 12000
rect 13424 11936 13440 12000
rect 13504 11936 13520 12000
rect 13584 11936 13600 12000
rect 13664 11936 13680 12000
rect 13744 11936 13752 12000
rect 13352 10912 13752 11936
rect 13352 10848 13360 10912
rect 13424 10848 13440 10912
rect 13504 10848 13520 10912
rect 13584 10848 13600 10912
rect 13664 10848 13680 10912
rect 13744 10848 13752 10912
rect 13352 9824 13752 10848
rect 13352 9760 13360 9824
rect 13424 9760 13440 9824
rect 13504 9760 13520 9824
rect 13584 9760 13600 9824
rect 13664 9760 13680 9824
rect 13744 9760 13752 9824
rect 13352 8736 13752 9760
rect 13352 8672 13360 8736
rect 13424 8672 13440 8736
rect 13504 8672 13520 8736
rect 13584 8672 13600 8736
rect 13664 8672 13680 8736
rect 13744 8672 13752 8736
rect 13352 7648 13752 8672
rect 13352 7584 13360 7648
rect 13424 7584 13440 7648
rect 13504 7584 13520 7648
rect 13584 7584 13600 7648
rect 13664 7584 13680 7648
rect 13744 7584 13752 7648
rect 13352 6560 13752 7584
rect 14046 7445 14106 12683
rect 16352 12544 16752 13568
rect 16352 12480 16360 12544
rect 16424 12480 16440 12544
rect 16504 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16752 12544
rect 16352 11456 16752 12480
rect 16352 11392 16360 11456
rect 16424 11392 16440 11456
rect 16504 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16752 11456
rect 16352 10368 16752 11392
rect 16352 10304 16360 10368
rect 16424 10304 16440 10368
rect 16504 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16752 10368
rect 16352 9280 16752 10304
rect 16352 9216 16360 9280
rect 16424 9216 16440 9280
rect 16504 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16752 9280
rect 16352 8192 16752 9216
rect 16352 8128 16360 8192
rect 16424 8128 16440 8192
rect 16504 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16752 8192
rect 14043 7444 14109 7445
rect 14043 7380 14044 7444
rect 14108 7380 14109 7444
rect 14043 7379 14109 7380
rect 13859 7172 13925 7173
rect 13859 7108 13860 7172
rect 13924 7108 13925 7172
rect 13859 7107 13925 7108
rect 13352 6496 13360 6560
rect 13424 6496 13440 6560
rect 13504 6496 13520 6560
rect 13584 6496 13600 6560
rect 13664 6496 13680 6560
rect 13744 6496 13752 6560
rect 13352 5472 13752 6496
rect 13862 6221 13922 7107
rect 16352 7104 16752 8128
rect 16352 7040 16360 7104
rect 16424 7040 16440 7104
rect 16504 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16752 7104
rect 14779 7036 14845 7037
rect 14779 6972 14780 7036
rect 14844 6972 14845 7036
rect 14779 6971 14845 6972
rect 13859 6220 13925 6221
rect 13859 6156 13860 6220
rect 13924 6156 13925 6220
rect 13859 6155 13925 6156
rect 13352 5408 13360 5472
rect 13424 5408 13440 5472
rect 13504 5408 13520 5472
rect 13584 5408 13600 5472
rect 13664 5408 13680 5472
rect 13744 5408 13752 5472
rect 13352 4384 13752 5408
rect 13352 4320 13360 4384
rect 13424 4320 13440 4384
rect 13504 4320 13520 4384
rect 13584 4320 13600 4384
rect 13664 4320 13680 4384
rect 13744 4320 13752 4384
rect 13352 3296 13752 4320
rect 13352 3232 13360 3296
rect 13424 3232 13440 3296
rect 13504 3232 13520 3296
rect 13584 3232 13600 3296
rect 13664 3232 13680 3296
rect 13744 3232 13752 3296
rect 13352 2208 13752 3232
rect 14782 2685 14842 6971
rect 16352 6016 16752 7040
rect 16352 5952 16360 6016
rect 16424 5952 16440 6016
rect 16504 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16752 6016
rect 16352 4928 16752 5952
rect 16352 4864 16360 4928
rect 16424 4864 16440 4928
rect 16504 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16752 4928
rect 15147 4044 15213 4045
rect 15147 3980 15148 4044
rect 15212 3980 15213 4044
rect 15147 3979 15213 3980
rect 14779 2684 14845 2685
rect 14779 2620 14780 2684
rect 14844 2620 14845 2684
rect 14779 2619 14845 2620
rect 13352 2144 13360 2208
rect 13424 2144 13440 2208
rect 13504 2144 13520 2208
rect 13584 2144 13600 2208
rect 13664 2144 13680 2208
rect 13744 2144 13752 2208
rect 13123 2004 13189 2005
rect 13123 1940 13124 2004
rect 13188 1940 13189 2004
rect 13123 1939 13189 1940
rect 11283 1324 11349 1325
rect 11283 1260 11284 1324
rect 11348 1260 11349 1324
rect 11283 1259 11349 1260
rect 10352 512 10360 576
rect 10424 512 10440 576
rect 10504 512 10520 576
rect 10584 512 10600 576
rect 10664 512 10680 576
rect 10744 512 10752 576
rect 10352 496 10752 512
rect 13352 1120 13752 2144
rect 15150 1597 15210 3979
rect 16352 3840 16752 4864
rect 16352 3776 16360 3840
rect 16424 3776 16440 3840
rect 16504 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16752 3840
rect 16352 2752 16752 3776
rect 16352 2688 16360 2752
rect 16424 2688 16440 2752
rect 16504 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16752 2752
rect 16352 1664 16752 2688
rect 16352 1600 16360 1664
rect 16424 1600 16440 1664
rect 16504 1600 16520 1664
rect 16584 1600 16600 1664
rect 16664 1600 16680 1664
rect 16744 1600 16752 1664
rect 15147 1596 15213 1597
rect 15147 1532 15148 1596
rect 15212 1532 15213 1596
rect 15147 1531 15213 1532
rect 15150 1325 15210 1531
rect 15147 1324 15213 1325
rect 15147 1260 15148 1324
rect 15212 1260 15213 1324
rect 15147 1259 15213 1260
rect 13352 1056 13360 1120
rect 13424 1056 13440 1120
rect 13504 1056 13520 1120
rect 13584 1056 13600 1120
rect 13664 1056 13680 1120
rect 13744 1056 13752 1120
rect 13352 496 13752 1056
rect 16352 576 16752 1600
rect 16352 512 16360 576
rect 16424 512 16440 576
rect 16504 512 16520 576
rect 16584 512 16600 576
rect 16664 512 16680 576
rect 16744 512 16752 576
rect 16352 496 16752 512
use sky130_fd_sc_hd__buf_1  _0512_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3956 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3588 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4416 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0515_
timestamp 1704896540
transform 1 0 3772 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0516_
timestamp 1704896540
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0517_
timestamp 1704896540
transform 1 0 2300 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0518_
timestamp 1704896540
transform 1 0 5244 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0519_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0520_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4324 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0521_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5244 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0522_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4048 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0523_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4600 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0524_
timestamp 1704896540
transform 1 0 4508 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0525_
timestamp 1704896540
transform -1 0 4416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0526_
timestamp 1704896540
transform -1 0 4140 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0527_
timestamp 1704896540
transform 1 0 3128 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0528_
timestamp 1704896540
transform 1 0 3404 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0529_
timestamp 1704896540
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0530_
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4324 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0532_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4784 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0533_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0534_
timestamp 1704896540
transform 1 0 3128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0535_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3864 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0536_
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0537_
timestamp 1704896540
transform 1 0 5152 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _0538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0539_
timestamp 1704896540
transform -1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0540_
timestamp 1704896540
transform -1 0 11960 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0541_
timestamp 1704896540
transform 1 0 12236 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0542_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12144 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0543_
timestamp 1704896540
transform -1 0 11408 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0544_
timestamp 1704896540
transform 1 0 12788 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0545_
timestamp 1704896540
transform -1 0 11684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0546_
timestamp 1704896540
transform -1 0 11408 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0547_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12696 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1704896540
transform -1 0 16376 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0549_
timestamp 1704896540
transform -1 0 17296 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0550_
timestamp 1704896540
transform -1 0 16652 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0551_
timestamp 1704896540
transform 1 0 15088 0 1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1704896540
transform -1 0 17020 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0553_
timestamp 1704896540
transform 1 0 16652 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0554_
timestamp 1704896540
transform -1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0555_
timestamp 1704896540
transform -1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0556_
timestamp 1704896540
transform 1 0 6072 0 1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1704896540
transform 1 0 17020 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0558_
timestamp 1704896540
transform -1 0 17020 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0559_
timestamp 1704896540
transform -1 0 16928 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0560_
timestamp 1704896540
transform -1 0 17112 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0561_
timestamp 1704896540
transform -1 0 17204 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0562_
timestamp 1704896540
transform -1 0 13248 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0563_
timestamp 1704896540
transform -1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0564_
timestamp 1704896540
transform -1 0 12236 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0565_
timestamp 1704896540
transform 1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0566_
timestamp 1704896540
transform -1 0 9936 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0567_
timestamp 1704896540
transform -1 0 11960 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0568_
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0569_
timestamp 1704896540
transform -1 0 11500 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0570_
timestamp 1704896540
transform 1 0 9384 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0571_
timestamp 1704896540
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13156 0 -1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__nand2_1  _0573_
timestamp 1704896540
transform 1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16008 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0575_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16468 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0576_
timestamp 1704896540
transform 1 0 17020 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0577_
timestamp 1704896540
transform 1 0 16928 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0578_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16744 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12144 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0580_
timestamp 1704896540
transform 1 0 15272 0 1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _0581_
timestamp 1704896540
transform 1 0 15824 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0582_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15088 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0583_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12880 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0584_
timestamp 1704896540
transform -1 0 13340 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0585_
timestamp 1704896540
transform -1 0 3128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0586_
timestamp 1704896540
transform 1 0 9384 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14260 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0588_
timestamp 1704896540
transform 1 0 12696 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0589_
timestamp 1704896540
transform 1 0 13524 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0590_
timestamp 1704896540
transform -1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0591_
timestamp 1704896540
transform 1 0 13708 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0592_
timestamp 1704896540
transform -1 0 12512 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0593_
timestamp 1704896540
transform 1 0 16468 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16928 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0595_
timestamp 1704896540
transform 1 0 16284 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0596_
timestamp 1704896540
transform -1 0 16836 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0597_
timestamp 1704896540
transform -1 0 16744 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0598_
timestamp 1704896540
transform -1 0 15640 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0599_
timestamp 1704896540
transform -1 0 12880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0600_
timestamp 1704896540
transform -1 0 13432 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0601_
timestamp 1704896540
transform 1 0 8832 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0602_
timestamp 1704896540
transform 1 0 4416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0603_
timestamp 1704896540
transform 1 0 9200 0 1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_1  _0604_
timestamp 1704896540
transform -1 0 17112 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12696 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0606_
timestamp 1704896540
transform -1 0 11592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12696 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11776 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12052 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0611_
timestamp 1704896540
transform -1 0 16836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0612_
timestamp 1704896540
transform -1 0 12788 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0613_
timestamp 1704896540
transform 1 0 12052 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0614_
timestamp 1704896540
transform -1 0 12972 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0615_
timestamp 1704896540
transform -1 0 12972 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0616_
timestamp 1704896540
transform 1 0 12604 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0617_
timestamp 1704896540
transform 1 0 12880 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0618_
timestamp 1704896540
transform -1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0619_
timestamp 1704896540
transform -1 0 9752 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0620_
timestamp 1704896540
transform -1 0 14720 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _0621_
timestamp 1704896540
transform 1 0 9752 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _0622_
timestamp 1704896540
transform 1 0 11592 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0623_
timestamp 1704896540
transform 1 0 11868 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0624_
timestamp 1704896540
transform 1 0 12880 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0625_
timestamp 1704896540
transform 1 0 13156 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16744 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0627_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0628_
timestamp 1704896540
transform 1 0 15824 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0629_
timestamp 1704896540
transform 1 0 16100 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1704896540
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0631_
timestamp 1704896540
transform -1 0 17388 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0632_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17020 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0633_
timestamp 1704896540
transform -1 0 17388 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0634_
timestamp 1704896540
transform -1 0 17112 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0635_
timestamp 1704896540
transform 1 0 16652 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0636_
timestamp 1704896540
transform -1 0 17112 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0637_
timestamp 1704896540
transform 1 0 17112 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0638_
timestamp 1704896540
transform -1 0 14168 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0639_
timestamp 1704896540
transform 1 0 12604 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0640_
timestamp 1704896540
transform -1 0 10488 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0641_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11408 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11224 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1704896540
transform -1 0 15456 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0644_
timestamp 1704896540
transform -1 0 16560 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0645_
timestamp 1704896540
transform 1 0 15456 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0646_
timestamp 1704896540
transform 1 0 15180 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16100 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0648_
timestamp 1704896540
transform 1 0 17112 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1704896540
transform -1 0 14720 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0650_
timestamp 1704896540
transform -1 0 17112 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1704896540
transform -1 0 14444 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0652_
timestamp 1704896540
transform -1 0 12696 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0653_
timestamp 1704896540
transform -1 0 11776 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0654_
timestamp 1704896540
transform -1 0 10856 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0655_
timestamp 1704896540
transform -1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0656_
timestamp 1704896540
transform -1 0 8740 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0657_
timestamp 1704896540
transform -1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0658_
timestamp 1704896540
transform 1 0 6348 0 -1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_1  _0659_
timestamp 1704896540
transform -1 0 10396 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0660_
timestamp 1704896540
transform -1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0661_
timestamp 1704896540
transform 1 0 10948 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0662_
timestamp 1704896540
transform -1 0 10948 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0663_
timestamp 1704896540
transform 1 0 12236 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0664_
timestamp 1704896540
transform 1 0 10120 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0665_
timestamp 1704896540
transform 1 0 2668 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0666_
timestamp 1704896540
transform 1 0 4048 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0667_
timestamp 1704896540
transform 1 0 4324 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0668_
timestamp 1704896540
transform 1 0 5612 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0669_
timestamp 1704896540
transform 1 0 9016 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0670_
timestamp 1704896540
transform 1 0 5428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0671_
timestamp 1704896540
transform 1 0 6900 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0672_
timestamp 1704896540
transform 1 0 8004 0 -1 13600
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _0673_
timestamp 1704896540
transform -1 0 10120 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0674_
timestamp 1704896540
transform -1 0 10212 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0675_
timestamp 1704896540
transform 1 0 10948 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0676_
timestamp 1704896540
transform 1 0 11316 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0677_
timestamp 1704896540
transform 1 0 15088 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0678_
timestamp 1704896540
transform 1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0679_
timestamp 1704896540
transform -1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_2  _0680_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15548 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0681_
timestamp 1704896540
transform 1 0 4600 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0682_
timestamp 1704896540
transform 1 0 2484 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0683_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4600 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0684_
timestamp 1704896540
transform -1 0 4232 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1704896540
transform 1 0 4692 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1704896540
transform -1 0 9844 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0687_
timestamp 1704896540
transform -1 0 9568 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0688_
timestamp 1704896540
transform -1 0 10856 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0689_
timestamp 1704896540
transform 1 0 9660 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1704896540
transform 1 0 3956 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1704896540
transform -1 0 3956 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0692_
timestamp 1704896540
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0693_
timestamp 1704896540
transform 1 0 4600 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0694_
timestamp 1704896540
transform -1 0 10212 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0695_
timestamp 1704896540
transform 1 0 9384 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0696_
timestamp 1704896540
transform -1 0 6624 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1704896540
transform 1 0 2576 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0698_
timestamp 1704896540
transform -1 0 2484 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0699_
timestamp 1704896540
transform -1 0 3036 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0700_
timestamp 1704896540
transform -1 0 2208 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0701_
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _0702_
timestamp 1704896540
transform -1 0 4232 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0703_
timestamp 1704896540
transform 1 0 4232 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0704_
timestamp 1704896540
transform -1 0 4876 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0705_
timestamp 1704896540
transform -1 0 4324 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0707_
timestamp 1704896540
transform -1 0 4416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0708_
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0709_
timestamp 1704896540
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0710_
timestamp 1704896540
transform 1 0 6348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0711_
timestamp 1704896540
transform 1 0 6992 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0712_
timestamp 1704896540
transform 1 0 7636 0 -1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_1  _0713_
timestamp 1704896540
transform -1 0 2852 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0714_
timestamp 1704896540
transform 1 0 4048 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0715_
timestamp 1704896540
transform -1 0 12696 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _0716_
timestamp 1704896540
transform -1 0 7452 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0717_
timestamp 1704896540
transform -1 0 8280 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0718_
timestamp 1704896540
transform 1 0 10764 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0719_
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0720_
timestamp 1704896540
transform 1 0 2392 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0721_
timestamp 1704896540
transform -1 0 2760 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1704896540
transform 1 0 2116 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0723_
timestamp 1704896540
transform 1 0 1472 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0724_
timestamp 1704896540
transform 1 0 1564 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0725_
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0726_
timestamp 1704896540
transform 1 0 2024 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0727_
timestamp 1704896540
transform 1 0 2760 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0728_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0729_
timestamp 1704896540
transform -1 0 3772 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0730_
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0731_
timestamp 1704896540
transform -1 0 3864 0 -1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0732_
timestamp 1704896540
transform 1 0 4968 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0733_
timestamp 1704896540
transform -1 0 3864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0734_
timestamp 1704896540
transform 1 0 4048 0 -1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__o22a_1  _0735_
timestamp 1704896540
transform 1 0 7084 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0736_
timestamp 1704896540
transform 1 0 5336 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0737_
timestamp 1704896540
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0738_
timestamp 1704896540
transform 1 0 4968 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1704896540
transform -1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0740_
timestamp 1704896540
transform 1 0 1840 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0741_
timestamp 1704896540
transform 1 0 4692 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_2  _0742_
timestamp 1704896540
transform -1 0 4968 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0743_
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0744_
timestamp 1704896540
transform 1 0 1196 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0745_
timestamp 1704896540
transform -1 0 2760 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0746_
timestamp 1704896540
transform 1 0 2208 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0747_
timestamp 1704896540
transform 1 0 2576 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1704896540
transform -1 0 8648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0749_
timestamp 1704896540
transform 1 0 5060 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0750_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7084 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0751_
timestamp 1704896540
transform 1 0 5796 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0752_
timestamp 1704896540
transform -1 0 7176 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1704896540
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0755_
timestamp 1704896540
transform -1 0 1932 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0756_
timestamp 1704896540
transform 1 0 5888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0757_
timestamp 1704896540
transform 1 0 6348 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0758_
timestamp 1704896540
transform -1 0 7820 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0759_
timestamp 1704896540
transform 1 0 6900 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0760_
timestamp 1704896540
transform 1 0 8556 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0761_
timestamp 1704896540
transform 1 0 6072 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0762_
timestamp 1704896540
transform 1 0 13432 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0763_
timestamp 1704896540
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0764_
timestamp 1704896540
transform -1 0 13800 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1704896540
transform 1 0 16560 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0766_
timestamp 1704896540
transform -1 0 15180 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0767_
timestamp 1704896540
transform -1 0 16560 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0768_
timestamp 1704896540
transform 1 0 8924 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0769_
timestamp 1704896540
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0770_
timestamp 1704896540
transform -1 0 15732 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0771_
timestamp 1704896540
transform -1 0 12144 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0772_
timestamp 1704896540
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0773_
timestamp 1704896540
transform 1 0 13524 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0774_
timestamp 1704896540
transform -1 0 14904 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0775_
timestamp 1704896540
transform 1 0 14260 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0776_
timestamp 1704896540
transform 1 0 13708 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0777_
timestamp 1704896540
transform 1 0 13800 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0778_
timestamp 1704896540
transform 1 0 14720 0 -1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0779_
timestamp 1704896540
transform 1 0 14812 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0780_
timestamp 1704896540
transform -1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0781_
timestamp 1704896540
transform -1 0 8096 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0782_
timestamp 1704896540
transform 1 0 6164 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0783_
timestamp 1704896540
transform 1 0 13340 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0784_
timestamp 1704896540
transform 1 0 12144 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0785_
timestamp 1704896540
transform -1 0 13800 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0786_
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0787_
timestamp 1704896540
transform 1 0 12604 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0788_
timestamp 1704896540
transform 1 0 14812 0 -1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0789_
timestamp 1704896540
transform 1 0 13800 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0790_
timestamp 1704896540
transform -1 0 14168 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0791_
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0792_
timestamp 1704896540
transform -1 0 13432 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0793_
timestamp 1704896540
transform 1 0 13156 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0794_
timestamp 1704896540
transform -1 0 10764 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0795_
timestamp 1704896540
transform -1 0 12236 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0796_
timestamp 1704896540
transform 1 0 7268 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0797_
timestamp 1704896540
transform -1 0 11776 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0798_
timestamp 1704896540
transform 1 0 11040 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0799_
timestamp 1704896540
transform 1 0 10212 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0800_
timestamp 1704896540
transform -1 0 10304 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0801_
timestamp 1704896540
transform -1 0 8464 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0802_
timestamp 1704896540
transform 1 0 2760 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0803_
timestamp 1704896540
transform -1 0 9936 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0804_
timestamp 1704896540
transform 1 0 9476 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0805_
timestamp 1704896540
transform 1 0 9384 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0806_
timestamp 1704896540
transform 1 0 8832 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0807_
timestamp 1704896540
transform 1 0 7360 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0808_
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0809_
timestamp 1704896540
transform 1 0 7544 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0810_
timestamp 1704896540
transform -1 0 8188 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0811_
timestamp 1704896540
transform -1 0 8372 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0812_
timestamp 1704896540
transform 1 0 5336 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0813_
timestamp 1704896540
transform -1 0 5704 0 -1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0814_
timestamp 1704896540
transform -1 0 6348 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0815_
timestamp 1704896540
transform -1 0 6624 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0816_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5520 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0817_
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0818_
timestamp 1704896540
transform -1 0 12328 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0819_
timestamp 1704896540
transform -1 0 3956 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _0820_
timestamp 1704896540
transform 1 0 7820 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0821_
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0822_
timestamp 1704896540
transform -1 0 7544 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0823_
timestamp 1704896540
transform 1 0 7268 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0824_
timestamp 1704896540
transform -1 0 15180 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0825_
timestamp 1704896540
transform -1 0 14904 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1704896540
transform 1 0 10212 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0827_
timestamp 1704896540
transform -1 0 9752 0 -1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0828_
timestamp 1704896540
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0829_
timestamp 1704896540
transform -1 0 12604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0830_
timestamp 1704896540
transform 1 0 9936 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0831_
timestamp 1704896540
transform 1 0 12512 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0832_
timestamp 1704896540
transform 1 0 14260 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0833_
timestamp 1704896540
transform 1 0 14996 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0834_
timestamp 1704896540
transform -1 0 14720 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0835_
timestamp 1704896540
transform -1 0 15364 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0836_
timestamp 1704896540
transform -1 0 14996 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1704896540
transform -1 0 14628 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0838_
timestamp 1704896540
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0839_
timestamp 1704896540
transform -1 0 14996 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0840_
timestamp 1704896540
transform 1 0 14076 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0841_
timestamp 1704896540
transform -1 0 14812 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 1704896540
transform -1 0 14076 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0844_
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0845_
timestamp 1704896540
transform -1 0 14444 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0846_
timestamp 1704896540
transform -1 0 14260 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0847_
timestamp 1704896540
transform -1 0 14812 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0848_
timestamp 1704896540
transform -1 0 11040 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0849_
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1704896540
transform 1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0851_
timestamp 1704896540
transform -1 0 11500 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0852_
timestamp 1704896540
transform -1 0 12512 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0853_
timestamp 1704896540
transform -1 0 11684 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0854_
timestamp 1704896540
transform 1 0 11040 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0855_
timestamp 1704896540
transform -1 0 11500 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0856_
timestamp 1704896540
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0857_
timestamp 1704896540
transform 1 0 8924 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0858_
timestamp 1704896540
transform 1 0 4876 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0859_
timestamp 1704896540
transform -1 0 9660 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0860_
timestamp 1704896540
transform -1 0 10856 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0861_
timestamp 1704896540
transform -1 0 12604 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0862_
timestamp 1704896540
transform -1 0 7268 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0863_
timestamp 1704896540
transform -1 0 7728 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0864_
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0865_
timestamp 1704896540
transform 1 0 7176 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0866_
timestamp 1704896540
transform -1 0 7360 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0867_
timestamp 1704896540
transform -1 0 11500 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0868_
timestamp 1704896540
transform 1 0 5244 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0870_
timestamp 1704896540
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1704896540
transform -1 0 6624 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0872_
timestamp 1704896540
transform -1 0 6900 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0873_
timestamp 1704896540
transform 1 0 9108 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0874_
timestamp 1704896540
transform -1 0 9200 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0875_
timestamp 1704896540
transform -1 0 9752 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0876_
timestamp 1704896540
transform 1 0 8832 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1704896540
transform -1 0 9108 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0878_
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0880_
timestamp 1704896540
transform 1 0 6072 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0881_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10672 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1704896540
transform -1 0 14352 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0883_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0884_
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0885_
timestamp 1704896540
transform -1 0 3128 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0886_
timestamp 1704896540
transform 1 0 6072 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0887_
timestamp 1704896540
transform -1 0 7360 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1704896540
transform -1 0 7728 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0889_
timestamp 1704896540
transform -1 0 8648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0890_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0891_
timestamp 1704896540
transform 1 0 6808 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0892_
timestamp 1704896540
transform 1 0 6992 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _0893_
timestamp 1704896540
transform -1 0 8004 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _0894_
timestamp 1704896540
transform -1 0 8096 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0895_
timestamp 1704896540
transform -1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 1704896540
transform 1 0 2300 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 1704896540
transform 1 0 1656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0898_
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0900_
timestamp 1704896540
transform -1 0 17020 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0901_
timestamp 1704896540
transform 1 0 7912 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0902_
timestamp 1704896540
transform -1 0 9292 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0903_
timestamp 1704896540
transform 1 0 4508 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0904_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0905_
timestamp 1704896540
transform 1 0 5428 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0906_
timestamp 1704896540
transform 1 0 13984 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1704896540
transform 1 0 6900 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0908_
timestamp 1704896540
transform 1 0 8004 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1704896540
transform 1 0 14996 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0910_
timestamp 1704896540
transform 1 0 14352 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1704896540
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0912_
timestamp 1704896540
transform 1 0 5060 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0913_
timestamp 1704896540
transform -1 0 14628 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0914_
timestamp 1704896540
transform 1 0 8464 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0915_
timestamp 1704896540
transform -1 0 16008 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 1704896540
transform -1 0 13984 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1704896540
transform -1 0 13984 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0918_
timestamp 1704896540
transform 1 0 14628 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0919_
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0920_
timestamp 1704896540
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0921_
timestamp 1704896540
transform -1 0 13248 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0922_
timestamp 1704896540
transform -1 0 12328 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0923_
timestamp 1704896540
transform -1 0 11960 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0924_
timestamp 1704896540
transform -1 0 3680 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1704896540
transform 1 0 13800 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0926_
timestamp 1704896540
transform 1 0 13800 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0927_
timestamp 1704896540
transform -1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0928_
timestamp 1704896540
transform -1 0 2760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0929_
timestamp 1704896540
transform -1 0 3404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0930_
timestamp 1704896540
transform -1 0 3128 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0931_
timestamp 1704896540
transform 1 0 3404 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0932_
timestamp 1704896540
transform 1 0 2300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0933_
timestamp 1704896540
transform -1 0 3128 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0934_
timestamp 1704896540
transform -1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1704896540
transform -1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0936_
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1704896540
transform 1 0 1380 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0938_
timestamp 1704896540
transform -1 0 2300 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1704896540
transform 1 0 1196 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0940_
timestamp 1704896540
transform 1 0 13984 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1704896540
transform 1 0 17112 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0942_
timestamp 1704896540
transform -1 0 12972 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0943_
timestamp 1704896540
transform 1 0 12788 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1704896540
transform 1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0945_
timestamp 1704896540
transform 1 0 14260 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0946_
timestamp 1704896540
transform -1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6716 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0948_
timestamp 1704896540
transform -1 0 6072 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1704896540
transform -1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0950_
timestamp 1704896540
transform 1 0 4784 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_2  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0952_
timestamp 1704896540
transform -1 0 6256 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0953_
timestamp 1704896540
transform -1 0 4784 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0954_
timestamp 1704896540
transform -1 0 13892 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0955_
timestamp 1704896540
transform 1 0 13708 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0956_
timestamp 1704896540
transform -1 0 11316 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1704896540
transform -1 0 2668 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0958_
timestamp 1704896540
transform 1 0 12420 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0959_
timestamp 1704896540
transform -1 0 3864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0960_
timestamp 1704896540
transform 1 0 2484 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 1704896540
transform -1 0 3220 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1704896540
transform -1 0 2116 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0963_
timestamp 1704896540
transform -1 0 5152 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0964_
timestamp 1704896540
transform 1 0 2116 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0965_
timestamp 1704896540
transform 1 0 1472 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1704896540
transform -1 0 2208 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0967_
timestamp 1704896540
transform -1 0 2576 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0968_
timestamp 1704896540
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0969_
timestamp 1704896540
transform -1 0 3036 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0970_
timestamp 1704896540
transform -1 0 1932 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0971_
timestamp 1704896540
transform 1 0 1288 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0972_
timestamp 1704896540
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0973_
timestamp 1704896540
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0974_
timestamp 1704896540
transform -1 0 3128 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0975_
timestamp 1704896540
transform 1 0 2392 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0976_
timestamp 1704896540
transform 1 0 2484 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1704896540
transform -1 0 3128 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0978_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2484 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0979_
timestamp 1704896540
transform 1 0 1380 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0980_
timestamp 1704896540
transform 1 0 16100 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1704896540
transform 1 0 15732 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp 1704896540
transform -1 0 15640 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1704896540
transform -1 0 15732 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp 1704896540
transform 1 0 13524 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1704896540
transform -1 0 13800 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0986_
timestamp 1704896540
transform -1 0 12880 0 -1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0987_
timestamp 1704896540
transform 1 0 11868 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1704896540
transform -1 0 9384 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0989_
timestamp 1704896540
transform -1 0 12236 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1704896540
transform 1 0 13340 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0991_
timestamp 1704896540
transform 1 0 11040 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1704896540
transform -1 0 11500 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1704896540
transform 1 0 9936 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1704896540
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 1704896540
transform 1 0 7360 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1704896540
transform 1 0 4600 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0997_
timestamp 1704896540
transform 1 0 6256 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0998_
timestamp 1704896540
transform 1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0999_
timestamp 1704896540
transform -1 0 12604 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1704896540
transform -1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1001_
timestamp 1704896540
transform -1 0 14812 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1002_
timestamp 1704896540
transform 1 0 15456 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1003_
timestamp 1704896540
transform -1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1004_
timestamp 1704896540
transform 1 0 16100 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1704896540
transform 1 0 16560 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1006_
timestamp 1704896540
transform -1 0 13064 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1007_
timestamp 1704896540
transform 1 0 9108 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1704896540
transform -1 0 11408 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1009_
timestamp 1704896540
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1010_
timestamp 1704896540
transform 1 0 4784 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _1011_
timestamp 1704896540
transform -1 0 10488 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1012_
timestamp 1704896540
transform -1 0 11868 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1013_
timestamp 1704896540
transform 1 0 10028 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1014_
timestamp 1704896540
transform 1 0 10120 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1015_
timestamp 1704896540
transform -1 0 9660 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1016_
timestamp 1704896540
transform 1 0 9752 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1704896540
transform 1 0 8924 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1018_
timestamp 1704896540
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1019_
timestamp 1704896540
transform 1 0 6348 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1704896540
transform 1 0 6992 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1021_
timestamp 1704896540
transform 1 0 6624 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1022_
timestamp 1704896540
transform -1 0 6164 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1023_
timestamp 1704896540
transform 1 0 7268 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1024_
timestamp 1704896540
transform -1 0 6992 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1025_
timestamp 1704896540
transform 1 0 5796 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1026_
timestamp 1704896540
transform -1 0 6624 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1027_
timestamp 1704896540
transform 1 0 5888 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1704896540
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1029_
timestamp 1704896540
transform 1 0 6256 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1030_
timestamp 1704896540
transform 1 0 7636 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1031_
timestamp 1704896540
transform -1 0 7360 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1032_
timestamp 1704896540
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1033_
timestamp 1704896540
transform 1 0 6072 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1034_
timestamp 1704896540
transform 1 0 6256 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1035_
timestamp 1704896540
transform -1 0 7636 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1036_
timestamp 1704896540
transform 1 0 4600 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1704896540
transform 1 0 7820 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1038_
timestamp 1704896540
transform -1 0 9660 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1039_
timestamp 1704896540
transform -1 0 9660 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1704896540
transform 1 0 6716 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1041_
timestamp 1704896540
transform 1 0 4968 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _1042_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7820 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1043_
timestamp 1704896540
transform -1 0 8372 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1044_
timestamp 1704896540
transform -1 0 9200 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1045_
timestamp 1704896540
transform -1 0 9108 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1046_
timestamp 1704896540
transform -1 0 12604 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1047_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8096 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1048_
timestamp 1704896540
transform 1 0 7176 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1049_
timestamp 1704896540
transform 1 0 6072 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1050_
timestamp 1704896540
transform 1 0 5336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1051_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1012 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1704896540
transform 1 0 15272 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1704896540
transform 1 0 14536 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1704896540
transform 1 0 14352 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1704896540
transform 1 0 11408 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1704896540
transform 1 0 15824 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1704896540
transform 1 0 15824 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1704896540
transform 1 0 14260 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1704896540
transform 1 0 920 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1704896540
transform 1 0 3128 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1704896540
transform 1 0 1196 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1704896540
transform 1 0 14536 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1704896540
transform 1 0 15640 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1704896540
transform 1 0 13800 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1704896540
transform -1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1704896540
transform -1 0 12972 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1704896540
transform 1 0 11500 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1704896540
transform 1 0 9292 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1704896540
transform -1 0 4692 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1704896540
transform 1 0 14812 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1704896540
transform 1 0 15916 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10488 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1704896540
transform 1 0 1748 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1704896540
transform -1 0 2300 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1704896540
transform -1 0 4692 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1704896540
transform 1 0 2300 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1704896540
transform 1 0 2576 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1704896540
transform 1 0 4784 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 1704896540
transform 1 0 1472 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1704896540
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1091_
timestamp 1704896540
transform -1 0 6716 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1704896540
transform 1 0 6716 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1093_
timestamp 1704896540
transform -1 0 12788 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1704896540
transform -1 0 12604 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10304 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1704896540
transform -1 0 6256 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1704896540
transform -1 0 6440 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1704896540
transform 1 0 12420 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1704896540
transform 1 0 11316 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1748 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2944 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_37
timestamp 1704896540
transform 1 0 3956 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_45
timestamp 1704896540
transform 1 0 4692 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_61
timestamp 1704896540
transform 1 0 6164 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77
timestamp 1704896540
transform 1 0 7636 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_91
timestamp 1704896540
transform 1 0 8924 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_119
timestamp 1704896540
transform 1 0 11500 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_131
timestamp 1704896540
transform 1 0 12604 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1704896540
transform 1 0 13248 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_147
timestamp 1704896540
transform 1 0 14076 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1704896540
transform 1 0 15916 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_180
timestamp 1704896540
transform 1 0 17112 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 1704896540
transform 1 0 1380 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_13
timestamp 1704896540
transform 1 0 1748 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_21
timestamp 1704896540
transform 1 0 2484 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_42
timestamp 1704896540
transform 1 0 4416 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_85
timestamp 1704896540
transform 1 0 8372 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_89
timestamp 1704896540
transform 1 0 8740 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1704896540
transform 1 0 15824 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_180
timestamp 1704896540
transform 1 0 17112 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_14
timestamp 1704896540
transform 1 0 1840 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_55
timestamp 1704896540
transform 1 0 5612 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_59
timestamp 1704896540
transform 1 0 5980 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_114
timestamp 1704896540
transform 1 0 11040 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1472 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_22
timestamp 1704896540
transform 1 0 2576 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_26
timestamp 1704896540
transform 1 0 2944 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_41
timestamp 1704896540
transform 1 0 4324 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1704896540
transform 1 0 5428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_66
timestamp 1704896540
transform 1 0 6624 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_72
timestamp 1704896540
transform 1 0 7176 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_78
timestamp 1704896540
transform 1 0 7728 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_97
timestamp 1704896540
transform 1 0 9476 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1704896540
transform 1 0 10580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_120
timestamp 1704896540
transform 1 0 11592 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_126
timestamp 1704896540
transform 1 0 12144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_136 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13064 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_144
timestamp 1704896540
transform 1 0 13800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_157
timestamp 1704896540
transform 1 0 14996 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_174
timestamp 1704896540
transform 1 0 16560 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_9
timestamp 1704896540
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_20
timestamp 1704896540
transform 1 0 2392 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_33
timestamp 1704896540
transform 1 0 3588 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_47
timestamp 1704896540
transform 1 0 4876 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_69
timestamp 1704896540
transform 1 0 6900 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_93
timestamp 1704896540
transform 1 0 9108 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_103
timestamp 1704896540
transform 1 0 10028 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_115
timestamp 1704896540
transform 1 0 11132 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_121
timestamp 1704896540
transform 1 0 11684 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_129
timestamp 1704896540
transform 1 0 12420 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_159
timestamp 1704896540
transform 1 0 15180 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_170
timestamp 1704896540
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_11
timestamp 1704896540
transform 1 0 1564 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_36
timestamp 1704896540
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_48
timestamp 1704896540
transform 1 0 4968 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_66
timestamp 1704896540
transform 1 0 6624 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_74
timestamp 1704896540
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_84
timestamp 1704896540
transform 1 0 8280 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_90
timestamp 1704896540
transform 1 0 8832 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_96
timestamp 1704896540
transform 1 0 9384 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_119
timestamp 1704896540
transform 1 0 11500 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_132
timestamp 1704896540
transform 1 0 12696 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_164
timestamp 1704896540
transform 1 0 15640 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_182
timestamp 1704896540
transform 1 0 17296 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_45
timestamp 1704896540
transform 1 0 4692 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_51
timestamp 1704896540
transform 1 0 5244 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_66
timestamp 1704896540
transform 1 0 6624 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_78
timestamp 1704896540
transform 1 0 7728 0 1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9476 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_101
timestamp 1704896540
transform 1 0 9844 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_107
timestamp 1704896540
transform 1 0 10396 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_121
timestamp 1704896540
transform 1 0 11684 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_132
timestamp 1704896540
transform 1 0 12696 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_156
timestamp 1704896540
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_173
timestamp 1704896540
transform 1 0 16468 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_10
timestamp 1704896540
transform 1 0 1472 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_34
timestamp 1704896540
transform 1 0 3680 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_46
timestamp 1704896540
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_66
timestamp 1704896540
transform 1 0 6624 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_84
timestamp 1704896540
transform 1 0 8280 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_135
timestamp 1704896540
transform 1 0 12972 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_141
timestamp 1704896540
transform 1 0 13524 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_159
timestamp 1704896540
transform 1 0 15180 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16100 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_177
timestamp 1704896540
transform 1 0 16836 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_56
timestamp 1704896540
transform 1 0 5704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_60
timestamp 1704896540
transform 1 0 6072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_78
timestamp 1704896540
transform 1 0 7728 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_102
timestamp 1704896540
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_119
timestamp 1704896540
transform 1 0 11500 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_135
timestamp 1704896540
transform 1 0 12972 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_148
timestamp 1704896540
transform 1 0 14168 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_160
timestamp 1704896540
transform 1 0 15272 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_172
timestamp 1704896540
transform 1 0 16376 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_180
timestamp 1704896540
transform 1 0 17112 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_19
timestamp 1704896540
transform 1 0 2300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_28
timestamp 1704896540
transform 1 0 3128 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_48
timestamp 1704896540
transform 1 0 4968 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_66
timestamp 1704896540
transform 1 0 6624 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_75
timestamp 1704896540
transform 1 0 7452 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_87
timestamp 1704896540
transform 1 0 8556 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_107
timestamp 1704896540
transform 1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_121
timestamp 1704896540
transform 1 0 11684 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_146
timestamp 1704896540
transform 1 0 13984 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_152
timestamp 1704896540
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_172
timestamp 1704896540
transform 1 0 16376 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_181
timestamp 1704896540
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_21
timestamp 1704896540
transform 1 0 2484 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1704896540
transform 1 0 2852 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1704896540
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_94
timestamp 1704896540
transform 1 0 9200 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_106
timestamp 1704896540
transform 1 0 10304 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_120
timestamp 1704896540
transform 1 0 11592 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_126
timestamp 1704896540
transform 1 0 12144 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_130
timestamp 1704896540
transform 1 0 12512 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 1704896540
transform 1 0 12880 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_156
timestamp 1704896540
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_180
timestamp 1704896540
transform 1 0 17112 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_19
timestamp 1704896540
transform 1 0 2300 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_26
timestamp 1704896540
transform 1 0 2944 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_32
timestamp 1704896540
transform 1 0 3496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_48
timestamp 1704896540
transform 1 0 4968 0 -1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_76
timestamp 1704896540
transform 1 0 7544 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_88
timestamp 1704896540
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_103
timestamp 1704896540
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_122
timestamp 1704896540
transform 1 0 11776 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_134
timestamp 1704896540
transform 1 0 12880 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_142
timestamp 1704896540
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_147
timestamp 1704896540
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_159
timestamp 1704896540
transform 1 0 15180 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1704896540
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16100 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_175
timestamp 1704896540
transform 1 0 16652 0 -1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1704896540
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1704896540
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_47
timestamp 1704896540
transform 1 0 4876 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_51
timestamp 1704896540
transform 1 0 5244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_61
timestamp 1704896540
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_66
timestamp 1704896540
transform 1 0 6624 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_78
timestamp 1704896540
transform 1 0 7728 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_100
timestamp 1704896540
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_111
timestamp 1704896540
transform 1 0 10764 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_121
timestamp 1704896540
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_131
timestamp 1704896540
transform 1 0 12604 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_163
timestamp 1704896540
transform 1 0 15548 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_178
timestamp 1704896540
transform 1 0 16928 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_182
timestamp 1704896540
transform 1 0 17296 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_30
timestamp 1704896540
transform 1 0 3312 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_68
timestamp 1704896540
transform 1 0 6808 0 -1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_86
timestamp 1704896540
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_98
timestamp 1704896540
transform 1 0 9568 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_133
timestamp 1704896540
transform 1 0 12788 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_139
timestamp 1704896540
transform 1 0 13340 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_158
timestamp 1704896540
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1704896540
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_177
timestamp 1704896540
transform 1 0 16836 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1704896540
transform 1 0 2300 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_76
timestamp 1704896540
transform 1 0 7544 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_99
timestamp 1704896540
transform 1 0 9660 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_108
timestamp 1704896540
transform 1 0 10488 0 1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_122
timestamp 1704896540
transform 1 0 11776 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_134
timestamp 1704896540
transform 1 0 12880 0 1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_150
timestamp 1704896540
transform 1 0 14352 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_162
timestamp 1704896540
transform 1 0 15456 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_166
timestamp 1704896540
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_11
timestamp 1704896540
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_77
timestamp 1704896540
transform 1 0 7636 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_99
timestamp 1704896540
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_103
timestamp 1704896540
transform 1 0 10028 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_123
timestamp 1704896540
transform 1 0 11868 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_127
timestamp 1704896540
transform 1 0 12236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_131
timestamp 1704896540
transform 1 0 12604 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_160
timestamp 1704896540
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_164
timestamp 1704896540
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_182
timestamp 1704896540
transform 1 0 17296 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_25
timestamp 1704896540
transform 1 0 2852 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4324 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_70
timestamp 1704896540
transform 1 0 6992 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1704896540
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_96
timestamp 1704896540
transform 1 0 9384 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_134
timestamp 1704896540
transform 1 0 12880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_146
timestamp 1704896540
transform 1 0 13984 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_171
timestamp 1704896540
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_48
timestamp 1704896540
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_77
timestamp 1704896540
transform 1 0 7636 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_88
timestamp 1704896540
transform 1 0 8648 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_101
timestamp 1704896540
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_107
timestamp 1704896540
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1704896540
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_135
timestamp 1704896540
transform 1 0 12972 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_139
timestamp 1704896540
transform 1 0 13340 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_143
timestamp 1704896540
transform 1 0 13708 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_151
timestamp 1704896540
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_182
timestamp 1704896540
transform 1 0 17296 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_9
timestamp 1704896540
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_13
timestamp 1704896540
transform 1 0 1748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_25
timestamp 1704896540
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_42
timestamp 1704896540
transform 1 0 4416 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_51
timestamp 1704896540
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_68
timestamp 1704896540
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_80
timestamp 1704896540
transform 1 0 7912 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_106
timestamp 1704896540
transform 1 0 10304 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_118
timestamp 1704896540
transform 1 0 11408 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_130
timestamp 1704896540
transform 1 0 12512 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_146
timestamp 1704896540
transform 1 0 13984 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_165
timestamp 1704896540
transform 1 0 15732 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_178
timestamp 1704896540
transform 1 0 16928 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_182
timestamp 1704896540
transform 1 0 17296 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_11
timestamp 1704896540
transform 1 0 1564 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_21
timestamp 1704896540
transform 1 0 2484 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1704896540
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_60
timestamp 1704896540
transform 1 0 6072 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_66
timestamp 1704896540
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_82
timestamp 1704896540
transform 1 0 8096 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_99
timestamp 1704896540
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1704896540
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_149
timestamp 1704896540
transform 1 0 14260 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_153
timestamp 1704896540
transform 1 0 14628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_172
timestamp 1704896540
transform 1 0 16376 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_179
timestamp 1704896540
transform 1 0 17020 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_12
timestamp 1704896540
transform 1 0 1656 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_22
timestamp 1704896540
transform 1 0 2576 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_33
timestamp 1704896540
transform 1 0 3588 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_64
timestamp 1704896540
transform 1 0 6440 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_72
timestamp 1704896540
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1704896540
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_128
timestamp 1704896540
transform 1 0 12328 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1704896540
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_158
timestamp 1704896540
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_176
timestamp 1704896540
transform 1 0 16744 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_182
timestamp 1704896540
transform 1 0 17296 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_19
timestamp 1704896540
transform 1 0 2300 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_25
timestamp 1704896540
transform 1 0 2852 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_29
timestamp 1704896540
transform 1 0 3220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_88
timestamp 1704896540
transform 1 0 8648 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_100
timestamp 1704896540
transform 1 0 9752 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_117
timestamp 1704896540
transform 1 0 11316 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_134
timestamp 1704896540
transform 1 0 12880 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_142
timestamp 1704896540
transform 1 0 13616 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_7
timestamp 1704896540
transform 1 0 1196 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_15
timestamp 1704896540
transform 1 0 1932 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_45
timestamp 1704896540
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_72
timestamp 1704896540
transform 1 0 7176 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_89
timestamp 1704896540
transform 1 0 8740 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_118
timestamp 1704896540
transform 1 0 11408 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_127
timestamp 1704896540
transform 1 0 12236 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1704896540
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_154
timestamp 1704896540
transform 1 0 14720 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_165
timestamp 1704896540
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_182
timestamp 1704896540
transform 1 0 17296 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_34
timestamp 1704896540
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_41
timestamp 1704896540
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_60
timestamp 1704896540
transform 1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1704896540
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_116
timestamp 1704896540
transform 1 0 11224 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_15
timestamp 1704896540
transform 1 0 1932 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_21
timestamp 1704896540
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_57
timestamp 1704896540
transform 1 0 5796 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1704896540
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_88
timestamp 1704896540
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_93
timestamp 1704896540
transform 1 0 9108 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1704896540
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_173
timestamp 1704896540
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_181
timestamp 1704896540
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_17
timestamp 1704896540
transform 1 0 2116 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_37
timestamp 1704896540
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_67
timestamp 1704896540
transform 1 0 6716 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_95
timestamp 1704896540
transform 1 0 9292 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_100
timestamp 1704896540
transform 1 0 9752 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1704896540
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_116
timestamp 1704896540
transform 1 0 11224 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_120
timestamp 1704896540
transform 1 0 11592 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_136
timestamp 1704896540
transform 1 0 13064 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_142
timestamp 1704896540
transform 1 0 13616 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_147
timestamp 1704896540
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_181
timestamp 1704896540
transform 1 0 17204 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_19
timestamp 1704896540
transform 1 0 2300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_43
timestamp 1704896540
transform 1 0 4508 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_60
timestamp 1704896540
transform 1 0 6072 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_69
timestamp 1704896540
transform 1 0 6900 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_90
timestamp 1704896540
transform 1 0 8832 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_102
timestamp 1704896540
transform 1 0 9936 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_114
timestamp 1704896540
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1704896540
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_147
timestamp 1704896540
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_156
timestamp 1704896540
transform 1 0 14904 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_165
timestamp 1704896540
transform 1 0 15732 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_182
timestamp 1704896540
transform 1 0 17296 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_3
timestamp 1704896540
transform 1 0 828 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_31
timestamp 1704896540
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_63
timestamp 1704896540
transform 1 0 6348 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_67
timestamp 1704896540
transform 1 0 6716 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_82
timestamp 1704896540
transform 1 0 8096 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_90
timestamp 1704896540
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_95
timestamp 1704896540
transform 1 0 9292 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1704896540
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1704896540
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_119
timestamp 1704896540
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_142
timestamp 1704896540
transform 1 0 13616 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_158
timestamp 1704896540
transform 1 0 15088 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_175
timestamp 1704896540
transform 1 0 16652 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_182
timestamp 1704896540
transform 1 0 17296 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_3
timestamp 1704896540
transform 1 0 828 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_23
timestamp 1704896540
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_45
timestamp 1704896540
transform 1 0 4692 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_71
timestamp 1704896540
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_93
timestamp 1704896540
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_117
timestamp 1704896540
transform 1 0 11316 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_133
timestamp 1704896540
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_154
timestamp 1704896540
transform 1 0 14720 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_180
timestamp 1704896540
transform 1 0 17112 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_3
timestamp 1704896540
transform 1 0 828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_21
timestamp 1704896540
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_47
timestamp 1704896540
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1704896540
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_64
timestamp 1704896540
transform 1 0 6440 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_72
timestamp 1704896540
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1704896540
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_113
timestamp 1704896540
transform 1 0 10948 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_135
timestamp 1704896540
transform 1 0 12972 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_139
timestamp 1704896540
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1704896540
transform 1 0 15824 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_181
timestamp 1704896540
transform 1 0 17204 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_3
timestamp 1704896540
transform 1 0 828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_41
timestamp 1704896540
transform 1 0 4324 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_54
timestamp 1704896540
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_63
timestamp 1704896540
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_69
timestamp 1704896540
transform 1 0 6900 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_79
timestamp 1704896540
transform 1 0 7820 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_88
timestamp 1704896540
transform 1 0 8648 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_96
timestamp 1704896540
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_113
timestamp 1704896540
transform 1 0 10948 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_150
timestamp 1704896540
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_169
timestamp 1704896540
transform 1 0 16100 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_180
timestamp 1704896540
transform 1 0 17112 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3956 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 6164 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 13432 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1704896540
transform 1 0 16192 0 1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform -1 0 17204 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform 1 0 15548 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1704896540
transform 1 0 14076 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1704896540
transform 1 0 13800 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1704896540
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1704896540
transform -1 0 10120 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1704896540
transform 1 0 9568 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4324 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1704896540
transform 1 0 7084 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1704896540
transform -1 0 6164 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1704896540
transform -1 0 5428 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1704896540
transform -1 0 4692 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1704896540
transform -1 0 3956 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1704896540
transform -1 0 3588 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1704896540
transform -1 0 2944 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1748 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1704896540
transform -1 0 1196 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1704896540
transform -1 0 4968 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1704896540
transform 1 0 7912 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1704896540
transform -1 0 12052 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1704896540
transform -1 0 12604 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1704896540
transform -1 0 9752 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1704896540
transform 1 0 10304 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1704896540
transform -1 0 8280 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1704896540
transform 1 0 7268 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1704896540
transform -1 0 6900 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1704896540
transform -1 0 1656 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1704896540
transform 1 0 4968 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1704896540
transform -1 0 6348 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1704896540
transform -1 0 9108 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1704896540
transform -1 0 15088 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1704896540
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1704896540
transform 1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1704896540
transform 1 0 14812 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1704896540
transform 1 0 16100 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1704896540
transform 1 0 16100 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1704896540
transform 1 0 15364 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1704896540
transform -1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1704896540
transform 1 0 7452 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 17664 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 17664 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 17664 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 17664 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 17664 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 17664 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 17664 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 17664 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 17664 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 17664 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 17664 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 17664 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 17664 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 17664 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 17664 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp 1704896540
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 17664 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp 1704896540
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp 1704896540
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 17664 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp 1704896540
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 1704896540
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_68
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_69
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_70
timestamp 1704896540
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_71
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_72
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_73
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_74
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_75
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp 1704896540
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_78
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_79
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp 1704896540
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_87
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp 1704896540
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_92
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_93
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp 1704896540
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_96
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_97
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp 1704896540
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_102
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_103
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_105
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_106
timestamp 1704896540
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_108
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_109
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_111
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_112
timestamp 1704896540
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_113
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_114
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_115
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_116
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_117
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_118
timestamp 1704896540
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_119
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_120
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_121
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_122
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_123
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_124
timestamp 1704896540
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_125
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_126
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_127
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_128
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_129
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_130
timestamp 1704896540
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_131
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_132
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_133
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_134
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_135
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_136
timestamp 1704896540
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_137
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_138
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_139
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_140
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_141
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_142
timestamp 1704896540
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_143
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_144
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_145
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_146
timestamp 1704896540
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_147
timestamp 1704896540
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_148
timestamp 1704896540
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 1704896540
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 1704896540
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_151
timestamp 1704896540
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_152
timestamp 1704896540
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_153
timestamp 1704896540
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp 1704896540
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_155
timestamp 1704896540
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_156
timestamp 1704896540
transform 1 0 5704 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_157
timestamp 1704896540
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_158
timestamp 1704896540
transform 1 0 10856 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_159
timestamp 1704896540
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_160
timestamp 1704896540
transform 1 0 16008 0 1 16864
box -38 -48 130 592
<< labels >>
flabel metal4 s 4352 496 4752 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10352 496 10752 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16352 496 16752 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1352 496 1752 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7352 496 7752 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13352 496 13752 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 3698 17845 3754 18245 0 FreeSans 224 90 0 0 b6
port 2 nsew signal tristate
flabel metal2 s 7010 17845 7066 18245 0 FreeSans 224 90 0 0 b7
port 3 nsew signal tristate
flabel metal2 s 5722 0 5778 400 0 FreeSans 224 90 0 0 b[0]
port 4 nsew signal tristate
flabel metal2 s 4986 0 5042 400 0 FreeSans 224 90 0 0 b[1]
port 5 nsew signal tristate
flabel metal2 s 4250 0 4306 400 0 FreeSans 224 90 0 0 b[2]
port 6 nsew signal tristate
flabel metal2 s 3514 0 3570 400 0 FreeSans 224 90 0 0 b[3]
port 7 nsew signal tristate
flabel metal2 s 2778 0 2834 400 0 FreeSans 224 90 0 0 b[4]
port 8 nsew signal tristate
flabel metal2 s 2042 0 2098 400 0 FreeSans 224 90 0 0 b[5]
port 9 nsew signal tristate
flabel metal2 s 1306 0 1362 400 0 FreeSans 224 90 0 0 b[6]
port 10 nsew signal tristate
flabel metal2 s 570 0 626 400 0 FreeSans 224 90 0 0 b[7]
port 11 nsew signal tristate
flabel metal2 s 16946 17845 17002 18245 0 FreeSans 224 90 0 0 clk
port 12 nsew signal input
flabel metal2 s 4526 17845 4582 18245 0 FreeSans 224 90 0 0 g6
port 13 nsew signal tristate
flabel metal2 s 7838 17845 7894 18245 0 FreeSans 224 90 0 0 g7
port 14 nsew signal tristate
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 g[0]
port 15 nsew signal tristate
flabel metal2 s 10874 0 10930 400 0 FreeSans 224 90 0 0 g[1]
port 16 nsew signal tristate
flabel metal2 s 10138 0 10194 400 0 FreeSans 224 90 0 0 g[2]
port 17 nsew signal tristate
flabel metal2 s 9402 0 9458 400 0 FreeSans 224 90 0 0 g[3]
port 18 nsew signal tristate
flabel metal2 s 8666 0 8722 400 0 FreeSans 224 90 0 0 g[4]
port 19 nsew signal tristate
flabel metal2 s 7930 0 7986 400 0 FreeSans 224 90 0 0 g[5]
port 20 nsew signal tristate
flabel metal2 s 7194 0 7250 400 0 FreeSans 224 90 0 0 g[6]
port 21 nsew signal tristate
flabel metal2 s 6458 0 6514 400 0 FreeSans 224 90 0 0 g[7]
port 22 nsew signal tristate
flabel metal2 s 1214 17845 1270 18245 0 FreeSans 224 90 0 0 hblank
port 23 nsew signal tristate
flabel metal2 s 2870 17845 2926 18245 0 FreeSans 224 90 0 0 hsync
port 24 nsew signal tristate
flabel metal2 s 5354 17845 5410 18245 0 FreeSans 224 90 0 0 r6
port 25 nsew signal tristate
flabel metal2 s 8666 17845 8722 18245 0 FreeSans 224 90 0 0 r7
port 26 nsew signal tristate
flabel metal2 s 17498 0 17554 400 0 FreeSans 224 90 0 0 r[0]
port 27 nsew signal tristate
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 r[1]
port 28 nsew signal tristate
flabel metal2 s 16026 0 16082 400 0 FreeSans 224 90 0 0 r[2]
port 29 nsew signal tristate
flabel metal2 s 15290 0 15346 400 0 FreeSans 224 90 0 0 r[3]
port 30 nsew signal tristate
flabel metal2 s 14554 0 14610 400 0 FreeSans 224 90 0 0 r[4]
port 31 nsew signal tristate
flabel metal2 s 13818 0 13874 400 0 FreeSans 224 90 0 0 r[5]
port 32 nsew signal tristate
flabel metal2 s 13082 0 13138 400 0 FreeSans 224 90 0 0 r[6]
port 33 nsew signal tristate
flabel metal2 s 12346 0 12402 400 0 FreeSans 224 90 0 0 r[7]
port 34 nsew signal tristate
flabel metal2 s 16118 17845 16174 18245 0 FreeSans 224 90 0 0 rst_n
port 35 nsew signal input
flabel metal2 s 15290 17845 15346 18245 0 FreeSans 224 90 0 0 ui_in[0]
port 36 nsew signal input
flabel metal2 s 14462 17845 14518 18245 0 FreeSans 224 90 0 0 ui_in[1]
port 37 nsew signal input
flabel metal2 s 13634 17845 13690 18245 0 FreeSans 224 90 0 0 ui_in[2]
port 38 nsew signal input
flabel metal2 s 12806 17845 12862 18245 0 FreeSans 224 90 0 0 ui_in[3]
port 39 nsew signal input
flabel metal2 s 11978 17845 12034 18245 0 FreeSans 224 90 0 0 ui_in[4]
port 40 nsew signal input
flabel metal2 s 11150 17845 11206 18245 0 FreeSans 224 90 0 0 ui_in[5]
port 41 nsew signal input
flabel metal2 s 10322 17845 10378 18245 0 FreeSans 224 90 0 0 ui_in[6]
port 42 nsew signal input
flabel metal2 s 9494 17845 9550 18245 0 FreeSans 224 90 0 0 ui_in[7]
port 43 nsew signal input
flabel metal2 s 2042 17845 2098 18245 0 FreeSans 224 90 0 0 vblank
port 44 nsew signal tristate
flabel metal2 s 6182 17845 6238 18245 0 FreeSans 224 90 0 0 vsync
port 45 nsew signal tristate
rlabel metal1 9108 16864 9108 16864 0 VGND
rlabel metal1 9108 17408 9108 17408 0 VPWR
rlabel metal1 1513 16694 1513 16694 0 _0000_
rlabel metal2 16146 11458 16146 11458 0 _0001_
rlabel metal1 14750 12342 14750 12342 0 _0002_
rlabel metal2 15778 13668 15778 13668 0 _0003_
rlabel metal1 11822 11866 11822 11866 0 _0004_
rlabel metal1 2254 5882 2254 5882 0 _0005_
rlabel metal1 2070 5678 2070 5678 0 _0006_
rlabel via1 3537 4046 3537 4046 0 _0007_
rlabel metal1 1191 3978 1191 3978 0 _0008_
rlabel metal1 16647 12750 16647 12750 0 _0009_
rlabel metal1 15900 14858 15900 14858 0 _0010_
rlabel metal1 13987 14586 13987 14586 0 _0011_
rlabel via1 3537 12682 3537 12682 0 _0012_
rlabel metal1 1375 10098 1375 10098 0 _0013_
rlabel metal1 1288 11866 1288 11866 0 _0014_
rlabel metal1 1288 12954 1288 12954 0 _0015_
rlabel metal1 1659 14586 1659 14586 0 _0016_
rlabel metal1 3174 16150 3174 16150 0 _0017_
rlabel metal1 1472 15674 1472 15674 0 _0018_
rlabel metal1 15456 15334 15456 15334 0 _0019_
rlabel metal1 15732 15674 15732 15674 0 _0020_
rlabel metal1 14020 16626 14020 16626 0 _0021_
rlabel viali 9342 16626 9342 16626 0 _0022_
rlabel via1 12654 14858 12654 14858 0 _0023_
rlabel metal1 11720 16626 11720 16626 0 _0024_
rlabel metal1 9655 15946 9655 15946 0 _0025_
rlabel metal1 4523 15946 4523 15946 0 _0026_
rlabel metal1 14934 9418 14934 9418 0 _0027_
rlabel metal1 16698 8058 16698 8058 0 _0028_
rlabel metal2 10442 9758 10442 9758 0 _0029_
rlabel metal1 10902 9146 10902 9146 0 _0030_
rlabel via2 2622 9027 2622 9027 0 _0031_
rlabel metal1 6578 8806 6578 8806 0 _0032_
rlabel metal1 2384 8330 2384 8330 0 _0033_
rlabel metal1 4472 9010 4472 9010 0 _0034_
rlabel metal1 3859 10166 3859 10166 0 _0035_
rlabel via2 7038 10795 7038 10795 0 _0036_
rlabel metal1 5239 16014 5239 16014 0 _0037_
rlabel metal2 4324 13396 4324 13396 0 _0038_
rlabel metal1 5704 13838 5704 13838 0 _0039_
rlabel metal2 6762 11135 6762 11135 0 _0040_
rlabel metal2 4186 10676 4186 10676 0 _0041_
rlabel metal1 4646 7718 4646 7718 0 _0042_
rlabel metal1 2254 9622 2254 9622 0 _0043_
rlabel metal1 5520 10982 5520 10982 0 _0044_
rlabel metal1 3910 10234 3910 10234 0 _0045_
rlabel metal2 5290 9894 5290 9894 0 _0046_
rlabel metal1 4416 10778 4416 10778 0 _0047_
rlabel metal1 4738 11322 4738 11322 0 _0048_
rlabel metal1 4968 13158 4968 13158 0 _0049_
rlabel metal2 8602 14756 8602 14756 0 _0050_
rlabel metal2 3542 15164 3542 15164 0 _0051_
rlabel metal1 10074 13362 10074 13362 0 _0052_
rlabel metal1 6670 13804 6670 13804 0 _0053_
rlabel metal1 8832 13362 8832 13362 0 _0054_
rlabel metal1 4646 7242 4646 7242 0 _0055_
rlabel metal1 3956 13498 3956 13498 0 _0056_
rlabel metal1 4278 9418 4278 9418 0 _0057_
rlabel metal1 3634 14042 3634 14042 0 _0058_
rlabel metal1 4370 14892 4370 14892 0 _0059_
rlabel metal1 3818 14926 3818 14926 0 _0060_
rlabel metal1 5474 12682 5474 12682 0 _0061_
rlabel viali 12462 3570 12462 3570 0 _0062_
rlabel metal1 11914 14479 11914 14479 0 _0063_
rlabel metal2 12558 9248 12558 9248 0 _0064_
rlabel metal1 9545 2482 9545 2482 0 _0065_
rlabel metal1 12374 1938 12374 1938 0 _0066_
rlabel metal1 12926 1326 12926 1326 0 _0067_
rlabel metal2 7222 5372 7222 5372 0 _0068_
rlabel metal2 13800 2380 13800 2380 0 _0069_
rlabel metal1 12696 1870 12696 1870 0 _0070_
rlabel metal1 15824 5610 15824 5610 0 _0071_
rlabel metal1 16514 15402 16514 15402 0 _0072_
rlabel metal1 8234 6732 8234 6732 0 _0073_
rlabel metal2 7406 6052 7406 6052 0 _0074_
rlabel metal1 17066 7310 17066 7310 0 _0075_
rlabel metal1 12282 7276 12282 7276 0 _0076_
rlabel metal1 8786 7276 8786 7276 0 _0077_
rlabel metal1 5980 6358 5980 6358 0 _0078_
rlabel metal1 7636 6222 7636 6222 0 _0079_
rlabel metal2 17158 9418 17158 9418 0 _0080_
rlabel metal1 12374 9044 12374 9044 0 _0081_
rlabel metal1 12788 13906 12788 13906 0 _0082_
rlabel metal1 14858 4624 14858 4624 0 _0083_
rlabel metal1 17204 13702 17204 13702 0 _0084_
rlabel metal1 14536 13362 14536 13362 0 _0085_
rlabel metal1 8878 13940 8878 13940 0 _0086_
rlabel metal1 10856 14042 10856 14042 0 _0087_
rlabel metal1 13432 9554 13432 9554 0 _0088_
rlabel metal1 9890 13498 9890 13498 0 _0089_
rlabel metal1 10166 14450 10166 14450 0 _0090_
rlabel metal1 13110 13365 13110 13365 0 _0091_
rlabel metal1 11362 14790 11362 14790 0 _0092_
rlabel metal1 9246 14416 9246 14416 0 _0093_
rlabel metal1 13754 13464 13754 13464 0 _0094_
rlabel metal1 15042 13158 15042 13158 0 _0095_
rlabel metal1 16054 5746 16054 5746 0 _0096_
rlabel metal1 15410 4080 15410 4080 0 _0097_
rlabel metal1 16698 4658 16698 4658 0 _0098_
rlabel metal1 17204 8806 17204 8806 0 _0099_
rlabel metal2 16974 4794 16974 4794 0 _0100_
rlabel metal1 16514 3978 16514 3978 0 _0101_
rlabel metal2 12880 10948 12880 10948 0 _0102_
rlabel metal1 15870 3026 15870 3026 0 _0103_
rlabel metal1 15778 4046 15778 4046 0 _0104_
rlabel metal1 13524 918 13524 918 0 _0105_
rlabel metal1 13248 15674 13248 15674 0 _0106_
rlabel metal1 13662 16422 13662 16422 0 _0107_
rlabel metal1 9246 15572 9246 15572 0 _0108_
rlabel metal1 12466 16048 12466 16048 0 _0109_
rlabel metal2 15134 1037 15134 1037 0 _0110_
rlabel metal1 9338 15640 9338 15640 0 _0111_
rlabel metal1 13110 15946 13110 15946 0 _0112_
rlabel metal1 12880 1394 12880 1394 0 _0113_
rlabel metal1 10120 2550 10120 2550 0 _0114_
rlabel metal1 16376 10574 16376 10574 0 _0115_
rlabel metal1 16514 11220 16514 11220 0 _0116_
rlabel metal1 16790 4590 16790 4590 0 _0117_
rlabel metal1 16330 3502 16330 3502 0 _0118_
rlabel metal1 12006 2992 12006 2992 0 _0119_
rlabel metal1 14122 7922 14122 7922 0 _0120_
rlabel metal1 13340 6086 13340 6086 0 _0121_
rlabel metal1 13478 7854 13478 7854 0 _0122_
rlabel metal1 9246 13702 9246 13702 0 _0123_
rlabel metal1 5888 14790 5888 14790 0 _0124_
rlabel metal2 10994 13345 10994 13345 0 _0125_
rlabel metal1 13018 5678 13018 5678 0 _0126_
rlabel metal1 12190 5712 12190 5712 0 _0127_
rlabel metal2 11362 5270 11362 5270 0 _0128_
rlabel metal2 12558 4284 12558 4284 0 _0129_
rlabel metal2 11822 1870 11822 1870 0 _0130_
rlabel metal1 8970 2312 8970 2312 0 _0131_
rlabel metal1 14168 8398 14168 8398 0 _0132_
rlabel metal1 14030 10574 14030 10574 0 _0133_
rlabel via2 6578 4165 6578 4165 0 _0134_
rlabel metal1 7866 4556 7866 4556 0 _0135_
rlabel metal1 9246 11866 9246 11866 0 _0136_
rlabel metal1 12880 9010 12880 9010 0 _0137_
rlabel metal1 13018 8942 13018 8942 0 _0138_
rlabel metal1 10304 12750 10304 12750 0 _0139_
rlabel metal1 10258 12648 10258 12648 0 _0140_
rlabel metal1 13938 16082 13938 16082 0 _0141_
rlabel metal2 11960 12614 11960 12614 0 _0142_
rlabel metal1 11960 4794 11960 4794 0 _0143_
rlabel metal1 13018 1904 13018 1904 0 _0144_
rlabel metal1 13110 1904 13110 1904 0 _0145_
rlabel metal1 13478 1802 13478 1802 0 _0146_
rlabel metal1 17388 3026 17388 3026 0 _0147_
rlabel metal1 17066 1462 17066 1462 0 _0148_
rlabel metal2 16330 13804 16330 13804 0 _0149_
rlabel metal1 17158 2448 17158 2448 0 _0150_
rlabel metal1 16330 9146 16330 9146 0 _0151_
rlabel metal1 16882 11186 16882 11186 0 _0152_
rlabel metal1 17342 2516 17342 2516 0 _0153_
rlabel metal1 16284 2550 16284 2550 0 _0154_
rlabel metal2 16882 1530 16882 1530 0 _0155_
rlabel metal1 17250 1394 17250 1394 0 _0156_
rlabel metal1 16238 1326 16238 1326 0 _0157_
rlabel metal1 16192 2278 16192 2278 0 _0158_
rlabel metal1 13432 1870 13432 1870 0 _0159_
rlabel metal1 6302 1972 6302 1972 0 _0160_
rlabel metal1 10810 11594 10810 11594 0 _0161_
rlabel via3 12259 11084 12259 11084 0 _0162_
rlabel metal1 15870 10064 15870 10064 0 _0163_
rlabel metal1 15962 13158 15962 13158 0 _0164_
rlabel metal2 15410 2924 15410 2924 0 _0165_
rlabel metal1 15640 1530 15640 1530 0 _0166_
rlabel metal1 16560 1870 16560 1870 0 _0167_
rlabel metal1 17066 2074 17066 2074 0 _0168_
rlabel metal1 16146 1938 16146 1938 0 _0169_
rlabel metal1 14398 1836 14398 1836 0 _0170_
rlabel metal1 11316 1258 11316 1258 0 _0171_
rlabel metal1 11822 8398 11822 8398 0 _0172_
rlabel metal1 11868 8262 11868 8262 0 _0173_
rlabel metal1 10626 6868 10626 6868 0 _0174_
rlabel metal1 8326 13974 8326 13974 0 _0175_
rlabel metal1 8970 3672 8970 3672 0 _0176_
rlabel metal2 5658 13855 5658 13855 0 _0177_
rlabel metal1 11224 7922 11224 7922 0 _0178_
rlabel metal2 7360 5134 7360 5134 0 _0179_
rlabel metal1 11500 11526 11500 11526 0 _0180_
rlabel metal1 10948 5134 10948 5134 0 _0181_
rlabel metal2 10396 1326 10396 1326 0 _0182_
rlabel metal1 10856 1394 10856 1394 0 _0183_
rlabel metal1 4830 5678 4830 5678 0 _0184_
rlabel metal2 9614 4896 9614 4896 0 _0185_
rlabel metal1 5290 7854 5290 7854 0 _0186_
rlabel metal1 8464 7854 8464 7854 0 _0187_
rlabel viali 9890 4659 9890 4659 0 _0188_
rlabel metal1 5888 14518 5888 14518 0 _0189_
rlabel metal1 7912 13838 7912 13838 0 _0190_
rlabel metal1 8878 5678 8878 5678 0 _0191_
rlabel metal2 9522 5134 9522 5134 0 _0192_
rlabel metal2 9522 3604 9522 3604 0 _0193_
rlabel metal1 10580 15334 10580 15334 0 _0194_
rlabel metal1 10672 2278 10672 2278 0 _0195_
rlabel metal2 15502 2176 15502 2176 0 _0196_
rlabel metal1 15318 2448 15318 2448 0 _0197_
rlabel metal1 15778 1870 15778 1870 0 _0198_
rlabel metal2 15686 1581 15686 1581 0 _0199_
rlabel metal1 4094 7378 4094 7378 0 _0200_
rlabel metal1 3358 7310 3358 7310 0 _0201_
rlabel metal2 4278 7072 4278 7072 0 _0202_
rlabel metal1 4738 6868 4738 6868 0 _0203_
rlabel metal1 4140 3026 4140 3026 0 _0204_
rlabel metal1 8970 10132 8970 10132 0 _0205_
rlabel metal1 9292 11662 9292 11662 0 _0206_
rlabel metal1 10212 11118 10212 11118 0 _0207_
rlabel metal1 4324 2958 4324 2958 0 _0208_
rlabel metal2 4278 2652 4278 2652 0 _0209_
rlabel metal1 3956 2482 3956 2482 0 _0210_
rlabel metal1 4002 1360 4002 1360 0 _0211_
rlabel metal1 5198 1292 5198 1292 0 _0212_
rlabel via1 10074 1411 10074 1411 0 _0213_
rlabel metal2 5750 2652 5750 2652 0 _0214_
rlabel metal1 3128 9554 3128 9554 0 _0215_
rlabel metal1 1932 7310 1932 7310 0 _0216_
rlabel metal1 2162 7344 2162 7344 0 _0217_
rlabel metal1 2070 7820 2070 7820 0 _0218_
rlabel metal1 3634 6868 3634 6868 0 _0219_
rlabel metal1 3588 2482 3588 2482 0 _0220_
rlabel metal1 4646 2992 4646 2992 0 _0221_
rlabel viali 4370 1393 4370 1393 0 _0222_
rlabel metal1 4416 1734 4416 1734 0 _0223_
rlabel metal2 3450 1972 3450 1972 0 _0224_
rlabel metal1 3588 1326 3588 1326 0 _0225_
rlabel metal1 5796 1326 5796 1326 0 _0226_
rlabel metal2 6118 4046 6118 4046 0 _0227_
rlabel metal1 7314 2550 7314 2550 0 _0228_
rlabel viali 7682 4657 7682 4657 0 _0229_
rlabel metal2 8832 13396 8832 13396 0 _0230_
rlabel metal1 6394 4692 6394 4692 0 _0231_
rlabel metal1 5428 5270 5428 5270 0 _0232_
rlabel metal1 8510 4590 8510 4590 0 _0233_
rlabel metal1 8263 4658 8263 4658 0 _0234_
rlabel metal1 6440 1326 6440 1326 0 _0235_
rlabel metal1 8142 1428 8142 1428 0 _0236_
rlabel metal1 2392 2958 2392 2958 0 _0237_
rlabel metal1 2070 3604 2070 3604 0 _0238_
rlabel metal2 2162 3366 2162 3366 0 _0239_
rlabel metal1 2116 1870 2116 1870 0 _0240_
rlabel metal1 2024 1394 2024 1394 0 _0241_
rlabel metal1 2254 1734 2254 1734 0 _0242_
rlabel metal1 2576 1530 2576 1530 0 _0243_
rlabel metal2 2990 1564 2990 1564 0 _0244_
rlabel metal1 3404 2074 3404 2074 0 _0245_
rlabel metal1 2392 714 2392 714 0 _0246_
rlabel metal1 5014 2006 5014 2006 0 _0247_
rlabel via1 2622 5117 2622 5117 0 _0248_
rlabel metal1 5796 7718 5796 7718 0 _0249_
rlabel metal1 5060 14518 5060 14518 0 _0250_
rlabel metal2 5566 13333 5566 13333 0 _0251_
rlabel metal1 5842 4080 5842 4080 0 _0252_
rlabel metal2 5382 2958 5382 2958 0 _0253_
rlabel metal1 6026 2550 6026 2550 0 _0254_
rlabel metal1 2116 3706 2116 3706 0 _0255_
rlabel metal1 1656 1870 1656 1870 0 _0256_
rlabel metal1 5198 8330 5198 8330 0 _0257_
rlabel metal3 6302 2516 6302 2516 0 _0258_
rlabel metal1 1656 1938 1656 1938 0 _0259_
rlabel metal1 2530 1836 2530 1836 0 _0260_
rlabel metal2 2806 1462 2806 1462 0 _0261_
rlabel metal2 2530 1190 2530 1190 0 _0262_
rlabel metal1 3174 1530 3174 1530 0 _0263_
rlabel metal1 7084 17034 7084 17034 0 _0264_
rlabel metal1 5612 14994 5612 14994 0 _0265_
rlabel metal1 6946 16218 6946 16218 0 _0266_
rlabel metal1 6164 15674 6164 15674 0 _0267_
rlabel metal2 6578 16898 6578 16898 0 _0268_
rlabel metal1 8050 16048 8050 16048 0 _0269_
rlabel metal2 9246 7650 9246 7650 0 _0270_
rlabel metal1 1334 5100 1334 5100 0 _0271_
rlabel metal1 6026 7514 6026 7514 0 _0272_
rlabel metal2 7130 6528 7130 6528 0 _0273_
rlabel metal1 7084 5746 7084 5746 0 _0274_
rlabel metal1 6716 5542 6716 5542 0 _0275_
rlabel metal2 9062 2108 9062 2108 0 _0276_
rlabel metal1 13248 10234 13248 10234 0 _0277_
rlabel metal1 14720 8874 14720 8874 0 _0278_
rlabel metal2 15134 6290 15134 6290 0 _0279_
rlabel metal1 16514 6256 16514 6256 0 _0280_
rlabel metal1 8878 6256 8878 6256 0 _0281_
rlabel metal1 13018 6392 13018 6392 0 _0282_
rlabel metal1 10120 7310 10120 7310 0 _0283_
rlabel metal1 8050 6732 8050 6732 0 _0284_
rlabel metal1 14812 7922 14812 7922 0 _0285_
rlabel metal2 11730 13333 11730 13333 0 _0286_
rlabel metal1 7866 6766 7866 6766 0 _0287_
rlabel metal1 14674 6256 14674 6256 0 _0288_
rlabel metal1 14812 4114 14812 4114 0 _0289_
rlabel metal2 14214 3332 14214 3332 0 _0290_
rlabel metal1 14030 6732 14030 6732 0 _0291_
rlabel metal1 14904 2550 14904 2550 0 _0292_
rlabel via2 13846 3043 13846 3043 0 _0293_
rlabel metal1 9430 5134 9430 5134 0 _0294_
rlabel metal1 6256 5202 6256 5202 0 _0295_
rlabel metal1 8694 5304 8694 5304 0 _0296_
rlabel metal1 13294 3638 13294 3638 0 _0297_
rlabel metal1 8234 3536 8234 3536 0 _0298_
rlabel metal1 13984 3026 13984 3026 0 _0299_
rlabel metal1 13294 3026 13294 3026 0 _0300_
rlabel metal2 14030 3910 14030 3910 0 _0301_
rlabel metal2 13846 4658 13846 4658 0 _0302_
rlabel metal1 14076 4046 14076 4046 0 _0303_
rlabel metal1 12972 4114 12972 4114 0 _0304_
rlabel metal1 13570 1428 13570 1428 0 _0305_
rlabel metal1 7866 1258 7866 1258 0 _0306_
rlabel metal1 10350 7888 10350 7888 0 _0307_
rlabel metal1 7544 6834 7544 6834 0 _0308_
rlabel metal1 11132 6222 11132 6222 0 _0309_
rlabel metal2 11086 6596 11086 6596 0 _0310_
rlabel metal1 9936 986 9936 986 0 _0311_
rlabel metal1 9430 8364 9430 8364 0 _0312_
rlabel metal1 2346 11186 2346 11186 0 _0313_
rlabel metal1 9982 3604 9982 3604 0 _0314_
rlabel metal1 9890 3094 9890 3094 0 _0315_
rlabel metal2 9246 1700 9246 1700 0 _0316_
rlabel metal2 1748 4964 1748 4964 0 _0317_
rlabel metal1 8050 3604 8050 3604 0 _0318_
rlabel metal1 7774 3026 7774 3026 0 _0319_
rlabel metal1 7958 1462 7958 1462 0 _0320_
rlabel metal1 5704 7514 5704 7514 0 _0321_
rlabel metal1 1886 12784 1886 12784 0 _0322_
rlabel via1 6039 2958 6039 2958 0 _0323_
rlabel metal1 6256 2958 6256 2958 0 _0324_
rlabel metal1 5888 2822 5888 2822 0 _0325_
rlabel metal2 7866 714 7866 714 0 _0326_
rlabel metal3 5198 7276 5198 7276 0 _0327_
rlabel metal1 8602 6324 8602 6324 0 _0328_
rlabel metal1 7728 6426 7728 6426 0 _0329_
rlabel metal1 7774 1394 7774 1394 0 _0330_
rlabel metal1 14536 3502 14536 3502 0 _0331_
rlabel metal2 14490 4012 14490 4012 0 _0332_
rlabel metal1 9936 6766 9936 6766 0 _0333_
rlabel metal2 10534 7361 10534 7361 0 _0334_
rlabel metal1 10994 7718 10994 7718 0 _0335_
rlabel metal2 13846 7820 13846 7820 0 _0336_
rlabel metal1 13708 8398 13708 8398 0 _0337_
rlabel metal1 13524 7922 13524 7922 0 _0338_
rlabel metal1 15134 7310 15134 7310 0 _0339_
rlabel metal2 14214 3604 14214 3604 0 _0340_
rlabel metal1 14812 986 14812 986 0 _0341_
rlabel metal1 14628 2414 14628 2414 0 _0342_
rlabel metal2 14260 2652 14260 2652 0 _0343_
rlabel metal1 14858 7310 14858 7310 0 _0344_
rlabel metal3 14697 2652 14697 2652 0 _0345_
rlabel metal1 14352 986 14352 986 0 _0346_
rlabel metal2 13938 4148 13938 4148 0 _0347_
rlabel metal2 14030 6970 14030 6970 0 _0348_
rlabel metal1 14260 7310 14260 7310 0 _0349_
rlabel metal1 13478 4658 13478 4658 0 _0350_
rlabel metal2 14306 4012 14306 4012 0 _0351_
rlabel metal1 9614 2006 9614 2006 0 _0352_
rlabel metal1 6486 3060 6486 3060 0 _0353_
rlabel metal1 11362 7412 11362 7412 0 _0354_
rlabel metal1 11178 7378 11178 7378 0 _0355_
rlabel metal1 11592 7922 11592 7922 0 _0356_
rlabel metal1 11592 7378 11592 7378 0 _0357_
rlabel metal1 11132 986 11132 986 0 _0358_
rlabel metal1 10534 3604 10534 3604 0 _0359_
rlabel metal1 10626 3468 10626 3468 0 _0360_
rlabel metal1 6256 5338 6256 5338 0 _0361_
rlabel metal1 10304 3570 10304 3570 0 _0362_
rlabel metal1 12052 1190 12052 1190 0 _0363_
rlabel metal2 7038 1700 7038 1700 0 _0364_
rlabel metal1 7222 1938 7222 1938 0 _0365_
rlabel metal1 7176 4046 7176 4046 0 _0366_
rlabel metal1 7038 1802 7038 1802 0 _0367_
rlabel metal2 8970 1360 8970 1360 0 _0368_
rlabel metal1 6578 2890 6578 2890 0 _0369_
rlabel viali 6674 3026 6674 3026 0 _0370_
rlabel metal1 6348 4046 6348 4046 0 _0371_
rlabel metal2 6394 3434 6394 3434 0 _0372_
rlabel metal1 9522 1836 9522 1836 0 _0373_
rlabel metal2 9522 7106 9522 7106 0 _0374_
rlabel metal1 9522 7174 9522 7174 0 _0375_
rlabel metal2 8878 2074 8878 2074 0 _0376_
rlabel metal1 8556 1870 8556 1870 0 _0377_
rlabel metal1 10810 13498 10810 13498 0 _0378_
rlabel metal1 6946 13702 6946 13702 0 _0379_
rlabel metal1 9890 14824 9890 14824 0 _0380_
rlabel metal2 8602 15232 8602 15232 0 _0381_
rlabel viali 8418 14931 8418 14931 0 _0382_
rlabel metal1 8280 15538 8280 15538 0 _0383_
rlabel metal2 4922 15334 4922 15334 0 _0384_
rlabel metal1 6578 15334 6578 15334 0 _0385_
rlabel metal1 7590 15572 7590 15572 0 _0386_
rlabel metal2 7314 16694 7314 16694 0 _0387_
rlabel metal1 7038 12750 7038 12750 0 _0388_
rlabel metal1 6946 14518 6946 14518 0 _0389_
rlabel metal1 7498 14586 7498 14586 0 _0390_
rlabel metal1 7636 15130 7636 15130 0 _0391_
rlabel metal2 7222 14331 7222 14331 0 _0392_
rlabel metal1 8004 15674 8004 15674 0 _0393_
rlabel metal1 7590 16150 7590 16150 0 _0394_
rlabel metal1 1886 17068 1886 17068 0 _0395_
rlabel metal1 7084 10506 7084 10506 0 _0396_
rlabel metal1 7360 9962 7360 9962 0 _0397_
rlabel metal1 16652 10166 16652 10166 0 _0398_
rlabel metal1 5658 10098 5658 10098 0 _0399_
rlabel metal1 7958 11050 7958 11050 0 _0400_
rlabel metal1 4968 10234 4968 10234 0 _0401_
rlabel metal1 5428 10234 5428 10234 0 _0402_
rlabel via2 6394 10659 6394 10659 0 _0403_
rlabel metal1 15134 10710 15134 10710 0 _0404_
rlabel metal1 7958 9010 7958 9010 0 _0405_
rlabel metal3 5336 7820 5336 7820 0 _0406_
rlabel metal1 14766 10540 14766 10540 0 _0407_
rlabel metal1 15640 10778 15640 10778 0 _0408_
rlabel metal2 14398 11577 14398 11577 0 _0409_
rlabel metal1 13984 11526 13984 11526 0 _0410_
rlabel metal1 14122 9520 14122 9520 0 _0411_
rlabel metal1 14812 11322 14812 11322 0 _0412_
rlabel metal1 13386 10778 13386 10778 0 _0413_
rlabel metal1 14214 11594 14214 11594 0 _0414_
rlabel metal1 14214 11866 14214 11866 0 _0415_
rlabel metal1 12466 11560 12466 11560 0 _0416_
rlabel metal1 11914 11628 11914 11628 0 _0417_
rlabel metal1 2530 5712 2530 5712 0 _0418_
rlabel metal1 13938 12750 13938 12750 0 _0419_
rlabel metal2 9568 10132 9568 10132 0 _0420_
rlabel metal1 2714 5780 2714 5780 0 _0421_
rlabel metal2 3082 5270 3082 5270 0 _0422_
rlabel metal1 3174 5338 3174 5338 0 _0423_
rlabel metal1 1426 5168 1426 5168 0 _0424_
rlabel metal1 3450 4692 3450 4692 0 _0425_
rlabel metal1 1426 4998 1426 4998 0 _0426_
rlabel metal1 1518 5338 1518 5338 0 _0427_
rlabel metal1 1916 5066 1916 5066 0 _0428_
rlabel metal1 1426 4692 1426 4692 0 _0429_
rlabel metal1 15962 12682 15962 12682 0 _0430_
rlabel via2 5290 13821 5290 13821 0 _0431_
rlabel metal1 12742 14314 12742 14314 0 _0432_
rlabel metal2 15042 16286 15042 16286 0 _0433_
rlabel metal1 15180 14926 15180 14926 0 _0434_
rlabel metal1 5566 13940 5566 13940 0 _0435_
rlabel metal1 5014 13872 5014 13872 0 _0436_
rlabel metal1 3726 13770 3726 13770 0 _0437_
rlabel metal1 4784 13838 4784 13838 0 _0438_
rlabel metal1 5888 12274 5888 12274 0 _0439_
rlabel metal2 5106 12585 5106 12585 0 _0440_
rlabel metal1 2254 11764 2254 11764 0 _0441_
rlabel metal1 13708 14042 13708 14042 0 _0442_
rlabel via1 2622 14365 2622 14365 0 _0443_
rlabel via1 1970 11526 1970 11526 0 _0444_
rlabel via2 12558 12835 12558 12835 0 _0445_
rlabel metal1 3634 12376 3634 12376 0 _0446_
rlabel metal2 3036 12308 3036 12308 0 _0447_
rlabel metal1 2070 11322 2070 11322 0 _0448_
rlabel via1 6775 9418 6775 9418 0 _0449_
rlabel metal1 1518 10540 1518 10540 0 _0450_
rlabel metal1 1702 11662 1702 11662 0 _0451_
rlabel metal1 1426 11628 1426 11628 0 _0452_
rlabel metal1 1702 14246 1702 14246 0 _0453_
rlabel metal1 1334 12716 1334 12716 0 _0454_
rlabel metal1 1748 14518 1748 14518 0 _0455_
rlabel metal1 2622 15402 2622 15402 0 _0456_
rlabel metal2 2898 14960 2898 14960 0 _0457_
rlabel metal1 3082 15504 3082 15504 0 _0458_
rlabel metal1 1610 15572 1610 15572 0 _0459_
rlabel metal1 16054 15538 16054 15538 0 _0460_
rlabel metal1 15548 15538 15548 15538 0 _0461_
rlabel metal1 13432 16218 13432 16218 0 _0462_
rlabel metal1 12558 15436 12558 15436 0 _0463_
rlabel metal1 9154 17068 9154 17068 0 _0464_
rlabel metal1 13570 15572 13570 15572 0 _0465_
rlabel metal1 11178 16626 11178 16626 0 _0466_
rlabel metal1 9936 16626 9936 16626 0 _0467_
rlabel metal1 4830 16660 4830 16660 0 _0468_
rlabel metal1 5934 8976 5934 8976 0 _0469_
rlabel metal1 13800 10506 13800 10506 0 _0470_
rlabel metal1 15410 7956 15410 7956 0 _0471_
rlabel metal1 14720 9146 14720 9146 0 _0472_
rlabel metal1 16100 7718 16100 7718 0 _0473_
rlabel metal1 15832 8058 15832 8058 0 _0474_
rlabel metal1 16652 7922 16652 7922 0 _0475_
rlabel metal1 12535 10438 12535 10438 0 _0476_
rlabel metal2 7360 9894 7360 9894 0 _0477_
rlabel metal1 10810 9078 10810 9078 0 _0478_
rlabel metal1 10350 10132 10350 10132 0 _0479_
rlabel metal1 6808 9350 6808 9350 0 _0480_
rlabel metal2 8142 8194 8142 8194 0 _0481_
rlabel viali 10176 9010 10176 9010 0 _0482_
rlabel metal1 9430 8602 9430 8602 0 _0483_
rlabel metal2 9798 8772 9798 8772 0 _0484_
rlabel metal1 7314 8602 7314 8602 0 _0485_
rlabel metal1 6900 8058 6900 8058 0 _0486_
rlabel metal1 6854 9044 6854 9044 0 _0487_
rlabel metal1 6210 8602 6210 8602 0 _0488_
rlabel metal1 6854 8466 6854 8466 0 _0489_
rlabel metal1 6026 8432 6026 8432 0 _0490_
rlabel metal2 6210 9248 6210 9248 0 _0491_
rlabel metal1 7406 8942 7406 8942 0 _0492_
rlabel metal1 6992 9146 6992 9146 0 _0493_
rlabel metal1 7866 10744 7866 10744 0 _0494_
rlabel metal1 6670 10234 6670 10234 0 _0495_
rlabel metal1 7038 10030 7038 10030 0 _0496_
rlabel metal1 6946 9894 6946 9894 0 _0497_
rlabel metal2 5290 7582 5290 7582 0 _0498_
rlabel metal1 8050 11288 8050 11288 0 _0499_
rlabel metal1 9430 11322 9430 11322 0 _0500_
rlabel metal2 8326 12121 8326 12121 0 _0501_
rlabel metal1 7222 11016 7222 11016 0 _0502_
rlabel metal1 6210 9622 6210 9622 0 _0503_
rlabel metal1 7498 12206 7498 12206 0 _0504_
rlabel via2 7958 12427 7958 12427 0 _0505_
rlabel metal1 8878 11322 8878 11322 0 _0506_
rlabel metal1 8372 11866 8372 11866 0 _0507_
rlabel metal1 11638 9350 11638 9350 0 _0508_
rlabel metal1 7958 11866 7958 11866 0 _0509_
rlabel metal1 6992 12274 6992 12274 0 _0510_
rlabel metal1 6026 12954 6026 12954 0 _0511_
rlabel metal1 3910 17306 3910 17306 0 b6
rlabel metal1 7176 17306 7176 17306 0 b7
rlabel metal2 5750 398 5750 398 0 b[0]
rlabel metal2 5014 398 5014 398 0 b[1]
rlabel metal2 4278 500 4278 500 0 b[2]
rlabel metal2 3542 398 3542 398 0 b[3]
rlabel metal2 2806 500 2806 500 0 b[4]
rlabel metal2 2070 636 2070 636 0 b[5]
rlabel metal2 1334 500 1334 500 0 b[6]
rlabel metal2 598 500 598 500 0 b[7]
rlabel metal1 10580 10574 10580 10574 0 clk
rlabel metal2 11362 11662 11362 11662 0 clknet_0_clk
rlabel metal1 1380 4046 1380 4046 0 clknet_2_0__leaf_clk
rlabel metal1 3450 12750 3450 12750 0 clknet_2_1__leaf_clk
rlabel metal1 15548 12750 15548 12750 0 clknet_2_2__leaf_clk
rlabel metal1 9614 16660 9614 16660 0 clknet_2_3__leaf_clk
rlabel metal1 15042 16422 15042 16422 0 divider\[0\]
rlabel metal2 9522 14144 9522 14144 0 divider\[1\]
rlabel metal1 4646 17306 4646 17306 0 g6
rlabel metal1 8004 17306 8004 17306 0 g7
rlabel metal2 11638 772 11638 772 0 g[0]
rlabel metal2 10902 398 10902 398 0 g[1]
rlabel metal2 10166 500 10166 500 0 g[2]
rlabel metal2 9430 636 9430 636 0 g[3]
rlabel metal2 8694 398 8694 398 0 g[4]
rlabel metal2 7958 398 7958 398 0 g[5]
rlabel metal2 7222 500 7222 500 0 g[6]
rlabel metal2 6486 398 6486 398 0 g[7]
rlabel metal1 17020 15538 17020 15538 0 gate
rlabel metal2 1242 17588 1242 17588 0 hblank
rlabel metal1 4094 17238 4094 17238 0 hsync
rlabel metal1 12742 14892 12742 14892 0 mode\[0\]
rlabel metal1 12926 16524 12926 16524 0 mode\[1\]
rlabel metal1 10764 16218 10764 16218 0 mode\[2\]
rlabel metal1 13846 14892 13846 14892 0 net1
rlabel metal1 1748 1394 1748 1394 0 net10
rlabel metal1 1288 1394 1288 1394 0 net11
rlabel metal2 12834 714 12834 714 0 net12
rlabel metal2 5382 986 5382 986 0 net13
rlabel metal2 12558 799 12558 799 0 net14
rlabel metal1 4048 782 4048 782 0 net15
rlabel metal1 3542 748 3542 748 0 net16
rlabel metal1 2898 816 2898 816 0 net17
rlabel metal1 1702 782 1702 782 0 net18
rlabel metal2 1150 986 1150 986 0 net19
rlabel metal1 16284 16626 16284 16626 0 net2
rlabel via2 5842 2635 5842 2635 0 net20
rlabel metal1 6946 1462 6946 1462 0 net21
rlabel metal1 12240 1462 12240 1462 0 net22
rlabel metal2 12466 1088 12466 1088 0 net23
rlabel metal1 12926 952 12926 952 0 net24
rlabel metal1 10350 714 10350 714 0 net25
rlabel metal1 8234 816 8234 816 0 net26
rlabel metal2 8510 1054 8510 1054 0 net27
rlabel metal1 7314 748 7314 748 0 net28
rlabel metal1 6808 782 6808 782 0 net29
rlabel metal1 15410 15946 15410 15946 0 net3
rlabel metal1 1518 17136 1518 17136 0 net30
rlabel metal1 3818 17034 3818 17034 0 net31
rlabel metal3 9223 2380 9223 2380 0 net32
rlabel metal2 8602 1785 8602 1785 0 net33
rlabel metal1 15180 986 15180 986 0 net34
rlabel metal1 14766 680 14766 680 0 net35
rlabel metal1 14996 1258 14996 1258 0 net36
rlabel metal1 14766 408 14766 408 0 net37
rlabel metal1 15640 1462 15640 1462 0 net38
rlabel metal1 16238 306 16238 306 0 net39
rlabel metal1 14628 16014 14628 16014 0 net4
rlabel metal1 15502 748 15502 748 0 net40
rlabel metal1 13478 782 13478 782 0 net41
rlabel metal1 2944 16626 2944 16626 0 net42
rlabel metal2 6394 16864 6394 16864 0 net43
rlabel metal1 2990 17034 2990 17034 0 net44
rlabel metal1 10304 16762 10304 16762 0 net45
rlabel metal2 6578 13804 6578 13804 0 net46
rlabel metal1 11546 17204 11546 17204 0 net47
rlabel metal1 13110 17000 13110 17000 0 net5
rlabel metal2 12834 16354 12834 16354 0 net6
rlabel metal1 13294 17238 13294 17238 0 net7
rlabel metal1 10212 16626 10212 16626 0 net8
rlabel metal1 9246 16014 9246 16014 0 net9
rlabel metal1 5658 17306 5658 17306 0 r6
rlabel metal1 8786 17306 8786 17306 0 r7
rlabel metal2 17526 1350 17526 1350 0 r[0]
rlabel metal1 16698 2822 16698 2822 0 r[1]
rlabel metal2 16054 755 16054 755 0 r[2]
rlabel metal2 15318 942 15318 942 0 r[3]
rlabel metal2 14582 415 14582 415 0 r[4]
rlabel metal2 13846 415 13846 415 0 r[5]
rlabel metal2 13110 415 13110 415 0 r[6]
rlabel metal1 13018 680 13018 680 0 r[7]
rlabel viali 16338 5746 16338 5746 0 rampc\[0\]
rlabel viali 15594 11185 15594 11185 0 rampc\[1\]
rlabel metal1 16422 13838 16422 13838 0 rampc\[2\]
rlabel metal1 13202 11662 13202 11662 0 rampc\[3\]
rlabel metal1 2484 6834 2484 6834 0 rampc\[4\]
rlabel metal1 2254 6188 2254 6188 0 rampc\[5\]
rlabel metal1 2622 3604 2622 3604 0 rampc\[6\]
rlabel metal1 2024 3910 2024 3910 0 rampc\[7\]
rlabel metal1 15916 16966 15916 16966 0 registered
rlabel metal1 16192 17170 16192 17170 0 rst_n
rlabel metal1 17158 16660 17158 16660 0 ui_in[0]
rlabel metal1 15778 16694 15778 16694 0 ui_in[1]
rlabel metal1 15042 16626 15042 16626 0 ui_in[2]
rlabel metal1 14214 17102 14214 17102 0 ui_in[3]
rlabel metal1 13202 17068 13202 17068 0 ui_in[4]
rlabel metal1 13708 17102 13708 17102 0 ui_in[5]
rlabel metal1 10120 17102 10120 17102 0 ui_in[6]
rlabel metal1 9660 17102 9660 17102 0 ui_in[7]
rlabel metal2 2070 17588 2070 17588 0 vblank
rlabel metal1 17066 12954 17066 12954 0 vga_sync.hpos\[0\]
rlabel metal1 17112 13838 17112 13838 0 vga_sync.hpos\[1\]
rlabel metal1 15824 14450 15824 14450 0 vga_sync.hpos\[2\]
rlabel metal1 9890 13294 9890 13294 0 vga_sync.hpos\[3\]
rlabel metal1 2714 8024 2714 8024 0 vga_sync.hpos\[4\]
rlabel metal1 2254 7888 2254 7888 0 vga_sync.hpos\[5\]
rlabel metal1 2438 4046 2438 4046 0 vga_sync.hpos\[6\]
rlabel metal1 4830 15606 4830 15606 0 vga_sync.hpos\[7\]
rlabel metal1 4416 16422 4416 16422 0 vga_sync.hpos\[8\]
rlabel metal1 3174 15606 3174 15606 0 vga_sync.hpos\[9\]
rlabel metal2 3312 15878 3312 15878 0 vga_sync.mode
rlabel metal1 17066 9078 17066 9078 0 vga_sync.o_vpos\[0\]
rlabel metal1 16514 9452 16514 9452 0 vga_sync.o_vpos\[1\]
rlabel metal1 15410 10132 15410 10132 0 vga_sync.o_vpos\[2\]
rlabel metal2 9798 9894 9798 9894 0 vga_sync.o_vpos\[3\]
rlabel metal1 4232 9486 4232 9486 0 vga_sync.o_vpos\[4\]
rlabel metal1 4922 9486 4922 9486 0 vga_sync.o_vpos\[5\]
rlabel metal1 1702 2924 1702 2924 0 vga_sync.o_vpos\[6\]
rlabel metal1 3818 9520 3818 9520 0 vga_sync.o_vpos\[7\]
rlabel metal1 4922 10030 4922 10030 0 vga_sync.o_vpos\[8\]
rlabel metal1 5290 11152 5290 11152 0 vga_sync.o_vpos\[9\]
rlabel metal2 6210 15436 6210 15436 0 vga_sync.vsync
rlabel metal1 7314 17238 7314 17238 0 vsync
<< properties >>
string FIXED_BBOX 0 0 18261 18245
<< end >>
