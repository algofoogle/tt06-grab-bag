magic
tech sky130A
magscale 1 2
timestamp 1713544590
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 545 163 735 203
rect 1 27 735 163
rect 30 -17 64 27
rect 545 21 735 27
<< scnmos >>
rect 79 53 109 137
rect 267 53 297 137
rect 358 53 388 137
rect 442 53 472 137
rect 526 53 556 137
rect 624 47 654 177
<< scpmoshvt >>
rect 79 297 109 381
rect 267 297 297 381
rect 362 297 392 381
rect 435 297 465 381
rect 526 297 556 381
rect 624 297 654 497
<< ndiff >>
rect 571 137 624 177
rect 27 117 79 137
rect 27 83 35 117
rect 69 83 79 117
rect 27 53 79 83
rect 109 117 161 137
rect 109 83 119 117
rect 153 83 161 117
rect 109 53 161 83
rect 215 117 267 137
rect 215 83 223 117
rect 257 83 267 117
rect 215 53 267 83
rect 297 111 358 137
rect 297 77 313 111
rect 347 77 358 111
rect 297 53 358 77
rect 388 97 442 137
rect 388 63 398 97
rect 432 63 442 97
rect 388 53 442 63
rect 472 111 526 137
rect 472 77 482 111
rect 516 77 526 111
rect 472 53 526 77
rect 556 97 624 137
rect 556 63 576 97
rect 610 63 624 97
rect 556 53 624 63
rect 571 47 624 53
rect 654 135 709 177
rect 654 101 664 135
rect 698 101 709 135
rect 654 47 709 101
<< pdiff >>
rect 571 485 624 497
rect 571 451 579 485
rect 613 451 624 485
rect 571 417 624 451
rect 571 383 579 417
rect 613 383 624 417
rect 571 381 624 383
rect 27 361 79 381
rect 27 327 35 361
rect 69 327 79 361
rect 27 297 79 327
rect 109 361 161 381
rect 109 327 119 361
rect 153 327 161 361
rect 109 297 161 327
rect 215 354 267 381
rect 215 320 223 354
rect 257 320 267 354
rect 215 297 267 320
rect 297 297 362 381
rect 392 297 435 381
rect 465 297 526 381
rect 556 297 624 381
rect 654 454 709 497
rect 654 420 664 454
rect 698 420 709 454
rect 654 386 709 420
rect 654 352 664 386
rect 698 352 709 386
rect 654 297 709 352
<< ndiffc >>
rect 35 83 69 117
rect 119 83 153 117
rect 223 83 257 117
rect 313 77 347 111
rect 398 63 432 97
rect 482 77 516 111
rect 576 63 610 97
rect 664 101 698 135
<< pdiffc >>
rect 579 451 613 485
rect 579 383 613 417
rect 35 327 69 361
rect 119 327 153 361
rect 223 320 257 354
rect 664 420 698 454
rect 664 352 698 386
<< poly >>
rect 624 497 654 523
rect 426 473 492 483
rect 426 439 442 473
rect 476 439 492 473
rect 426 433 492 439
rect 427 431 491 433
rect 428 429 490 431
rect 79 381 109 407
rect 267 381 297 407
rect 362 381 392 407
rect 435 381 465 429
rect 526 381 556 407
rect 79 265 109 297
rect 267 265 297 297
rect 362 265 392 297
rect 21 249 109 265
rect 21 215 35 249
rect 69 215 109 249
rect 21 199 109 215
rect 206 249 297 265
rect 206 215 216 249
rect 250 215 297 249
rect 206 199 297 215
rect 339 249 393 265
rect 339 215 349 249
rect 383 215 393 249
rect 339 199 393 215
rect 79 137 109 199
rect 267 137 297 199
rect 358 137 388 199
rect 435 182 465 297
rect 526 265 556 297
rect 624 265 654 297
rect 511 249 565 265
rect 511 215 521 249
rect 555 215 565 249
rect 511 199 565 215
rect 607 249 661 265
rect 607 215 617 249
rect 651 215 661 249
rect 607 199 661 215
rect 435 152 472 182
rect 442 137 472 152
rect 526 137 556 199
rect 624 177 654 199
rect 79 27 109 53
rect 267 27 297 53
rect 358 27 388 53
rect 442 27 472 53
rect 526 27 556 53
rect 624 21 654 47
<< polycont >>
rect 442 439 476 473
rect 35 215 69 249
rect 216 215 250 249
rect 349 215 383 249
rect 521 215 555 249
rect 617 215 651 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 361 85 527
rect 566 485 622 527
rect 122 473 532 483
rect 122 439 442 473
rect 476 439 532 473
rect 122 425 532 439
rect 566 451 579 485
rect 613 451 622 485
rect 566 417 622 451
rect 17 327 35 361
rect 69 327 85 361
rect 17 312 85 327
rect 119 361 167 384
rect 153 327 167 361
rect 119 265 167 327
rect 206 357 532 391
rect 566 383 579 417
rect 613 383 622 417
rect 566 367 622 383
rect 664 454 719 493
rect 698 420 719 454
rect 664 386 719 420
rect 206 354 270 357
rect 206 320 223 354
rect 257 320 270 354
rect 498 333 532 357
rect 698 352 719 386
rect 206 299 270 320
rect 17 249 85 265
rect 17 215 35 249
rect 69 215 85 249
rect 17 151 85 215
rect 119 249 250 265
rect 119 215 216 249
rect 119 199 250 215
rect 304 249 452 323
rect 498 299 630 333
rect 664 299 719 352
rect 596 265 630 299
rect 304 215 349 249
rect 383 215 452 249
rect 304 199 452 215
rect 486 249 562 265
rect 486 215 521 249
rect 555 215 562 249
rect 486 199 562 215
rect 596 249 651 265
rect 596 215 617 249
rect 596 199 651 215
rect 119 117 168 199
rect 596 165 630 199
rect 313 131 630 165
rect 685 152 719 299
rect 664 135 719 152
rect 17 83 35 117
rect 69 83 85 117
rect 17 17 85 83
rect 153 83 168 117
rect 119 61 168 83
rect 207 83 223 117
rect 257 83 273 117
rect 207 17 273 83
rect 313 111 347 131
rect 482 111 516 131
rect 313 61 347 77
rect 382 63 398 97
rect 432 63 448 97
rect 382 17 448 63
rect 698 101 719 135
rect 482 61 516 77
rect 550 63 576 97
rect 610 63 626 97
rect 664 83 719 101
rect 550 17 626 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 122 425 156 459 0 FreeSans 400 0 0 0 B
port 6 nsew
flabel locali s 30 153 64 187 0 FreeSans 400 0 0 0 D_N
port 10 nsew
flabel locali s 305 425 339 459 0 FreeSans 400 0 0 0 B
port 6 nsew
flabel locali s 213 425 247 459 0 FreeSans 400 0 0 0 B
port 6 nsew
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 A
port 8 nsew
flabel locali s 673 357 707 391 0 FreeSans 200 0 0 0 X
port 9 nsew
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 C
port 7 nsew
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 C
port 7 nsew
flabel locali s 397 425 431 459 0 FreeSans 400 0 0 0 B
port 6 nsew
flabel locali s 397 289 431 323 0 FreeSans 400 0 0 0 C
port 7 nsew
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 D_N
port 10 nsew
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 C
port 7 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 or4b_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 339122
string GDS_FILE controller.gds
string GDS_START 331898
string path 0.000 0.000 3.680 0.000 
<< end >>
