** sch_path: /home/anton/projects/tt06-grab-bag/xschem/tb_r2rV2.sch
**.subckt tb_r2rV2
x1 a_int d7 d6 d5 d4 d3 d2 d1 d0 GND GND r2r
x2 out c_int GND tt06_analog_load
V1 d0 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 20ns 40ns)
V2 d1 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 40ns 80ns)
V3 d6 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 80ns 160ns)
V4 d2 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 160ns 320ns)
V5 d3 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 320ns 640ns)
V6 d4 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 640ns 1280ns)
V7 d5 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 1280ns 2560ns)
V8 d7 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 2560ns 5120ns)
x3 a_int_parax d7 d6 d5 d4 d3 d2 d1 d0 GND GND r2r_parax
x4 out_parax a_int_parax GND tt06_analog_load
V10 VCC GND 1.8
R4 out GND 1e6 m=1
V9 net1 GND pwl(0ns,0.15v 5ns,0.15v 3us,0.85v 3.002us,0.15v 3.15us,0.15v 3.152us,0.85v 6us,0.15v 7us,0.15v)
R5 b_int a_int 250k m=1
V11 NBIAS GND 1.1
R1 a_int VCC 50k m=1
R2 GND b_int 400k m=1
x5jo VCC net3 net2 b_int c_int GND j_opamp
I0 net3 GND 150u
R3 GND net2 300k m=1
R6 net2 c_int 50k m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/anton/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.tech/ngspice/sky130.lib.spice tt





* .options filetype=ascii
.options savecurrents
.control
  save all
  tran 2n 7u uic
  *set filetype=ascii
  write tb_r2rV2.raw
  quit
.endc
.end



**** end user architecture code
**.ends

* expanding   symbol:  r2r.sym # of pins=11
** sym_path: /home/anton/projects/tt06-grab-bag/xschem/r2r.sym
** sch_path: /home/anton/projects/tt06-grab-bag/xschem/r2r.sch
.subckt r2r aout d7 d6 d5 d4 d3 d2 d1 d0 GND VSUBS
*.ipin d0
*.ipin d1
*.ipin d2
*.ipin d3
*.ipin d4
*.ipin d5
*.ipin d6
*.ipin d7
*.iopin GND
*.iopin VSUBS
*.opin aout
XR1 d0 net1 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR2 d1 net2 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR3 d2 net3 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR4 d3 net4 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR5 d4 net5 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR6 d5 net6 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR7 d6 net7 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR8 d7 aout VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR9 GND net1 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR10 net1 net2 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR11 net2 net3 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR12 net3 net4 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR13 net4 net5 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR14 net5 net6 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR15 net6 net7 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR16 net7 aout VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
.ends


* expanding   symbol:  tt06_analog_load.sym # of pins=3
** sym_path: /home/anton/projects/tt06-grab-bag/xschem/tt06_analog_load.sym
** sch_path: /home/anton/projects/tt06-grab-bag/xschem/tt06_analog_load.sch
.subckt tt06_analog_load a_ext a_int GND
*.iopin a_int
*.iopin a_ext
*.iopin GND
R1 a_ext a_int 500 m=1
C1 a_int GND 2.5p m=1
C2 a_ext GND 2.5p m=1
.ends


* expanding   symbol:  j_opamp.sym # of pins=6
** sym_path: /home/anton/projects/tt06-grab-bag/xschem/j_opamp.sym
** sch_path: /home/anton/projects/tt06-grab-bag/xschem/j_opamp.sch
.subckt j_opamp vdd iref vin_n vin_p vout vss
*.iopin vdd
*.iopin vss
*.ipin vin_n
*.ipin vin_p
*.ipin iref
*.opin vout
XM1 vbn vin_n vp vp sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 voe1 vin_p vp vp sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vbn vbn vss vss sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 voe1 vbn vss vss sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 vp iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.75 W=5 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 vout iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.6 W=16 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 iref iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.75 W=5 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net1 vdd voe1 vss sky130_fd_pr__nfet_01v8 L=0.6 W=10 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 net1 vout sky130_fd_pr__cap_mim_m3_1 W=28 L=20 MF=1 m=1
XM6 vout voe1 vss vss sky130_fd_pr__nfet_01v8 L=0.6 W=10 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  r2r_parax.sym # of pins=11
** sym_path: /home/anton/projects/tt06-grab-bag/xschem/r2r.sym
.include /home/anton/projects/tt06-grab-bag/mag/r2r.sim.spice
.GLOBAL GND
.end
