magic
tech sky130A
magscale 1 2
timestamp 1713529744
<< metal1 >>
rect 6494 42746 6626 42752
rect 6494 29886 6626 42614
rect 5994 29754 6626 29886
rect 5994 4846 6126 29754
rect 6686 26488 6742 26494
rect 7514 26488 7570 26494
rect 8342 26488 8398 26494
rect 9170 26488 9226 26494
rect 9998 26488 10054 26494
rect 10826 26488 10882 26494
rect 11654 26488 11710 26494
rect 12482 26488 12538 26494
rect 14966 26488 15022 26494
rect 15794 26488 15850 26494
rect 16622 26488 16678 26494
rect 17450 26488 17506 26494
rect 18278 26488 18334 26494
rect 19106 26488 19162 26494
rect 23246 26488 23302 26494
rect 24074 26488 24130 26494
rect 24902 26488 24958 26494
rect 25730 26488 25786 26494
rect 6742 26432 7048 26488
rect 6686 26426 6742 26432
rect 6992 25992 7048 26432
rect 7570 26432 7848 26488
rect 7514 26426 7570 26432
rect 7792 25992 7848 26432
rect 8398 26432 8648 26488
rect 8342 26426 8398 26432
rect 8592 25992 8648 26432
rect 9226 26432 9448 26488
rect 9170 26426 9226 26432
rect 9392 26032 9448 26432
rect 10054 26432 10248 26488
rect 9998 26426 10054 26432
rect 10192 25992 10248 26432
rect 10882 26432 11048 26488
rect 10826 26426 10882 26432
rect 10992 26032 11048 26432
rect 11710 26432 11848 26488
rect 11654 26426 11710 26432
rect 11792 26032 11848 26432
rect 12116 26460 12316 26466
rect 12538 26432 12648 26488
rect 12482 26426 12538 26432
rect 12116 25966 12316 26260
rect 12592 25972 12648 26432
rect 12986 26460 13186 26466
rect 15022 26432 15248 26488
rect 14966 26426 15022 26432
rect 12986 25966 13186 26260
rect 15192 26032 15248 26432
rect 15850 26432 16048 26488
rect 15794 26426 15850 26432
rect 15992 26012 16048 26432
rect 16678 26432 16848 26488
rect 16622 26426 16678 26432
rect 16792 26032 16848 26432
rect 17506 26432 17648 26488
rect 17450 26426 17506 26432
rect 17592 26032 17648 26432
rect 18334 26432 18448 26488
rect 18278 26426 18334 26432
rect 18392 25992 18448 26432
rect 19162 26432 19268 26488
rect 19928 26432 19934 26488
rect 19990 26432 20068 26488
rect 19106 26426 19162 26432
rect 19212 25972 19268 26432
rect 20012 25992 20068 26432
rect 20316 26480 20516 26486
rect 20756 26432 20762 26488
rect 20818 26432 20824 26488
rect 21186 26480 21386 26486
rect 20316 25966 20516 26280
rect 20762 25992 20818 26432
rect 23302 26432 23448 26488
rect 23246 26426 23302 26432
rect 21186 25966 21386 26280
rect 23392 26052 23448 26432
rect 24130 26432 24248 26488
rect 24074 26426 24130 26432
rect 24192 26032 24248 26432
rect 24958 26432 25048 26488
rect 24902 26426 24958 26432
rect 24992 26012 25048 26432
rect 25786 26432 25900 26488
rect 26552 26432 26558 26488
rect 26614 26432 26620 26488
rect 27380 26432 27386 26488
rect 27442 26432 27448 26488
rect 28208 26432 28214 26488
rect 28270 26432 28276 26488
rect 28516 26480 28716 26486
rect 25730 26426 25786 26432
rect 25844 26052 25900 26432
rect 26558 26032 26614 26432
rect 27386 26032 27442 26432
rect 28214 25992 28270 26432
rect 28516 25966 28716 26280
rect 28976 26440 29042 26496
rect 29098 26440 29104 26496
rect 29386 26480 29586 26486
rect 28976 25970 29032 26440
rect 29386 25960 29586 26280
rect 6414 16293 6826 16466
rect 14472 16311 15088 16488
rect 6414 10506 6587 16293
rect 14472 10508 14649 16311
rect 22666 16306 23294 16494
rect 22666 10514 22854 16306
rect 28706 10514 28894 10520
rect 6414 10333 13147 10506
rect 12974 10086 13147 10333
rect 14472 10331 21409 10508
rect 12974 9913 20907 10086
rect 20734 9626 20907 9913
rect 21232 10068 21409 10331
rect 22666 10326 28706 10514
rect 28706 10320 28894 10326
rect 25332 10068 25509 10074
rect 21232 9891 25332 10068
rect 25332 9885 25509 9891
rect 24574 9626 24747 9632
rect 20734 9453 24574 9626
rect 24574 9447 24747 9453
rect 5994 4714 6866 4846
rect 4854 4400 4860 4600
rect 5060 4400 6610 4600
rect 6410 4223 6610 4400
rect 4554 3123 4560 3323
rect 4760 3123 5180 3323
rect 6734 3239 6866 4714
rect 6444 3107 6866 3239
rect 6754 2740 6760 2940
rect 6960 2740 6966 2940
rect 6760 2540 6960 2740
rect 6400 2340 7320 2540
rect 7120 1800 7320 2340
rect 7114 1600 7120 1800
rect 7320 1600 7326 1800
<< via1 >>
rect 6494 42614 6626 42746
rect 6686 26432 6742 26488
rect 7514 26432 7570 26488
rect 8342 26432 8398 26488
rect 9170 26432 9226 26488
rect 9998 26432 10054 26488
rect 10826 26432 10882 26488
rect 11654 26432 11710 26488
rect 12116 26260 12316 26460
rect 12482 26432 12538 26488
rect 12986 26260 13186 26460
rect 14966 26432 15022 26488
rect 15794 26432 15850 26488
rect 16622 26432 16678 26488
rect 17450 26432 17506 26488
rect 18278 26432 18334 26488
rect 19106 26432 19162 26488
rect 19934 26432 19990 26488
rect 20316 26280 20516 26480
rect 20762 26432 20818 26488
rect 21186 26280 21386 26480
rect 23246 26432 23302 26488
rect 24074 26432 24130 26488
rect 24902 26432 24958 26488
rect 25730 26432 25786 26488
rect 26558 26432 26614 26488
rect 27386 26432 27442 26488
rect 28214 26432 28270 26488
rect 28516 26280 28716 26480
rect 29042 26440 29098 26496
rect 29386 26280 29586 26480
rect 28706 10326 28894 10514
rect 25332 9891 25509 10068
rect 24574 9453 24747 9626
rect 4860 4400 5060 4600
rect 4560 3123 4760 3323
rect 6760 2740 6960 2940
rect 7120 1600 7320 1800
<< metal2 >>
rect 10366 44488 10426 44490
rect 10359 44432 10368 44488
rect 10424 44432 10433 44488
rect 11102 44464 11162 44466
rect 11838 44464 11898 44466
rect 12574 44464 12634 44466
rect 13310 44464 13370 44466
rect 14046 44464 14106 44466
rect 14782 44464 14842 44466
rect 15518 44464 15578 44466
rect 16254 44464 16314 44466
rect 16990 44464 17050 44466
rect 17726 44464 17786 44466
rect 10366 44274 10426 44432
rect 11095 44408 11104 44464
rect 11160 44408 11169 44464
rect 11831 44408 11840 44464
rect 11896 44408 11905 44464
rect 12567 44408 12576 44464
rect 12632 44408 12641 44464
rect 13303 44408 13312 44464
rect 13368 44408 13377 44464
rect 14039 44408 14048 44464
rect 14104 44408 14113 44464
rect 14775 44408 14784 44464
rect 14840 44408 14849 44464
rect 15511 44408 15520 44464
rect 15576 44408 15585 44464
rect 16247 44408 16256 44464
rect 16312 44408 16321 44464
rect 16983 44408 16992 44464
rect 17048 44408 17057 44464
rect 17719 44408 17728 44464
rect 17784 44408 17793 44464
rect 10366 43214 10434 44274
rect 11102 43388 11162 44408
rect 11838 43388 11898 44408
rect 12574 43388 12634 44408
rect 13310 43388 13370 44408
rect 14046 43388 14106 44408
rect 14782 43388 14842 44408
rect 15518 43388 15578 44408
rect 16254 43388 16314 44408
rect 16990 43388 17050 44408
rect 17726 43388 17786 44408
rect 24350 44264 24410 44266
rect 25086 44264 25146 44266
rect 25822 44264 25882 44266
rect 26558 44264 26618 44266
rect 27294 44264 27354 44266
rect 28030 44264 28090 44266
rect 28766 44264 28826 44266
rect 29502 44264 29562 44266
rect 24343 44208 24352 44264
rect 24408 44208 24417 44264
rect 25079 44208 25088 44264
rect 25144 44208 25153 44264
rect 25815 44208 25824 44264
rect 25880 44208 25889 44264
rect 26551 44208 26560 44264
rect 26616 44208 26625 44264
rect 27287 44208 27296 44264
rect 27352 44208 27361 44264
rect 28023 44208 28032 44264
rect 28088 44208 28097 44264
rect 28759 44208 28768 44264
rect 28824 44208 28833 44264
rect 29495 44208 29504 44264
rect 29560 44208 29569 44264
rect 24350 43388 24410 44208
rect 25086 43388 25146 44208
rect 25822 43388 25882 44208
rect 26558 43388 26618 44208
rect 27294 43388 27354 44208
rect 28030 43388 28090 44208
rect 28766 43388 28826 44208
rect 29502 43388 29562 44208
rect 6786 43146 10434 43214
rect 6494 43026 6626 43035
rect 6494 42746 6626 42894
rect 6488 42614 6494 42746
rect 6626 42614 6632 42746
rect 6786 29540 6854 43146
rect 6280 29340 6920 29540
rect 6280 17120 6480 29340
rect 6686 26488 6742 27794
rect 7514 26488 7570 27794
rect 8342 26488 8398 27794
rect 9170 26488 9226 27794
rect 9998 26488 10054 27808
rect 10826 26488 10882 27794
rect 11654 26488 11710 27794
rect 12116 26880 12316 26889
rect 6680 26432 6686 26488
rect 6742 26432 6748 26488
rect 7508 26432 7514 26488
rect 7570 26432 7576 26488
rect 8336 26432 8342 26488
rect 8398 26432 8404 26488
rect 9164 26432 9170 26488
rect 9226 26432 9232 26488
rect 9992 26432 9998 26488
rect 10054 26432 10060 26488
rect 10820 26432 10826 26488
rect 10882 26432 10888 26488
rect 11648 26432 11654 26488
rect 11710 26432 11716 26488
rect 12116 26460 12316 26680
rect 12482 26488 12538 27794
rect 12986 26880 13186 26889
rect 12110 26260 12116 26460
rect 12316 26260 12322 26460
rect 12476 26432 12482 26488
rect 12538 26432 12544 26488
rect 12986 26460 13186 26680
rect 14966 26488 15022 27794
rect 15794 26488 15850 27794
rect 16622 26488 16678 27794
rect 17450 26488 17506 27794
rect 18278 26488 18334 27794
rect 19106 26488 19162 27794
rect 19934 26488 19990 27794
rect 12980 26260 12986 26460
rect 13186 26260 13192 26460
rect 14960 26432 14966 26488
rect 15022 26432 15028 26488
rect 15788 26432 15794 26488
rect 15850 26432 15856 26488
rect 16616 26432 16622 26488
rect 16678 26432 16684 26488
rect 17444 26432 17450 26488
rect 17506 26432 17512 26488
rect 18272 26432 18278 26488
rect 18334 26432 18340 26488
rect 19100 26432 19106 26488
rect 19162 26432 19168 26488
rect 20316 26880 20516 26889
rect 20316 26480 20516 26680
rect 20762 26488 20818 27794
rect 19934 26426 19990 26432
rect 20310 26280 20316 26480
rect 20516 26280 20522 26480
rect 21186 26880 21386 26889
rect 21186 26480 21386 26680
rect 23246 26488 23302 27794
rect 24074 26488 24130 27794
rect 24902 26488 24958 27794
rect 25730 26488 25786 27794
rect 26558 26488 26614 27794
rect 20762 26426 20818 26432
rect 21180 26280 21186 26480
rect 21386 26280 21392 26480
rect 23240 26432 23246 26488
rect 23302 26432 23308 26488
rect 24068 26432 24074 26488
rect 24130 26432 24136 26488
rect 24896 26432 24902 26488
rect 24958 26432 24964 26488
rect 25724 26432 25730 26488
rect 25786 26432 25792 26488
rect 26558 26426 26614 26432
rect 27386 26488 27442 27794
rect 27386 26426 27442 26432
rect 28214 26488 28270 27794
rect 28516 26880 28716 26889
rect 28516 26480 28716 26680
rect 29042 26496 29098 27794
rect 28214 26426 28270 26432
rect 28510 26280 28516 26480
rect 28716 26280 28722 26480
rect 29386 26880 29586 26889
rect 29386 26480 29586 26680
rect 29042 26434 29098 26440
rect 29380 26280 29386 26480
rect 29586 26280 29592 26480
rect 6040 16920 6480 17120
rect 6040 5000 6240 16920
rect 29391 10514 29569 10518
rect 28700 10326 28706 10514
rect 28894 10509 29574 10514
rect 28894 10331 29391 10509
rect 29569 10331 29574 10509
rect 28894 10326 29574 10331
rect 29391 10322 29569 10326
rect 26057 10068 26224 10072
rect 25326 9891 25332 10068
rect 25509 10063 26229 10068
rect 25509 9896 26057 10063
rect 26224 9896 26229 10063
rect 25509 9891 26229 9896
rect 26057 9887 26224 9891
rect 25319 9626 25482 9630
rect 24568 9453 24574 9626
rect 24747 9621 25487 9626
rect 24747 9458 25319 9621
rect 25482 9458 25487 9621
rect 24747 9453 25487 9458
rect 25319 9449 25482 9453
rect 6040 4800 6960 5000
rect 4860 4600 5060 4606
rect 4091 4400 4100 4600
rect 4300 4400 4860 4600
rect 4860 4394 5060 4400
rect 4560 3323 4760 3329
rect 4091 3123 4100 3323
rect 4300 3123 4560 3323
rect 4560 3117 4760 3123
rect 6760 2940 6960 4800
rect 6760 2734 6960 2740
rect 7120 1800 7320 1806
rect 7120 1535 7320 1600
rect 7116 1345 7125 1535
rect 7315 1345 7324 1535
rect 7120 1340 7320 1345
<< via2 >>
rect 10368 44432 10424 44488
rect 11104 44408 11160 44464
rect 11840 44408 11896 44464
rect 12576 44408 12632 44464
rect 13312 44408 13368 44464
rect 14048 44408 14104 44464
rect 14784 44408 14840 44464
rect 15520 44408 15576 44464
rect 16256 44408 16312 44464
rect 16992 44408 17048 44464
rect 17728 44408 17784 44464
rect 24352 44208 24408 44264
rect 25088 44208 25144 44264
rect 25824 44208 25880 44264
rect 26560 44208 26616 44264
rect 27296 44208 27352 44264
rect 28032 44208 28088 44264
rect 28768 44208 28824 44264
rect 29504 44208 29560 44264
rect 6494 42894 6626 43026
rect 12116 26680 12316 26880
rect 12986 26680 13186 26880
rect 20316 26680 20516 26880
rect 21186 26680 21386 26880
rect 28516 26680 28716 26880
rect 29386 26680 29586 26880
rect 29391 10331 29569 10509
rect 26057 9896 26224 10063
rect 25319 9458 25482 9621
rect 4100 4400 4300 4600
rect 4100 3123 4300 3323
rect 7125 1345 7315 1535
<< metal3 >>
rect 6494 44781 6626 44806
rect 18432 44789 18528 44795
rect 6494 44700 18432 44781
rect 6270 44459 6370 44460
rect 6265 44361 6271 44459
rect 6369 44361 6375 44459
rect 6270 44210 6370 44361
rect 4124 44110 4130 44210
rect 4230 44110 6370 44210
rect 1861 43680 1939 43685
rect 1860 43679 2520 43680
rect 1860 43601 1861 43679
rect 1939 43601 2520 43679
rect 1860 43600 2520 43601
rect 2600 43600 2606 43680
rect 1861 43595 1939 43600
rect 6494 43031 6626 44700
rect 18432 44687 18528 44693
rect 10358 44568 10364 44632
rect 10428 44568 10434 44632
rect 10366 44493 10426 44568
rect 11094 44554 11100 44618
rect 11164 44554 11170 44618
rect 11830 44554 11836 44618
rect 11900 44554 11906 44618
rect 12566 44554 12572 44618
rect 12636 44554 12642 44618
rect 13302 44554 13308 44618
rect 13372 44554 13378 44618
rect 14038 44554 14044 44618
rect 14108 44554 14114 44618
rect 14774 44554 14780 44618
rect 14844 44554 14850 44618
rect 15510 44554 15516 44618
rect 15580 44554 15586 44618
rect 16246 44554 16252 44618
rect 16316 44554 16322 44618
rect 16982 44554 16988 44618
rect 17052 44554 17058 44618
rect 17718 44554 17724 44618
rect 17788 44554 17794 44618
rect 24342 44554 24348 44618
rect 24412 44554 24418 44618
rect 25078 44554 25084 44618
rect 25148 44554 25154 44618
rect 25814 44554 25820 44618
rect 25884 44554 25890 44618
rect 26550 44554 26556 44618
rect 26620 44554 26626 44618
rect 27286 44554 27292 44618
rect 27356 44554 27362 44618
rect 28022 44554 28028 44618
rect 28092 44554 28098 44618
rect 28758 44554 28764 44618
rect 28828 44554 28834 44618
rect 29494 44554 29500 44618
rect 29564 44554 29570 44618
rect 10363 44488 10429 44493
rect 10363 44432 10368 44488
rect 10424 44432 10429 44488
rect 11102 44469 11162 44554
rect 11838 44469 11898 44554
rect 12574 44469 12634 44554
rect 13310 44469 13370 44554
rect 14046 44469 14106 44554
rect 14782 44469 14842 44554
rect 15518 44469 15578 44554
rect 16254 44469 16314 44554
rect 16990 44469 17050 44554
rect 17726 44469 17786 44554
rect 10363 44427 10429 44432
rect 11099 44464 11165 44469
rect 11099 44408 11104 44464
rect 11160 44408 11165 44464
rect 11099 44403 11165 44408
rect 11835 44464 11901 44469
rect 11835 44408 11840 44464
rect 11896 44408 11901 44464
rect 11835 44403 11901 44408
rect 12571 44464 12637 44469
rect 12571 44408 12576 44464
rect 12632 44408 12637 44464
rect 12571 44403 12637 44408
rect 13307 44464 13373 44469
rect 13307 44408 13312 44464
rect 13368 44408 13373 44464
rect 13307 44403 13373 44408
rect 14043 44464 14109 44469
rect 14043 44408 14048 44464
rect 14104 44408 14109 44464
rect 14043 44403 14109 44408
rect 14779 44464 14845 44469
rect 14779 44408 14784 44464
rect 14840 44408 14845 44464
rect 14779 44403 14845 44408
rect 15515 44464 15581 44469
rect 15515 44408 15520 44464
rect 15576 44408 15581 44464
rect 15515 44403 15581 44408
rect 16251 44464 16317 44469
rect 16251 44408 16256 44464
rect 16312 44408 16317 44464
rect 16251 44403 16317 44408
rect 16987 44464 17053 44469
rect 16987 44408 16992 44464
rect 17048 44408 17053 44464
rect 16987 44403 17053 44408
rect 17723 44464 17789 44469
rect 17723 44408 17728 44464
rect 17784 44408 17789 44464
rect 17723 44403 17789 44408
rect 11102 44320 11162 44403
rect 11838 44320 11898 44403
rect 12574 44320 12634 44403
rect 13310 44320 13370 44403
rect 14046 44320 14106 44403
rect 14782 44320 14842 44403
rect 15518 44320 15578 44403
rect 16254 44320 16314 44403
rect 16990 44320 17050 44403
rect 17726 44320 17786 44403
rect 24350 44269 24410 44554
rect 25086 44269 25146 44554
rect 25822 44269 25882 44554
rect 26558 44269 26618 44554
rect 27294 44269 27354 44554
rect 28030 44269 28090 44554
rect 28766 44269 28826 44554
rect 29502 44269 29562 44554
rect 24347 44264 24413 44269
rect 24347 44208 24352 44264
rect 24408 44208 24413 44264
rect 24347 44203 24413 44208
rect 25083 44264 25149 44269
rect 25083 44208 25088 44264
rect 25144 44208 25149 44264
rect 25083 44203 25149 44208
rect 25819 44264 25885 44269
rect 25819 44208 25824 44264
rect 25880 44208 25885 44264
rect 25819 44203 25885 44208
rect 26555 44264 26621 44269
rect 26555 44208 26560 44264
rect 26616 44208 26621 44264
rect 26555 44203 26621 44208
rect 27291 44264 27357 44269
rect 27291 44208 27296 44264
rect 27352 44208 27357 44264
rect 27291 44203 27357 44208
rect 28027 44264 28093 44269
rect 28027 44208 28032 44264
rect 28088 44208 28093 44264
rect 28027 44203 28093 44208
rect 28763 44264 28829 44269
rect 28763 44208 28768 44264
rect 28824 44208 28829 44264
rect 28763 44203 28829 44208
rect 29499 44264 29565 44269
rect 29499 44208 29504 44264
rect 29560 44208 29565 44264
rect 29499 44203 29565 44208
rect 19188 44141 19268 44146
rect 19039 44140 19269 44141
rect 19039 44060 19188 44140
rect 19268 44060 19269 44140
rect 19039 44059 19269 44060
rect 19188 44054 19268 44059
rect 19925 43981 20004 43986
rect 19040 43980 20005 43981
rect 19040 43901 19925 43980
rect 20004 43901 20005 43980
rect 19040 43900 20005 43901
rect 19925 43895 20004 43900
rect 20662 43820 20739 43825
rect 19041 43819 20740 43820
rect 19041 43742 20662 43819
rect 20739 43742 20740 43819
rect 19041 43741 20740 43742
rect 20662 43736 20739 43741
rect 21397 43660 21475 43665
rect 19040 43659 21476 43660
rect 19040 43581 21397 43659
rect 21475 43581 21476 43659
rect 19040 43580 21476 43581
rect 21397 43575 21475 43580
rect 6489 43026 6631 43031
rect 6489 42894 6494 43026
rect 6626 42894 6631 43026
rect 6489 42889 6631 42894
rect 30964 42339 31044 42340
rect 30959 42261 30965 42339
rect 31043 42261 31049 42339
rect 30964 41722 31044 42261
rect 30304 41642 31044 41722
rect 30804 41201 30876 41202
rect 30799 41131 30805 41201
rect 30875 41131 30881 41201
rect 30804 40620 30876 41131
rect 30294 40548 30876 40620
rect 2531 26930 2829 26935
rect 2530 26929 29970 26930
rect 2530 26631 2531 26929
rect 2829 26880 29970 26929
rect 2829 26680 12116 26880
rect 12316 26680 12986 26880
rect 13186 26680 20316 26880
rect 20516 26680 21186 26880
rect 21386 26680 28516 26880
rect 28716 26680 29386 26880
rect 29586 26680 29970 26880
rect 2829 26631 29970 26680
rect 2530 26630 29970 26631
rect 2531 26625 2829 26630
rect 31279 10514 31465 10519
rect 29386 10513 31466 10514
rect 29386 10509 31279 10513
rect 29386 10331 29391 10509
rect 29569 10331 31279 10509
rect 29386 10327 31279 10331
rect 31465 10327 31466 10513
rect 29386 10326 31466 10327
rect 31279 10321 31465 10326
rect 26869 10068 27044 10073
rect 26052 10067 27045 10068
rect 26052 10063 26869 10067
rect 26052 9896 26057 10063
rect 26224 9896 26869 10063
rect 26052 9892 26869 9896
rect 27044 9892 27045 10067
rect 26052 9891 27045 9892
rect 26869 9886 27044 9891
rect 26134 9626 26305 9631
rect 25314 9625 26306 9626
rect 25314 9621 26134 9625
rect 25314 9458 25319 9621
rect 25482 9458 26134 9621
rect 25314 9454 26134 9458
rect 26305 9454 26306 9625
rect 25314 9453 26306 9454
rect 26134 9448 26305 9453
rect 4095 4600 4305 4605
rect 3414 4400 3420 4600
rect 3620 4400 4100 4600
rect 4300 4400 4305 4600
rect 4095 4395 4305 4400
rect 4095 3323 4305 3328
rect 1174 3123 1180 3323
rect 1380 3123 4100 3323
rect 4300 3123 4305 3323
rect 4095 3118 4305 3123
rect 7120 1535 7320 1540
rect 7120 1345 7125 1535
rect 7315 1345 7320 1535
rect 7120 1340 7320 1345
rect 7120 1134 7320 1140
<< via3 >>
rect 6271 44361 6369 44459
rect 4130 44110 4230 44210
rect 1861 43601 1939 43679
rect 2520 43600 2600 43680
rect 18432 44693 18528 44789
rect 10364 44568 10428 44632
rect 11100 44554 11164 44618
rect 11836 44554 11900 44618
rect 12572 44554 12636 44618
rect 13308 44554 13372 44618
rect 14044 44554 14108 44618
rect 14780 44554 14844 44618
rect 15516 44554 15580 44618
rect 16252 44554 16316 44618
rect 16988 44554 17052 44618
rect 17724 44554 17788 44618
rect 24348 44554 24412 44618
rect 25084 44554 25148 44618
rect 25820 44554 25884 44618
rect 26556 44554 26620 44618
rect 27292 44554 27356 44618
rect 28028 44554 28092 44618
rect 28764 44554 28828 44618
rect 29500 44554 29564 44618
rect 19188 44060 19268 44140
rect 19925 43901 20004 43980
rect 20662 43742 20739 43819
rect 21397 43581 21475 43659
rect 30965 42261 31043 42339
rect 30805 41131 30875 41201
rect 2531 26631 2829 26929
rect 31279 10327 31465 10513
rect 26869 9892 27044 10067
rect 26134 9454 26305 9625
rect 3420 4400 3620 4600
rect 1180 3123 1380 3323
rect 7120 1140 7320 1340
<< metal4 >>
rect 200 44080 500 44152
rect 798 44080 858 45152
rect 1534 44460 1594 45152
rect 2270 44460 2330 45152
rect 3006 44460 3066 45152
rect 3742 44460 3802 45152
rect 4478 44460 4538 45152
rect 5214 44460 5274 45152
rect 5950 44460 6010 45152
rect 6686 44460 6746 45152
rect 7422 44460 7482 45152
rect 8158 44460 8218 45152
rect 8894 44460 8954 45152
rect 9630 44460 9690 45152
rect 10366 44633 10426 45152
rect 10363 44632 10429 44633
rect 10363 44568 10364 44632
rect 10428 44568 10429 44632
rect 11102 44619 11162 45152
rect 11838 44619 11898 45152
rect 12574 44619 12634 45152
rect 13310 44619 13370 45152
rect 14046 44619 14106 45152
rect 14782 44619 14842 45152
rect 15518 44619 15578 45152
rect 16254 44619 16314 45152
rect 16990 44619 17050 45152
rect 17726 44619 17786 45152
rect 18462 44908 18522 45152
rect 18432 44790 18528 44908
rect 18431 44789 18529 44790
rect 18431 44693 18432 44789
rect 18528 44693 18529 44789
rect 18431 44692 18529 44693
rect 10363 44567 10429 44568
rect 11099 44618 11165 44619
rect 11099 44554 11100 44618
rect 11164 44554 11165 44618
rect 11099 44553 11165 44554
rect 11835 44618 11901 44619
rect 11835 44554 11836 44618
rect 11900 44554 11901 44618
rect 11835 44553 11901 44554
rect 12571 44618 12637 44619
rect 12571 44554 12572 44618
rect 12636 44554 12637 44618
rect 12571 44553 12637 44554
rect 13307 44618 13373 44619
rect 13307 44554 13308 44618
rect 13372 44554 13373 44618
rect 13307 44553 13373 44554
rect 14043 44618 14109 44619
rect 14043 44554 14044 44618
rect 14108 44554 14109 44618
rect 14043 44553 14109 44554
rect 14779 44618 14845 44619
rect 14779 44554 14780 44618
rect 14844 44554 14845 44618
rect 14779 44553 14845 44554
rect 15515 44618 15581 44619
rect 15515 44554 15516 44618
rect 15580 44554 15581 44618
rect 15515 44553 15581 44554
rect 16251 44618 16317 44619
rect 16251 44554 16252 44618
rect 16316 44554 16317 44618
rect 16251 44553 16317 44554
rect 16987 44618 17053 44619
rect 16987 44554 16988 44618
rect 17052 44554 17053 44618
rect 16987 44553 17053 44554
rect 17723 44618 17789 44619
rect 17723 44554 17724 44618
rect 17788 44554 17789 44618
rect 17723 44553 17789 44554
rect 11102 44540 11162 44553
rect 11838 44540 11898 44553
rect 12574 44540 12634 44553
rect 13310 44540 13370 44553
rect 14046 44540 14106 44553
rect 14782 44540 14842 44553
rect 15518 44540 15578 44553
rect 16254 44540 16314 44553
rect 16990 44540 17050 44553
rect 1480 44438 3802 44460
rect 1480 44210 3800 44438
rect 4440 44360 6020 44460
rect 6270 44459 9740 44460
rect 6270 44361 6271 44459
rect 6369 44361 9740 44459
rect 6270 44360 9740 44361
rect 4129 44210 4231 44211
rect 1480 44110 4130 44210
rect 4230 44110 4231 44210
rect 200 44000 860 44080
rect 200 43680 500 44000
rect 1480 43920 3800 44110
rect 4129 44109 4231 44110
rect 4440 43920 4600 44360
rect 19198 44141 19258 45152
rect 19187 44140 19269 44141
rect 19187 44060 19188 44140
rect 19268 44060 19269 44140
rect 19187 44059 19269 44060
rect 19198 44040 19258 44059
rect 19934 43981 19994 45152
rect 19924 43980 20005 43981
rect 200 43679 1940 43680
rect 200 43601 1861 43679
rect 1939 43601 1940 43679
rect 200 43600 1940 43601
rect 200 3323 500 43600
rect 2100 26930 2400 43920
rect 2519 43680 2601 43681
rect 4480 43680 4560 43920
rect 19924 43901 19925 43980
rect 20004 43901 20005 43980
rect 19924 43900 20005 43901
rect 19934 43880 19994 43900
rect 20670 43820 20730 45152
rect 20661 43819 20740 43820
rect 20661 43742 20662 43819
rect 20739 43742 20740 43819
rect 20661 43741 20740 43742
rect 20670 43720 20730 43741
rect 2519 43600 2520 43680
rect 2600 43600 4560 43680
rect 21406 43660 21466 45152
rect 22142 44854 22202 45152
rect 22878 44854 22938 45152
rect 23614 44854 23674 45152
rect 24350 44619 24410 45152
rect 25086 44619 25146 45152
rect 25822 44619 25882 45152
rect 26558 44619 26618 45152
rect 27294 44619 27354 45152
rect 28030 44619 28090 45152
rect 28766 44619 28826 45152
rect 29502 44619 29562 45152
rect 24347 44618 24413 44619
rect 24347 44554 24348 44618
rect 24412 44554 24413 44618
rect 24347 44553 24413 44554
rect 25083 44618 25149 44619
rect 25083 44554 25084 44618
rect 25148 44554 25149 44618
rect 25083 44553 25149 44554
rect 25819 44618 25885 44619
rect 25819 44554 25820 44618
rect 25884 44554 25885 44618
rect 25819 44553 25885 44554
rect 26555 44618 26621 44619
rect 26555 44554 26556 44618
rect 26620 44554 26621 44618
rect 26555 44553 26621 44554
rect 27291 44618 27357 44619
rect 27291 44554 27292 44618
rect 27356 44554 27357 44618
rect 27291 44553 27357 44554
rect 28027 44618 28093 44619
rect 28027 44554 28028 44618
rect 28092 44554 28093 44618
rect 28027 44553 28093 44554
rect 28763 44618 28829 44619
rect 28763 44554 28764 44618
rect 28828 44554 28829 44618
rect 28763 44553 28829 44554
rect 29499 44618 29565 44619
rect 29499 44554 29500 44618
rect 29564 44554 29565 44618
rect 29499 44553 29565 44554
rect 30238 44256 30298 45152
rect 30238 44196 30600 44256
rect 21396 43659 21476 43660
rect 2519 43599 2601 43600
rect 21396 43581 21397 43659
rect 21475 43581 21476 43659
rect 21396 43580 21476 43581
rect 21406 43560 21466 43580
rect 30540 42024 30600 44196
rect 30974 42340 31034 45152
rect 31710 44952 31770 45152
rect 30964 42339 31044 42340
rect 30964 42261 30965 42339
rect 31043 42261 31044 42339
rect 30964 42260 31044 42261
rect 30540 41964 30870 42024
rect 30810 41202 30870 41964
rect 30804 41201 30876 41202
rect 30804 41131 30805 41201
rect 30875 41131 30876 41201
rect 30804 41130 30876 41131
rect 2100 26929 2830 26930
rect 2100 26631 2531 26929
rect 2829 26631 2830 26929
rect 2100 26630 2830 26631
rect 2100 4600 2400 26630
rect 31278 10513 31466 10514
rect 31278 10327 31279 10513
rect 31465 10327 31466 10513
rect 26868 10067 27045 10068
rect 26868 9892 26869 10067
rect 27044 9892 27045 10067
rect 26133 9625 26306 9626
rect 26133 9454 26134 9625
rect 26305 9454 26306 9625
rect 3419 4600 3621 4601
rect 2100 4400 3420 4600
rect 3620 4400 3621 4600
rect 1179 3323 1381 3324
rect 200 3123 1180 3323
rect 1380 3123 1381 3323
rect 200 1000 500 3123
rect 1179 3122 1381 3123
rect 2100 1000 2400 4400
rect 3419 4399 3621 4400
rect 7119 1340 7321 1341
rect 7119 1140 7120 1340
rect 7320 1140 7321 1340
rect 7119 1139 7321 1140
rect 7120 760 7320 1139
rect 26133 827 26306 9454
rect 7120 560 9380 760
rect 22454 654 26306 827
rect 26868 772 27045 9892
rect 31278 846 31466 10327
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 560
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 654
rect 26896 0 27016 772
rect 31312 0 31432 846
use controller  controller_0
timestamp 1713497815
transform 1 0 6668 0 1 27738
box 14 0 24000 16000
use inverter  inverter_0
timestamp 1712241802
transform 1 0 5390 0 1 1613
box -410 547 1220 2810
use r2r  r2r_blue
timestamp 1713380768
transform 0 1 12386 -1 0 25766
box -400 -5786 14766 800
use r2r  r2r_green
timestamp 1713380768
transform 0 1 20586 -1 0 25766
box -400 -5786 14766 800
use r2r  r2r_red
timestamp 1713380768
transform 0 1 28786 -1 0 25766
box -400 -5786 14766 800
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 2100 1000 2400 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
