magic
tech sky130A
magscale 1 2
timestamp 1713392524
<< metal1 >>
rect 29432 44410 29632 44420
rect 29432 44350 29502 44410
rect 29562 44350 29632 44410
rect 17660 43260 17860 43266
rect 17660 42060 17860 43060
rect 17660 41860 28980 42060
rect 29180 41860 29186 42060
rect 10894 41380 10900 41580
rect 11100 41380 24766 41580
rect 18496 41268 18696 41274
rect 18496 40714 18696 41068
rect 19296 41268 19496 41274
rect 19296 40714 19496 41068
rect 20096 41268 20296 41274
rect 20096 40714 20296 41068
rect 20896 41268 21096 41274
rect 20896 40714 21096 41068
rect 21696 41268 21896 41274
rect 21696 40714 21896 41068
rect 22496 41268 22696 41274
rect 22496 40714 22696 41068
rect 23296 41268 23496 41274
rect 23296 40714 23496 41068
rect 23696 40714 23896 41380
rect 24096 41268 24296 41274
rect 24096 40714 24296 41068
rect 24566 40714 24766 41380
rect 17340 31054 18380 31254
rect 17340 25060 17540 31054
rect 17340 24860 27020 25060
rect 26820 7980 27020 24860
rect 26820 7774 27020 7780
rect 29432 7686 29632 44350
rect 29860 42060 30060 42066
rect 30060 41860 31060 42060
rect 29860 41854 30060 41860
rect 29432 7486 30410 7686
rect 29432 7480 29632 7486
rect 11598 7037 11604 7237
rect 11804 7037 30116 7237
rect 2102 5937 2108 6137
rect 2308 5937 28688 6137
rect 30204 6090 30404 7486
rect 29920 5892 30404 6090
rect 29916 3982 30116 5357
rect 30860 4040 31060 41860
rect 30800 3982 31060 4040
rect 29916 3782 31060 3982
rect 29916 2070 30116 3782
rect 30580 3780 31060 3782
rect 31270 2070 31470 2076
rect 29916 1870 31270 2070
rect 31270 1864 31470 1870
<< via1 >>
rect 29502 44350 29562 44410
rect 17660 43060 17860 43260
rect 28980 41860 29180 42060
rect 10900 41380 11100 41580
rect 18496 41068 18696 41268
rect 19296 41068 19496 41268
rect 20096 41068 20296 41268
rect 20896 41068 21096 41268
rect 21696 41068 21896 41268
rect 22496 41068 22696 41268
rect 23296 41068 23496 41268
rect 24096 41068 24296 41268
rect 26820 7780 27020 7980
rect 29860 41860 30060 42060
rect 11604 7037 11804 7237
rect 2108 5937 2308 6137
rect 31270 1870 31470 2070
<< metal2 >>
rect 29502 44590 29562 44592
rect 29495 44534 29504 44590
rect 29560 44534 29569 44590
rect 29502 44410 29562 44534
rect 29502 44344 29562 44350
rect 17660 43700 17860 43709
rect 17660 43260 17860 43500
rect 17654 43060 17660 43260
rect 17860 43060 17866 43260
rect 18496 42380 18696 42389
rect 10900 41580 11100 41586
rect 10611 41380 10620 41580
rect 10820 41380 10900 41580
rect 10900 41374 11100 41380
rect 18496 41268 18696 42180
rect 19296 42380 19496 42389
rect 19296 41268 19496 42180
rect 20096 42380 20296 42389
rect 20096 41268 20296 42180
rect 20896 42380 21096 42389
rect 20896 41268 21096 42180
rect 21696 42380 21896 42389
rect 21696 41268 21896 42180
rect 22496 42380 22696 42389
rect 22496 41268 22696 42180
rect 23296 42380 23496 42389
rect 23296 41268 23496 42180
rect 24096 42380 24296 42389
rect 24096 41268 24296 42180
rect 28980 42060 29180 42066
rect 29180 41860 29860 42060
rect 30060 41860 30066 42060
rect 28980 41854 29180 41860
rect 18490 41068 18496 41268
rect 18696 41068 18702 41268
rect 19290 41068 19296 41268
rect 19496 41068 19502 41268
rect 20090 41068 20096 41268
rect 20296 41068 20302 41268
rect 20890 41068 20896 41268
rect 21096 41068 21102 41268
rect 21690 41068 21696 41268
rect 21896 41068 21902 41268
rect 22490 41068 22496 41268
rect 22696 41068 22702 41268
rect 23290 41068 23296 41268
rect 23496 41068 23502 41268
rect 24090 41068 24096 41268
rect 24296 41068 24302 41268
rect 26814 7780 26820 7980
rect 27020 7780 27026 7980
rect 11604 7237 11804 7243
rect 11147 7037 11156 7237
rect 11356 7037 11604 7237
rect 11604 7031 11804 7037
rect 2108 6137 2308 6143
rect 1611 5937 1620 6137
rect 1820 5937 2108 6137
rect 2108 5931 2308 5937
rect 26820 1620 27020 7780
rect 31264 1870 31270 2070
rect 31470 1870 31476 2070
rect 31270 1660 31470 1870
rect 31270 1451 31470 1460
rect 26820 1411 27020 1420
<< via2 >>
rect 29504 44534 29560 44590
rect 17660 43500 17860 43700
rect 18496 42180 18696 42380
rect 10620 41380 10820 41580
rect 19296 42180 19496 42380
rect 20096 42180 20296 42380
rect 20896 42180 21096 42380
rect 21696 42180 21896 42380
rect 22496 42180 22696 42380
rect 23296 42180 23496 42380
rect 24096 42180 24296 42380
rect 11156 7037 11356 7237
rect 1620 5937 1820 6137
rect 26820 1420 27020 1620
rect 31270 1460 31470 1660
<< metal3 >>
rect 29494 44752 29500 44816
rect 29564 44752 29570 44816
rect 29502 44595 29562 44752
rect 29499 44590 29565 44595
rect 29499 44534 29504 44590
rect 29560 44534 29565 44590
rect 29499 44529 29565 44534
rect 17660 44090 17860 44096
rect 17660 43705 17860 43890
rect 17655 43700 17865 43705
rect 17655 43500 17660 43700
rect 17860 43500 17865 43700
rect 17655 43495 17865 43500
rect 18496 42860 18696 42866
rect 18496 42385 18696 42660
rect 19296 42860 19496 42866
rect 19296 42385 19496 42660
rect 20096 42860 20296 42866
rect 20096 42385 20296 42660
rect 20896 42860 21096 42866
rect 20896 42385 21096 42660
rect 21696 42860 21896 42866
rect 21696 42385 21896 42660
rect 22496 42860 22696 42866
rect 22496 42385 22696 42660
rect 23296 42860 23496 42866
rect 23296 42385 23496 42660
rect 24096 42860 24296 42866
rect 24096 42385 24296 42660
rect 18491 42380 18701 42385
rect 18491 42180 18496 42380
rect 18696 42180 18701 42380
rect 18491 42175 18701 42180
rect 19291 42380 19501 42385
rect 19291 42180 19296 42380
rect 19496 42180 19501 42380
rect 19291 42175 19501 42180
rect 20091 42380 20301 42385
rect 20091 42180 20096 42380
rect 20296 42180 20301 42380
rect 20091 42175 20301 42180
rect 20891 42380 21101 42385
rect 20891 42180 20896 42380
rect 21096 42180 21101 42380
rect 20891 42175 21101 42180
rect 21691 42380 21901 42385
rect 21691 42180 21696 42380
rect 21896 42180 21901 42380
rect 21691 42175 21901 42180
rect 22491 42380 22701 42385
rect 22491 42180 22496 42380
rect 22696 42180 22701 42380
rect 22491 42175 22701 42180
rect 23291 42380 23501 42385
rect 23291 42180 23296 42380
rect 23496 42180 23501 42380
rect 23291 42175 23501 42180
rect 24091 42380 24301 42385
rect 24091 42180 24096 42380
rect 24296 42180 24301 42380
rect 24091 42175 24301 42180
rect 10615 41580 10825 41585
rect 10374 41380 10380 41580
rect 10580 41380 10620 41580
rect 10820 41380 10825 41580
rect 10615 41375 10825 41380
rect 11151 7237 11361 7242
rect 10664 7037 10670 7237
rect 10870 7037 11156 7237
rect 11356 7037 11361 7237
rect 11151 7032 11361 7037
rect 1615 6137 1825 6142
rect 1078 5937 1084 6137
rect 1284 5937 1620 6137
rect 1820 5937 1825 6137
rect 1615 5932 1825 5937
rect 31265 1660 31475 1665
rect 26815 1620 27025 1625
rect 26815 1420 26820 1620
rect 27020 1420 27025 1620
rect 31265 1460 31270 1660
rect 31470 1460 31475 1660
rect 31265 1455 31475 1460
rect 26815 1415 27025 1420
rect 26820 1140 27020 1415
rect 31270 1240 31470 1455
rect 31270 1034 31470 1040
rect 26820 934 27020 940
<< via3 >>
rect 29500 44752 29564 44816
rect 17660 43890 17860 44090
rect 18496 42660 18696 42860
rect 19296 42660 19496 42860
rect 20096 42660 20296 42860
rect 20896 42660 21096 42860
rect 21696 42660 21896 42860
rect 22496 42660 22696 42860
rect 23296 42660 23496 42860
rect 24096 42660 24296 42860
rect 10380 41380 10580 41580
rect 10670 7037 10870 7237
rect 1084 5937 1284 6137
rect 26820 940 27020 1140
rect 31270 1040 31470 1240
<< metal4 >>
rect 798 44438 858 45152
rect 1534 44438 1594 45152
rect 2270 44438 2330 45152
rect 3006 44438 3066 45152
rect 3742 44438 3802 45152
rect 4478 44438 4538 45152
rect 5214 44438 5274 45152
rect 5950 44438 6010 45152
rect 6686 44438 6746 45152
rect 7422 44438 7482 45152
rect 8158 44438 8218 45152
rect 8894 44438 8954 45152
rect 9630 44438 9690 45152
rect 10366 44438 10426 45152
rect 11102 44438 11162 45152
rect 11838 44438 11898 45152
rect 12574 44438 12634 45152
rect 13310 44438 13370 45152
rect 14046 44438 14106 45152
rect 14782 44438 14842 45152
rect 15518 44438 15578 45152
rect 16254 44438 16314 45152
rect 16990 44438 17050 45152
rect 17726 44620 17786 45152
rect 200 6137 500 44152
rect 748 43926 17168 44438
rect 17660 44091 17860 44620
rect 18462 44150 18522 45152
rect 19198 44150 19258 45152
rect 19934 44150 19994 45152
rect 20670 44150 20730 45152
rect 21406 44150 21466 45152
rect 22142 44150 22202 45152
rect 22878 44150 22938 45152
rect 23614 44150 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44817 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29499 44816 29565 44817
rect 29499 44752 29500 44816
rect 29564 44752 29565 44816
rect 29499 44751 29565 44752
rect 17659 44090 17861 44091
rect 18462 44090 18630 44150
rect 19198 44090 19430 44150
rect 19934 44090 20230 44150
rect 20670 44090 21030 44150
rect 21406 44090 21830 44150
rect 22142 44090 22630 44150
rect 22878 44090 23430 44150
rect 23614 44090 24230 44150
rect 9800 41580 10100 43926
rect 17659 43890 17660 44090
rect 17860 43890 17861 44090
rect 17659 43889 17861 43890
rect 18570 43380 18630 44090
rect 19370 43380 19430 44090
rect 20170 43380 20230 44090
rect 20970 43380 21030 44090
rect 21770 43380 21830 44090
rect 22570 43380 22630 44090
rect 23370 43380 23430 44090
rect 24170 43380 24230 44090
rect 18496 42861 18696 43380
rect 19296 42861 19496 43380
rect 20096 42861 20296 43380
rect 20896 42861 21096 43380
rect 21696 42861 21896 43380
rect 22496 42861 22696 43380
rect 23296 42861 23496 43380
rect 24096 42861 24296 43380
rect 18495 42860 18697 42861
rect 18495 42660 18496 42860
rect 18696 42660 18697 42860
rect 18495 42659 18697 42660
rect 19295 42860 19497 42861
rect 19295 42660 19296 42860
rect 19496 42660 19497 42860
rect 19295 42659 19497 42660
rect 20095 42860 20297 42861
rect 20095 42660 20096 42860
rect 20296 42660 20297 42860
rect 20095 42659 20297 42660
rect 20895 42860 21097 42861
rect 20895 42660 20896 42860
rect 21096 42660 21097 42860
rect 20895 42659 21097 42660
rect 21695 42860 21897 42861
rect 21695 42660 21696 42860
rect 21896 42660 21897 42860
rect 21695 42659 21897 42660
rect 22495 42860 22697 42861
rect 22495 42660 22496 42860
rect 22696 42660 22697 42860
rect 22495 42659 22697 42660
rect 23295 42860 23497 42861
rect 23295 42660 23296 42860
rect 23496 42660 23497 42860
rect 23295 42659 23497 42660
rect 24095 42860 24297 42861
rect 24095 42660 24096 42860
rect 24296 42660 24297 42860
rect 24095 42659 24297 42660
rect 10379 41580 10581 41581
rect 9800 41380 10380 41580
rect 10580 41380 10581 41580
rect 9800 7237 10100 41380
rect 10379 41379 10581 41380
rect 10669 7237 10871 7238
rect 9800 7037 10670 7237
rect 10870 7037 10871 7237
rect 1083 6137 1285 6138
rect 200 5937 1084 6137
rect 1284 5937 1285 6137
rect 200 1000 500 5937
rect 1083 5936 1285 5937
rect 9800 1000 10100 7037
rect 10669 7036 10871 7037
rect 31269 1240 31471 1241
rect 26819 1140 27021 1141
rect 26819 940 26820 1140
rect 27020 940 27021 1140
rect 31269 1040 31270 1240
rect 31470 1040 31471 1240
rect 31269 1039 31471 1040
rect 26819 939 27021 940
rect 26820 580 27020 939
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 580
rect 31286 496 31455 1039
rect 31312 0 31432 496
use inverter  inverter_0
timestamp 1712241802
transform 1 0 28896 0 1 4427
box -410 547 1220 2810
use r2r  r2r_0
timestamp 1713380768
transform 0 1 23966 -1 0 40514
box -400 -5786 14766 800
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
