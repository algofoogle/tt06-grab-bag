magic
tech sky130A
magscale 1 2
timestamp 1713538698
<< metal1 >>
rect 6494 42738 6626 42752
rect 6494 42622 6502 42738
rect 6618 42622 6626 42738
rect 6494 29886 6626 42622
rect 5994 29754 6626 29886
rect 5994 4846 6126 29754
rect 28976 26494 29104 26496
rect 6686 26488 6742 26494
rect 7514 26488 7570 26494
rect 8342 26488 8398 26494
rect 9170 26488 9226 26494
rect 9998 26488 10054 26494
rect 10826 26488 10882 26494
rect 11654 26488 11710 26494
rect 12482 26488 12538 26494
rect 14966 26488 15022 26494
rect 15794 26488 15850 26494
rect 16622 26488 16678 26494
rect 17450 26488 17506 26494
rect 18278 26488 18334 26494
rect 19106 26488 19162 26494
rect 23246 26488 23302 26494
rect 24074 26488 24130 26494
rect 24902 26488 24958 26494
rect 25730 26488 25786 26494
rect 6686 26486 7048 26488
rect 6686 26434 6688 26486
rect 6740 26434 7048 26486
rect 6686 26432 7048 26434
rect 6686 26426 6742 26432
rect 6992 25992 7048 26432
rect 7514 26486 7848 26488
rect 7514 26434 7516 26486
rect 7568 26434 7848 26486
rect 7514 26432 7848 26434
rect 7514 26426 7570 26432
rect 7792 25992 7848 26432
rect 8342 26486 8648 26488
rect 8342 26434 8344 26486
rect 8396 26434 8648 26486
rect 8342 26432 8648 26434
rect 8342 26426 8398 26432
rect 8592 25992 8648 26432
rect 9170 26486 9448 26488
rect 9170 26434 9172 26486
rect 9224 26434 9448 26486
rect 9170 26432 9448 26434
rect 9170 26426 9226 26432
rect 9392 26032 9448 26432
rect 9998 26486 10248 26488
rect 9998 26434 10000 26486
rect 10052 26434 10248 26486
rect 9998 26432 10248 26434
rect 9998 26426 10054 26432
rect 10192 25992 10248 26432
rect 10826 26486 11048 26488
rect 10826 26434 10828 26486
rect 10880 26434 11048 26486
rect 10826 26432 11048 26434
rect 10826 26426 10882 26432
rect 10992 26032 11048 26432
rect 11654 26486 11848 26488
rect 11654 26434 11656 26486
rect 11708 26434 11848 26486
rect 12482 26486 12648 26488
rect 11654 26432 11848 26434
rect 11654 26426 11710 26432
rect 11792 26032 11848 26432
rect 12116 26450 12316 26466
rect 12116 26270 12126 26450
rect 12306 26270 12316 26450
rect 12482 26434 12484 26486
rect 12536 26434 12648 26486
rect 14966 26486 15248 26488
rect 12482 26432 12648 26434
rect 12482 26426 12538 26432
rect 12116 25966 12316 26270
rect 12592 25972 12648 26432
rect 12986 26450 13186 26466
rect 12986 26270 12996 26450
rect 13176 26270 13186 26450
rect 14966 26434 14968 26486
rect 15020 26434 15248 26486
rect 14966 26432 15248 26434
rect 14966 26426 15022 26432
rect 12986 25966 13186 26270
rect 15192 26032 15248 26432
rect 15794 26486 16048 26488
rect 15794 26434 15796 26486
rect 15848 26434 16048 26486
rect 15794 26432 16048 26434
rect 15794 26426 15850 26432
rect 15992 26012 16048 26432
rect 16622 26486 16848 26488
rect 16622 26434 16624 26486
rect 16676 26434 16848 26486
rect 16622 26432 16848 26434
rect 16622 26426 16678 26432
rect 16792 26032 16848 26432
rect 17450 26486 17648 26488
rect 17450 26434 17452 26486
rect 17504 26434 17648 26486
rect 17450 26432 17648 26434
rect 17450 26426 17506 26432
rect 17592 26032 17648 26432
rect 18278 26486 18448 26488
rect 18278 26434 18280 26486
rect 18332 26434 18448 26486
rect 18278 26432 18448 26434
rect 18278 26426 18334 26432
rect 18392 25992 18448 26432
rect 19106 26486 19268 26488
rect 19106 26434 19108 26486
rect 19160 26434 19268 26486
rect 19106 26432 19268 26434
rect 19928 26486 20068 26488
rect 20756 26486 20824 26488
rect 23246 26486 23448 26488
rect 19928 26434 19936 26486
rect 19988 26434 20068 26486
rect 19928 26432 20068 26434
rect 19106 26426 19162 26432
rect 19212 25972 19268 26432
rect 20012 25992 20068 26432
rect 20316 26470 20516 26486
rect 20316 26290 20326 26470
rect 20506 26290 20516 26470
rect 20756 26434 20764 26486
rect 20816 26434 20824 26486
rect 20756 26432 20824 26434
rect 21186 26470 21386 26486
rect 20316 25966 20516 26290
rect 20762 25992 20818 26432
rect 21186 26290 21196 26470
rect 21376 26290 21386 26470
rect 23246 26434 23248 26486
rect 23300 26434 23448 26486
rect 23246 26432 23448 26434
rect 23246 26426 23302 26432
rect 21186 25966 21386 26290
rect 23392 26052 23448 26432
rect 24074 26486 24248 26488
rect 24074 26434 24076 26486
rect 24128 26434 24248 26486
rect 24074 26432 24248 26434
rect 24074 26426 24130 26432
rect 24192 26032 24248 26432
rect 24902 26486 25048 26488
rect 24902 26434 24904 26486
rect 24956 26434 25048 26486
rect 24902 26432 25048 26434
rect 24902 26426 24958 26432
rect 24992 26012 25048 26432
rect 25730 26486 25900 26488
rect 25730 26434 25732 26486
rect 25784 26434 25900 26486
rect 25730 26432 25900 26434
rect 26552 26486 26620 26488
rect 26552 26434 26560 26486
rect 26612 26434 26620 26486
rect 26552 26432 26620 26434
rect 27380 26486 27448 26488
rect 27380 26434 27388 26486
rect 27440 26434 27448 26486
rect 27380 26432 27448 26434
rect 28208 26486 28276 26488
rect 28208 26434 28216 26486
rect 28268 26434 28276 26486
rect 28208 26432 28276 26434
rect 28516 26470 28716 26486
rect 25730 26426 25786 26432
rect 25844 26052 25900 26432
rect 26558 26032 26614 26432
rect 27386 26032 27442 26432
rect 28214 25992 28270 26432
rect 28516 26290 28526 26470
rect 28706 26290 28716 26470
rect 28516 25966 28716 26290
rect 28976 26442 29044 26494
rect 29096 26442 29104 26494
rect 28976 26440 29104 26442
rect 29386 26470 29586 26486
rect 28976 25970 29032 26440
rect 29386 26290 29396 26470
rect 29576 26290 29586 26470
rect 29386 25960 29586 26290
rect 6414 16293 6826 16466
rect 14472 16311 15088 16488
rect 6414 10506 6587 16293
rect 14472 10508 14649 16311
rect 22666 16306 23294 16494
rect 22666 10514 22854 16306
rect 28706 10514 28894 10520
rect 22666 10510 28894 10514
rect 6414 10333 13147 10506
rect 12974 10086 13147 10333
rect 14472 10331 21409 10508
rect 12974 9913 20907 10086
rect 20734 9626 20907 9913
rect 21232 10068 21409 10331
rect 22666 10330 28710 10510
rect 28890 10330 28894 10510
rect 22666 10326 28894 10330
rect 28706 10320 28894 10326
rect 25332 10068 25509 10074
rect 21232 10037 25509 10068
rect 21232 9921 25362 10037
rect 25478 9921 25509 10037
rect 21232 9891 25509 9921
rect 25332 9885 25509 9891
rect 24574 9626 24747 9632
rect 20734 9597 24747 9626
rect 20734 9481 24602 9597
rect 24718 9481 24747 9597
rect 20734 9453 24747 9481
rect 24574 9447 24747 9453
rect 5994 4714 6866 4846
rect 4854 4590 6610 4600
rect 4854 4410 4870 4590
rect 5050 4410 6610 4590
rect 4854 4400 6610 4410
rect 6410 4223 6610 4400
rect 4554 3313 5180 3323
rect 4554 3133 4570 3313
rect 4750 3133 5180 3313
rect 6734 3239 6866 4714
rect 4554 3123 5180 3133
rect 6444 3107 6866 3239
rect 6754 2930 6966 2940
rect 6754 2750 6770 2930
rect 6950 2750 6966 2930
rect 6754 2740 6966 2750
rect 6760 2540 6960 2740
rect 6400 2340 7320 2540
rect 7120 1800 7320 2340
rect 7114 1790 7326 1800
rect 7114 1610 7130 1790
rect 7310 1610 7326 1790
rect 7114 1600 7326 1610
<< via1 >>
rect 6502 42622 6618 42738
rect 6688 26434 6740 26486
rect 7516 26434 7568 26486
rect 8344 26434 8396 26486
rect 9172 26434 9224 26486
rect 10000 26434 10052 26486
rect 10828 26434 10880 26486
rect 11656 26434 11708 26486
rect 12126 26270 12306 26450
rect 12484 26434 12536 26486
rect 12996 26270 13176 26450
rect 14968 26434 15020 26486
rect 15796 26434 15848 26486
rect 16624 26434 16676 26486
rect 17452 26434 17504 26486
rect 18280 26434 18332 26486
rect 19108 26434 19160 26486
rect 19936 26434 19988 26486
rect 20326 26290 20506 26470
rect 20764 26434 20816 26486
rect 21196 26290 21376 26470
rect 23248 26434 23300 26486
rect 24076 26434 24128 26486
rect 24904 26434 24956 26486
rect 25732 26434 25784 26486
rect 26560 26434 26612 26486
rect 27388 26434 27440 26486
rect 28216 26434 28268 26486
rect 28526 26290 28706 26470
rect 29044 26442 29096 26494
rect 29396 26290 29576 26470
rect 28710 10330 28890 10510
rect 25362 9921 25478 10037
rect 24602 9481 24718 9597
rect 4870 4410 5050 4590
rect 4570 3133 4750 3313
rect 6770 2750 6950 2930
rect 7130 1610 7310 1790
<< metal2 >>
rect 10366 44488 10426 44490
rect 10359 44432 10368 44488
rect 10424 44432 10433 44488
rect 11102 44464 11162 44466
rect 11838 44464 11898 44466
rect 12574 44464 12634 44466
rect 13310 44464 13370 44466
rect 14046 44464 14106 44466
rect 14782 44464 14842 44466
rect 15518 44464 15578 44466
rect 16254 44464 16314 44466
rect 16990 44464 17050 44466
rect 17726 44464 17786 44466
rect 10366 44274 10426 44432
rect 11095 44408 11104 44464
rect 11160 44408 11169 44464
rect 11831 44408 11840 44464
rect 11896 44408 11905 44464
rect 12567 44408 12576 44464
rect 12632 44408 12641 44464
rect 13303 44408 13312 44464
rect 13368 44408 13377 44464
rect 14039 44408 14048 44464
rect 14104 44408 14113 44464
rect 14775 44408 14784 44464
rect 14840 44408 14849 44464
rect 15511 44408 15520 44464
rect 15576 44408 15585 44464
rect 16247 44408 16256 44464
rect 16312 44408 16321 44464
rect 16983 44408 16992 44464
rect 17048 44408 17057 44464
rect 17719 44408 17728 44464
rect 17784 44408 17793 44464
rect 10366 43214 10434 44274
rect 11102 43388 11162 44408
rect 11838 43388 11898 44408
rect 12574 43388 12634 44408
rect 13310 43388 13370 44408
rect 14046 43388 14106 44408
rect 14782 43388 14842 44408
rect 15518 43388 15578 44408
rect 16254 43388 16314 44408
rect 16990 43388 17050 44408
rect 17726 43388 17786 44408
rect 24350 44264 24410 44266
rect 25086 44264 25146 44266
rect 25822 44264 25882 44266
rect 26558 44264 26618 44266
rect 27294 44264 27354 44266
rect 28030 44264 28090 44266
rect 28766 44264 28826 44266
rect 29502 44264 29562 44266
rect 24343 44208 24352 44264
rect 24408 44208 24417 44264
rect 25079 44208 25088 44264
rect 25144 44208 25153 44264
rect 25815 44208 25824 44264
rect 25880 44208 25889 44264
rect 26551 44208 26560 44264
rect 26616 44208 26625 44264
rect 27287 44208 27296 44264
rect 27352 44208 27361 44264
rect 28023 44208 28032 44264
rect 28088 44208 28097 44264
rect 28759 44208 28768 44264
rect 28824 44208 28833 44264
rect 29495 44208 29504 44264
rect 29560 44208 29569 44264
rect 24350 43388 24410 44208
rect 25086 43388 25146 44208
rect 25822 43388 25882 44208
rect 26558 43388 26618 44208
rect 27294 43388 27354 44208
rect 28030 43388 28090 44208
rect 28766 43388 28826 44208
rect 29502 43388 29562 44208
rect 6786 43146 10434 43214
rect 6494 42988 6626 43035
rect 6494 42932 6532 42988
rect 6588 42932 6626 42988
rect 6494 42746 6626 42932
rect 6488 42738 6632 42746
rect 6488 42622 6502 42738
rect 6618 42622 6632 42738
rect 6488 42614 6632 42622
rect 6786 29540 6854 43146
rect 6280 29340 6920 29540
rect 6280 17120 6480 29340
rect 6686 26488 6742 27794
rect 7514 26488 7570 27794
rect 8342 26488 8398 27794
rect 9170 26488 9226 27794
rect 9998 26488 10054 27808
rect 10826 26488 10882 27794
rect 11654 26488 11710 27794
rect 12116 26848 12316 26889
rect 12116 26712 12148 26848
rect 12284 26712 12316 26848
rect 6680 26486 6748 26488
rect 6680 26434 6688 26486
rect 6740 26434 6748 26486
rect 6680 26432 6748 26434
rect 7508 26486 7576 26488
rect 7508 26434 7516 26486
rect 7568 26434 7576 26486
rect 7508 26432 7576 26434
rect 8336 26486 8404 26488
rect 8336 26434 8344 26486
rect 8396 26434 8404 26486
rect 8336 26432 8404 26434
rect 9164 26486 9232 26488
rect 9164 26434 9172 26486
rect 9224 26434 9232 26486
rect 9164 26432 9232 26434
rect 9992 26486 10060 26488
rect 9992 26434 10000 26486
rect 10052 26434 10060 26486
rect 9992 26432 10060 26434
rect 10820 26486 10888 26488
rect 10820 26434 10828 26486
rect 10880 26434 10888 26486
rect 10820 26432 10888 26434
rect 11648 26486 11716 26488
rect 11648 26434 11656 26486
rect 11708 26434 11716 26486
rect 12116 26460 12316 26712
rect 12482 26488 12538 27794
rect 12986 26848 13186 26889
rect 12986 26712 13018 26848
rect 13154 26712 13186 26848
rect 12476 26486 12544 26488
rect 11648 26432 11716 26434
rect 12110 26450 12322 26460
rect 12110 26270 12126 26450
rect 12306 26270 12322 26450
rect 12476 26434 12484 26486
rect 12536 26434 12544 26486
rect 12986 26460 13186 26712
rect 14966 26488 15022 27794
rect 15794 26488 15850 27794
rect 16622 26488 16678 27794
rect 17450 26488 17506 27794
rect 18278 26488 18334 27794
rect 19106 26488 19162 27794
rect 14960 26486 15028 26488
rect 12476 26432 12544 26434
rect 12980 26450 13192 26460
rect 12110 26260 12322 26270
rect 12980 26270 12996 26450
rect 13176 26270 13192 26450
rect 14960 26434 14968 26486
rect 15020 26434 15028 26486
rect 14960 26432 15028 26434
rect 15788 26486 15856 26488
rect 15788 26434 15796 26486
rect 15848 26434 15856 26486
rect 15788 26432 15856 26434
rect 16616 26486 16684 26488
rect 16616 26434 16624 26486
rect 16676 26434 16684 26486
rect 16616 26432 16684 26434
rect 17444 26486 17512 26488
rect 17444 26434 17452 26486
rect 17504 26434 17512 26486
rect 17444 26432 17512 26434
rect 18272 26486 18340 26488
rect 18272 26434 18280 26486
rect 18332 26434 18340 26486
rect 18272 26432 18340 26434
rect 19100 26486 19168 26488
rect 19100 26434 19108 26486
rect 19160 26434 19168 26486
rect 19100 26432 19168 26434
rect 19934 26486 19990 27794
rect 19934 26434 19936 26486
rect 19988 26434 19990 26486
rect 20316 26848 20516 26889
rect 20316 26712 20348 26848
rect 20484 26712 20516 26848
rect 20316 26480 20516 26712
rect 20762 26486 20818 27794
rect 19934 26426 19990 26434
rect 20310 26470 20522 26480
rect 20310 26290 20326 26470
rect 20506 26290 20522 26470
rect 20762 26434 20764 26486
rect 20816 26434 20818 26486
rect 21186 26848 21386 26889
rect 21186 26712 21218 26848
rect 21354 26712 21386 26848
rect 21186 26480 21386 26712
rect 23246 26488 23302 27794
rect 24074 26488 24130 27794
rect 24902 26488 24958 27794
rect 25730 26488 25786 27794
rect 23240 26486 23308 26488
rect 20762 26426 20818 26434
rect 21180 26470 21392 26480
rect 20310 26280 20522 26290
rect 21180 26290 21196 26470
rect 21376 26290 21392 26470
rect 23240 26434 23248 26486
rect 23300 26434 23308 26486
rect 23240 26432 23308 26434
rect 24068 26486 24136 26488
rect 24068 26434 24076 26486
rect 24128 26434 24136 26486
rect 24068 26432 24136 26434
rect 24896 26486 24964 26488
rect 24896 26434 24904 26486
rect 24956 26434 24964 26486
rect 24896 26432 24964 26434
rect 25724 26486 25792 26488
rect 25724 26434 25732 26486
rect 25784 26434 25792 26486
rect 25724 26432 25792 26434
rect 26558 26486 26614 27794
rect 26558 26434 26560 26486
rect 26612 26434 26614 26486
rect 26558 26426 26614 26434
rect 27386 26486 27442 27794
rect 27386 26434 27388 26486
rect 27440 26434 27442 26486
rect 27386 26426 27442 26434
rect 28214 26486 28270 27794
rect 28214 26434 28216 26486
rect 28268 26434 28270 26486
rect 28516 26848 28716 26889
rect 28516 26712 28548 26848
rect 28684 26712 28716 26848
rect 28516 26480 28716 26712
rect 29042 26494 29098 27794
rect 28214 26426 28270 26434
rect 28510 26470 28722 26480
rect 21180 26280 21392 26290
rect 28510 26290 28526 26470
rect 28706 26290 28722 26470
rect 29042 26442 29044 26494
rect 29096 26442 29098 26494
rect 29386 26848 29586 26889
rect 29386 26712 29418 26848
rect 29554 26712 29586 26848
rect 29386 26480 29586 26712
rect 29042 26434 29098 26442
rect 29380 26470 29592 26480
rect 28510 26280 28722 26290
rect 29380 26290 29396 26470
rect 29576 26290 29592 26470
rect 29380 26280 29592 26290
rect 12980 26260 13192 26270
rect 6040 16920 6480 17120
rect 6040 5000 6240 16920
rect 29391 10514 29569 10518
rect 28700 10510 29574 10514
rect 28700 10330 28710 10510
rect 28890 10488 29574 10510
rect 28890 10352 29412 10488
rect 29548 10352 29574 10488
rect 28890 10330 29574 10352
rect 28700 10326 29574 10330
rect 29391 10322 29569 10326
rect 26057 10068 26224 10072
rect 25326 10047 26229 10068
rect 25326 10037 26072 10047
rect 25326 9921 25362 10037
rect 25478 9921 26072 10037
rect 25326 9911 26072 9921
rect 26208 9911 26229 10047
rect 25326 9891 26229 9911
rect 26057 9887 26224 9891
rect 25319 9626 25482 9630
rect 24568 9607 25487 9626
rect 24568 9597 25332 9607
rect 24568 9481 24602 9597
rect 24718 9481 25332 9597
rect 24568 9471 25332 9481
rect 25468 9471 25487 9607
rect 24568 9453 25487 9471
rect 25319 9449 25482 9453
rect 6040 4800 6960 5000
rect 4860 4600 5060 4606
rect 4091 4590 5060 4600
rect 4091 4568 4870 4590
rect 4091 4432 4132 4568
rect 4268 4432 4870 4568
rect 4091 4410 4870 4432
rect 5050 4410 5060 4590
rect 4091 4400 5060 4410
rect 4860 4394 5060 4400
rect 4560 3323 4760 3329
rect 4091 3313 4760 3323
rect 4091 3291 4570 3313
rect 4091 3155 4132 3291
rect 4268 3155 4570 3291
rect 4091 3133 4570 3155
rect 4750 3133 4760 3313
rect 4091 3123 4760 3133
rect 4560 3117 4760 3123
rect 6760 2930 6960 4800
rect 6760 2750 6770 2930
rect 6950 2750 6960 2930
rect 6760 2734 6960 2750
rect 7120 1790 7320 1806
rect 7120 1610 7130 1790
rect 7310 1610 7320 1790
rect 7120 1535 7320 1610
rect 7116 1508 7324 1535
rect 7116 1372 7152 1508
rect 7288 1372 7324 1508
rect 7116 1345 7324 1372
rect 7120 1340 7320 1345
<< via2 >>
rect 10368 44432 10424 44488
rect 11104 44408 11160 44464
rect 11840 44408 11896 44464
rect 12576 44408 12632 44464
rect 13312 44408 13368 44464
rect 14048 44408 14104 44464
rect 14784 44408 14840 44464
rect 15520 44408 15576 44464
rect 16256 44408 16312 44464
rect 16992 44408 17048 44464
rect 17728 44408 17784 44464
rect 24352 44208 24408 44264
rect 25088 44208 25144 44264
rect 25824 44208 25880 44264
rect 26560 44208 26616 44264
rect 27296 44208 27352 44264
rect 28032 44208 28088 44264
rect 28768 44208 28824 44264
rect 29504 44208 29560 44264
rect 6532 42932 6588 42988
rect 12148 26712 12284 26848
rect 13018 26712 13154 26848
rect 20348 26712 20484 26848
rect 21218 26712 21354 26848
rect 28548 26712 28684 26848
rect 29418 26712 29554 26848
rect 29412 10352 29548 10488
rect 26072 9911 26208 10047
rect 25332 9471 25468 9607
rect 4132 4432 4268 4568
rect 4132 3155 4268 3291
rect 7152 1372 7288 1508
<< metal3 >>
rect 6494 44781 6626 44806
rect 18432 44781 18528 44795
rect 6494 44773 18528 44781
rect 6494 44709 18448 44773
rect 18512 44709 18528 44773
rect 6494 44700 18528 44709
rect 6270 44459 6370 44460
rect 6265 44442 6375 44459
rect 6265 44378 6288 44442
rect 6352 44378 6375 44442
rect 6265 44361 6375 44378
rect 6270 44210 6370 44361
rect 4124 44192 6370 44210
rect 4124 44128 4148 44192
rect 4212 44128 6370 44192
rect 4124 44110 6370 44128
rect 1861 43680 1939 43685
rect 1860 43672 2606 43680
rect 1860 43608 1868 43672
rect 1932 43608 2528 43672
rect 2592 43608 2606 43672
rect 1860 43600 2606 43608
rect 1861 43595 1939 43600
rect 6494 43031 6626 44700
rect 18432 44687 18528 44700
rect 10358 44568 10364 44632
rect 10428 44568 10434 44632
rect 10366 44493 10426 44568
rect 11094 44554 11100 44618
rect 11164 44554 11170 44618
rect 11830 44554 11836 44618
rect 11900 44554 11906 44618
rect 12566 44554 12572 44618
rect 12636 44554 12642 44618
rect 13302 44554 13308 44618
rect 13372 44554 13378 44618
rect 14038 44554 14044 44618
rect 14108 44554 14114 44618
rect 14774 44554 14780 44618
rect 14844 44554 14850 44618
rect 15510 44554 15516 44618
rect 15580 44554 15586 44618
rect 16246 44554 16252 44618
rect 16316 44554 16322 44618
rect 16982 44554 16988 44618
rect 17052 44554 17058 44618
rect 17718 44554 17724 44618
rect 17788 44554 17794 44618
rect 24342 44554 24348 44618
rect 24412 44554 24418 44618
rect 25078 44554 25084 44618
rect 25148 44554 25154 44618
rect 25814 44554 25820 44618
rect 25884 44554 25890 44618
rect 26550 44554 26556 44618
rect 26620 44554 26626 44618
rect 27286 44554 27292 44618
rect 27356 44554 27362 44618
rect 28022 44554 28028 44618
rect 28092 44554 28098 44618
rect 28758 44554 28764 44618
rect 28828 44554 28834 44618
rect 29494 44554 29500 44618
rect 29564 44554 29570 44618
rect 10363 44488 10429 44493
rect 10363 44432 10368 44488
rect 10424 44432 10429 44488
rect 11102 44469 11162 44554
rect 11838 44469 11898 44554
rect 12574 44469 12634 44554
rect 13310 44469 13370 44554
rect 14046 44469 14106 44554
rect 14782 44469 14842 44554
rect 15518 44469 15578 44554
rect 16254 44469 16314 44554
rect 16990 44469 17050 44554
rect 17726 44469 17786 44554
rect 10363 44427 10429 44432
rect 11099 44464 11165 44469
rect 11099 44408 11104 44464
rect 11160 44408 11165 44464
rect 11099 44403 11165 44408
rect 11835 44464 11901 44469
rect 11835 44408 11840 44464
rect 11896 44408 11901 44464
rect 11835 44403 11901 44408
rect 12571 44464 12637 44469
rect 12571 44408 12576 44464
rect 12632 44408 12637 44464
rect 12571 44403 12637 44408
rect 13307 44464 13373 44469
rect 13307 44408 13312 44464
rect 13368 44408 13373 44464
rect 13307 44403 13373 44408
rect 14043 44464 14109 44469
rect 14043 44408 14048 44464
rect 14104 44408 14109 44464
rect 14043 44403 14109 44408
rect 14779 44464 14845 44469
rect 14779 44408 14784 44464
rect 14840 44408 14845 44464
rect 14779 44403 14845 44408
rect 15515 44464 15581 44469
rect 15515 44408 15520 44464
rect 15576 44408 15581 44464
rect 15515 44403 15581 44408
rect 16251 44464 16317 44469
rect 16251 44408 16256 44464
rect 16312 44408 16317 44464
rect 16251 44403 16317 44408
rect 16987 44464 17053 44469
rect 16987 44408 16992 44464
rect 17048 44408 17053 44464
rect 16987 44403 17053 44408
rect 17723 44464 17789 44469
rect 17723 44408 17728 44464
rect 17784 44408 17789 44464
rect 17723 44403 17789 44408
rect 11102 44320 11162 44403
rect 11838 44320 11898 44403
rect 12574 44320 12634 44403
rect 13310 44320 13370 44403
rect 14046 44320 14106 44403
rect 14782 44320 14842 44403
rect 15518 44320 15578 44403
rect 16254 44320 16314 44403
rect 16990 44320 17050 44403
rect 17726 44320 17786 44403
rect 24350 44269 24410 44554
rect 25086 44269 25146 44554
rect 25822 44269 25882 44554
rect 26558 44269 26618 44554
rect 27294 44269 27354 44554
rect 28030 44269 28090 44554
rect 28766 44269 28826 44554
rect 29502 44269 29562 44554
rect 24347 44264 24413 44269
rect 24347 44208 24352 44264
rect 24408 44208 24413 44264
rect 24347 44203 24413 44208
rect 25083 44264 25149 44269
rect 25083 44208 25088 44264
rect 25144 44208 25149 44264
rect 25083 44203 25149 44208
rect 25819 44264 25885 44269
rect 25819 44208 25824 44264
rect 25880 44208 25885 44264
rect 25819 44203 25885 44208
rect 26555 44264 26621 44269
rect 26555 44208 26560 44264
rect 26616 44208 26621 44264
rect 26555 44203 26621 44208
rect 27291 44264 27357 44269
rect 27291 44208 27296 44264
rect 27352 44208 27357 44264
rect 27291 44203 27357 44208
rect 28027 44264 28093 44269
rect 28027 44208 28032 44264
rect 28088 44208 28093 44264
rect 28027 44203 28093 44208
rect 28763 44264 28829 44269
rect 28763 44208 28768 44264
rect 28824 44208 28829 44264
rect 28763 44203 28829 44208
rect 29499 44264 29565 44269
rect 29499 44208 29504 44264
rect 29560 44208 29565 44264
rect 29499 44203 29565 44208
rect 19188 44141 19268 44146
rect 19039 44132 19269 44141
rect 19039 44068 19196 44132
rect 19260 44068 19269 44132
rect 19039 44059 19269 44068
rect 19188 44054 19268 44059
rect 19925 43981 20004 43986
rect 19040 43972 20005 43981
rect 19040 43908 19932 43972
rect 19996 43908 20005 43972
rect 19040 43900 20005 43908
rect 19925 43895 20004 43900
rect 20662 43820 20739 43825
rect 19041 43812 20740 43820
rect 19041 43748 20668 43812
rect 20732 43748 20740 43812
rect 19041 43741 20740 43748
rect 20662 43736 20739 43741
rect 21397 43660 21475 43665
rect 19040 43652 21476 43660
rect 19040 43588 21404 43652
rect 21468 43588 21476 43652
rect 19040 43580 21476 43588
rect 21397 43575 21475 43580
rect 6489 42988 6631 43031
rect 6489 42932 6532 42988
rect 6588 42932 6631 42988
rect 6489 42889 6631 42932
rect 30964 42339 31044 42340
rect 30959 42332 31049 42339
rect 30959 42268 30972 42332
rect 31036 42268 31049 42332
rect 30959 42261 31049 42268
rect 30964 41722 31044 42261
rect 30304 41642 31044 41722
rect 30804 41201 30876 41202
rect 30799 41198 30881 41201
rect 30799 41134 30808 41198
rect 30872 41134 30881 41198
rect 30799 41131 30881 41134
rect 30804 40620 30876 41131
rect 30294 40548 30876 40620
rect 8595 27532 9005 27539
rect 691 27490 989 27495
rect 8595 27490 8608 27532
rect 690 27452 8608 27490
rect 690 27228 728 27452
rect 952 27228 8608 27452
rect 690 27190 8608 27228
rect 691 27185 989 27190
rect 8595 27148 8608 27190
rect 8992 27490 9005 27532
rect 14015 27532 14425 27539
rect 14015 27490 14028 27532
rect 8992 27190 14028 27490
rect 8992 27148 9005 27190
rect 8595 27141 9005 27148
rect 14015 27148 14028 27190
rect 14412 27490 14425 27532
rect 19355 27532 19765 27539
rect 19355 27490 19368 27532
rect 14412 27190 19368 27490
rect 14412 27148 14425 27190
rect 14015 27141 14425 27148
rect 19355 27148 19368 27190
rect 19752 27490 19765 27532
rect 26015 27532 26425 27539
rect 26015 27490 26028 27532
rect 19752 27190 26028 27490
rect 19752 27148 19765 27190
rect 19355 27141 19765 27148
rect 26015 27148 26028 27190
rect 26412 27490 26425 27532
rect 26412 27190 27170 27490
rect 26412 27148 26425 27190
rect 26015 27141 26425 27148
rect 11015 26952 11425 26959
rect 2531 26930 2829 26935
rect 11015 26930 11028 26952
rect 2530 26892 11028 26930
rect 2530 26668 2568 26892
rect 2792 26668 11028 26892
rect 2530 26630 11028 26668
rect 2531 26625 2829 26630
rect 11015 26568 11028 26630
rect 11412 26930 11425 26952
rect 16855 26952 17265 26959
rect 16855 26930 16868 26952
rect 11412 26848 16868 26930
rect 11412 26712 12148 26848
rect 12284 26712 13018 26848
rect 13154 26712 16868 26848
rect 11412 26630 16868 26712
rect 11412 26568 11425 26630
rect 11015 26561 11425 26568
rect 16855 26568 16868 26630
rect 17252 26930 17265 26952
rect 22435 26952 22845 26959
rect 22435 26930 22448 26952
rect 17252 26848 22448 26930
rect 17252 26712 20348 26848
rect 20484 26712 21218 26848
rect 21354 26712 22448 26848
rect 17252 26630 22448 26712
rect 17252 26568 17265 26630
rect 16855 26561 17265 26568
rect 22435 26568 22448 26630
rect 22832 26930 22845 26952
rect 29555 26952 29965 26959
rect 29555 26930 29568 26952
rect 22832 26848 29568 26930
rect 22832 26712 28548 26848
rect 28684 26712 29418 26848
rect 29554 26712 29568 26848
rect 22832 26630 29568 26712
rect 22832 26568 22845 26630
rect 22435 26561 22845 26568
rect 29555 26568 29568 26630
rect 29952 26930 29965 26952
rect 29952 26630 29970 26930
rect 29952 26568 29965 26630
rect 29555 26561 29965 26568
rect 31279 10514 31465 10519
rect 29386 10492 31466 10514
rect 29386 10488 31300 10492
rect 29386 10352 29412 10488
rect 29548 10352 31300 10488
rect 29386 10348 31300 10352
rect 31444 10348 31466 10492
rect 29386 10326 31466 10348
rect 31279 10321 31465 10326
rect 26869 10068 27044 10073
rect 26052 10051 27045 10068
rect 26052 10047 26884 10051
rect 26052 9911 26072 10047
rect 26208 9911 26884 10047
rect 26052 9907 26884 9911
rect 27028 9907 27045 10051
rect 26052 9891 27045 9907
rect 26869 9886 27044 9891
rect 26134 9626 26305 9631
rect 25314 9611 26306 9626
rect 25314 9607 26147 9611
rect 25314 9471 25332 9607
rect 25468 9471 26147 9607
rect 25314 9467 26147 9471
rect 26291 9467 26306 9611
rect 25314 9453 26306 9467
rect 26134 9448 26305 9453
rect 4095 4600 4305 4605
rect 3414 4572 4305 4600
rect 3414 4428 3448 4572
rect 3592 4568 4305 4572
rect 3592 4432 4132 4568
rect 4268 4432 4305 4568
rect 3592 4428 4305 4432
rect 3414 4400 4305 4428
rect 4095 4395 4305 4400
rect 4095 3323 4305 3328
rect 1174 3295 4305 3323
rect 1174 3151 1208 3295
rect 1352 3291 4305 3295
rect 1352 3155 4132 3291
rect 4268 3155 4305 3291
rect 1352 3151 4305 3155
rect 1174 3123 4305 3151
rect 4095 3118 4305 3123
rect 7120 1508 7320 1540
rect 7120 1372 7152 1508
rect 7288 1372 7320 1508
rect 7120 1312 7320 1372
rect 7120 1168 7148 1312
rect 7292 1168 7320 1312
rect 7120 1134 7320 1168
<< via3 >>
rect 18448 44709 18512 44773
rect 6288 44378 6352 44442
rect 4148 44128 4212 44192
rect 1868 43608 1932 43672
rect 2528 43608 2592 43672
rect 10364 44568 10428 44632
rect 11100 44554 11164 44618
rect 11836 44554 11900 44618
rect 12572 44554 12636 44618
rect 13308 44554 13372 44618
rect 14044 44554 14108 44618
rect 14780 44554 14844 44618
rect 15516 44554 15580 44618
rect 16252 44554 16316 44618
rect 16988 44554 17052 44618
rect 17724 44554 17788 44618
rect 24348 44554 24412 44618
rect 25084 44554 25148 44618
rect 25820 44554 25884 44618
rect 26556 44554 26620 44618
rect 27292 44554 27356 44618
rect 28028 44554 28092 44618
rect 28764 44554 28828 44618
rect 29500 44554 29564 44618
rect 19196 44068 19260 44132
rect 19932 43908 19996 43972
rect 20668 43748 20732 43812
rect 21404 43588 21468 43652
rect 30972 42268 31036 42332
rect 30808 41134 30872 41198
rect 728 27228 952 27452
rect 8608 27148 8992 27532
rect 14028 27148 14412 27532
rect 19368 27148 19752 27532
rect 26028 27148 26412 27532
rect 2568 26668 2792 26892
rect 11028 26568 11412 26952
rect 16868 26568 17252 26952
rect 22448 26568 22832 26952
rect 29568 26568 29952 26952
rect 31300 10348 31444 10492
rect 26884 9907 27028 10051
rect 26147 9467 26291 9611
rect 3448 4428 3592 4572
rect 1208 3151 1352 3295
rect 7148 1168 7292 1312
<< metal4 >>
rect 798 44160 858 45152
rect 1534 44460 1594 45152
rect 2270 44460 2330 45152
rect 3006 44460 3066 45152
rect 3742 44460 3802 45152
rect 4478 44460 4538 45152
rect 5214 44460 5274 45152
rect 5950 44460 6010 45152
rect 6686 44460 6746 45152
rect 7422 44460 7482 45152
rect 8158 44460 8218 45152
rect 8894 44460 8954 45152
rect 9630 44460 9690 45152
rect 10366 44633 10426 45152
rect 10363 44632 10429 44633
rect 10363 44568 10364 44632
rect 10428 44568 10429 44632
rect 11102 44619 11162 45152
rect 11838 44619 11898 45152
rect 12574 44619 12634 45152
rect 13310 44619 13370 45152
rect 14046 44619 14106 45152
rect 14782 44619 14842 45152
rect 15518 44619 15578 45152
rect 16254 44619 16314 45152
rect 16990 44619 17050 45152
rect 17726 44619 17786 45152
rect 18462 44908 18522 45152
rect 18432 44790 18528 44908
rect 18431 44773 18529 44790
rect 18431 44709 18448 44773
rect 18512 44709 18529 44773
rect 18431 44692 18529 44709
rect 10363 44567 10429 44568
rect 11099 44618 11165 44619
rect 11099 44554 11100 44618
rect 11164 44554 11165 44618
rect 11099 44553 11165 44554
rect 11835 44618 11901 44619
rect 11835 44554 11836 44618
rect 11900 44554 11901 44618
rect 11835 44553 11901 44554
rect 12571 44618 12637 44619
rect 12571 44554 12572 44618
rect 12636 44554 12637 44618
rect 12571 44553 12637 44554
rect 13307 44618 13373 44619
rect 13307 44554 13308 44618
rect 13372 44554 13373 44618
rect 13307 44553 13373 44554
rect 14043 44618 14109 44619
rect 14043 44554 14044 44618
rect 14108 44554 14109 44618
rect 14043 44553 14109 44554
rect 14779 44618 14845 44619
rect 14779 44554 14780 44618
rect 14844 44554 14845 44618
rect 14779 44553 14845 44554
rect 15515 44618 15581 44619
rect 15515 44554 15516 44618
rect 15580 44554 15581 44618
rect 15515 44553 15581 44554
rect 16251 44618 16317 44619
rect 16251 44554 16252 44618
rect 16316 44554 16317 44618
rect 16251 44553 16317 44554
rect 16987 44618 17053 44619
rect 16987 44554 16988 44618
rect 17052 44554 17053 44618
rect 16987 44553 17053 44554
rect 17723 44618 17789 44619
rect 17723 44554 17724 44618
rect 17788 44554 17789 44618
rect 17723 44553 17789 44554
rect 11102 44540 11162 44553
rect 11838 44540 11898 44553
rect 12574 44540 12634 44553
rect 13310 44540 13370 44553
rect 14046 44540 14106 44553
rect 14782 44540 14842 44553
rect 15518 44540 15578 44553
rect 16254 44540 16314 44553
rect 16990 44540 17050 44553
rect 1480 44438 3802 44460
rect 1480 44210 3800 44438
rect 4440 44360 6020 44460
rect 6270 44442 9740 44460
rect 6270 44378 6288 44442
rect 6352 44378 9740 44442
rect 6270 44360 9740 44378
rect 4129 44210 4231 44211
rect 1480 44192 4231 44210
rect 1480 44160 4148 44192
rect 200 43680 500 44152
rect 798 44128 4148 44160
rect 4212 44128 4231 44192
rect 798 44110 4231 44128
rect 798 44100 3800 44110
rect 4129 44109 4231 44110
rect 1480 43920 3800 44100
rect 4440 43920 4600 44360
rect 19198 44141 19258 45152
rect 19187 44132 19269 44141
rect 19187 44068 19196 44132
rect 19260 44068 19269 44132
rect 19187 44059 19269 44068
rect 19198 44040 19258 44059
rect 19934 43981 19994 45152
rect 19924 43972 20005 43981
rect 200 43672 1940 43680
rect 200 43608 1868 43672
rect 1932 43608 1940 43672
rect 200 43600 1940 43608
rect 200 27490 500 43600
rect 200 27452 990 27490
rect 200 27228 728 27452
rect 952 27228 990 27452
rect 200 27190 990 27228
rect 200 3323 500 27190
rect 2100 26930 2400 43920
rect 2519 43680 2601 43681
rect 4480 43680 4560 43920
rect 19924 43908 19932 43972
rect 19996 43908 20005 43972
rect 19924 43900 20005 43908
rect 19934 43880 19994 43900
rect 20670 43820 20730 45152
rect 20661 43812 20740 43820
rect 20661 43748 20668 43812
rect 20732 43748 20740 43812
rect 20661 43741 20740 43748
rect 20670 43720 20730 43741
rect 2519 43672 4560 43680
rect 2519 43608 2528 43672
rect 2592 43608 4560 43672
rect 21406 43660 21466 45152
rect 22142 44854 22202 45152
rect 22878 44854 22938 45152
rect 23614 44854 23674 45152
rect 24350 44619 24410 45152
rect 25086 44619 25146 45152
rect 25822 44619 25882 45152
rect 26558 44619 26618 45152
rect 27294 44619 27354 45152
rect 28030 44619 28090 45152
rect 28766 44619 28826 45152
rect 29502 44619 29562 45152
rect 24347 44618 24413 44619
rect 24347 44554 24348 44618
rect 24412 44554 24413 44618
rect 24347 44553 24413 44554
rect 25083 44618 25149 44619
rect 25083 44554 25084 44618
rect 25148 44554 25149 44618
rect 25083 44553 25149 44554
rect 25819 44618 25885 44619
rect 25819 44554 25820 44618
rect 25884 44554 25885 44618
rect 25819 44553 25885 44554
rect 26555 44618 26621 44619
rect 26555 44554 26556 44618
rect 26620 44554 26621 44618
rect 26555 44553 26621 44554
rect 27291 44618 27357 44619
rect 27291 44554 27292 44618
rect 27356 44554 27357 44618
rect 27291 44553 27357 44554
rect 28027 44618 28093 44619
rect 28027 44554 28028 44618
rect 28092 44554 28093 44618
rect 28027 44553 28093 44554
rect 28763 44618 28829 44619
rect 28763 44554 28764 44618
rect 28828 44554 28829 44618
rect 28763 44553 28829 44554
rect 29499 44618 29565 44619
rect 29499 44554 29500 44618
rect 29564 44554 29565 44618
rect 29499 44553 29565 44554
rect 30238 44256 30298 45152
rect 30238 44196 30600 44256
rect 2519 43600 4560 43608
rect 21396 43652 21476 43660
rect 2519 43599 2601 43600
rect 21396 43588 21404 43652
rect 21468 43588 21476 43652
rect 21396 43580 21476 43588
rect 21406 43560 21466 43580
rect 30540 42024 30600 44196
rect 30974 42340 31034 45152
rect 31710 44952 31770 45152
rect 30964 42332 31044 42340
rect 30964 42268 30972 42332
rect 31036 42268 31044 42332
rect 30964 42260 31044 42268
rect 30540 41964 30870 42024
rect 30810 41202 30870 41964
rect 30804 41198 30876 41202
rect 30804 41134 30808 41198
rect 30872 41134 30876 41198
rect 30804 41130 30876 41134
rect 8020 28240 9000 28640
rect 8600 27532 9000 28240
rect 8600 27148 8608 27532
rect 8992 27148 9000 27532
rect 8600 27140 9000 27148
rect 11020 26952 11420 28714
rect 14020 27532 14420 28634
rect 14020 27148 14028 27532
rect 14412 27148 14420 27532
rect 14020 27140 14420 27148
rect 16860 28400 17520 28800
rect 2100 26892 2830 26930
rect 2100 26668 2568 26892
rect 2792 26668 2830 26892
rect 2100 26630 2830 26668
rect 2100 4600 2400 26630
rect 11020 26568 11028 26952
rect 11412 26568 11420 26952
rect 11020 26560 11420 26568
rect 16860 26952 17260 28400
rect 19360 28234 20420 28634
rect 22440 28314 23420 28714
rect 19360 27532 19760 28234
rect 19360 27148 19368 27532
rect 19752 27148 19760 27532
rect 19360 27140 19760 27148
rect 16860 26568 16868 26952
rect 17252 26568 17260 26952
rect 16860 26560 17260 26568
rect 22440 26952 22840 28314
rect 26020 27532 26420 28634
rect 29020 28314 29960 28714
rect 26020 27148 26028 27532
rect 26412 27148 26420 27532
rect 26020 27140 26420 27148
rect 22440 26568 22448 26952
rect 22832 26568 22840 26952
rect 22440 26560 22840 26568
rect 29560 26952 29960 28314
rect 29560 26568 29568 26952
rect 29952 26568 29960 26952
rect 29560 26560 29960 26568
rect 31278 10492 31466 10514
rect 31278 10348 31300 10492
rect 31444 10348 31466 10492
rect 26868 10051 27045 10068
rect 26868 9907 26884 10051
rect 27028 9907 27045 10051
rect 26133 9611 26306 9626
rect 26133 9467 26147 9611
rect 26291 9467 26306 9611
rect 3419 4600 3621 4601
rect 2100 4572 3621 4600
rect 2100 4428 3448 4572
rect 3592 4428 3621 4572
rect 2100 4400 3621 4428
rect 1179 3323 1381 3324
rect 200 3295 1381 3323
rect 200 3151 1208 3295
rect 1352 3151 1381 3295
rect 200 3123 1381 3151
rect 200 1000 500 3123
rect 1179 3122 1381 3123
rect 2100 1000 2400 4400
rect 3419 4399 3621 4400
rect 7119 1312 7321 1341
rect 7119 1168 7148 1312
rect 7292 1168 7321 1312
rect 7119 1139 7321 1168
rect 7120 760 7320 1139
rect 26133 827 26306 9467
rect 7120 720 17980 760
rect 7120 600 18184 720
rect 22454 654 26306 827
rect 26868 772 27045 9907
rect 31278 846 31466 10348
rect 7120 560 17980 600
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 280
rect 13648 0 13768 200
rect 18064 0 18184 600
rect 22480 0 22600 654
rect 26896 0 27016 772
rect 31312 0 31432 846
use inverter  inverter_0
timestamp 1713537803
transform 1 0 5390 0 1 1613
box -410 547 1220 2810
use r2r  r2r_blue
timestamp 1713537803
transform 0 1 12386 -1 0 25766
box -400 -5786 14766 800
use r2r  r2r_green
timestamp 1713537803
transform 0 1 20586 -1 0 25766
box -400 -5786 14766 800
use r2r  r2r_red
timestamp 1713537803
transform 0 1 28786 -1 0 25766
box -400 -5786 14766 800
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 600 90 0 0 clk
port 1 nsew
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 600 90 0 0 ena
port 2 nsew
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 600 90 0 0 rst_n
port 3 nsew
flabel metal4 s 31312 0 31432 200 0 FreeSans 1200 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26896 0 27016 200 0 FreeSans 1200 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 22480 0 22600 200 0 FreeSans 1200 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 18064 0 18184 200 0 FreeSans 1200 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 13648 0 13768 200 0 FreeSans 1200 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 9232 0 9352 200 0 FreeSans 1200 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 4816 0 4936 200 0 FreeSans 1200 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 400 0 520 200 0 FreeSans 1200 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 600 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 600 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 600 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 600 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 600 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 600 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 600 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 600 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 600 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 600 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 600 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 600 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 600 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 600 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 600 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 600 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 600 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 600 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 798 44952 858 45152 0 FreeSans 600 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 600 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 600 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 600 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 600 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 600 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 600 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 600 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 600 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 600 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 600 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 200 1000 500 44152 1 FreeSans 3 0 0 0 VPWR
port 52 nsew
flabel metal4 s 2100 1000 2400 44152 1 FreeSans 3 0 0 0 VGND
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
string GDS_END 2390302
string GDS_FILE /home/anton/projects/tt06-grab-bag/gds/tt_um_algofoogle_tt06_grab_bag.gds
string GDS_START 2316714
<< end >>
