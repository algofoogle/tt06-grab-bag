** sch_path: /home/anton/projects/tt06-grab-bag/xschem/tb_r2r.sch
**.subckt tb_r2r
x1 a_int d7 d6 d5 d4 d3 d2 d1 d0 GND GND r2r
x2 out net1 GND tt06_analog_load
V1 d0 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 20ns 40ns)
V2 d1 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 40ns 80ns)
V3 d2 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 80ns 160ns)
V4 d3 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 160ns 320ns)
V5 d4 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 320ns 640ns)
V6 d5 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 640ns 1280ns)
V7 d6 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 1280ns 2560ns)
V8 d7 GND pulse(0V 1.8V 0ns 0.5ns 0.5ns 2560ns 5120ns)
x3 a_int_parax d7 d6 d5 d4 d3 d2 d1 d0 GND GND r2r_parax
x4 out_parax a_int_parax GND tt06_analog_load
V10 VCC GND 1.8
R1 net1 GND 100k m=1
XM1 VCC b_int net1 net1 sky130_fd_pr__nfet_01v8 L=0.15 W=40 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R2 b_int a_int 150k m=1
R3 VCC b_int 200k m=1
R4 out GND 200k m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/anton/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.tech/ngspice/sky130.lib.spice tt





* .options filetype=ascii
.options savecurrents
.control
  save all
  tran 2n 5.5u uic
  write tb_r2r.raw
  quit
.endc
.end



**** end user architecture code
**.ends

* expanding   symbol:  r2r.sym # of pins=11
** sym_path: /home/anton/projects/tt06-grab-bag/xschem/r2r.sym
** sch_path: /home/anton/projects/tt06-grab-bag/xschem/r2r.sch
.subckt r2r aout d7 d6 d5 d4 d3 d2 d1 d0 GND VSUBS
*.ipin d0
*.ipin d1
*.ipin d2
*.ipin d3
*.ipin d4
*.ipin d5
*.ipin d6
*.ipin d7
*.iopin GND
*.iopin VSUBS
*.opin aout
XR1 d0 net1 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR2 d1 net2 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR3 d2 net3 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR4 d3 net4 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR5 d4 net5 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR6 d5 net6 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR7 d6 net7 VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR8 d7 aout VSUBS sky130_fd_pr__res_high_po_0p69 L=39.9 mult=1 m=1
XR9 GND net1 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR10 net1 net2 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR11 net2 net3 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR12 net3 net4 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR13 net4 net5 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR14 net5 net6 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR15 net6 net7 VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
XR16 net7 aout VSUBS sky130_fd_pr__res_high_po_0p69 L=19.55 mult=1 m=1
.ends


* expanding   symbol:  tt06_analog_load.sym # of pins=3
** sym_path: /home/anton/projects/tt06-grab-bag/xschem/tt06_analog_load.sym
** sch_path: /home/anton/projects/tt06-grab-bag/xschem/tt06_analog_load.sch
.subckt tt06_analog_load a_ext a_int GND
*.iopin a_int
*.iopin a_ext
*.iopin GND
R1 a_ext a_int 500 m=1
C1 a_int GND 2.5p m=1
C2 a_ext GND 2.5p m=1
.ends


* expanding   symbol:  r2r_parax.sym # of pins=11
** sym_path: /home/anton/projects/tt06-grab-bag/xschem/r2r.sym
.include /home/anton/projects/tt06-grab-bag/mag/r2r.sim.spice
.GLOBAL GND
.end
