magic
tech sky130A
magscale 1 2
timestamp 1713537803
<< locali >>
rect 4772 431 4932 448
rect 4772 397 4799 431
rect 4833 397 4871 431
rect 4905 397 4932 431
rect 4772 380 4932 397
rect 14586 361 14658 362
rect 14586 327 14605 361
rect 14639 327 14658 361
rect 14586 289 14658 327
rect 14586 255 14605 289
rect 14639 255 14658 289
rect 14586 217 14658 255
rect 14586 183 14605 217
rect 14639 183 14658 217
rect 14586 145 14658 183
rect 14586 111 14605 145
rect 14639 111 14658 145
rect 14586 110 14658 111
rect 4772 71 4932 88
rect 4772 37 4799 71
rect 4833 37 4871 71
rect 4905 37 4932 71
rect 4772 20 4932 37
rect 4772 -369 4932 -352
rect 4772 -403 4799 -369
rect 4833 -403 4871 -369
rect 4905 -403 4932 -369
rect 4772 -420 4932 -403
rect 14586 -439 14658 -438
rect 14586 -473 14605 -439
rect 14639 -473 14658 -439
rect 14586 -511 14658 -473
rect 14586 -545 14605 -511
rect 14639 -545 14658 -511
rect 14586 -583 14658 -545
rect 14586 -617 14605 -583
rect 14639 -617 14658 -583
rect 14586 -655 14658 -617
rect 14586 -689 14605 -655
rect 14639 -689 14658 -655
rect 14586 -690 14658 -689
rect 4772 -729 4932 -712
rect 4772 -763 4799 -729
rect 4833 -763 4871 -729
rect 4905 -763 4932 -729
rect 4772 -780 4932 -763
rect 4772 -1169 4932 -1152
rect 4772 -1203 4799 -1169
rect 4833 -1203 4871 -1169
rect 4905 -1203 4932 -1169
rect 4772 -1220 4932 -1203
rect 14586 -1239 14658 -1238
rect 14586 -1273 14605 -1239
rect 14639 -1273 14658 -1239
rect 14586 -1311 14658 -1273
rect 14586 -1345 14605 -1311
rect 14639 -1345 14658 -1311
rect 14586 -1383 14658 -1345
rect 14586 -1417 14605 -1383
rect 14639 -1417 14658 -1383
rect 14586 -1455 14658 -1417
rect 14586 -1489 14605 -1455
rect 14639 -1489 14658 -1455
rect 14586 -1490 14658 -1489
rect 4772 -1529 4932 -1512
rect 4772 -1563 4799 -1529
rect 4833 -1563 4871 -1529
rect 4905 -1563 4932 -1529
rect 4772 -1580 4932 -1563
rect 4772 -1969 4932 -1952
rect 4772 -2003 4799 -1969
rect 4833 -2003 4871 -1969
rect 4905 -2003 4932 -1969
rect 4772 -2020 4932 -2003
rect 14586 -2039 14658 -2038
rect 14586 -2073 14605 -2039
rect 14639 -2073 14658 -2039
rect 14586 -2111 14658 -2073
rect 14586 -2145 14605 -2111
rect 14639 -2145 14658 -2111
rect 14586 -2183 14658 -2145
rect 14586 -2217 14605 -2183
rect 14639 -2217 14658 -2183
rect 14586 -2255 14658 -2217
rect 14586 -2289 14605 -2255
rect 14639 -2289 14658 -2255
rect 14586 -2290 14658 -2289
rect 4772 -2329 4932 -2312
rect 4772 -2363 4799 -2329
rect 4833 -2363 4871 -2329
rect 4905 -2363 4932 -2329
rect 4772 -2380 4932 -2363
rect 4772 -2769 4932 -2752
rect 4772 -2803 4799 -2769
rect 4833 -2803 4871 -2769
rect 4905 -2803 4932 -2769
rect 4772 -2820 4932 -2803
rect 14586 -2839 14658 -2838
rect 14586 -2873 14605 -2839
rect 14639 -2873 14658 -2839
rect 14586 -2911 14658 -2873
rect 14586 -2945 14605 -2911
rect 14639 -2945 14658 -2911
rect 14586 -2983 14658 -2945
rect 14586 -3017 14605 -2983
rect 14639 -3017 14658 -2983
rect 14586 -3055 14658 -3017
rect 14586 -3089 14605 -3055
rect 14639 -3089 14658 -3055
rect 14586 -3090 14658 -3089
rect 4772 -3129 4932 -3112
rect 4772 -3163 4799 -3129
rect 4833 -3163 4871 -3129
rect 4905 -3163 4932 -3129
rect 4772 -3180 4932 -3163
rect 4772 -3569 4932 -3552
rect 4772 -3603 4799 -3569
rect 4833 -3603 4871 -3569
rect 4905 -3603 4932 -3569
rect 4772 -3620 4932 -3603
rect 14586 -3639 14658 -3638
rect 14586 -3673 14605 -3639
rect 14639 -3673 14658 -3639
rect 14586 -3711 14658 -3673
rect 14586 -3745 14605 -3711
rect 14639 -3745 14658 -3711
rect 14586 -3783 14658 -3745
rect 14586 -3817 14605 -3783
rect 14639 -3817 14658 -3783
rect 14586 -3855 14658 -3817
rect 14586 -3889 14605 -3855
rect 14639 -3889 14658 -3855
rect 14586 -3890 14658 -3889
rect 4772 -3929 4932 -3912
rect 4772 -3963 4799 -3929
rect 4833 -3963 4871 -3929
rect 4905 -3963 4932 -3929
rect 4772 -3980 4932 -3963
rect 4772 -4369 4932 -4352
rect 4772 -4403 4799 -4369
rect 4833 -4403 4871 -4369
rect 4905 -4403 4932 -4369
rect 4772 -4420 4932 -4403
rect 14586 -4439 14658 -4438
rect 14586 -4473 14605 -4439
rect 14639 -4473 14658 -4439
rect 14586 -4511 14658 -4473
rect 14586 -4545 14605 -4511
rect 14639 -4545 14658 -4511
rect 14586 -4583 14658 -4545
rect 14586 -4617 14605 -4583
rect 14639 -4617 14658 -4583
rect 14586 -4655 14658 -4617
rect 14586 -4689 14605 -4655
rect 14639 -4689 14658 -4655
rect 14586 -4690 14658 -4689
rect 4772 -4729 4932 -4712
rect 4772 -4763 4799 -4729
rect 4833 -4763 4871 -4729
rect 4905 -4763 4932 -4729
rect 4772 -4780 4932 -4763
rect 4772 -5169 4932 -5152
rect 4772 -5203 4799 -5169
rect 4833 -5203 4871 -5169
rect 4905 -5203 4932 -5169
rect 4772 -5220 4932 -5203
rect 14586 -5239 14658 -5238
rect 14586 -5273 14605 -5239
rect 14639 -5273 14658 -5239
rect 14586 -5311 14658 -5273
rect 14586 -5345 14605 -5311
rect 14639 -5345 14658 -5311
rect 14586 -5383 14658 -5345
rect 14586 -5417 14605 -5383
rect 14639 -5417 14658 -5383
rect 14586 -5455 14658 -5417
rect 14586 -5489 14605 -5455
rect 14639 -5489 14658 -5455
rect 14586 -5490 14658 -5489
rect 4772 -5529 4932 -5512
rect 4772 -5563 4799 -5529
rect 4833 -5563 4871 -5529
rect 4905 -5563 4932 -5529
rect 4772 -5580 4932 -5563
<< viali >>
rect 4799 397 4833 431
rect 4871 397 4905 431
rect 14605 327 14639 361
rect 14605 255 14639 289
rect 14605 183 14639 217
rect 14605 111 14639 145
rect 4799 37 4833 71
rect 4871 37 4905 71
rect 4799 -403 4833 -369
rect 4871 -403 4905 -369
rect 14605 -473 14639 -439
rect 14605 -545 14639 -511
rect 14605 -617 14639 -583
rect 14605 -689 14639 -655
rect 4799 -763 4833 -729
rect 4871 -763 4905 -729
rect 4799 -1203 4833 -1169
rect 4871 -1203 4905 -1169
rect 14605 -1273 14639 -1239
rect 14605 -1345 14639 -1311
rect 14605 -1417 14639 -1383
rect 14605 -1489 14639 -1455
rect 4799 -1563 4833 -1529
rect 4871 -1563 4905 -1529
rect 4799 -2003 4833 -1969
rect 4871 -2003 4905 -1969
rect 14605 -2073 14639 -2039
rect 14605 -2145 14639 -2111
rect 14605 -2217 14639 -2183
rect 14605 -2289 14639 -2255
rect 4799 -2363 4833 -2329
rect 4871 -2363 4905 -2329
rect 4799 -2803 4833 -2769
rect 4871 -2803 4905 -2769
rect 14605 -2873 14639 -2839
rect 14605 -2945 14639 -2911
rect 14605 -3017 14639 -2983
rect 14605 -3089 14639 -3055
rect 4799 -3163 4833 -3129
rect 4871 -3163 4905 -3129
rect 4799 -3603 4833 -3569
rect 4871 -3603 4905 -3569
rect 14605 -3673 14639 -3639
rect 14605 -3745 14639 -3711
rect 14605 -3817 14639 -3783
rect 14605 -3889 14639 -3855
rect 4799 -3963 4833 -3929
rect 4871 -3963 4905 -3929
rect 4799 -4403 4833 -4369
rect 4871 -4403 4905 -4369
rect 14605 -4473 14639 -4439
rect 14605 -4545 14639 -4511
rect 14605 -4617 14639 -4583
rect 14605 -4689 14639 -4655
rect 4799 -4763 4833 -4729
rect 4871 -4763 4905 -4729
rect 4799 -5203 4833 -5169
rect 4871 -5203 4905 -5169
rect 14605 -5273 14639 -5239
rect 14605 -5345 14639 -5311
rect 14605 -5417 14639 -5383
rect 14605 -5489 14639 -5455
rect 4799 -5563 4833 -5529
rect 4871 -5563 4905 -5529
<< metal1 >>
rect -400 600 14380 800
rect 4750 431 4950 496
rect 4750 397 4799 431
rect 4833 397 4871 431
rect 4905 397 4950 431
rect -400 130 500 330
rect 4750 71 4950 397
rect 9880 330 10080 336
rect 8636 130 10080 330
rect 4750 37 4799 71
rect 4833 37 4871 71
rect 4905 37 4950 71
rect 4750 -66 4950 37
rect 9880 -60 10080 130
rect 14180 118 14380 600
rect 14560 361 14760 398
rect 14560 327 14605 361
rect 14639 327 14760 361
rect 14560 289 14760 327
rect 14560 255 14605 289
rect 14639 255 14760 289
rect 14560 217 14760 255
rect 14560 183 14605 217
rect 14639 183 14760 217
rect 14560 145 14760 183
rect 14560 111 14605 145
rect 14639 111 14760 145
rect 4744 -70 4956 -66
rect -400 -76 4956 -70
rect -400 -256 4760 -76
rect 4940 -256 4956 -76
rect -400 -266 4956 -256
rect 9880 -260 14378 -60
rect -400 -270 4950 -266
rect 4750 -369 4950 -270
rect 4750 -403 4799 -369
rect 4833 -403 4871 -369
rect 4905 -403 4950 -369
rect -400 -670 500 -470
rect 4750 -729 4950 -403
rect 9880 -470 10080 -464
rect 8636 -670 10080 -470
rect 4750 -763 4799 -729
rect 4833 -763 4871 -729
rect 4905 -763 4950 -729
rect 4750 -1169 4950 -763
rect 9880 -860 10080 -670
rect 14178 -688 14378 -260
rect 14560 -76 14760 111
rect 14560 -256 14570 -76
rect 14750 -256 14760 -76
rect 14560 -439 14760 -256
rect 14560 -473 14605 -439
rect 14639 -473 14760 -439
rect 14560 -511 14760 -473
rect 14560 -545 14605 -511
rect 14639 -545 14760 -511
rect 14560 -583 14760 -545
rect 14560 -617 14605 -583
rect 14639 -617 14760 -583
rect 14560 -655 14760 -617
rect 14560 -689 14605 -655
rect 14639 -689 14760 -655
rect 9880 -1060 14378 -860
rect 4750 -1203 4799 -1169
rect 4833 -1203 4871 -1169
rect 4905 -1203 4950 -1169
rect -400 -1470 500 -1270
rect 4750 -1529 4950 -1203
rect 9880 -1270 10080 -1264
rect 8636 -1470 10080 -1270
rect 4750 -1563 4799 -1529
rect 4833 -1563 4871 -1529
rect 4905 -1563 4950 -1529
rect 4750 -1969 4950 -1563
rect 9880 -1660 10080 -1470
rect 14178 -1488 14378 -1060
rect 14560 -1239 14760 -689
rect 14560 -1273 14605 -1239
rect 14639 -1273 14760 -1239
rect 14560 -1311 14760 -1273
rect 14560 -1345 14605 -1311
rect 14639 -1345 14760 -1311
rect 14560 -1383 14760 -1345
rect 14560 -1417 14605 -1383
rect 14639 -1417 14760 -1383
rect 14560 -1455 14760 -1417
rect 14560 -1489 14605 -1455
rect 14639 -1489 14760 -1455
rect 9880 -1860 14378 -1660
rect 4750 -2003 4799 -1969
rect 4833 -2003 4871 -1969
rect 4905 -2003 4950 -1969
rect -400 -2270 500 -2070
rect 4750 -2329 4950 -2003
rect 9880 -2070 10080 -2064
rect 8636 -2270 10080 -2070
rect 4750 -2363 4799 -2329
rect 4833 -2363 4871 -2329
rect 4905 -2363 4950 -2329
rect 4750 -2769 4950 -2363
rect 9880 -2460 10080 -2270
rect 14178 -2288 14378 -1860
rect 14560 -2039 14760 -1489
rect 14560 -2073 14605 -2039
rect 14639 -2073 14760 -2039
rect 14560 -2111 14760 -2073
rect 14560 -2145 14605 -2111
rect 14639 -2145 14760 -2111
rect 14560 -2183 14760 -2145
rect 14560 -2217 14605 -2183
rect 14639 -2217 14760 -2183
rect 14560 -2255 14760 -2217
rect 14560 -2289 14605 -2255
rect 14639 -2289 14760 -2255
rect 9880 -2660 14378 -2460
rect 4750 -2803 4799 -2769
rect 4833 -2803 4871 -2769
rect 4905 -2803 4950 -2769
rect -400 -3070 500 -2870
rect 4750 -3129 4950 -2803
rect 9880 -2870 10080 -2864
rect 8636 -3070 10080 -2870
rect 4750 -3163 4799 -3129
rect 4833 -3163 4871 -3129
rect 4905 -3163 4950 -3129
rect 4750 -3569 4950 -3163
rect 9880 -3260 10080 -3070
rect 14178 -3088 14378 -2660
rect 14560 -2839 14760 -2289
rect 14560 -2873 14605 -2839
rect 14639 -2873 14760 -2839
rect 14560 -2911 14760 -2873
rect 14560 -2945 14605 -2911
rect 14639 -2945 14760 -2911
rect 14560 -2983 14760 -2945
rect 14560 -3017 14605 -2983
rect 14639 -3017 14760 -2983
rect 14560 -3055 14760 -3017
rect 14560 -3089 14605 -3055
rect 14639 -3089 14760 -3055
rect 9880 -3460 14378 -3260
rect 4750 -3603 4799 -3569
rect 4833 -3603 4871 -3569
rect 4905 -3603 4950 -3569
rect -400 -3870 500 -3670
rect 4750 -3929 4950 -3603
rect 9880 -3670 10080 -3664
rect 8636 -3870 10080 -3670
rect 4750 -3963 4799 -3929
rect 4833 -3963 4871 -3929
rect 4905 -3963 4950 -3929
rect 4750 -4369 4950 -3963
rect 9880 -4060 10080 -3870
rect 14178 -3888 14378 -3460
rect 14560 -3639 14760 -3089
rect 14560 -3673 14605 -3639
rect 14639 -3673 14760 -3639
rect 14560 -3711 14760 -3673
rect 14560 -3745 14605 -3711
rect 14639 -3745 14760 -3711
rect 14560 -3783 14760 -3745
rect 14560 -3817 14605 -3783
rect 14639 -3817 14760 -3783
rect 14560 -3855 14760 -3817
rect 14560 -3889 14605 -3855
rect 14639 -3889 14760 -3855
rect 9880 -4260 14378 -4060
rect 4750 -4403 4799 -4369
rect 4833 -4403 4871 -4369
rect 4905 -4403 4950 -4369
rect -400 -4670 500 -4470
rect 4750 -4729 4950 -4403
rect 9880 -4470 10080 -4464
rect 8636 -4670 10080 -4470
rect 4750 -4763 4799 -4729
rect 4833 -4763 4871 -4729
rect 4905 -4763 4950 -4729
rect 4750 -5169 4950 -4763
rect 9880 -4860 10080 -4670
rect 14178 -4688 14378 -4260
rect 14560 -4439 14760 -3889
rect 14560 -4473 14605 -4439
rect 14639 -4473 14760 -4439
rect 14560 -4511 14760 -4473
rect 14560 -4545 14605 -4511
rect 14639 -4545 14760 -4511
rect 14560 -4583 14760 -4545
rect 14560 -4617 14605 -4583
rect 14639 -4617 14760 -4583
rect 14560 -4655 14760 -4617
rect 14560 -4689 14605 -4655
rect 14639 -4689 14760 -4655
rect 9880 -5060 14378 -4860
rect 4750 -5203 4799 -5169
rect 4833 -5203 4871 -5169
rect 4905 -5203 4950 -5169
rect -400 -5470 500 -5270
rect 4750 -5529 4950 -5203
rect 8636 -5470 10080 -5270
rect 4750 -5563 4799 -5529
rect 4833 -5563 4871 -5529
rect 4905 -5563 4950 -5529
rect 4750 -5606 4950 -5563
rect 9260 -5786 9460 -5470
rect 14178 -5488 14378 -5060
rect 14560 -5239 14760 -4689
rect 14560 -5273 14605 -5239
rect 14639 -5273 14760 -5239
rect 14560 -5311 14760 -5273
rect 14560 -5345 14605 -5311
rect 14639 -5345 14760 -5311
rect 14560 -5383 14760 -5345
rect 14560 -5417 14605 -5383
rect 14639 -5417 14760 -5383
rect 14560 -5455 14760 -5417
rect 14560 -5489 14605 -5455
rect 14639 -5489 14760 -5455
rect 14560 -5590 14760 -5489
<< via1 >>
rect 4760 -256 4940 -76
rect 14570 -256 14750 -76
<< metal2 >>
rect 4750 -66 4950 -60
rect 4750 -76 14766 -66
rect 4750 -256 4760 -76
rect 4940 -256 14570 -76
rect 14750 -256 14766 -76
rect 4750 -266 14766 -256
rect 4750 -272 4950 -266
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR1
timestamp 1713537803
transform 0 1 4572 -1 0 235
box -225 -4562 225 4562
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR2
timestamp 1713537803
transform 0 1 4572 -1 0 -565
box -225 -4562 225 4562
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR3
timestamp 1713537803
transform 0 1 4572 -1 0 -1365
box -225 -4562 225 4562
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR4
timestamp 1713537803
transform 0 1 4572 -1 0 -2165
box -225 -4562 225 4562
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR5
timestamp 1713537803
transform 0 1 4572 -1 0 -2965
box -225 -4562 225 4562
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR6
timestamp 1713537803
transform 0 1 4572 -1 0 -3765
box -225 -4562 225 4562
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR7
timestamp 1713537803
transform 0 1 4572 -1 0 -4565
box -225 -4562 225 4562
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR8
timestamp 1713537803
transform 0 1 4572 -1 0 -5365
box -225 -4562 225 4562
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR9
timestamp 1713537803
transform 0 1 12137 -1 0 235
box -225 -2527 225 2527
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR10
timestamp 1713537803
transform 0 1 12137 -1 0 -565
box -225 -2527 225 2527
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR11
timestamp 1713537803
transform 0 1 12137 -1 0 -1365
box -225 -2527 225 2527
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR12
timestamp 1713537803
transform 0 1 12137 -1 0 -2165
box -225 -2527 225 2527
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR13
timestamp 1713537803
transform 0 1 12137 -1 0 -2965
box -225 -2527 225 2527
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR14
timestamp 1713537803
transform 0 1 12137 -1 0 -3765
box -225 -2527 225 2527
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR15
timestamp 1713537803
transform 0 1 12137 -1 0 -4565
box -225 -2527 225 2527
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR16
timestamp 1713537803
transform 0 1 12137 -1 0 -5365
box -225 -2527 225 2527
<< labels >>
flabel metal1 s 9260 -5786 9460 -5586 0 FreeSans 320 0 0 0 aout
port 1 nsew
flabel metal1 s -400 -5470 -200 -5270 0 FreeSans 320 0 0 0 d7
port 2 nsew
flabel metal1 s -400 -4670 -200 -4470 0 FreeSans 320 0 0 0 d6
port 3 nsew
flabel metal1 s -400 -3870 -200 -3670 0 FreeSans 320 0 0 0 d5
port 4 nsew
flabel metal1 s -400 -3070 -200 -2870 0 FreeSans 320 0 0 0 d4
port 5 nsew
flabel metal1 s -400 -2270 -200 -2070 0 FreeSans 320 0 0 0 d3
port 6 nsew
flabel metal1 s -400 -1470 -200 -1270 0 FreeSans 320 0 0 0 d2
port 7 nsew
flabel metal1 s -400 -670 -200 -470 0 FreeSans 320 0 0 0 d1
port 8 nsew
flabel metal1 s -400 130 -200 330 0 FreeSans 320 0 0 0 d0
port 9 nsew
flabel metal1 s -400 600 -200 800 0 FreeSans 320 0 0 0 GND
port 10 nsew
flabel metal1 s -400 -270 -200 -70 0 FreeSans 320 0 0 0 VSUBS
port 11 nsew
<< properties >>
string GDS_END 45798
string GDS_FILE /home/anton/projects/tt06-grab-bag/gds/tt_um_algofoogle_tt06_grab_bag.gds
string GDS_START 32528
<< end >>
