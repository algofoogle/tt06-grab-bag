magic
tech sky130A
magscale 1 2
timestamp 1713537803
<< locali >>
rect 850 1893 910 1920
rect 850 1859 863 1893
rect 897 1859 910 1893
rect 850 1821 910 1859
rect 850 1787 863 1821
rect 897 1787 910 1821
rect 850 1760 910 1787
rect -30 1663 30 1680
rect -30 1629 -17 1663
rect 17 1629 30 1663
rect -30 1591 30 1629
rect -30 1557 -17 1591
rect 17 1557 30 1591
rect -30 1540 30 1557
<< viali >>
rect 863 1859 897 1893
rect 863 1787 897 1821
rect -17 1629 17 1663
rect -17 1557 17 1591
<< metal1 >>
rect 130 2400 750 2460
rect 690 2060 750 2400
rect 930 2060 990 2066
rect 670 2056 990 2060
rect 670 2004 934 2056
rect 986 2004 990 2056
rect 670 2000 990 2004
rect 930 1994 990 2000
rect 1020 1940 1220 2810
rect 740 1893 1220 1940
rect 740 1859 863 1893
rect 897 1859 1220 1893
rect 740 1821 1220 1859
rect 740 1787 863 1821
rect 897 1787 1220 1821
rect -410 1663 140 1710
rect -410 1629 -17 1663
rect 17 1629 140 1663
rect -410 1591 140 1629
rect -410 1557 -17 1591
rect 17 1557 140 1591
rect -410 1510 140 1557
rect 180 1510 700 1760
rect 740 1740 1220 1787
rect 930 1590 990 1596
rect 1020 1590 1220 1660
rect 930 1586 1220 1590
rect 930 1534 934 1586
rect 986 1534 1220 1586
rect 930 1530 1220 1534
rect 930 1524 990 1530
rect 420 860 480 1510
rect 1020 1460 1220 1530
rect 930 1140 990 1146
rect 670 1136 990 1140
rect 670 1084 934 1136
rect 986 1084 990 1136
rect 670 1080 990 1084
rect 590 860 650 866
rect 420 856 650 860
rect 420 804 594 856
rect 646 804 650 856
rect 420 800 650 804
rect 590 794 650 800
rect 690 730 750 1080
rect 930 1074 990 1080
rect 1020 860 1220 930
rect 794 856 1220 860
rect 794 804 804 856
rect 856 804 1220 856
rect 794 800 1220 804
rect 1020 730 1220 800
rect 120 670 750 730
<< via1 >>
rect 934 2004 986 2056
rect 934 1534 986 1586
rect 934 1084 986 1136
rect 594 804 646 856
rect 804 804 856 856
<< metal2 >>
rect 924 2056 996 2060
rect 924 2004 934 2056
rect 986 2004 996 2056
rect 924 2000 996 2004
rect 930 1590 990 2000
rect 924 1586 996 1590
rect 924 1534 934 1586
rect 986 1534 996 1586
rect 924 1530 996 1534
rect 930 1140 990 1530
rect 924 1136 996 1140
rect 924 1084 934 1136
rect 986 1084 996 1136
rect 924 1080 996 1084
rect 800 860 860 866
rect 584 856 860 860
rect 584 804 594 856
rect 646 804 804 856
rect 856 804 860 856
rect 584 800 860 804
rect 800 794 860 800
use sky130_fd_pr__pfet_01v8_UGACMG  XM1
timestamp 1713537803
transform 1 0 158 0 1 1566
box -211 -1019 211 1019
use sky130_fd_pr__nfet_01v8_PWNS5P  XM2
timestamp 1713537803
transform 1 0 721 0 1 1570
box -201 -600 201 600
<< labels >>
flabel metal1 s -410 1510 -210 1710 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 s 1020 2610 1220 2810 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 s 1020 1460 1220 1660 0 FreeSans 1600 0 0 0 A
port 3 nsew
flabel metal1 s 1020 730 1220 930 0 FreeSans 1600 0 0 0 Y
port 4 nsew
<< properties >>
string GDS_END 67878
string GDS_FILE /home/anton/projects/tt06-grab-bag/gds/tt_um_algofoogle_tt06_grab_bag.gds
string GDS_START 64338
<< end >>
