magic
tech sky130A
magscale 1 2
timestamp 1712241802
<< viali >>
rect 850 1760 910 1920
rect -30 1540 30 1680
<< metal1 >>
rect 130 2400 750 2460
rect 690 2060 750 2400
rect 930 2060 990 2066
rect 670 2000 930 2060
rect 930 1994 990 2000
rect 1020 1940 1220 2810
rect 740 1920 1220 1940
rect 740 1760 850 1920
rect 910 1760 1220 1920
rect -410 1680 140 1710
rect -410 1540 -30 1680
rect 30 1540 140 1680
rect -410 1510 140 1540
rect 180 1510 700 1760
rect 740 1740 1220 1760
rect 930 1590 990 1596
rect 1020 1590 1220 1660
rect 990 1530 1220 1590
rect 930 1524 990 1530
rect 420 860 480 1510
rect 1020 1460 1220 1530
rect 930 1140 990 1146
rect 670 1080 930 1140
rect 590 860 650 866
rect 420 800 590 860
rect 590 794 650 800
rect 690 730 750 1080
rect 930 1074 990 1080
rect 1020 860 1220 930
rect 794 800 800 860
rect 860 800 1220 860
rect 1020 730 1220 800
rect 120 670 750 730
<< via1 >>
rect 930 2000 990 2060
rect 930 1530 990 1590
rect 930 1080 990 1140
rect 590 800 650 860
rect 800 800 860 860
<< metal2 >>
rect 924 2000 930 2060
rect 990 2000 996 2060
rect 930 1590 990 2000
rect 924 1530 930 1590
rect 990 1530 996 1590
rect 930 1140 990 1530
rect 924 1080 930 1140
rect 990 1080 996 1140
rect 800 860 860 866
rect 584 800 590 860
rect 650 800 800 860
rect 800 794 860 800
use sky130_fd_pr__pfet_01v8_UGACMG  XM1
timestamp 1712240008
transform 1 0 158 0 1 1566
box -211 -1019 211 1019
use sky130_fd_pr__nfet_01v8_PWNS5P  XM2
timestamp 1712240008
transform 1 0 721 0 1 1570
box -211 -610 211 610
<< labels >>
flabel metal1 -410 1510 -210 1710 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 1020 1460 1220 1660 0 FreeSans 1280 0 0 0 A
port 2 nsew
flabel metal1 1020 730 1220 930 0 FreeSans 1280 0 0 0 Y
port 3 nsew
flabel metal1 1020 2610 1220 2810 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
<< end >>
