`default_nettype none

// just a stub to keep the Tiny Tapeout tools happy

module tt_um_algofoogle_tt06_grab_bag(
    input  wire       VGND,
    input  wire       VPWR,
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    inout  wire [7:0] ua, // analog pins
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    wire Y; // Inverter output -- goes to multiple places.
    assign uo_out[0] = Y;
    assign ua[0] = Y;

    inverter inverter(
        .VDD    (VPWR),
        .VSS    (VGND),
        .A      (ui_in[0]),
        .Y      (Y)
    );

    // Tie other digital outputs to VGND, so they don't float:
    assign uo_out[7:1] = {7{VGND}};
    assign uio_out[7:0] = {8{VGND}};
    assign uio_oe[7:0] = {8{VGND}};

endmodule

