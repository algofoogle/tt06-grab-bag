magic
tech sky130A
magscale 1 2
timestamp 1713380768
<< viali >>
rect 4772 380 4932 448
rect 14586 110 14658 362
rect 4772 20 4932 88
rect 4772 -420 4932 -352
rect 14586 -690 14658 -438
rect 4772 -780 4932 -712
rect 4772 -1220 4932 -1152
rect 14586 -1490 14658 -1238
rect 4772 -1580 4932 -1512
rect 4772 -2020 4932 -1952
rect 14586 -2290 14658 -2038
rect 4772 -2380 4932 -2312
rect 4772 -2820 4932 -2752
rect 14586 -3090 14658 -2838
rect 4772 -3180 4932 -3112
rect 4772 -3620 4932 -3552
rect 14586 -3890 14658 -3638
rect 4772 -3980 4932 -3912
rect 4772 -4420 4932 -4352
rect 14586 -4690 14658 -4438
rect 4772 -4780 4932 -4712
rect 4772 -5220 4932 -5152
rect 14586 -5490 14658 -5238
rect 4772 -5580 4932 -5512
<< metal1 >>
rect -400 600 14380 800
rect 4750 448 4950 496
rect 4750 380 4772 448
rect 4932 380 4950 448
rect -400 130 500 330
rect 4750 88 4950 380
rect 9880 330 10080 336
rect 8636 130 10080 330
rect 4750 20 4772 88
rect 4932 20 4950 88
rect 4750 -66 4950 20
rect 9880 -60 10080 130
rect 14180 118 14380 600
rect 14560 362 14760 398
rect 14560 110 14586 362
rect 14658 110 14760 362
rect 4744 -70 4750 -66
rect -400 -266 4750 -70
rect 4950 -266 4956 -66
rect 9880 -260 14378 -60
rect -400 -270 4950 -266
rect 4750 -352 4950 -270
rect 4750 -420 4772 -352
rect 4932 -420 4950 -352
rect -400 -670 500 -470
rect 4750 -712 4950 -420
rect 9880 -470 10080 -464
rect 8636 -670 10080 -470
rect 4750 -780 4772 -712
rect 4932 -780 4950 -712
rect 4750 -1152 4950 -780
rect 9880 -860 10080 -670
rect 14178 -688 14378 -260
rect 14560 -66 14760 110
rect 14560 -438 14760 -266
rect 14560 -690 14586 -438
rect 14658 -690 14760 -438
rect 9880 -1060 14378 -860
rect 4750 -1220 4772 -1152
rect 4932 -1220 4950 -1152
rect -400 -1470 500 -1270
rect 4750 -1512 4950 -1220
rect 9880 -1270 10080 -1264
rect 8636 -1470 10080 -1270
rect 4750 -1580 4772 -1512
rect 4932 -1580 4950 -1512
rect 4750 -1952 4950 -1580
rect 9880 -1660 10080 -1470
rect 14178 -1488 14378 -1060
rect 14560 -1238 14760 -690
rect 14560 -1490 14586 -1238
rect 14658 -1490 14760 -1238
rect 9880 -1860 14378 -1660
rect 4750 -2020 4772 -1952
rect 4932 -2020 4950 -1952
rect -400 -2270 500 -2070
rect 4750 -2312 4950 -2020
rect 9880 -2070 10080 -2064
rect 8636 -2270 10080 -2070
rect 4750 -2380 4772 -2312
rect 4932 -2380 4950 -2312
rect 4750 -2752 4950 -2380
rect 9880 -2460 10080 -2270
rect 14178 -2288 14378 -1860
rect 14560 -2038 14760 -1490
rect 14560 -2290 14586 -2038
rect 14658 -2290 14760 -2038
rect 9880 -2660 14378 -2460
rect 4750 -2820 4772 -2752
rect 4932 -2820 4950 -2752
rect -400 -3070 500 -2870
rect 4750 -3112 4950 -2820
rect 9880 -2870 10080 -2864
rect 8636 -3070 10080 -2870
rect 4750 -3180 4772 -3112
rect 4932 -3180 4950 -3112
rect 4750 -3552 4950 -3180
rect 9880 -3260 10080 -3070
rect 14178 -3088 14378 -2660
rect 14560 -2838 14760 -2290
rect 14560 -3090 14586 -2838
rect 14658 -3090 14760 -2838
rect 9880 -3460 14378 -3260
rect 4750 -3620 4772 -3552
rect 4932 -3620 4950 -3552
rect -400 -3870 500 -3670
rect 4750 -3912 4950 -3620
rect 9880 -3670 10080 -3664
rect 8636 -3870 10080 -3670
rect 4750 -3980 4772 -3912
rect 4932 -3980 4950 -3912
rect 4750 -4352 4950 -3980
rect 9880 -4060 10080 -3870
rect 14178 -3888 14378 -3460
rect 14560 -3638 14760 -3090
rect 14560 -3890 14586 -3638
rect 14658 -3890 14760 -3638
rect 9880 -4260 14378 -4060
rect 4750 -4420 4772 -4352
rect 4932 -4420 4950 -4352
rect -400 -4670 500 -4470
rect 4750 -4712 4950 -4420
rect 9880 -4470 10080 -4464
rect 8636 -4670 10080 -4470
rect 4750 -4780 4772 -4712
rect 4932 -4780 4950 -4712
rect 4750 -5152 4950 -4780
rect 9880 -4860 10080 -4670
rect 14178 -4688 14378 -4260
rect 14560 -4438 14760 -3890
rect 14560 -4690 14586 -4438
rect 14658 -4690 14760 -4438
rect 9880 -5060 14378 -4860
rect 4750 -5220 4772 -5152
rect 4932 -5220 4950 -5152
rect -400 -5470 500 -5270
rect 4750 -5512 4950 -5220
rect 8636 -5470 10080 -5270
rect 4750 -5580 4772 -5512
rect 4932 -5580 4950 -5512
rect 4750 -5606 4950 -5580
rect 9260 -5786 9460 -5470
rect 14178 -5488 14378 -5060
rect 14560 -5238 14760 -4690
rect 14560 -5490 14586 -5238
rect 14658 -5490 14760 -5238
rect 14560 -5590 14760 -5490
<< via1 >>
rect 4750 -266 4950 -66
rect 14560 -266 14760 -66
<< metal2 >>
rect 4750 -66 4950 -60
rect 4950 -266 14560 -66
rect 14760 -266 14766 -66
rect 4750 -272 4950 -266
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR1
timestamp 1713376360
transform 0 1 4572 -1 0 235
box -235 -4572 235 4572
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR2
timestamp 1713376360
transform 0 1 4572 -1 0 -565
box -235 -4572 235 4572
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR3
timestamp 1713376360
transform 0 1 4572 -1 0 -1365
box -235 -4572 235 4572
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR4
timestamp 1713376360
transform 0 1 4572 -1 0 -2165
box -235 -4572 235 4572
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR5
timestamp 1713376360
transform 0 1 4572 -1 0 -2965
box -235 -4572 235 4572
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR6
timestamp 1713376360
transform 0 1 4572 -1 0 -3765
box -235 -4572 235 4572
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR7
timestamp 1713376360
transform 0 1 4572 -1 0 -4565
box -235 -4572 235 4572
use sky130_fd_pr__res_high_po_0p69_5ANSK2  XR8
timestamp 1713376360
transform 0 1 4572 -1 0 -5365
box -235 -4572 235 4572
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR9
timestamp 1713376360
transform 0 1 12137 -1 0 235
box -235 -2537 235 2537
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR10
timestamp 1713376360
transform 0 1 12137 -1 0 -565
box -235 -2537 235 2537
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR11
timestamp 1713376360
transform 0 1 12137 -1 0 -1365
box -235 -2537 235 2537
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR12
timestamp 1713376360
transform 0 1 12137 -1 0 -2165
box -235 -2537 235 2537
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR13
timestamp 1713376360
transform 0 1 12137 -1 0 -2965
box -235 -2537 235 2537
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR14
timestamp 1713376360
transform 0 1 12137 -1 0 -3765
box -235 -2537 235 2537
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR15
timestamp 1713376360
transform 0 1 12137 -1 0 -4565
box -235 -2537 235 2537
use sky130_fd_pr__res_high_po_0p69_5G96UM  XR16
timestamp 1713376360
transform 0 1 12137 -1 0 -5365
box -235 -2537 235 2537
<< labels >>
flabel metal1 -400 130 -200 330 0 FreeSans 256 0 0 0 {d\[0\]}
port 8 nsew
flabel metal1 -400 -670 -200 -470 0 FreeSans 256 0 0 0 {d\[1\]}
port 7 nsew
flabel metal1 -400 -1470 -200 -1270 0 FreeSans 256 0 0 0 {d\[2\]}
port 6 nsew
flabel metal1 -400 -2270 -200 -2070 0 FreeSans 256 0 0 0 {d\[3\]}
port 5 nsew
flabel metal1 -400 -3070 -200 -2870 0 FreeSans 256 0 0 0 {d\[4\]}
port 4 nsew
flabel metal1 -400 -3870 -200 -3670 0 FreeSans 256 0 0 0 {d\[5\]}
port 3 nsew
flabel metal1 -400 -4670 -200 -4470 0 FreeSans 256 0 0 0 {d\[6\]}
port 2 nsew
flabel metal1 -400 -5470 -200 -5270 0 FreeSans 256 0 0 0 {d\[7\]}
port 1 nsew
flabel metal1 -400 600 -200 800 0 FreeSans 256 0 0 0 GND
port 9 nsew
flabel metal1 -400 -270 -200 -70 0 FreeSans 256 0 0 0 VSUBS
port 10 nsew
flabel metal1 9260 -5786 9460 -5586 0 FreeSans 256 0 0 0 aout
port 0 nsew
<< end >>
