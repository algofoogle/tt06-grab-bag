magic
tech sky130A
magscale 1 2
timestamp 1713545776
<< viali >>
rect 4629 15113 4663 15147
rect 5181 15113 5215 15147
rect 6193 15113 6227 15147
rect 6653 15113 6687 15147
rect 7573 15113 7607 15147
rect 8493 15113 8527 15147
rect 9137 15113 9171 15147
rect 9597 15113 9631 15147
rect 10517 15113 10551 15147
rect 11069 15113 11103 15147
rect 21465 15113 21499 15147
rect 16129 15045 16163 15079
rect 21281 15045 21315 15079
rect 22201 15045 22235 15079
rect 22845 15045 22879 15079
rect 16589 14977 16623 15011
rect 16681 14977 16715 15011
rect 2329 14909 2363 14943
rect 4813 14909 4847 14943
rect 6009 14909 6043 14943
rect 7757 14909 7791 14943
rect 7849 14909 7883 14943
rect 8033 14909 8067 14943
rect 8953 14909 8987 14943
rect 10701 14909 10735 14943
rect 13185 14909 13219 14943
rect 13553 14909 13587 14943
rect 13829 14909 13863 14943
rect 17785 14909 17819 14943
rect 18705 14909 18739 14943
rect 19441 14909 19475 14943
rect 20085 14909 20119 14943
rect 20361 14909 20395 14943
rect 20913 14909 20947 14943
rect 21741 14909 21775 14943
rect 22017 14909 22051 14943
rect 22385 14909 22419 14943
rect 23029 14909 23063 14943
rect 5457 14841 5491 14875
rect 6929 14841 6963 14875
rect 8769 14841 8803 14875
rect 9873 14841 9907 14875
rect 11345 14841 11379 14875
rect 16497 14841 16531 14875
rect 2973 14773 3007 14807
rect 7941 14773 7975 14807
rect 13093 14773 13127 14807
rect 17969 14773 18003 14807
rect 18889 14773 18923 14807
rect 19257 14773 19291 14807
rect 19901 14773 19935 14807
rect 20177 14773 20211 14807
rect 20729 14773 20763 14807
rect 21833 14773 21867 14807
rect 2237 14569 2271 14603
rect 2421 14569 2455 14603
rect 5641 14569 5675 14603
rect 6193 14569 6227 14603
rect 6745 14569 6779 14603
rect 10241 14569 10275 14603
rect 10425 14569 10459 14603
rect 11069 14569 11103 14603
rect 16589 14569 16623 14603
rect 16957 14569 16991 14603
rect 18061 14569 18095 14603
rect 18429 14569 18463 14603
rect 21097 14569 21131 14603
rect 21557 14569 21591 14603
rect 23029 14569 23063 14603
rect 6101 14501 6135 14535
rect 10977 14501 11011 14535
rect 21894 14501 21928 14535
rect 1124 14433 1158 14467
rect 2513 14433 2547 14467
rect 2605 14433 2639 14467
rect 2872 14433 2906 14467
rect 4261 14433 4295 14467
rect 4528 14433 4562 14467
rect 6561 14433 6595 14467
rect 6653 14433 6687 14467
rect 6837 14433 6871 14467
rect 7113 14433 7147 14467
rect 7573 14433 7607 14467
rect 8217 14433 8251 14467
rect 9505 14433 9539 14467
rect 10333 14433 10367 14467
rect 10609 14433 10643 14467
rect 12081 14433 12115 14467
rect 12357 14433 12391 14467
rect 12613 14433 12647 14467
rect 13829 14433 13863 14467
rect 14096 14433 14130 14467
rect 15669 14433 15703 14467
rect 16497 14433 16531 14467
rect 17141 14433 17175 14467
rect 17693 14433 17727 14467
rect 19165 14433 19199 14467
rect 19257 14433 19291 14467
rect 19717 14433 19751 14467
rect 19984 14433 20018 14467
rect 21373 14433 21407 14467
rect 21649 14433 21683 14467
rect 857 14365 891 14399
rect 7665 14365 7699 14399
rect 8125 14365 8159 14399
rect 9321 14365 9355 14399
rect 9689 14365 9723 14399
rect 9781 14365 9815 14399
rect 11345 14365 11379 14399
rect 15485 14365 15519 14399
rect 15945 14365 15979 14399
rect 16773 14365 16807 14399
rect 17417 14365 17451 14399
rect 17969 14365 18003 14399
rect 18521 14365 18555 14399
rect 18705 14365 18739 14399
rect 18981 14365 19015 14399
rect 6929 14297 6963 14331
rect 7941 14297 7975 14331
rect 10057 14297 10091 14331
rect 12265 14297 12299 14331
rect 15853 14297 15887 14331
rect 17509 14297 17543 14331
rect 3985 14229 4019 14263
rect 6377 14229 6411 14263
rect 8493 14229 8527 14263
rect 10793 14229 10827 14263
rect 11253 14229 11287 14263
rect 11345 14229 11379 14263
rect 13737 14229 13771 14263
rect 15209 14229 15243 14263
rect 16129 14229 16163 14263
rect 17325 14229 17359 14263
rect 17877 14229 17911 14263
rect 19625 14229 19659 14263
rect 1869 14025 1903 14059
rect 2881 14025 2915 14059
rect 7849 14025 7883 14059
rect 8493 14025 8527 14059
rect 9045 14025 9079 14059
rect 9781 14025 9815 14059
rect 10977 14025 11011 14059
rect 14565 14025 14599 14059
rect 16313 14025 16347 14059
rect 17601 14025 17635 14059
rect 18245 14025 18279 14059
rect 18889 14025 18923 14059
rect 20085 14025 20119 14059
rect 6377 13957 6411 13991
rect 10609 13957 10643 13991
rect 11437 13957 11471 13991
rect 13737 13957 13771 13991
rect 8861 13889 8895 13923
rect 10333 13889 10367 13923
rect 11069 13889 11103 13923
rect 15393 13889 15427 13923
rect 15669 13889 15703 13923
rect 16773 13889 16807 13923
rect 16957 13889 16991 13923
rect 18337 13889 18371 13923
rect 19441 13889 19475 13923
rect 19625 13889 19659 13923
rect 20637 13889 20671 13923
rect 1869 13821 1903 13855
rect 2053 13821 2087 13855
rect 2145 13821 2179 13855
rect 2329 13821 2363 13855
rect 2697 13821 2731 13855
rect 6285 13821 6319 13855
rect 7849 13821 7883 13855
rect 8033 13821 8067 13855
rect 8401 13821 8435 13855
rect 8677 13821 8711 13855
rect 8953 13821 8987 13855
rect 10241 13821 10275 13855
rect 10701 13821 10735 13855
rect 10885 13821 10919 13855
rect 11161 13821 11195 13855
rect 11529 13821 11563 13855
rect 11713 13821 11747 13855
rect 13093 13821 13127 13855
rect 13185 13821 13219 13855
rect 13277 13821 13311 13855
rect 13829 13821 13863 13855
rect 14013 13821 14047 13855
rect 14749 13821 14783 13855
rect 17325 13821 17359 13855
rect 17417 13821 17451 13855
rect 17877 13821 17911 13855
rect 18061 13821 18095 13855
rect 18889 13821 18923 13855
rect 19073 13821 19107 13855
rect 19717 13821 19751 13855
rect 20821 13821 20855 13855
rect 6040 13753 6074 13787
rect 6561 13753 6595 13787
rect 9413 13753 9447 13787
rect 9597 13753 9631 13787
rect 2513 13685 2547 13719
rect 4905 13685 4939 13719
rect 11621 13685 11655 13719
rect 16681 13685 16715 13719
rect 17141 13685 17175 13719
rect 18705 13685 18739 13719
rect 7849 13481 7883 13515
rect 17877 13481 17911 13515
rect 18429 13481 18463 13515
rect 18521 13481 18555 13515
rect 18889 13481 18923 13515
rect 19165 13481 19199 13515
rect 21557 13481 21591 13515
rect 1869 13413 1903 13447
rect 2085 13413 2119 13447
rect 2596 13413 2630 13447
rect 10425 13413 10459 13447
rect 16129 13413 16163 13447
rect 21894 13413 21928 13447
rect 2329 13345 2363 13379
rect 6285 13345 6319 13379
rect 6377 13345 6411 13379
rect 7665 13345 7699 13379
rect 7849 13345 7883 13379
rect 8769 13345 8803 13379
rect 10149 13345 10183 13379
rect 10333 13345 10367 13379
rect 10609 13345 10643 13379
rect 11161 13345 11195 13379
rect 16313 13345 16347 13379
rect 16865 13345 16899 13379
rect 17141 13345 17175 13379
rect 17785 13345 17819 13379
rect 18061 13345 18095 13379
rect 19257 13345 19291 13379
rect 19993 13345 20027 13379
rect 21373 13345 21407 13379
rect 11069 13277 11103 13311
rect 11713 13277 11747 13311
rect 16589 13277 16623 13311
rect 18337 13277 18371 13311
rect 21649 13277 21683 13311
rect 11437 13209 11471 13243
rect 16497 13209 16531 13243
rect 2053 13141 2087 13175
rect 2237 13141 2271 13175
rect 3709 13141 3743 13175
rect 6101 13141 6135 13175
rect 6469 13141 6503 13175
rect 8953 13141 8987 13175
rect 10241 13141 10275 13175
rect 10793 13141 10827 13175
rect 16681 13141 16715 13175
rect 17049 13141 17083 13175
rect 17601 13141 17635 13175
rect 20177 13141 20211 13175
rect 23029 13141 23063 13175
rect 1685 12937 1719 12971
rect 1869 12937 1903 12971
rect 2329 12937 2363 12971
rect 3341 12937 3375 12971
rect 5917 12937 5951 12971
rect 9229 12937 9263 12971
rect 13645 12937 13679 12971
rect 16589 12937 16623 12971
rect 18429 12937 18463 12971
rect 21649 12937 21683 12971
rect 1317 12869 1351 12903
rect 6285 12869 6319 12903
rect 12909 12869 12943 12903
rect 19625 12869 19659 12903
rect 3525 12801 3559 12835
rect 5181 12801 5215 12835
rect 5365 12801 5399 12835
rect 9597 12801 9631 12835
rect 10609 12801 10643 12835
rect 10885 12801 10919 12835
rect 11069 12801 11103 12835
rect 11253 12801 11287 12835
rect 13277 12801 13311 12835
rect 13369 12801 13403 12835
rect 13829 12801 13863 12835
rect 14197 12801 14231 12835
rect 19533 12801 19567 12835
rect 22201 12801 22235 12835
rect 1225 12733 1259 12767
rect 1409 12733 1443 12767
rect 1961 12733 1995 12767
rect 2145 12733 2179 12767
rect 2421 12733 2455 12767
rect 2605 12733 2639 12767
rect 2697 12733 2731 12767
rect 2835 12733 2869 12767
rect 3249 12733 3283 12767
rect 3433 12733 3467 12767
rect 5457 12733 5491 12767
rect 6101 12733 6135 12767
rect 6193 12733 6227 12767
rect 6377 12733 6411 12767
rect 6561 12733 6595 12767
rect 6745 12733 6779 12767
rect 6837 12733 6871 12767
rect 9413 12733 9447 12767
rect 9689 12733 9723 12767
rect 10793 12733 10827 12767
rect 10977 12733 11011 12767
rect 11437 12733 11471 12767
rect 11621 12733 11655 12767
rect 11713 12733 11747 12767
rect 13093 12733 13127 12767
rect 13921 12733 13955 12767
rect 14289 12733 14323 12767
rect 14473 12733 14507 12767
rect 16405 12733 16439 12767
rect 16681 12733 16715 12767
rect 18245 12733 18279 12767
rect 18521 12733 18555 12767
rect 19257 12733 19291 12767
rect 19809 12733 19843 12767
rect 20177 12733 20211 12767
rect 20444 12733 20478 12767
rect 22109 12733 22143 12767
rect 23029 12733 23063 12767
rect 1501 12665 1535 12699
rect 3781 12665 3815 12699
rect 6653 12665 6687 12699
rect 7104 12665 7138 12699
rect 22017 12665 22051 12699
rect 1701 12597 1735 12631
rect 3065 12597 3099 12631
rect 4905 12597 4939 12631
rect 5825 12597 5859 12631
rect 8217 12597 8251 12631
rect 14657 12597 14691 12631
rect 16221 12597 16255 12631
rect 18061 12597 18095 12631
rect 21557 12597 21591 12631
rect 22845 12597 22879 12631
rect 2053 12393 2087 12427
rect 7481 12393 7515 12427
rect 12173 12393 12207 12427
rect 14013 12393 14047 12427
rect 1869 12325 1903 12359
rect 2789 12325 2823 12359
rect 17242 12325 17276 12359
rect 1685 12257 1719 12291
rect 1961 12257 1995 12291
rect 2329 12257 2363 12291
rect 2513 12257 2547 12291
rect 3341 12257 3375 12291
rect 4445 12257 4479 12291
rect 4813 12257 4847 12291
rect 5181 12257 5215 12291
rect 5457 12257 5491 12291
rect 7665 12257 7699 12291
rect 8024 12257 8058 12291
rect 9689 12257 9723 12291
rect 10609 12257 10643 12291
rect 10793 12257 10827 12291
rect 10969 12257 11003 12291
rect 11437 12257 11471 12291
rect 12357 12257 12391 12291
rect 12449 12257 12483 12291
rect 12541 12257 12575 12291
rect 13001 12257 13035 12291
rect 13461 12257 13495 12291
rect 13645 12257 13679 12291
rect 13737 12257 13771 12291
rect 13853 12257 13887 12291
rect 15761 12257 15795 12291
rect 17509 12257 17543 12291
rect 18429 12257 18463 12291
rect 18613 12257 18647 12291
rect 19818 12257 19852 12291
rect 20085 12257 20119 12291
rect 2237 12189 2271 12223
rect 2421 12189 2455 12223
rect 3065 12189 3099 12223
rect 5825 12189 5859 12223
rect 6101 12189 6135 12223
rect 7757 12189 7791 12223
rect 9505 12189 9539 12223
rect 9965 12189 9999 12223
rect 12633 12189 12667 12223
rect 12909 12189 12943 12223
rect 13369 12189 13403 12223
rect 1777 12121 1811 12155
rect 5273 12121 5307 12155
rect 5365 12121 5399 12155
rect 9873 12121 9907 12155
rect 11161 12121 11195 12155
rect 2881 12053 2915 12087
rect 4629 12053 4663 12087
rect 4997 12053 5031 12087
rect 5641 12053 5675 12087
rect 9137 12053 9171 12087
rect 10701 12053 10735 12087
rect 11345 12053 11379 12087
rect 15945 12053 15979 12087
rect 16129 12053 16163 12087
rect 18521 12053 18555 12087
rect 18705 12053 18739 12087
rect 2145 11849 2179 11883
rect 4629 11849 4663 11883
rect 5273 11849 5307 11883
rect 11253 11849 11287 11883
rect 13553 11849 13587 11883
rect 14473 11849 14507 11883
rect 16221 11849 16255 11883
rect 17417 11849 17451 11883
rect 18337 11849 18371 11883
rect 18705 11849 18739 11883
rect 4537 11781 4571 11815
rect 14289 11781 14323 11815
rect 5549 11713 5583 11747
rect 5733 11713 5767 11747
rect 10885 11713 10919 11747
rect 10977 11713 11011 11747
rect 11437 11713 11471 11747
rect 11621 11713 11655 11747
rect 15301 11713 15335 11747
rect 16865 11713 16899 11747
rect 21189 11713 21223 11747
rect 1593 11645 1627 11679
rect 1777 11645 1811 11679
rect 2329 11645 2363 11679
rect 2513 11645 2547 11679
rect 3249 11645 3283 11679
rect 3525 11645 3559 11679
rect 4353 11645 4387 11679
rect 4813 11645 4847 11679
rect 5089 11645 5123 11679
rect 5457 11645 5491 11679
rect 5641 11645 5675 11679
rect 6193 11645 6227 11679
rect 10517 11645 10551 11679
rect 10793 11645 10827 11679
rect 11069 11645 11103 11679
rect 11529 11645 11563 11679
rect 11713 11645 11747 11679
rect 13737 11645 13771 11679
rect 13829 11645 13863 11679
rect 14105 11645 14139 11679
rect 14197 11645 14231 11679
rect 14933 11645 14967 11679
rect 15117 11645 15151 11679
rect 15393 11645 15427 11679
rect 15945 11645 15979 11679
rect 16589 11645 16623 11679
rect 18153 11645 18187 11679
rect 18981 11645 19015 11679
rect 19073 11645 19107 11679
rect 19165 11645 19199 11679
rect 19349 11645 19383 11679
rect 20821 11645 20855 11679
rect 6653 11577 6687 11611
rect 10149 11577 10183 11611
rect 10333 11577 10367 11611
rect 13921 11577 13955 11611
rect 14657 11577 14691 11611
rect 17325 11577 17359 11611
rect 21434 11577 21468 11611
rect 1685 11509 1719 11543
rect 4905 11509 4939 11543
rect 6101 11509 6135 11543
rect 6745 11509 6779 11543
rect 10609 11509 10643 11543
rect 14457 11509 14491 11543
rect 15025 11509 15059 11543
rect 16129 11509 16163 11543
rect 16681 11509 16715 11543
rect 21005 11509 21039 11543
rect 22569 11509 22603 11543
rect 5549 11305 5583 11339
rect 6009 11305 6043 11339
rect 7113 11305 7147 11339
rect 7941 11305 7975 11339
rect 8762 11305 8796 11339
rect 10609 11305 10643 11339
rect 11069 11305 11103 11339
rect 14105 11305 14139 11339
rect 14289 11305 14323 11339
rect 18889 11305 18923 11339
rect 20269 11305 20303 11339
rect 6285 11237 6319 11271
rect 6745 11237 6779 11271
rect 8125 11237 8159 11271
rect 8677 11237 8711 11271
rect 15669 11237 15703 11271
rect 15853 11237 15887 11271
rect 18521 11237 18555 11271
rect 20177 11237 20211 11271
rect 21526 11237 21560 11271
rect 1492 11169 1526 11203
rect 3433 11169 3467 11203
rect 3985 11169 4019 11203
rect 4353 11169 4387 11203
rect 4813 11169 4847 11203
rect 5273 11169 5307 11203
rect 5365 11169 5399 11203
rect 6377 11169 6411 11203
rect 8585 11169 8619 11203
rect 8861 11169 8895 11203
rect 9505 11169 9539 11203
rect 10425 11169 10459 11203
rect 11253 11169 11287 11203
rect 11621 11169 11655 11203
rect 13093 11169 13127 11203
rect 14013 11169 14047 11203
rect 14197 11169 14231 11203
rect 14473 11169 14507 11203
rect 16129 11169 16163 11203
rect 17601 11169 17635 11203
rect 17877 11169 17911 11203
rect 18061 11169 18095 11203
rect 18429 11169 18463 11203
rect 18705 11169 18739 11203
rect 20913 11169 20947 11203
rect 21097 11169 21131 11203
rect 21281 11169 21315 11203
rect 1225 11101 1259 11135
rect 4629 11101 4663 11135
rect 8493 11101 8527 11135
rect 11529 11101 11563 11135
rect 11897 11101 11931 11135
rect 13369 11101 13403 11135
rect 15117 11101 15151 11135
rect 15393 11101 15427 11135
rect 16221 11101 16255 11135
rect 17325 11101 17359 11135
rect 17969 11101 18003 11135
rect 18153 11101 18187 11135
rect 18337 11101 18371 11135
rect 19993 11101 20027 11135
rect 20729 11101 20763 11135
rect 2605 11033 2639 11067
rect 3893 11033 3927 11067
rect 5181 11033 5215 11067
rect 7297 11033 7331 11067
rect 11437 11033 11471 11067
rect 20637 11033 20671 11067
rect 3249 10965 3283 10999
rect 4077 10965 4111 10999
rect 4445 10965 4479 10999
rect 4537 10965 4571 10999
rect 8125 10965 8159 10999
rect 9321 10965 9355 10999
rect 15485 10965 15519 10999
rect 22661 10965 22695 10999
rect 1869 10761 1903 10795
rect 3985 10761 4019 10795
rect 6745 10761 6779 10795
rect 8401 10761 8435 10795
rect 9045 10761 9079 10795
rect 10885 10761 10919 10795
rect 11713 10761 11747 10795
rect 12725 10761 12759 10795
rect 14381 10761 14415 10795
rect 16313 10761 16347 10795
rect 17325 10761 17359 10795
rect 18889 10761 18923 10795
rect 19625 10761 19659 10795
rect 19901 10761 19935 10795
rect 20269 10761 20303 10795
rect 20913 10761 20947 10795
rect 9137 10693 9171 10727
rect 12081 10693 12115 10727
rect 12449 10693 12483 10727
rect 13553 10693 13587 10727
rect 14933 10693 14967 10727
rect 17601 10693 17635 10727
rect 1777 10625 1811 10659
rect 4905 10625 4939 10659
rect 5273 10625 5307 10659
rect 6285 10625 6319 10659
rect 8953 10625 8987 10659
rect 11345 10625 11379 10659
rect 15393 10625 15427 10659
rect 16681 10625 16715 10659
rect 21557 10625 21591 10659
rect 1961 10557 1995 10591
rect 2053 10557 2087 10591
rect 3985 10557 4019 10591
rect 4353 10557 4387 10591
rect 4445 10557 4479 10591
rect 4629 10557 4663 10591
rect 4813 10557 4847 10591
rect 5641 10557 5675 10591
rect 6561 10557 6595 10591
rect 8631 10557 8665 10591
rect 8769 10557 8803 10591
rect 8861 10557 8895 10591
rect 9228 10535 9262 10569
rect 9505 10557 9539 10591
rect 11069 10557 11103 10591
rect 11253 10557 11287 10591
rect 11437 10557 11471 10591
rect 11621 10557 11655 10591
rect 11897 10557 11931 10591
rect 12173 10557 12207 10591
rect 12633 10557 12667 10591
rect 13001 10557 13035 10591
rect 13093 10557 13127 10591
rect 13185 10557 13219 10591
rect 13369 10557 13403 10591
rect 13737 10557 13771 10591
rect 13921 10557 13955 10591
rect 14013 10557 14047 10591
rect 14105 10557 14139 10591
rect 14289 10547 14323 10581
rect 14562 10557 14596 10591
rect 15025 10557 15059 10591
rect 15117 10557 15151 10591
rect 15301 10557 15335 10591
rect 15669 10557 15703 10591
rect 16497 10557 16531 10591
rect 16589 10557 16623 10591
rect 16773 10557 16807 10591
rect 17141 10557 17175 10591
rect 17417 10557 17451 10591
rect 19073 10557 19107 10591
rect 19165 10557 19199 10591
rect 19441 10557 19475 10591
rect 20177 10557 20211 10591
rect 20729 10557 20763 10591
rect 21833 10557 21867 10591
rect 22201 10557 22235 10591
rect 19855 10523 19889 10557
rect 5181 10489 5215 10523
rect 6837 10489 6871 10523
rect 19257 10489 19291 10523
rect 20085 10489 20119 10523
rect 21925 10489 21959 10523
rect 22109 10489 22143 10523
rect 3801 10421 3835 10455
rect 5089 10421 5123 10455
rect 5457 10421 5491 10455
rect 9321 10421 9355 10455
rect 14565 10421 14599 10455
rect 15301 10421 15335 10455
rect 19717 10421 19751 10455
rect 22017 10421 22051 10455
rect 1869 10217 1903 10251
rect 2329 10217 2363 10251
rect 8217 10217 8251 10251
rect 11621 10217 11655 10251
rect 16681 10217 16715 10251
rect 17233 10217 17267 10251
rect 18981 10217 19015 10251
rect 21557 10217 21591 10251
rect 22201 10217 22235 10251
rect 2697 10149 2731 10183
rect 3233 10149 3267 10183
rect 3433 10149 3467 10183
rect 8585 10149 8619 10183
rect 10793 10149 10827 10183
rect 13277 10149 13311 10183
rect 13553 10149 13587 10183
rect 21373 10149 21407 10183
rect 8355 10115 8389 10149
rect 1593 10081 1627 10115
rect 1685 10081 1719 10115
rect 1961 10081 1995 10115
rect 2145 10081 2179 10115
rect 2237 10081 2271 10115
rect 2513 10081 2547 10115
rect 2605 10081 2639 10115
rect 2835 10081 2869 10115
rect 4629 10081 4663 10115
rect 4813 10081 4847 10115
rect 5365 10081 5399 10115
rect 7849 10081 7883 10115
rect 8677 10081 8711 10115
rect 9229 10081 9263 10115
rect 10241 10081 10275 10115
rect 10517 10081 10551 10115
rect 10609 10081 10643 10115
rect 10977 10081 11011 10115
rect 11161 10081 11195 10115
rect 11253 10081 11287 10115
rect 11365 10081 11399 10115
rect 13093 10081 13127 10115
rect 13369 10081 13403 10115
rect 13461 10081 13495 10115
rect 13645 10081 13679 10115
rect 14841 10081 14875 10115
rect 16865 10081 16899 10115
rect 17095 10081 17129 10115
rect 17509 10081 17543 10115
rect 19533 10081 19567 10115
rect 20453 10081 20487 10115
rect 21281 10081 21315 10115
rect 21925 10081 21959 10115
rect 22385 10081 22419 10115
rect 2973 10013 3007 10047
rect 8769 10013 8803 10047
rect 8953 10013 8987 10047
rect 16957 10013 16991 10047
rect 17325 10013 17359 10047
rect 19349 10013 19383 10047
rect 20269 10013 20303 10047
rect 21741 10013 21775 10047
rect 21833 10013 21867 10047
rect 22017 10013 22051 10047
rect 22569 10013 22603 10047
rect 1961 9945 1995 9979
rect 3065 9945 3099 9979
rect 9045 9945 9079 9979
rect 13093 9945 13127 9979
rect 1409 9877 1443 9911
rect 3249 9877 3283 9911
rect 4721 9877 4755 9911
rect 5549 9877 5583 9911
rect 6561 9877 6595 9911
rect 8401 9877 8435 9911
rect 8861 9877 8895 9911
rect 10333 9877 10367 9911
rect 14657 9877 14691 9911
rect 20637 9877 20671 9911
rect 2513 9673 2547 9707
rect 3249 9673 3283 9707
rect 3433 9673 3467 9707
rect 16773 9673 16807 9707
rect 17417 9673 17451 9707
rect 18889 9673 18923 9707
rect 19073 9673 19107 9707
rect 19809 9673 19843 9707
rect 21189 9673 21223 9707
rect 21741 9673 21775 9707
rect 22569 9673 22603 9707
rect 2789 9605 2823 9639
rect 5457 9605 5491 9639
rect 8217 9605 8251 9639
rect 13783 9605 13817 9639
rect 19993 9605 20027 9639
rect 22385 9605 22419 9639
rect 5181 9537 5215 9571
rect 12541 9537 12575 9571
rect 13553 9537 13587 9571
rect 15301 9537 15335 9571
rect 15669 9537 15703 9571
rect 19165 9537 19199 9571
rect 19533 9537 19567 9571
rect 21281 9537 21315 9571
rect 22293 9537 22327 9571
rect 2697 9469 2731 9503
rect 2881 9469 2915 9503
rect 2973 9469 3007 9503
rect 3433 9469 3467 9503
rect 3525 9469 3559 9503
rect 4997 9469 5031 9503
rect 5089 9469 5123 9503
rect 5273 9469 5307 9503
rect 6469 9469 6503 9503
rect 7944 9447 7978 9481
rect 8033 9469 8067 9503
rect 8401 9469 8435 9503
rect 8657 9469 8691 9503
rect 11069 9469 11103 9503
rect 12265 9469 12299 9503
rect 15025 9469 15059 9503
rect 15393 9469 15427 9503
rect 16405 9469 16439 9503
rect 16589 9469 16623 9503
rect 16773 9469 16807 9503
rect 17141 9469 17175 9503
rect 18245 9469 18279 9503
rect 19349 9469 19383 9503
rect 19855 9435 19889 9469
rect 20085 9445 20119 9479
rect 21005 9469 21039 9503
rect 21097 9469 21131 9503
rect 21431 9469 21465 9503
rect 21557 9469 21591 9503
rect 21833 9469 21867 9503
rect 21925 9469 21959 9503
rect 22017 9469 22051 9503
rect 3709 9401 3743 9435
rect 5733 9401 5767 9435
rect 6009 9401 6043 9435
rect 6101 9401 6135 9435
rect 8217 9401 8251 9435
rect 17969 9401 18003 9435
rect 18061 9401 18095 9435
rect 18705 9401 18739 9435
rect 19625 9401 19659 9435
rect 22753 9401 22787 9435
rect 6837 9333 6871 9367
rect 7021 9333 7055 9367
rect 9781 9333 9815 9367
rect 10885 9333 10919 9367
rect 17601 9333 17635 9367
rect 17693 9333 17727 9367
rect 17785 9333 17819 9367
rect 18429 9333 18463 9367
rect 18905 9333 18939 9367
rect 20269 9333 20303 9367
rect 20729 9333 20763 9367
rect 22543 9333 22577 9367
rect 2237 9129 2271 9163
rect 3893 9129 3927 9163
rect 5365 9129 5399 9163
rect 9137 9129 9171 9163
rect 9505 9129 9539 9163
rect 13369 9129 13403 9163
rect 18061 9129 18095 9163
rect 20177 9129 20211 9163
rect 21833 9129 21867 9163
rect 11713 9061 11747 9095
rect 16221 9061 16255 9095
rect 17693 9061 17727 9095
rect 17893 9061 17927 9095
rect 1961 8993 1995 9027
rect 2145 8993 2179 9027
rect 2237 8993 2271 9027
rect 2329 8993 2363 9027
rect 2513 8993 2547 9027
rect 2973 8993 3007 9027
rect 3065 8993 3099 9027
rect 3249 8993 3283 9027
rect 3525 8993 3559 9027
rect 3985 8993 4019 9027
rect 4077 8993 4111 9027
rect 4997 8993 5031 9027
rect 5181 8993 5215 9027
rect 6193 8993 6227 9027
rect 8861 8993 8895 9027
rect 9321 8993 9355 9027
rect 9597 8993 9631 9027
rect 9873 8993 9907 9027
rect 10333 8993 10367 9027
rect 10977 8993 11011 9027
rect 11161 8993 11195 9027
rect 11253 8993 11287 9027
rect 11345 8993 11379 9027
rect 11897 8993 11931 9027
rect 11989 8993 12023 9027
rect 12265 8993 12299 9027
rect 12541 8993 12575 9027
rect 12633 8993 12667 9027
rect 12817 8993 12851 9027
rect 12909 8993 12943 9027
rect 13185 8993 13219 9027
rect 13645 8993 13679 9027
rect 13783 8993 13817 9027
rect 13927 8993 13961 9027
rect 14025 8995 14059 9029
rect 14197 8993 14231 9027
rect 14473 8993 14507 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 15301 8993 15335 9027
rect 16773 8977 16807 9011
rect 17049 8993 17083 9027
rect 18337 8993 18371 9027
rect 18797 8993 18831 9027
rect 19257 8993 19291 9027
rect 19625 8993 19659 9027
rect 19809 8993 19843 9027
rect 19901 8993 19935 9027
rect 20361 8993 20395 9027
rect 21360 8993 21394 9027
rect 21649 8993 21683 9027
rect 22109 8993 22143 9027
rect 2697 8925 2731 8959
rect 3617 8925 3651 8959
rect 9689 8925 9723 8959
rect 10057 8925 10091 8959
rect 13001 8925 13035 8959
rect 15025 8925 15059 8959
rect 17325 8925 17359 8959
rect 4353 8857 4387 8891
rect 10241 8857 10275 8891
rect 16957 8857 16991 8891
rect 18521 8857 18555 8891
rect 18981 8857 19015 8891
rect 19073 8857 19107 8891
rect 19993 8857 20027 8891
rect 21465 8857 21499 8891
rect 21557 8857 21591 8891
rect 21925 8857 21959 8891
rect 2789 8789 2823 8823
rect 3157 8789 3191 8823
rect 3709 8789 3743 8823
rect 3985 8789 4019 8823
rect 6009 8789 6043 8823
rect 9045 8789 9079 8823
rect 11621 8789 11655 8823
rect 12173 8789 12207 8823
rect 12357 8789 12391 8823
rect 13461 8789 13495 8823
rect 14289 8789 14323 8823
rect 14841 8789 14875 8823
rect 16313 8789 16347 8823
rect 17417 8789 17451 8823
rect 17601 8789 17635 8823
rect 17877 8789 17911 8823
rect 19809 8789 19843 8823
rect 2697 8585 2731 8619
rect 3249 8585 3283 8619
rect 11437 8585 11471 8619
rect 13277 8585 13311 8619
rect 16313 8585 16347 8619
rect 16865 8585 16899 8619
rect 17325 8585 17359 8619
rect 17601 8585 17635 8619
rect 19901 8585 19935 8619
rect 20361 8585 20395 8619
rect 20637 8585 20671 8619
rect 21373 8585 21407 8619
rect 21649 8585 21683 8619
rect 2421 8517 2455 8551
rect 2881 8517 2915 8551
rect 7205 8517 7239 8551
rect 15945 8517 15979 8551
rect 20453 8517 20487 8551
rect 22753 8517 22787 8551
rect 8677 8449 8711 8483
rect 13369 8449 13403 8483
rect 15117 8449 15151 8483
rect 15209 8449 15243 8483
rect 19073 8449 19107 8483
rect 20269 8449 20303 8483
rect 20821 8449 20855 8483
rect 21281 8449 21315 8483
rect 22017 8449 22051 8483
rect 2237 8381 2271 8415
rect 2513 8381 2547 8415
rect 3065 8381 3099 8415
rect 3433 8381 3467 8415
rect 3525 8381 3559 8415
rect 4721 8381 4755 8415
rect 6193 8381 6227 8415
rect 6285 8381 6319 8415
rect 11161 8381 11195 8415
rect 11253 8381 11287 8415
rect 11529 8381 11563 8415
rect 11621 8381 11655 8415
rect 11713 8381 11747 8415
rect 11897 8381 11931 8415
rect 12357 8381 12391 8415
rect 13093 8381 13127 8415
rect 14841 8381 14875 8415
rect 15301 8381 15335 8415
rect 15485 8381 15519 8415
rect 15761 8381 15795 8415
rect 16221 8381 16255 8415
rect 16497 8381 16531 8415
rect 16589 8381 16623 8415
rect 17049 8381 17083 8415
rect 17141 8381 17175 8415
rect 17417 8381 17451 8415
rect 18889 8381 18923 8415
rect 19441 8381 19475 8415
rect 19625 8381 19659 8415
rect 20085 8381 20119 8415
rect 20637 8381 20671 8415
rect 20913 8381 20947 8415
rect 21465 8381 21499 8415
rect 21741 8381 21775 8415
rect 22661 8381 22695 8415
rect 22845 8381 22879 8415
rect 2789 8313 2823 8347
rect 2973 8313 3007 8347
rect 3249 8313 3283 8347
rect 5917 8313 5951 8347
rect 6653 8313 6687 8347
rect 9229 8313 9263 8347
rect 10977 8313 11011 8347
rect 12909 8313 12943 8347
rect 15669 8313 15703 8347
rect 16865 8313 16899 8347
rect 20361 8313 20395 8347
rect 21189 8313 21223 8347
rect 3709 8245 3743 8279
rect 4905 8245 4939 8279
rect 7021 8245 7055 8279
rect 12081 8245 12115 8279
rect 12173 8245 12207 8279
rect 16037 8245 16071 8279
rect 16773 8245 16807 8279
rect 18705 8245 18739 8279
rect 19533 8245 19567 8279
rect 2237 8041 2271 8075
rect 3433 8041 3467 8075
rect 3893 8041 3927 8075
rect 5181 8041 5215 8075
rect 6009 8041 6043 8075
rect 7113 8041 7147 8075
rect 11161 8041 11195 8075
rect 12449 8041 12483 8075
rect 15577 8041 15611 8075
rect 17233 8041 17267 8075
rect 20361 8041 20395 8075
rect 20821 8041 20855 8075
rect 17325 7973 17359 8007
rect 20729 7973 20763 8007
rect 1124 7905 1158 7939
rect 2789 7905 2823 7939
rect 3249 7905 3283 7939
rect 3709 7905 3743 7939
rect 4077 7905 4111 7939
rect 4997 7905 5031 7939
rect 5273 7905 5307 7939
rect 6278 7905 6312 7939
rect 6365 7905 6399 7939
rect 6745 7905 6779 7939
rect 9321 7905 9355 7939
rect 9597 7905 9631 7939
rect 11345 7905 11379 7939
rect 11621 7905 11655 7939
rect 11713 7905 11747 7939
rect 11897 7905 11931 7939
rect 13737 7905 13771 7939
rect 13829 7905 13863 7939
rect 14013 7905 14047 7939
rect 14105 7905 14139 7939
rect 14197 7905 14231 7939
rect 14381 7905 14415 7939
rect 14657 7905 14691 7939
rect 14841 7905 14875 7939
rect 15301 7905 15335 7939
rect 15393 7905 15427 7939
rect 16865 7905 16899 7939
rect 16957 7905 16991 7939
rect 17049 7905 17083 7939
rect 19717 7905 19751 7939
rect 20177 7905 20211 7939
rect 21629 7905 21663 7939
rect 857 7837 891 7871
rect 3065 7837 3099 7871
rect 8861 7837 8895 7871
rect 11529 7837 11563 7871
rect 14565 7837 14599 7871
rect 16773 7837 16807 7871
rect 19993 7837 20027 7871
rect 20453 7837 20487 7871
rect 20938 7837 20972 7871
rect 21373 7837 21407 7871
rect 3617 7769 3651 7803
rect 15117 7769 15151 7803
rect 3249 7701 3283 7735
rect 5457 7701 5491 7735
rect 7297 7701 7331 7735
rect 15025 7701 15059 7735
rect 18797 7701 18831 7735
rect 19441 7701 19475 7735
rect 19993 7701 20027 7735
rect 21097 7701 21131 7735
rect 22753 7701 22787 7735
rect 1409 7497 1443 7531
rect 3249 7497 3283 7531
rect 3709 7497 3743 7531
rect 15485 7497 15519 7531
rect 17601 7497 17635 7531
rect 20361 7497 20395 7531
rect 20821 7497 20855 7531
rect 3985 7429 4019 7463
rect 4169 7429 4203 7463
rect 17417 7429 17451 7463
rect 21005 7429 21039 7463
rect 3065 7361 3099 7395
rect 13369 7361 13403 7395
rect 13829 7361 13863 7395
rect 13921 7361 13955 7395
rect 14473 7361 14507 7395
rect 16221 7361 16255 7395
rect 16497 7361 16531 7395
rect 17785 7361 17819 7395
rect 18981 7361 19015 7395
rect 1409 7293 1443 7327
rect 1593 7293 1627 7327
rect 2789 7293 2823 7327
rect 3433 7293 3467 7327
rect 3525 7293 3559 7327
rect 3709 7293 3743 7327
rect 3801 7293 3835 7327
rect 4721 7293 4755 7327
rect 5181 7293 5215 7327
rect 7481 7293 7515 7327
rect 9965 7293 9999 7327
rect 10149 7293 10183 7327
rect 10333 7293 10367 7327
rect 10793 7293 10827 7327
rect 10885 7293 10919 7327
rect 11069 7293 11103 7327
rect 11161 7293 11195 7327
rect 11253 7293 11287 7327
rect 11713 7293 11747 7327
rect 11805 7293 11839 7327
rect 11897 7293 11931 7327
rect 11989 7293 12023 7327
rect 13093 7293 13127 7327
rect 13553 7293 13587 7327
rect 13737 7293 13771 7327
rect 14105 7293 14139 7327
rect 14565 7293 14599 7327
rect 14657 7293 14691 7327
rect 14749 7293 14783 7327
rect 15209 7293 15243 7327
rect 15301 7293 15335 7327
rect 15577 7293 15611 7327
rect 17141 7293 17175 7327
rect 17509 7293 17543 7327
rect 17969 7293 18003 7327
rect 18153 7293 18187 7327
rect 18337 7293 18371 7327
rect 18705 7293 18739 7327
rect 18797 7293 18831 7327
rect 18889 7293 18923 7327
rect 20637 7293 20671 7327
rect 21097 7293 21131 7327
rect 5089 7225 5123 7259
rect 10425 7225 10459 7259
rect 10609 7225 10643 7259
rect 15025 7225 15059 7259
rect 17417 7225 17451 7259
rect 17785 7225 17819 7259
rect 18245 7225 18279 7259
rect 19226 7225 19260 7259
rect 4353 7157 4387 7191
rect 5457 7157 5491 7191
rect 6193 7157 6227 7191
rect 11529 7157 11563 7191
rect 12173 7157 12207 7191
rect 14289 7157 14323 7191
rect 14933 7157 14967 7191
rect 17233 7157 17267 7191
rect 18521 7157 18555 7191
rect 1777 6953 1811 6987
rect 2421 6953 2455 6987
rect 3341 6953 3375 6987
rect 3617 6953 3651 6987
rect 3801 6953 3835 6987
rect 7389 6953 7423 6987
rect 14013 6953 14047 6987
rect 21281 6953 21315 6987
rect 2589 6885 2623 6919
rect 2789 6885 2823 6919
rect 6285 6885 6319 6919
rect 2053 6817 2087 6851
rect 2881 6817 2915 6851
rect 3157 6817 3191 6851
rect 3341 6817 3375 6851
rect 3433 6817 3467 6851
rect 3985 6817 4019 6851
rect 4169 6817 4203 6851
rect 4629 6817 4663 6851
rect 6561 6817 6595 6851
rect 6653 6817 6687 6851
rect 7021 6817 7055 6851
rect 7849 6817 7883 6851
rect 8392 6817 8426 6851
rect 10609 6817 10643 6851
rect 10793 6817 10827 6851
rect 10977 6817 11011 6851
rect 11161 6817 11195 6851
rect 11253 6817 11287 6851
rect 11345 6817 11379 6851
rect 11529 6817 11563 6851
rect 12265 6817 12299 6851
rect 13277 6817 13311 6851
rect 13461 6817 13495 6851
rect 13829 6817 13863 6851
rect 14105 6817 14139 6851
rect 14289 6817 14323 6851
rect 14565 6817 14599 6851
rect 14841 6817 14875 6851
rect 16589 6817 16623 6851
rect 17325 6817 17359 6851
rect 17509 6817 17543 6851
rect 17601 6817 17635 6851
rect 21097 6817 21131 6851
rect 21557 6817 21591 6851
rect 21741 6817 21775 6851
rect 22017 6817 22051 6851
rect 1777 6749 1811 6783
rect 8125 6749 8159 6783
rect 11989 6749 12023 6783
rect 12081 6749 12115 6783
rect 12173 6749 12207 6783
rect 13553 6749 13587 6783
rect 13645 6749 13679 6783
rect 4445 6681 4479 6715
rect 7573 6681 7607 6715
rect 9505 6681 9539 6715
rect 10701 6681 10735 6715
rect 16773 6681 16807 6715
rect 17325 6681 17359 6715
rect 1961 6613 1995 6647
rect 2605 6613 2639 6647
rect 3065 6613 3099 6647
rect 4353 6613 4387 6647
rect 8033 6613 8067 6647
rect 11713 6613 11747 6647
rect 11805 6613 11839 6647
rect 14197 6613 14231 6647
rect 14657 6613 14691 6647
rect 15025 6613 15059 6647
rect 20913 6613 20947 6647
rect 21649 6613 21683 6647
rect 21833 6613 21867 6647
rect 2237 6409 2271 6443
rect 2605 6409 2639 6443
rect 2789 6409 2823 6443
rect 8585 6409 8619 6443
rect 20913 6409 20947 6443
rect 22845 6409 22879 6443
rect 1593 6341 1627 6375
rect 8953 6341 8987 6375
rect 13921 6341 13955 6375
rect 1777 6273 1811 6307
rect 11161 6273 11195 6307
rect 11253 6273 11287 6307
rect 11345 6273 11379 6307
rect 11712 6273 11746 6307
rect 11897 6273 11931 6307
rect 15301 6273 15335 6307
rect 21005 6273 21039 6307
rect 21465 6273 21499 6307
rect 1501 6205 1535 6239
rect 1961 6205 1995 6239
rect 2053 6205 2087 6239
rect 2329 6205 2363 6239
rect 2513 6205 2547 6239
rect 5549 6205 5583 6239
rect 6285 6205 6319 6239
rect 6377 6205 6411 6239
rect 11069 6205 11103 6239
rect 11620 6205 11654 6239
rect 11815 6205 11849 6239
rect 13737 6205 13771 6239
rect 14013 6205 14047 6239
rect 14841 6205 14875 6239
rect 15025 6205 15059 6239
rect 15209 6205 15243 6239
rect 15393 6205 15427 6239
rect 15485 6205 15519 6239
rect 16129 6205 16163 6239
rect 16405 6205 16439 6239
rect 17969 6205 18003 6239
rect 18153 6205 18187 6239
rect 18705 6205 18739 6239
rect 19073 6205 19107 6239
rect 21189 6205 21223 6239
rect 1777 6137 1811 6171
rect 2973 6137 3007 6171
rect 6009 6137 6043 6171
rect 6745 6137 6779 6171
rect 12173 6137 12207 6171
rect 12357 6137 12391 6171
rect 14933 6137 14967 6171
rect 15761 6137 15795 6171
rect 15945 6137 15979 6171
rect 18061 6137 18095 6171
rect 18889 6137 18923 6171
rect 18981 6137 19015 6171
rect 20913 6137 20947 6171
rect 21710 6137 21744 6171
rect 2421 6069 2455 6103
rect 2763 6069 2797 6103
rect 5733 6069 5767 6103
rect 7113 6069 7147 6103
rect 7297 6069 7331 6103
rect 8401 6069 8435 6103
rect 8585 6069 8619 6103
rect 10885 6069 10919 6103
rect 12081 6069 12115 6103
rect 12541 6069 12575 6103
rect 13553 6069 13587 6103
rect 15669 6069 15703 6103
rect 16221 6069 16255 6103
rect 19257 6069 19291 6103
rect 21373 6069 21407 6103
rect 8125 5865 8159 5899
rect 8401 5865 8435 5899
rect 8493 5865 8527 5899
rect 11621 5865 11655 5899
rect 15485 5865 15519 5899
rect 17693 5865 17727 5899
rect 18889 5865 18923 5899
rect 21097 5865 21131 5899
rect 22109 5865 22143 5899
rect 2053 5797 2087 5831
rect 8033 5797 8067 5831
rect 18521 5797 18555 5831
rect 19073 5797 19107 5831
rect 19962 5797 19996 5831
rect 2329 5729 2363 5763
rect 2585 5729 2619 5763
rect 5825 5729 5859 5763
rect 6081 5729 6115 5763
rect 7573 5729 7607 5763
rect 7849 5729 7883 5763
rect 8217 5729 8251 5763
rect 8677 5729 8711 5763
rect 9137 5729 9171 5763
rect 10793 5729 10827 5763
rect 10977 5729 11011 5763
rect 11161 5729 11195 5763
rect 11253 5729 11287 5763
rect 11345 5729 11379 5763
rect 12265 5729 12299 5763
rect 12449 5729 12483 5763
rect 12725 5729 12759 5763
rect 12909 5729 12943 5763
rect 13277 5729 13311 5763
rect 13461 5729 13495 5763
rect 13737 5729 13771 5763
rect 15393 5729 15427 5763
rect 15669 5729 15703 5763
rect 17049 5729 17083 5763
rect 17141 5729 17175 5763
rect 17601 5729 17635 5763
rect 17785 5729 17819 5763
rect 18061 5729 18095 5763
rect 18337 5729 18371 5763
rect 18613 5729 18647 5763
rect 18705 5729 18739 5763
rect 18981 5729 19015 5763
rect 19165 5729 19199 5763
rect 19717 5729 19751 5763
rect 21557 5729 21591 5763
rect 21925 5729 21959 5763
rect 22201 5729 22235 5763
rect 1685 5661 1719 5695
rect 5089 5661 5123 5695
rect 5181 5661 5215 5695
rect 5273 5661 5307 5695
rect 5365 5661 5399 5695
rect 8769 5661 8803 5695
rect 8861 5661 8895 5695
rect 8953 5661 8987 5695
rect 9229 5661 9263 5695
rect 12187 5661 12221 5695
rect 12357 5661 12391 5695
rect 13001 5661 13035 5695
rect 13093 5661 13127 5695
rect 14013 5661 14047 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 21465 5661 21499 5695
rect 7757 5593 7791 5627
rect 13553 5593 13587 5627
rect 22385 5593 22419 5627
rect 2053 5525 2087 5559
rect 2237 5525 2271 5559
rect 3709 5525 3743 5559
rect 4905 5525 4939 5559
rect 7205 5525 7239 5559
rect 10609 5525 10643 5559
rect 12633 5525 12667 5559
rect 13921 5525 13955 5559
rect 15209 5525 15243 5559
rect 16865 5525 16899 5559
rect 17325 5525 17359 5559
rect 21925 5525 21959 5559
rect 5365 5321 5399 5355
rect 6607 5321 6641 5355
rect 12357 5321 12391 5355
rect 18521 5321 18555 5355
rect 21097 5321 21131 5355
rect 21465 5321 21499 5355
rect 22017 5321 22051 5355
rect 2145 5253 2179 5287
rect 18889 5253 18923 5287
rect 1961 5185 1995 5219
rect 4813 5185 4847 5219
rect 5733 5185 5767 5219
rect 6377 5185 6411 5219
rect 7665 5185 7699 5219
rect 11069 5185 11103 5219
rect 11713 5185 11747 5219
rect 15485 5185 15519 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 18153 5185 18187 5219
rect 21557 5185 21591 5219
rect 2237 5117 2271 5151
rect 2513 5117 2547 5151
rect 4537 5117 4571 5151
rect 5181 5117 5215 5151
rect 5457 5117 5491 5151
rect 7573 5117 7607 5151
rect 8401 5117 8435 5151
rect 8677 5117 8711 5151
rect 10333 5117 10367 5151
rect 10701 5117 10735 5151
rect 10793 5117 10827 5151
rect 10977 5117 11011 5151
rect 11161 5117 11195 5151
rect 11345 5117 11379 5151
rect 11805 5117 11839 5151
rect 11897 5117 11931 5151
rect 11989 5117 12023 5151
rect 12633 5117 12667 5151
rect 12725 5117 12759 5151
rect 12817 5117 12851 5151
rect 13001 5117 13035 5151
rect 13553 5117 13587 5151
rect 13829 5117 13863 5151
rect 14933 5117 14967 5151
rect 15209 5117 15243 5151
rect 15301 5117 15335 5151
rect 15577 5117 15611 5151
rect 17693 5117 17727 5151
rect 18337 5117 18371 5151
rect 18705 5117 18739 5151
rect 18889 5117 18923 5151
rect 21373 5117 21407 5151
rect 21465 5117 21499 5151
rect 21741 5117 21775 5151
rect 21925 5117 21959 5151
rect 22109 5107 22143 5141
rect 8493 5049 8527 5083
rect 10517 5049 10551 5083
rect 1961 4981 1995 5015
rect 2329 4981 2363 5015
rect 7941 4981 7975 5015
rect 8861 4981 8895 5015
rect 11529 4981 11563 5015
rect 12173 4981 12207 5015
rect 14749 4981 14783 5015
rect 15025 4981 15059 5015
rect 15669 4981 15703 5015
rect 16313 4981 16347 5015
rect 17877 4981 17911 5015
rect 2697 4777 2731 4811
rect 3433 4777 3467 4811
rect 5549 4777 5583 4811
rect 7757 4777 7791 4811
rect 11897 4777 11931 4811
rect 13553 4777 13587 4811
rect 16865 4777 16899 4811
rect 18521 4777 18555 4811
rect 21097 4777 21131 4811
rect 22661 4777 22695 4811
rect 1584 4709 1618 4743
rect 18061 4709 18095 4743
rect 20637 4709 20671 4743
rect 1317 4641 1351 4675
rect 3617 4641 3651 4675
rect 4813 4641 4847 4675
rect 5365 4641 5399 4675
rect 5825 4641 5859 4675
rect 6929 4641 6963 4675
rect 7389 4641 7423 4675
rect 7573 4641 7607 4675
rect 10609 4641 10643 4675
rect 11713 4641 11747 4675
rect 11897 4641 11931 4675
rect 13093 4641 13127 4675
rect 13737 4641 13771 4675
rect 13829 4641 13863 4675
rect 14105 4641 14139 4675
rect 14381 4641 14415 4675
rect 15209 4641 15243 4675
rect 15393 4641 15427 4675
rect 15577 4641 15611 4675
rect 15761 4641 15795 4675
rect 16129 4641 16163 4675
rect 16313 4641 16347 4675
rect 16405 4641 16439 4675
rect 16497 4641 16531 4675
rect 16681 4641 16715 4675
rect 18337 4641 18371 4675
rect 19073 4641 19107 4675
rect 19533 4641 19567 4675
rect 19625 4641 19659 4675
rect 20913 4641 20947 4675
rect 21281 4641 21315 4675
rect 21537 4641 21571 4675
rect 3709 4573 3743 4607
rect 3985 4573 4019 4607
rect 4629 4573 4663 4607
rect 5917 4573 5951 4607
rect 7021 4573 7055 4607
rect 12817 4573 12851 4607
rect 12909 4573 12943 4607
rect 14013 4573 14047 4607
rect 15485 4573 15519 4607
rect 18245 4573 18279 4607
rect 19809 4573 19843 4607
rect 20821 4573 20855 4607
rect 7297 4505 7331 4539
rect 10793 4505 10827 4539
rect 20269 4505 20303 4539
rect 4997 4437 5031 4471
rect 13277 4437 13311 4471
rect 14197 4437 14231 4471
rect 15945 4437 15979 4471
rect 18337 4437 18371 4471
rect 18889 4437 18923 4471
rect 19717 4437 19751 4471
rect 20729 4437 20763 4471
rect 2697 4233 2731 4267
rect 18337 4233 18371 4267
rect 22017 4233 22051 4267
rect 21649 4165 21683 4199
rect 22569 4165 22603 4199
rect 4353 4097 4387 4131
rect 4629 4097 4663 4131
rect 7665 4097 7699 4131
rect 13369 4097 13403 4131
rect 13829 4097 13863 4131
rect 13921 4097 13955 4131
rect 14381 4097 14415 4131
rect 14473 4097 14507 4131
rect 15669 4097 15703 4131
rect 16037 4097 16071 4131
rect 18705 4097 18739 4131
rect 1777 4029 1811 4063
rect 2053 4029 2087 4063
rect 2329 4029 2363 4063
rect 2513 4029 2547 4063
rect 4261 4029 4295 4063
rect 4997 4029 5031 4063
rect 5089 4029 5123 4063
rect 5273 4029 5307 4063
rect 7849 4029 7883 4063
rect 8401 4029 8435 4063
rect 8493 4029 8527 4063
rect 8585 4029 8619 4063
rect 9137 4029 9171 4063
rect 12725 4029 12759 4063
rect 12909 4029 12943 4063
rect 13001 4029 13035 4063
rect 13093 4029 13127 4063
rect 13553 4029 13587 4063
rect 13737 4029 13771 4063
rect 14105 4029 14139 4063
rect 14657 4029 14691 4063
rect 15209 4029 15243 4063
rect 15393 4029 15427 4063
rect 15577 4029 15611 4063
rect 15761 4029 15795 4063
rect 15945 4019 15979 4053
rect 16129 4029 16163 4063
rect 16313 4029 16347 4063
rect 18521 4029 18555 4063
rect 18981 4029 19015 4063
rect 19901 4029 19935 4063
rect 20085 4029 20119 4063
rect 20177 4029 20211 4063
rect 20269 4029 20303 4063
rect 20637 4029 20671 4063
rect 20821 4029 20855 4063
rect 20913 4029 20947 4063
rect 21005 4029 21039 4063
rect 21557 4029 21591 4063
rect 21833 4029 21867 4063
rect 22109 4029 22143 4063
rect 22477 4029 22511 4063
rect 22753 4029 22787 4063
rect 5457 3961 5491 3995
rect 10149 3961 10183 3995
rect 14289 3961 14323 3995
rect 20545 3961 20579 3995
rect 1875 3893 1909 3927
rect 1961 3893 1995 3927
rect 8033 3893 8067 3927
rect 14841 3893 14875 3927
rect 16497 3893 16531 3927
rect 21281 3893 21315 3927
rect 21373 3893 21407 3927
rect 22293 3893 22327 3927
rect 2329 3689 2363 3723
rect 3617 3689 3651 3723
rect 6377 3689 6411 3723
rect 9045 3689 9079 3723
rect 10057 3689 10091 3723
rect 13093 3689 13127 3723
rect 18613 3689 18647 3723
rect 19191 3689 19225 3723
rect 19993 3689 20027 3723
rect 22661 3689 22695 3723
rect 2789 3621 2823 3655
rect 2973 3621 3007 3655
rect 4752 3621 4786 3655
rect 6561 3621 6595 3655
rect 11973 3621 12007 3655
rect 12173 3621 12207 3655
rect 18061 3621 18095 3655
rect 18981 3621 19015 3655
rect 21526 3621 21560 3655
rect 949 3553 983 3587
rect 1216 3553 1250 3587
rect 4997 3553 5031 3587
rect 5457 3553 5491 3587
rect 6469 3553 6503 3587
rect 6745 3553 6779 3587
rect 7021 3553 7055 3587
rect 7665 3553 7699 3587
rect 7941 3553 7975 3587
rect 8125 3553 8159 3587
rect 8217 3553 8251 3587
rect 8585 3553 8619 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 9413 3553 9447 3587
rect 9781 3553 9815 3587
rect 10333 3553 10367 3587
rect 10609 3553 10643 3587
rect 10793 3553 10827 3587
rect 12265 3553 12299 3587
rect 13277 3553 13311 3587
rect 13369 3553 13403 3587
rect 13627 3553 13661 3587
rect 13737 3553 13771 3587
rect 13921 3553 13955 3587
rect 15117 3553 15151 3587
rect 15301 3553 15335 3587
rect 15393 3553 15427 3587
rect 15485 3553 15519 3587
rect 16129 3553 16163 3587
rect 16313 3553 16347 3587
rect 17325 3553 17359 3587
rect 17509 3553 17543 3587
rect 18153 3553 18187 3587
rect 18245 3553 18279 3587
rect 18705 3553 18739 3587
rect 19625 3553 19659 3587
rect 19809 3553 19843 3587
rect 20269 3553 20303 3587
rect 21281 3553 21315 3587
rect 5365 3485 5399 3519
rect 6009 3485 6043 3519
rect 6193 3485 6227 3519
rect 8033 3485 8067 3519
rect 8677 3485 8711 3519
rect 8769 3485 8803 3519
rect 8861 3485 8895 3519
rect 9873 3485 9907 3519
rect 9965 3485 9999 3519
rect 10241 3485 10275 3519
rect 11621 3485 11655 3519
rect 5089 3417 5123 3451
rect 10701 3417 10735 3451
rect 11253 3417 11287 3451
rect 12449 3417 12483 3451
rect 6929 3349 6963 3383
rect 7849 3349 7883 3383
rect 8401 3349 8435 3383
rect 10517 3349 10551 3383
rect 11161 3349 11195 3383
rect 11805 3349 11839 3383
rect 11989 3349 12023 3383
rect 13553 3349 13587 3383
rect 13829 3349 13863 3383
rect 15761 3349 15795 3383
rect 16221 3349 16255 3383
rect 17325 3349 17359 3383
rect 18429 3349 18463 3383
rect 19165 3349 19199 3383
rect 19349 3349 19383 3383
rect 20085 3349 20119 3383
rect 1409 3145 1443 3179
rect 2789 3145 2823 3179
rect 3249 3145 3283 3179
rect 6561 3145 6595 3179
rect 12725 3145 12759 3179
rect 13369 3145 13403 3179
rect 15301 3145 15335 3179
rect 19717 3145 19751 3179
rect 2421 3077 2455 3111
rect 19901 3077 19935 3111
rect 10793 3009 10827 3043
rect 13645 3009 13679 3043
rect 13737 3009 13771 3043
rect 13921 3009 13955 3043
rect 14473 3009 14507 3043
rect 14565 3009 14599 3043
rect 14657 3009 14691 3043
rect 15761 3009 15795 3043
rect 16221 3009 16255 3043
rect 16313 3009 16347 3043
rect 16405 3009 16439 3043
rect 1593 2941 1627 2975
rect 1961 2941 1995 2975
rect 2329 2941 2363 2975
rect 2513 2941 2547 2975
rect 3433 2941 3467 2975
rect 3617 2941 3651 2975
rect 6929 2941 6963 2975
rect 7665 2941 7699 2975
rect 8953 2941 8987 2975
rect 9229 2941 9263 2975
rect 9321 2941 9355 2975
rect 9432 2941 9466 2975
rect 9597 2941 9631 2975
rect 9965 2941 9999 2975
rect 10149 2941 10183 2975
rect 10517 2941 10551 2975
rect 12909 2941 12943 2975
rect 13829 2941 13863 2975
rect 14381 2941 14415 2975
rect 15025 2941 15059 2975
rect 15485 2941 15519 2975
rect 15577 2941 15611 2975
rect 15669 2941 15703 2975
rect 16129 2941 16163 2975
rect 16589 2941 16623 2975
rect 16957 2941 16991 2975
rect 17141 2941 17175 2975
rect 18797 2941 18831 2975
rect 18981 2941 19015 2975
rect 19349 2941 19383 2975
rect 21097 2941 21131 2975
rect 2743 2907 2777 2941
rect 2973 2873 3007 2907
rect 7849 2873 7883 2907
rect 13001 2873 13035 2907
rect 13185 2873 13219 2907
rect 14841 2873 14875 2907
rect 15209 2873 15243 2907
rect 16681 2873 16715 2907
rect 19717 2873 19751 2907
rect 19993 2873 20027 2907
rect 20177 2873 20211 2907
rect 20361 2873 20395 2907
rect 1777 2805 1811 2839
rect 2605 2805 2639 2839
rect 6377 2805 6411 2839
rect 6561 2805 6595 2839
rect 7481 2805 7515 2839
rect 9137 2805 9171 2839
rect 9781 2805 9815 2839
rect 10333 2805 10367 2839
rect 14105 2805 14139 2839
rect 14197 2805 14231 2839
rect 15945 2805 15979 2839
rect 18797 2805 18831 2839
rect 21281 2805 21315 2839
rect 2513 2601 2547 2635
rect 9781 2601 9815 2635
rect 22845 2601 22879 2635
rect 1400 2533 1434 2567
rect 9505 2533 9539 2567
rect 9689 2533 9723 2567
rect 13553 2533 13587 2567
rect 19625 2533 19659 2567
rect 21710 2533 21744 2567
rect 1133 2465 1167 2499
rect 2881 2465 2915 2499
rect 3157 2465 3191 2499
rect 3985 2465 4019 2499
rect 9781 2465 9815 2499
rect 9965 2465 9999 2499
rect 10149 2465 10183 2499
rect 10241 2465 10275 2499
rect 11253 2465 11287 2499
rect 11345 2465 11379 2499
rect 11621 2465 11655 2499
rect 13185 2449 13219 2483
rect 14289 2465 14323 2499
rect 16313 2465 16347 2499
rect 16589 2465 16623 2499
rect 16773 2465 16807 2499
rect 18245 2465 18279 2499
rect 18889 2465 18923 2499
rect 19073 2465 19107 2499
rect 19349 2465 19383 2499
rect 19717 2465 19751 2499
rect 19901 2465 19935 2499
rect 21465 2465 21499 2499
rect 4445 2397 4479 2431
rect 4721 2397 4755 2431
rect 10333 2397 10367 2431
rect 11069 2397 11103 2431
rect 11161 2397 11195 2431
rect 11897 2397 11931 2431
rect 14013 2397 14047 2431
rect 16129 2397 16163 2431
rect 16497 2397 16531 2431
rect 19257 2397 19291 2431
rect 19441 2397 19475 2431
rect 19625 2397 19659 2431
rect 10057 2329 10091 2363
rect 13829 2329 13863 2363
rect 16405 2329 16439 2363
rect 3801 2261 3835 2295
rect 11529 2261 11563 2295
rect 13001 2261 13035 2295
rect 14105 2261 14139 2295
rect 18337 2261 18371 2295
rect 19901 2261 19935 2295
rect 6101 2057 6135 2091
rect 8953 2057 8987 2091
rect 9413 2057 9447 2091
rect 18889 2057 18923 2091
rect 21741 2057 21775 2091
rect 1685 1989 1719 2023
rect 6745 1989 6779 2023
rect 7205 1989 7239 2023
rect 18061 1989 18095 2023
rect 3801 1921 3835 1955
rect 4169 1921 4203 1955
rect 4721 1921 4755 1955
rect 4905 1921 4939 1955
rect 5365 1921 5399 1955
rect 7481 1921 7515 1955
rect 7849 1921 7883 1955
rect 7941 1921 7975 1955
rect 8493 1921 8527 1955
rect 8585 1921 8619 1955
rect 9045 1921 9079 1955
rect 10425 1921 10459 1955
rect 10609 1921 10643 1955
rect 12357 1921 12391 1955
rect 16313 1921 16347 1955
rect 16405 1921 16439 1955
rect 16957 1921 16991 1955
rect 20729 1921 20763 1955
rect 21281 1921 21315 1955
rect 21649 1921 21683 1955
rect 1593 1853 1627 1887
rect 1869 1853 1903 1887
rect 3985 1853 4019 1887
rect 4261 1853 4295 1887
rect 4537 1853 4571 1887
rect 4997 1853 5031 1887
rect 5457 1853 5491 1887
rect 5917 1853 5951 1887
rect 6561 1853 6595 1887
rect 7113 1853 7147 1887
rect 7297 1853 7331 1887
rect 7389 1853 7423 1887
rect 7573 1853 7607 1887
rect 7757 1853 7791 1887
rect 8033 1853 8067 1887
rect 8677 1853 8711 1887
rect 8769 1853 8803 1887
rect 9229 1853 9263 1887
rect 9597 1853 9631 1887
rect 9781 1853 9815 1887
rect 9965 1853 9999 1887
rect 10517 1853 10551 1887
rect 10701 1853 10735 1887
rect 11161 1853 11195 1887
rect 11253 1853 11287 1887
rect 11345 1853 11379 1887
rect 11529 1853 11563 1887
rect 12265 1853 12299 1887
rect 12449 1853 12483 1887
rect 15669 1853 15703 1887
rect 15761 1853 15795 1887
rect 15853 1853 15887 1887
rect 16037 1853 16071 1887
rect 16221 1853 16255 1887
rect 16497 1853 16531 1887
rect 17141 1853 17175 1887
rect 17409 1855 17443 1889
rect 17601 1853 17635 1887
rect 17877 1853 17911 1887
rect 18061 1853 18095 1887
rect 19165 1853 19199 1887
rect 20913 1853 20947 1887
rect 21189 1853 21223 1887
rect 21465 1853 21499 1887
rect 21925 1853 21959 1887
rect 22209 1847 22243 1881
rect 4353 1785 4387 1819
rect 5595 1785 5629 1819
rect 5733 1785 5767 1819
rect 5825 1785 5859 1819
rect 13277 1785 13311 1819
rect 13737 1785 13771 1819
rect 14565 1785 14599 1819
rect 17325 1785 17359 1819
rect 18429 1785 18463 1819
rect 1409 1717 1443 1751
rect 8217 1717 8251 1751
rect 10241 1717 10275 1751
rect 10885 1717 10919 1751
rect 13185 1717 13219 1751
rect 13645 1717 13679 1751
rect 14657 1717 14691 1751
rect 15393 1717 15427 1751
rect 16681 1717 16715 1751
rect 17417 1717 17451 1751
rect 18705 1717 18739 1751
rect 21097 1717 21131 1751
rect 22109 1717 22143 1751
rect 4537 1513 4571 1547
rect 7757 1513 7791 1547
rect 9045 1513 9079 1547
rect 22661 1513 22695 1547
rect 1961 1445 1995 1479
rect 2504 1445 2538 1479
rect 18061 1445 18095 1479
rect 22109 1445 22143 1479
rect 1225 1377 1259 1411
rect 3893 1377 3927 1411
rect 4353 1377 4387 1411
rect 4997 1377 5031 1411
rect 6377 1377 6411 1411
rect 6469 1377 6503 1411
rect 6653 1377 6687 1411
rect 6929 1377 6963 1411
rect 7113 1377 7147 1411
rect 7205 1377 7239 1411
rect 7389 1377 7423 1411
rect 7941 1377 7975 1411
rect 8217 1377 8251 1411
rect 8585 1377 8619 1411
rect 9229 1377 9263 1411
rect 9413 1377 9447 1411
rect 9505 1377 9539 1411
rect 9965 1377 9999 1411
rect 10149 1377 10183 1411
rect 10425 1377 10459 1411
rect 10609 1377 10643 1411
rect 11345 1377 11379 1411
rect 11437 1377 11471 1411
rect 11529 1377 11563 1411
rect 11713 1377 11747 1411
rect 12265 1377 12299 1411
rect 12449 1377 12483 1411
rect 13185 1377 13219 1411
rect 13737 1377 13771 1411
rect 13921 1377 13955 1411
rect 14289 1377 14323 1411
rect 14565 1377 14599 1411
rect 14749 1377 14783 1411
rect 14933 1377 14967 1411
rect 15209 1377 15243 1411
rect 15577 1377 15611 1411
rect 15761 1377 15795 1411
rect 16221 1377 16255 1411
rect 16405 1377 16439 1411
rect 16773 1377 16807 1411
rect 16957 1377 16991 1411
rect 17233 1377 17267 1411
rect 17601 1377 17635 1411
rect 17785 1377 17819 1411
rect 19973 1377 20007 1411
rect 22477 1377 22511 1411
rect 2237 1309 2271 1343
rect 3985 1309 4019 1343
rect 4261 1309 4295 1343
rect 4905 1309 4939 1343
rect 7297 1309 7331 1343
rect 8125 1309 8159 1343
rect 8861 1309 8895 1343
rect 10241 1309 10275 1343
rect 10333 1309 10367 1343
rect 12173 1309 12207 1343
rect 13461 1309 13495 1343
rect 14013 1309 14047 1343
rect 14841 1309 14875 1343
rect 15485 1309 15519 1343
rect 16129 1309 16163 1343
rect 16681 1309 16715 1343
rect 17509 1309 17543 1343
rect 18889 1309 18923 1343
rect 19717 1309 19751 1343
rect 21557 1309 21591 1343
rect 1777 1241 1811 1275
rect 3617 1241 3651 1275
rect 5365 1241 5399 1275
rect 8033 1241 8067 1275
rect 11069 1241 11103 1275
rect 14105 1241 14139 1275
rect 15393 1241 15427 1275
rect 17141 1241 17175 1275
rect 21097 1241 21131 1275
rect 949 1173 983 1207
rect 7113 1173 7147 1207
rect 8401 1173 8435 1207
rect 8769 1173 8803 1207
rect 9781 1173 9815 1207
rect 10793 1173 10827 1207
rect 12633 1173 12667 1207
rect 13001 1173 13035 1207
rect 13369 1173 13403 1207
rect 13553 1173 13587 1207
rect 14381 1173 14415 1207
rect 15117 1173 15151 1207
rect 15945 1173 15979 1207
rect 16589 1173 16623 1207
rect 17417 1173 17451 1207
rect 17969 1173 18003 1207
rect 2789 969 2823 1003
rect 11713 969 11747 1003
rect 16221 969 16255 1003
rect 18797 969 18831 1003
rect 9045 901 9079 935
rect 1409 833 1443 867
rect 11621 833 11655 867
rect 18705 833 18739 867
rect 21373 833 21407 867
rect 22109 833 22143 867
rect 1225 765 1259 799
rect 3525 765 3559 799
rect 4537 765 4571 799
rect 5365 765 5399 799
rect 6193 765 6227 799
rect 8677 765 8711 799
rect 8861 765 8895 799
rect 9229 765 9263 799
rect 9781 765 9815 799
rect 10057 765 10091 799
rect 11069 765 11103 799
rect 11897 765 11931 799
rect 12081 765 12115 799
rect 12173 765 12207 799
rect 12817 765 12851 799
rect 13553 765 13587 799
rect 14473 765 14507 799
rect 16129 765 16163 799
rect 16405 765 16439 799
rect 16681 765 16715 799
rect 17509 765 17543 799
rect 18245 765 18279 799
rect 18981 765 19015 799
rect 19993 765 20027 799
rect 20821 765 20855 799
rect 22201 765 22235 799
rect 22569 765 22603 799
rect 1676 697 1710 731
rect 3617 697 3651 731
rect 3985 697 4019 731
rect 19165 697 19199 731
rect 19349 697 19383 731
rect 1041 629 1075 663
rect 3341 629 3375 663
rect 4353 629 4387 663
rect 5181 629 5215 663
rect 6009 629 6043 663
rect 8493 629 8527 663
rect 9413 629 9447 663
rect 9597 629 9631 663
rect 10241 629 10275 663
rect 11161 629 11195 663
rect 12357 629 12391 663
rect 12633 629 12667 663
rect 13737 629 13771 663
rect 14289 629 14323 663
rect 16589 629 16623 663
rect 16865 629 16899 663
rect 17693 629 17727 663
rect 18429 629 18463 663
rect 19441 629 19475 663
rect 20177 629 20211 663
rect 21005 629 21039 663
rect 22753 629 22787 663
<< metal1 >>
rect 16206 15416 16212 15428
rect 6564 15388 16212 15416
rect 6564 15360 6592 15388
rect 16206 15376 16212 15388
rect 16264 15376 16270 15428
rect 17218 15376 17224 15428
rect 17276 15416 17282 15428
rect 17276 15388 22324 15416
rect 17276 15376 17282 15388
rect 22296 15360 22324 15388
rect 6546 15308 6552 15360
rect 6604 15308 6610 15360
rect 6730 15308 6736 15360
rect 6788 15348 6794 15360
rect 14458 15348 14464 15360
rect 6788 15320 14464 15348
rect 6788 15308 6794 15320
rect 14458 15308 14464 15320
rect 14516 15308 14522 15360
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 18046 15348 18052 15360
rect 14792 15320 18052 15348
rect 14792 15308 14798 15320
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 22278 15308 22284 15360
rect 22336 15308 22342 15360
rect 552 15258 23368 15280
rect 552 15206 1366 15258
rect 1418 15206 1430 15258
rect 1482 15206 1494 15258
rect 1546 15206 1558 15258
rect 1610 15206 1622 15258
rect 1674 15206 1686 15258
rect 1738 15206 7366 15258
rect 7418 15206 7430 15258
rect 7482 15206 7494 15258
rect 7546 15206 7558 15258
rect 7610 15206 7622 15258
rect 7674 15206 7686 15258
rect 7738 15206 13366 15258
rect 13418 15206 13430 15258
rect 13482 15206 13494 15258
rect 13546 15206 13558 15258
rect 13610 15206 13622 15258
rect 13674 15206 13686 15258
rect 13738 15206 19366 15258
rect 19418 15206 19430 15258
rect 19482 15206 19494 15258
rect 19546 15206 19558 15258
rect 19610 15206 19622 15258
rect 19674 15206 19686 15258
rect 19738 15206 23368 15258
rect 552 15184 23368 15206
rect 4614 15104 4620 15156
rect 4672 15104 4678 15156
rect 5166 15104 5172 15156
rect 5224 15104 5230 15156
rect 6178 15104 6184 15156
rect 6236 15104 6242 15156
rect 6638 15104 6644 15156
rect 6696 15104 6702 15156
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 7561 15147 7619 15153
rect 7561 15144 7573 15147
rect 7340 15116 7573 15144
rect 7340 15104 7346 15116
rect 7561 15113 7573 15116
rect 7607 15113 7619 15147
rect 7561 15107 7619 15113
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 8481 15147 8539 15153
rect 8481 15144 8493 15147
rect 8168 15116 8493 15144
rect 8168 15104 8174 15116
rect 8481 15113 8493 15116
rect 8527 15113 8539 15147
rect 8481 15107 8539 15113
rect 9122 15104 9128 15156
rect 9180 15104 9186 15156
rect 9582 15104 9588 15156
rect 9640 15104 9646 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 10505 15147 10563 15153
rect 10505 15144 10517 15147
rect 10376 15116 10517 15144
rect 10376 15104 10382 15116
rect 10505 15113 10517 15116
rect 10551 15113 10563 15147
rect 10505 15107 10563 15113
rect 11054 15104 11060 15156
rect 11112 15104 11118 15156
rect 14458 15104 14464 15156
rect 14516 15144 14522 15156
rect 14516 15116 16252 15144
rect 14516 15104 14522 15116
rect 16117 15079 16175 15085
rect 16117 15076 16129 15079
rect 7116 15048 16129 15076
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 2317 14943 2375 14949
rect 2317 14940 2329 14943
rect 2280 14912 2329 14940
rect 2280 14900 2286 14912
rect 2317 14909 2329 14912
rect 2363 14909 2375 14943
rect 2317 14903 2375 14909
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14909 4859 14943
rect 4801 14903 4859 14909
rect 4816 14872 4844 14903
rect 4890 14900 4896 14952
rect 4948 14940 4954 14952
rect 5997 14943 6055 14949
rect 5997 14940 6009 14943
rect 4948 14912 6009 14940
rect 4948 14900 4954 14912
rect 5997 14909 6009 14912
rect 6043 14909 6055 14943
rect 5997 14903 6055 14909
rect 5445 14875 5503 14881
rect 4816 14844 5212 14872
rect 5184 14816 5212 14844
rect 5445 14841 5457 14875
rect 5491 14872 5503 14875
rect 6730 14872 6736 14884
rect 5491 14844 6736 14872
rect 5491 14841 5503 14844
rect 5445 14835 5503 14841
rect 6730 14832 6736 14844
rect 6788 14832 6794 14884
rect 6914 14832 6920 14884
rect 6972 14832 6978 14884
rect 7116 14816 7144 15048
rect 16117 15045 16129 15048
rect 16163 15045 16175 15079
rect 16117 15039 16175 15045
rect 7650 14968 7656 15020
rect 7708 15008 7714 15020
rect 16224 15008 16252 15116
rect 18598 15104 18604 15156
rect 18656 15144 18662 15156
rect 21453 15147 21511 15153
rect 21453 15144 21465 15147
rect 18656 15116 21465 15144
rect 18656 15104 18662 15116
rect 21453 15113 21465 15116
rect 21499 15144 21511 15147
rect 21499 15116 23336 15144
rect 21499 15113 21511 15116
rect 21453 15107 21511 15113
rect 17034 15076 17040 15088
rect 16684 15048 17040 15076
rect 16684 15017 16712 15048
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 17310 15036 17316 15088
rect 17368 15076 17374 15088
rect 21269 15079 21327 15085
rect 21269 15076 21281 15079
rect 17368 15048 21281 15076
rect 17368 15036 17374 15048
rect 21269 15045 21281 15048
rect 21315 15045 21327 15079
rect 21269 15039 21327 15045
rect 22189 15079 22247 15085
rect 22189 15045 22201 15079
rect 22235 15045 22247 15079
rect 22189 15039 22247 15045
rect 16577 15011 16635 15017
rect 16577 15008 16589 15011
rect 7708 14980 16068 15008
rect 16224 14980 16589 15008
rect 7708 14968 7714 14980
rect 7745 14943 7803 14949
rect 7745 14909 7757 14943
rect 7791 14909 7803 14943
rect 7745 14903 7803 14909
rect 7760 14872 7788 14903
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8570 14940 8576 14952
rect 8067 14912 8576 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 8938 14900 8944 14952
rect 8996 14900 9002 14952
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 10192 14912 10701 14940
rect 10192 14900 10198 14912
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14909 13231 14943
rect 13173 14903 13231 14909
rect 8662 14872 8668 14884
rect 7760 14844 8668 14872
rect 8662 14832 8668 14844
rect 8720 14832 8726 14884
rect 8757 14875 8815 14881
rect 8757 14841 8769 14875
rect 8803 14872 8815 14875
rect 9490 14872 9496 14884
rect 8803 14844 9496 14872
rect 8803 14841 8815 14844
rect 8757 14835 8815 14841
rect 9490 14832 9496 14844
rect 9548 14832 9554 14884
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 9861 14875 9919 14881
rect 9861 14872 9873 14875
rect 9732 14844 9873 14872
rect 9732 14832 9738 14844
rect 9861 14841 9873 14844
rect 9907 14841 9919 14875
rect 9861 14835 9919 14841
rect 11333 14875 11391 14881
rect 11333 14841 11345 14875
rect 11379 14872 11391 14875
rect 11974 14872 11980 14884
rect 11379 14844 11980 14872
rect 11379 14841 11391 14844
rect 11333 14835 11391 14841
rect 11974 14832 11980 14844
rect 12032 14832 12038 14884
rect 13188 14872 13216 14903
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13320 14912 13553 14940
rect 13320 14900 13326 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14909 13875 14943
rect 16040 14940 16068 14980
rect 16577 14977 16589 14980
rect 16623 14977 16635 15011
rect 16577 14971 16635 14977
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 22204 15008 22232 15039
rect 22278 15036 22284 15088
rect 22336 15076 22342 15088
rect 22833 15079 22891 15085
rect 22833 15076 22845 15079
rect 22336 15048 22845 15076
rect 22336 15036 22342 15048
rect 22833 15045 22845 15048
rect 22879 15045 22891 15079
rect 22833 15039 22891 15045
rect 16816 14980 22232 15008
rect 16816 14968 16822 14980
rect 16850 14940 16856 14952
rect 16040 14912 16856 14940
rect 13817 14903 13875 14909
rect 13832 14872 13860 14903
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 17678 14900 17684 14952
rect 17736 14940 17742 14952
rect 17773 14943 17831 14949
rect 17773 14940 17785 14943
rect 17736 14912 17785 14940
rect 17736 14900 17742 14912
rect 17773 14909 17785 14912
rect 17819 14909 17831 14943
rect 17773 14903 17831 14909
rect 18414 14900 18420 14952
rect 18472 14940 18478 14952
rect 18693 14943 18751 14949
rect 18693 14940 18705 14943
rect 18472 14912 18705 14940
rect 18472 14900 18478 14912
rect 18693 14909 18705 14912
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 19150 14900 19156 14952
rect 19208 14940 19214 14952
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 19208 14912 19441 14940
rect 19208 14900 19214 14912
rect 19429 14909 19441 14912
rect 19475 14909 19487 14943
rect 19429 14903 19487 14909
rect 20070 14900 20076 14952
rect 20128 14900 20134 14952
rect 20162 14900 20168 14952
rect 20220 14940 20226 14952
rect 20349 14943 20407 14949
rect 20349 14940 20361 14943
rect 20220 14912 20361 14940
rect 20220 14900 20226 14912
rect 20349 14909 20361 14912
rect 20395 14909 20407 14943
rect 20349 14903 20407 14909
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20680 14912 20913 14940
rect 20680 14900 20686 14912
rect 20901 14909 20913 14912
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 21358 14900 21364 14952
rect 21416 14900 21422 14952
rect 21450 14900 21456 14952
rect 21508 14940 21514 14952
rect 21729 14943 21787 14949
rect 21729 14940 21741 14943
rect 21508 14912 21741 14940
rect 21508 14900 21514 14912
rect 21729 14909 21741 14912
rect 21775 14909 21787 14943
rect 21729 14903 21787 14909
rect 22005 14943 22063 14949
rect 22005 14909 22017 14943
rect 22051 14909 22063 14943
rect 22005 14903 22063 14909
rect 13188 14844 13860 14872
rect 13832 14816 13860 14844
rect 16485 14875 16543 14881
rect 16485 14841 16497 14875
rect 16531 14872 16543 14875
rect 18230 14872 18236 14884
rect 16531 14844 18236 14872
rect 16531 14841 16543 14844
rect 16485 14835 16543 14841
rect 18230 14832 18236 14844
rect 18288 14872 18294 14884
rect 21376 14872 21404 14900
rect 22020 14872 22048 14903
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 22152 14912 22385 14940
rect 22152 14900 22158 14912
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 22830 14900 22836 14952
rect 22888 14940 22894 14952
rect 23017 14943 23075 14949
rect 23017 14940 23029 14943
rect 22888 14912 23029 14940
rect 22888 14900 22894 14912
rect 23017 14909 23029 14912
rect 23063 14909 23075 14943
rect 23017 14903 23075 14909
rect 18288 14844 20760 14872
rect 21376 14844 22048 14872
rect 18288 14832 18294 14844
rect 2498 14764 2504 14816
rect 2556 14804 2562 14816
rect 2961 14807 3019 14813
rect 2961 14804 2973 14807
rect 2556 14776 2973 14804
rect 2556 14764 2562 14776
rect 2961 14773 2973 14776
rect 3007 14773 3019 14807
rect 2961 14767 3019 14773
rect 5166 14764 5172 14816
rect 5224 14764 5230 14816
rect 7098 14764 7104 14816
rect 7156 14764 7162 14816
rect 7926 14764 7932 14816
rect 7984 14764 7990 14816
rect 11882 14764 11888 14816
rect 11940 14804 11946 14816
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 11940 14776 13093 14804
rect 11940 14764 11946 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13081 14767 13139 14773
rect 13814 14764 13820 14816
rect 13872 14764 13878 14816
rect 17957 14807 18015 14813
rect 17957 14773 17969 14807
rect 18003 14804 18015 14807
rect 18506 14804 18512 14816
rect 18003 14776 18512 14804
rect 18003 14773 18015 14776
rect 17957 14767 18015 14773
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 18874 14764 18880 14816
rect 18932 14764 18938 14816
rect 19242 14764 19248 14816
rect 19300 14764 19306 14816
rect 19889 14807 19947 14813
rect 19889 14773 19901 14807
rect 19935 14804 19947 14807
rect 19978 14804 19984 14816
rect 19935 14776 19984 14804
rect 19935 14773 19947 14776
rect 19889 14767 19947 14773
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 20162 14764 20168 14816
rect 20220 14764 20226 14816
rect 20732 14813 20760 14844
rect 20717 14807 20775 14813
rect 20717 14773 20729 14807
rect 20763 14773 20775 14807
rect 20717 14767 20775 14773
rect 21542 14764 21548 14816
rect 21600 14804 21606 14816
rect 21821 14807 21879 14813
rect 21821 14804 21833 14807
rect 21600 14776 21833 14804
rect 21600 14764 21606 14776
rect 21821 14773 21833 14776
rect 21867 14773 21879 14807
rect 23308 14804 23336 15116
rect 23308 14776 23428 14804
rect 21821 14767 21879 14773
rect 552 14714 23368 14736
rect 552 14662 4366 14714
rect 4418 14662 4430 14714
rect 4482 14662 4494 14714
rect 4546 14662 4558 14714
rect 4610 14662 4622 14714
rect 4674 14662 4686 14714
rect 4738 14662 10366 14714
rect 10418 14662 10430 14714
rect 10482 14662 10494 14714
rect 10546 14662 10558 14714
rect 10610 14662 10622 14714
rect 10674 14662 10686 14714
rect 10738 14662 16366 14714
rect 16418 14662 16430 14714
rect 16482 14662 16494 14714
rect 16546 14662 16558 14714
rect 16610 14662 16622 14714
rect 16674 14662 16686 14714
rect 16738 14662 22366 14714
rect 22418 14662 22430 14714
rect 22482 14662 22494 14714
rect 22546 14662 22558 14714
rect 22610 14662 22622 14714
rect 22674 14662 22686 14714
rect 22738 14662 23368 14714
rect 552 14640 23368 14662
rect 2222 14560 2228 14612
rect 2280 14560 2286 14612
rect 2406 14560 2412 14612
rect 2464 14600 2470 14612
rect 4890 14600 4896 14612
rect 2464 14572 4896 14600
rect 2464 14560 2470 14572
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 5629 14603 5687 14609
rect 5629 14569 5641 14603
rect 5675 14569 5687 14603
rect 5629 14563 5687 14569
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 6638 14600 6644 14612
rect 6227 14572 6644 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 5644 14532 5672 14563
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 6733 14603 6791 14609
rect 6733 14569 6745 14603
rect 6779 14600 6791 14603
rect 7650 14600 7656 14612
rect 6779 14572 7656 14600
rect 6779 14569 6791 14572
rect 6733 14563 6791 14569
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 7926 14560 7932 14612
rect 7984 14560 7990 14612
rect 8938 14560 8944 14612
rect 8996 14560 9002 14612
rect 10229 14603 10287 14609
rect 10229 14569 10241 14603
rect 10275 14600 10287 14603
rect 10413 14603 10471 14609
rect 10275 14572 10364 14600
rect 10275 14569 10287 14572
rect 10229 14563 10287 14569
rect 6086 14532 6092 14544
rect 2608 14504 4292 14532
rect 5644 14504 6092 14532
rect 1112 14467 1170 14473
rect 1112 14433 1124 14467
rect 1158 14464 1170 14467
rect 1158 14436 1900 14464
rect 1158 14433 1170 14436
rect 1112 14427 1170 14433
rect 845 14399 903 14405
rect 845 14365 857 14399
rect 891 14365 903 14399
rect 845 14359 903 14365
rect 860 14260 888 14359
rect 1872 14272 1900 14436
rect 2498 14424 2504 14476
rect 2556 14424 2562 14476
rect 2608 14473 2636 14504
rect 2866 14473 2872 14476
rect 2593 14467 2651 14473
rect 2593 14433 2605 14467
rect 2639 14433 2651 14467
rect 2593 14427 2651 14433
rect 2860 14427 2872 14473
rect 2866 14424 2872 14427
rect 2924 14424 2930 14476
rect 4264 14473 4292 14504
rect 6086 14492 6092 14504
rect 6144 14492 6150 14544
rect 7944 14532 7972 14560
rect 7944 14504 8156 14532
rect 4249 14467 4307 14473
rect 4249 14433 4261 14467
rect 4295 14464 4307 14467
rect 4338 14464 4344 14476
rect 4295 14436 4344 14464
rect 4295 14433 4307 14436
rect 4249 14427 4307 14433
rect 4338 14424 4344 14436
rect 4396 14424 4402 14476
rect 4516 14467 4574 14473
rect 4516 14433 4528 14467
rect 4562 14464 4574 14467
rect 4562 14436 5304 14464
rect 4562 14433 4574 14436
rect 4516 14427 4574 14433
rect 5276 14328 5304 14436
rect 5350 14424 5356 14476
rect 5408 14424 5414 14476
rect 6546 14424 6552 14476
rect 6604 14424 6610 14476
rect 6641 14467 6699 14473
rect 6641 14433 6653 14467
rect 6687 14433 6699 14467
rect 6641 14427 6699 14433
rect 5368 14396 5396 14424
rect 6656 14396 6684 14427
rect 6730 14424 6736 14476
rect 6788 14464 6794 14476
rect 6825 14467 6883 14473
rect 6825 14464 6837 14467
rect 6788 14436 6837 14464
rect 6788 14424 6794 14436
rect 6825 14433 6837 14436
rect 6871 14433 6883 14467
rect 6825 14427 6883 14433
rect 7098 14424 7104 14476
rect 7156 14424 7162 14476
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14464 7619 14467
rect 8018 14464 8024 14476
rect 7607 14436 8024 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8128 14405 8156 14504
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14464 8263 14467
rect 8754 14464 8760 14476
rect 8251 14436 8760 14464
rect 8251 14433 8263 14436
rect 8205 14427 8263 14433
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 5368 14368 6684 14396
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14365 8171 14399
rect 8956 14396 8984 14560
rect 10336 14532 10364 14572
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10686 14600 10692 14612
rect 10459 14572 10692 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10686 14560 10692 14572
rect 10744 14600 10750 14612
rect 11057 14603 11115 14609
rect 11057 14600 11069 14603
rect 10744 14572 11069 14600
rect 10744 14560 10750 14572
rect 11057 14569 11069 14572
rect 11103 14569 11115 14603
rect 14734 14600 14740 14612
rect 11057 14563 11115 14569
rect 12084 14572 14740 14600
rect 10965 14535 11023 14541
rect 10965 14532 10977 14535
rect 10336 14504 10977 14532
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 9140 14436 9505 14464
rect 9140 14408 9168 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 10336 14473 10364 14504
rect 10965 14501 10977 14504
rect 11011 14501 11023 14535
rect 10965 14495 11023 14501
rect 12084 14473 12112 14572
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16577 14603 16635 14609
rect 16577 14600 16589 14603
rect 15804 14572 16589 14600
rect 15804 14560 15810 14572
rect 16577 14569 16589 14572
rect 16623 14569 16635 14603
rect 16577 14563 16635 14569
rect 16942 14560 16948 14612
rect 17000 14560 17006 14612
rect 18046 14560 18052 14612
rect 18104 14560 18110 14612
rect 18414 14560 18420 14612
rect 18472 14600 18478 14612
rect 19242 14600 19248 14612
rect 18472 14572 19248 14600
rect 18472 14560 18478 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 21085 14603 21143 14609
rect 21085 14569 21097 14603
rect 21131 14600 21143 14603
rect 21450 14600 21456 14612
rect 21131 14572 21456 14600
rect 21131 14569 21143 14572
rect 21085 14563 21143 14569
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 21545 14603 21603 14609
rect 21545 14569 21557 14603
rect 21591 14600 21603 14603
rect 23017 14603 23075 14609
rect 21591 14572 21772 14600
rect 21591 14569 21603 14572
rect 21545 14563 21603 14569
rect 17402 14532 17408 14544
rect 12360 14504 13860 14532
rect 12360 14473 12388 14504
rect 13832 14473 13860 14504
rect 14844 14504 17408 14532
rect 10321 14467 10379 14473
rect 10321 14464 10333 14467
rect 10284 14436 10333 14464
rect 10284 14424 10290 14436
rect 10321 14433 10333 14436
rect 10367 14433 10379 14467
rect 10321 14427 10379 14433
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14433 10655 14467
rect 10597 14427 10655 14433
rect 12069 14467 12127 14473
rect 12069 14433 12081 14467
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14433 12403 14467
rect 12601 14467 12659 14473
rect 12601 14464 12613 14467
rect 12345 14427 12403 14433
rect 12452 14436 12613 14464
rect 8113 14359 8171 14365
rect 8404 14368 8984 14396
rect 6917 14331 6975 14337
rect 6917 14328 6929 14331
rect 5276 14300 6929 14328
rect 6917 14297 6929 14300
rect 6963 14297 6975 14331
rect 6917 14291 6975 14297
rect 1026 14260 1032 14272
rect 860 14232 1032 14260
rect 1026 14220 1032 14232
rect 1084 14220 1090 14272
rect 1854 14220 1860 14272
rect 1912 14220 1918 14272
rect 3973 14263 4031 14269
rect 3973 14229 3985 14263
rect 4019 14260 4031 14263
rect 4246 14260 4252 14272
rect 4019 14232 4252 14260
rect 4019 14229 4031 14232
rect 3973 14223 4031 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 6178 14220 6184 14272
rect 6236 14260 6242 14272
rect 6365 14263 6423 14269
rect 6365 14260 6377 14263
rect 6236 14232 6377 14260
rect 6236 14220 6242 14232
rect 6365 14229 6377 14232
rect 6411 14229 6423 14263
rect 7668 14260 7696 14359
rect 7929 14331 7987 14337
rect 7929 14297 7941 14331
rect 7975 14328 7987 14331
rect 8404 14328 8432 14368
rect 9122 14356 9128 14408
rect 9180 14356 9186 14408
rect 9306 14356 9312 14408
rect 9364 14356 9370 14408
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 9723 14368 9781 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 9769 14365 9781 14368
rect 9815 14396 9827 14399
rect 10612 14396 10640 14427
rect 11333 14399 11391 14405
rect 11333 14396 11345 14399
rect 9815 14368 11345 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 11333 14365 11345 14368
rect 11379 14365 11391 14399
rect 12452 14396 12480 14436
rect 12601 14433 12613 14436
rect 12647 14433 12659 14467
rect 12601 14427 12659 14433
rect 13817 14467 13875 14473
rect 13817 14433 13829 14467
rect 13863 14433 13875 14467
rect 13817 14427 13875 14433
rect 14084 14467 14142 14473
rect 14084 14433 14096 14467
rect 14130 14464 14142 14467
rect 14550 14464 14556 14476
rect 14130 14436 14556 14464
rect 14130 14433 14142 14436
rect 14084 14427 14142 14433
rect 11333 14359 11391 14365
rect 12268 14368 12480 14396
rect 7975 14300 8432 14328
rect 7975 14297 7987 14300
rect 7929 14291 7987 14297
rect 10042 14288 10048 14340
rect 10100 14288 10106 14340
rect 12268 14337 12296 14368
rect 12253 14331 12311 14337
rect 12253 14297 12265 14331
rect 12299 14297 12311 14331
rect 12253 14291 12311 14297
rect 8110 14260 8116 14272
rect 7668 14232 8116 14260
rect 6365 14223 6423 14229
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 8481 14263 8539 14269
rect 8481 14229 8493 14263
rect 8527 14260 8539 14263
rect 9306 14260 9312 14272
rect 8527 14232 9312 14260
rect 8527 14229 8539 14232
rect 8481 14223 8539 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 10778 14220 10784 14272
rect 10836 14220 10842 14272
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 11241 14263 11299 14269
rect 11241 14260 11253 14263
rect 10928 14232 11253 14260
rect 10928 14220 10934 14232
rect 11241 14229 11253 14232
rect 11287 14229 11299 14263
rect 11241 14223 11299 14229
rect 11330 14220 11336 14272
rect 11388 14220 11394 14272
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13725 14263 13783 14269
rect 13725 14260 13737 14263
rect 13320 14232 13737 14260
rect 13320 14220 13326 14232
rect 13725 14229 13737 14232
rect 13771 14229 13783 14263
rect 13832 14260 13860 14427
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 14844 14260 14872 14504
rect 17402 14492 17408 14504
rect 17460 14532 17466 14544
rect 21744 14532 21772 14572
rect 23017 14569 23029 14603
rect 23063 14600 23075 14603
rect 23400 14600 23428 14776
rect 23063 14572 23428 14600
rect 23063 14569 23075 14572
rect 23017 14563 23075 14569
rect 21882 14535 21940 14541
rect 21882 14532 21894 14535
rect 17460 14504 21680 14532
rect 21744 14504 21894 14532
rect 17460 14492 17466 14504
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14464 15715 14467
rect 15703 14436 16436 14464
rect 15703 14433 15715 14436
rect 15657 14427 15715 14433
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 15473 14399 15531 14405
rect 15473 14396 15485 14399
rect 15252 14368 15485 14396
rect 15252 14356 15258 14368
rect 15473 14365 15485 14368
rect 15519 14365 15531 14399
rect 15473 14359 15531 14365
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14396 15991 14399
rect 16298 14396 16304 14408
rect 15979 14368 16304 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 16408 14396 16436 14436
rect 16482 14424 16488 14476
rect 16540 14424 16546 14476
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 16592 14436 17141 14464
rect 16592 14396 16620 14436
rect 17129 14433 17141 14436
rect 17175 14464 17187 14467
rect 17586 14464 17592 14476
rect 17175 14436 17592 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17586 14424 17592 14436
rect 17644 14464 17650 14476
rect 17681 14467 17739 14473
rect 17681 14464 17693 14467
rect 17644 14436 17693 14464
rect 17644 14424 17650 14436
rect 17681 14433 17693 14436
rect 17727 14433 17739 14467
rect 18230 14464 18236 14476
rect 17681 14427 17739 14433
rect 17880 14436 18236 14464
rect 16408 14368 16620 14396
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 17034 14396 17040 14408
rect 16807 14368 17040 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 17034 14356 17040 14368
rect 17092 14356 17098 14408
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14396 17463 14399
rect 17880 14396 17908 14436
rect 18230 14424 18236 14436
rect 18288 14424 18294 14476
rect 18598 14424 18604 14476
rect 18656 14464 18662 14476
rect 19720 14473 19748 14504
rect 19978 14473 19984 14476
rect 19153 14467 19211 14473
rect 19153 14464 19165 14467
rect 18656 14436 19165 14464
rect 18656 14424 18662 14436
rect 19153 14433 19165 14436
rect 19199 14433 19211 14467
rect 19153 14427 19211 14433
rect 19245 14467 19303 14473
rect 19245 14433 19257 14467
rect 19291 14433 19303 14467
rect 19245 14427 19303 14433
rect 19705 14467 19763 14473
rect 19705 14433 19717 14467
rect 19751 14433 19763 14467
rect 19972 14464 19984 14473
rect 19939 14436 19984 14464
rect 19705 14427 19763 14433
rect 19972 14427 19984 14436
rect 17451 14368 17908 14396
rect 17451 14365 17463 14368
rect 17405 14359 17463 14365
rect 17954 14356 17960 14408
rect 18012 14356 18018 14408
rect 18509 14399 18567 14405
rect 18509 14396 18521 14399
rect 18432 14368 18521 14396
rect 15838 14288 15844 14340
rect 15896 14288 15902 14340
rect 17126 14288 17132 14340
rect 17184 14288 17190 14340
rect 17494 14288 17500 14340
rect 17552 14288 17558 14340
rect 13832 14232 14872 14260
rect 15197 14263 15255 14269
rect 13725 14223 13783 14229
rect 15197 14229 15209 14263
rect 15243 14260 15255 14263
rect 15378 14260 15384 14272
rect 15243 14232 15384 14260
rect 15243 14229 15255 14232
rect 15197 14223 15255 14229
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 16114 14220 16120 14272
rect 16172 14220 16178 14272
rect 17144 14260 17172 14288
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 17144 14232 17325 14260
rect 17313 14229 17325 14232
rect 17359 14260 17371 14263
rect 17862 14260 17868 14272
rect 17359 14232 17868 14260
rect 17359 14229 17371 14232
rect 17313 14223 17371 14229
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 18432 14260 18460 14368
rect 18509 14365 18521 14368
rect 18555 14365 18567 14399
rect 18509 14359 18567 14365
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 18782 14396 18788 14408
rect 18739 14368 18788 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 18782 14356 18788 14368
rect 18840 14396 18846 14408
rect 18969 14399 19027 14405
rect 18969 14396 18981 14399
rect 18840 14368 18981 14396
rect 18840 14356 18846 14368
rect 18969 14365 18981 14368
rect 19015 14365 19027 14399
rect 19260 14396 19288 14427
rect 19978 14424 19984 14427
rect 20036 14424 20042 14476
rect 21652 14473 21680 14504
rect 21882 14501 21894 14504
rect 21928 14501 21940 14535
rect 21882 14495 21940 14501
rect 21361 14467 21419 14473
rect 21361 14464 21373 14467
rect 20732 14436 21373 14464
rect 18969 14359 19027 14365
rect 19168 14368 19288 14396
rect 18874 14288 18880 14340
rect 18932 14328 18938 14340
rect 19168 14328 19196 14368
rect 18932 14300 19196 14328
rect 18932 14288 18938 14300
rect 18598 14260 18604 14272
rect 18432 14232 18604 14260
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 19613 14263 19671 14269
rect 19613 14229 19625 14263
rect 19659 14260 19671 14263
rect 20732 14260 20760 14436
rect 21361 14433 21373 14436
rect 21407 14433 21419 14467
rect 21361 14427 21419 14433
rect 21637 14467 21695 14473
rect 21637 14433 21649 14467
rect 21683 14433 21695 14467
rect 21637 14427 21695 14433
rect 19659 14232 20760 14260
rect 19659 14229 19671 14232
rect 19613 14223 19671 14229
rect 552 14170 23368 14192
rect 552 14118 1366 14170
rect 1418 14118 1430 14170
rect 1482 14118 1494 14170
rect 1546 14118 1558 14170
rect 1610 14118 1622 14170
rect 1674 14118 1686 14170
rect 1738 14118 7366 14170
rect 7418 14118 7430 14170
rect 7482 14118 7494 14170
rect 7546 14118 7558 14170
rect 7610 14118 7622 14170
rect 7674 14118 7686 14170
rect 7738 14118 13366 14170
rect 13418 14118 13430 14170
rect 13482 14118 13494 14170
rect 13546 14118 13558 14170
rect 13610 14118 13622 14170
rect 13674 14118 13686 14170
rect 13738 14118 19366 14170
rect 19418 14118 19430 14170
rect 19482 14118 19494 14170
rect 19546 14118 19558 14170
rect 19610 14118 19622 14170
rect 19674 14118 19686 14170
rect 19738 14118 23368 14170
rect 552 14096 23368 14118
rect 1854 14016 1860 14068
rect 1912 14016 1918 14068
rect 2406 14016 2412 14068
rect 2464 14016 2470 14068
rect 2866 14016 2872 14068
rect 2924 14016 2930 14068
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 8481 14059 8539 14065
rect 8481 14056 8493 14059
rect 7892 14028 8493 14056
rect 7892 14016 7898 14028
rect 8481 14025 8493 14028
rect 8527 14025 8539 14059
rect 8481 14019 8539 14025
rect 8570 14016 8576 14068
rect 8628 14056 8634 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 8628 14028 9045 14056
rect 8628 14016 8634 14028
rect 9033 14025 9045 14028
rect 9079 14025 9091 14059
rect 9033 14019 9091 14025
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 10042 14056 10048 14068
rect 9815 14028 10048 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10870 14016 10876 14068
rect 10928 14016 10934 14068
rect 10965 14059 11023 14065
rect 10965 14025 10977 14059
rect 11011 14056 11023 14059
rect 11330 14056 11336 14068
rect 11011 14028 11336 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11532 14028 13124 14056
rect 2424 13920 2452 14016
rect 6270 13948 6276 14000
rect 6328 13988 6334 14000
rect 6365 13991 6423 13997
rect 6365 13988 6377 13991
rect 6328 13960 6377 13988
rect 6328 13948 6334 13960
rect 6365 13957 6377 13960
rect 6411 13988 6423 13991
rect 10502 13988 10508 14000
rect 6411 13960 10508 13988
rect 6411 13957 6423 13960
rect 6365 13951 6423 13957
rect 10502 13948 10508 13960
rect 10560 13948 10566 14000
rect 10597 13991 10655 13997
rect 10597 13957 10609 13991
rect 10643 13988 10655 13991
rect 10888 13988 10916 14016
rect 10643 13960 10916 13988
rect 10643 13957 10655 13960
rect 10597 13951 10655 13957
rect 2056 13892 2452 13920
rect 8849 13923 8907 13929
rect 1210 13812 1216 13864
rect 1268 13852 1274 13864
rect 2056 13861 2084 13892
rect 8849 13889 8861 13923
rect 8895 13920 8907 13923
rect 10321 13923 10379 13929
rect 8895 13892 9628 13920
rect 8895 13889 8907 13892
rect 8849 13883 8907 13889
rect 1857 13855 1915 13861
rect 1857 13852 1869 13855
rect 1268 13824 1869 13852
rect 1268 13812 1274 13824
rect 1857 13821 1869 13824
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 2130 13812 2136 13864
rect 2188 13812 2194 13864
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 1762 13744 1768 13796
rect 1820 13784 1826 13796
rect 2332 13784 2360 13815
rect 2682 13812 2688 13864
rect 2740 13812 2746 13864
rect 3878 13812 3884 13864
rect 3936 13852 3942 13864
rect 4338 13852 4344 13864
rect 3936 13824 4344 13852
rect 3936 13812 3942 13824
rect 4338 13812 4344 13824
rect 4396 13852 4402 13864
rect 6273 13855 6331 13861
rect 6273 13852 6285 13855
rect 4396 13824 6285 13852
rect 4396 13812 4402 13824
rect 6273 13821 6285 13824
rect 6319 13852 6331 13855
rect 6822 13852 6828 13864
rect 6319 13824 6828 13852
rect 6319 13821 6331 13824
rect 6273 13815 6331 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7742 13812 7748 13864
rect 7800 13852 7806 13864
rect 7837 13855 7895 13861
rect 7837 13852 7849 13855
rect 7800 13824 7849 13852
rect 7800 13812 7806 13824
rect 7837 13821 7849 13824
rect 7883 13821 7895 13855
rect 7837 13815 7895 13821
rect 8021 13855 8079 13861
rect 8021 13821 8033 13855
rect 8067 13852 8079 13855
rect 8202 13852 8208 13864
rect 8067 13824 8208 13852
rect 8067 13821 8079 13824
rect 8021 13815 8079 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8389 13855 8447 13861
rect 8389 13821 8401 13855
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 1820 13756 2360 13784
rect 6028 13787 6086 13793
rect 1820 13744 1826 13756
rect 6028 13753 6040 13787
rect 6074 13784 6086 13787
rect 6178 13784 6184 13796
rect 6074 13756 6184 13784
rect 6074 13753 6086 13756
rect 6028 13747 6086 13753
rect 6178 13744 6184 13756
rect 6236 13744 6242 13796
rect 6549 13787 6607 13793
rect 6549 13784 6561 13787
rect 6380 13756 6561 13784
rect 2501 13719 2559 13725
rect 2501 13685 2513 13719
rect 2547 13716 2559 13719
rect 2590 13716 2596 13728
rect 2547 13688 2596 13716
rect 2547 13685 2559 13688
rect 2501 13679 2559 13685
rect 2590 13676 2596 13688
rect 2648 13676 2654 13728
rect 4893 13719 4951 13725
rect 4893 13685 4905 13719
rect 4939 13716 4951 13719
rect 5534 13716 5540 13728
rect 4939 13688 5540 13716
rect 4939 13685 4951 13688
rect 4893 13679 4951 13685
rect 5534 13676 5540 13688
rect 5592 13716 5598 13728
rect 6380 13716 6408 13756
rect 6549 13753 6561 13756
rect 6595 13753 6607 13787
rect 6549 13747 6607 13753
rect 5592 13688 6408 13716
rect 8404 13716 8432 13815
rect 8570 13812 8576 13864
rect 8628 13852 8634 13864
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 8628 13824 8677 13852
rect 8628 13812 8634 13824
rect 8665 13821 8677 13824
rect 8711 13852 8723 13855
rect 8941 13855 8999 13861
rect 8941 13852 8953 13855
rect 8711 13824 8953 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 8941 13821 8953 13824
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 9180 13824 9260 13852
rect 9180 13812 9186 13824
rect 9232 13784 9260 13824
rect 9306 13812 9312 13864
rect 9364 13852 9370 13864
rect 9600 13852 9628 13892
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 10367 13892 10640 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 10229 13855 10287 13861
rect 10229 13852 10241 13855
rect 9364 13824 9536 13852
rect 9600 13824 10241 13852
rect 9364 13812 9370 13824
rect 9401 13787 9459 13793
rect 9401 13784 9413 13787
rect 9232 13756 9413 13784
rect 9401 13753 9413 13756
rect 9447 13753 9459 13787
rect 9508 13784 9536 13824
rect 10229 13821 10241 13824
rect 10275 13821 10287 13855
rect 10229 13815 10287 13821
rect 9585 13787 9643 13793
rect 9585 13784 9597 13787
rect 9508 13756 9597 13784
rect 9401 13747 9459 13753
rect 9585 13753 9597 13756
rect 9631 13753 9643 13787
rect 10612 13784 10640 13892
rect 10704 13861 10732 13960
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 11425 13991 11483 13997
rect 11425 13988 11437 13991
rect 11204 13960 11437 13988
rect 11204 13948 11210 13960
rect 11425 13957 11437 13960
rect 11471 13957 11483 13991
rect 11425 13951 11483 13957
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13920 11115 13923
rect 11532 13920 11560 14028
rect 11882 13948 11888 14000
rect 11940 13948 11946 14000
rect 11900 13920 11928 13948
rect 11103 13892 11560 13920
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 11532 13868 11560 13892
rect 11716 13892 11928 13920
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13821 10747 13855
rect 10689 13815 10747 13821
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10836 13824 10885 13852
rect 10836 13812 10842 13824
rect 10873 13821 10885 13824
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11422 13852 11428 13864
rect 11195 13824 11428 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 11532 13861 11566 13868
rect 11517 13855 11575 13861
rect 11517 13821 11529 13855
rect 11563 13821 11575 13855
rect 11517 13815 11575 13821
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 11716 13861 11744 13892
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11664 13824 11713 13852
rect 11664 13812 11670 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 12986 13852 12992 13864
rect 11701 13815 11759 13821
rect 11808 13824 12992 13852
rect 11808 13784 11836 13824
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13096 13861 13124 14028
rect 14550 14016 14556 14068
rect 14608 14016 14614 14068
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 16301 14059 16359 14065
rect 16301 14056 16313 14059
rect 16264 14028 16313 14056
rect 16264 14016 16270 14028
rect 16301 14025 16313 14028
rect 16347 14025 16359 14059
rect 16301 14019 16359 14025
rect 16850 14016 16856 14068
rect 16908 14016 16914 14068
rect 17586 14016 17592 14068
rect 17644 14016 17650 14068
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 18233 14059 18291 14065
rect 18233 14056 18245 14059
rect 17920 14028 18245 14056
rect 17920 14016 17926 14028
rect 18233 14025 18245 14028
rect 18279 14025 18291 14059
rect 18233 14019 18291 14025
rect 18414 14016 18420 14068
rect 18472 14016 18478 14068
rect 18598 14016 18604 14068
rect 18656 14056 18662 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 18656 14028 18889 14056
rect 18656 14016 18662 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 20070 14016 20076 14068
rect 20128 14016 20134 14068
rect 21450 14016 21456 14068
rect 21508 14016 21514 14068
rect 13725 13991 13783 13997
rect 13725 13957 13737 13991
rect 13771 13988 13783 13991
rect 14182 13988 14188 14000
rect 13771 13960 14188 13988
rect 13771 13957 13783 13960
rect 13725 13951 13783 13957
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 15378 13880 15384 13932
rect 15436 13880 15442 13932
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 15746 13920 15752 13932
rect 15703 13892 15752 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 15896 13892 16773 13920
rect 15896 13880 15902 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 10612 13756 11836 13784
rect 13096 13784 13124 13815
rect 13170 13812 13176 13864
rect 13228 13812 13234 13864
rect 13262 13812 13268 13864
rect 13320 13812 13326 13864
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14642 13852 14648 13864
rect 14047 13824 14648 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 14737 13855 14795 13861
rect 14737 13821 14749 13855
rect 14783 13852 14795 13855
rect 16114 13852 16120 13864
rect 14783 13824 16120 13852
rect 14783 13821 14795 13824
rect 14737 13815 14795 13821
rect 16114 13812 16120 13824
rect 16172 13812 16178 13864
rect 16868 13852 16896 14016
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13920 17003 13923
rect 17034 13920 17040 13932
rect 16991 13892 17040 13920
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 17034 13880 17040 13892
rect 17092 13920 17098 13932
rect 17604 13920 17632 14016
rect 18325 13923 18383 13929
rect 17092 13892 17540 13920
rect 17604 13892 18092 13920
rect 17092 13880 17098 13892
rect 17313 13855 17371 13861
rect 17313 13852 17325 13855
rect 16868 13824 17325 13852
rect 17313 13821 17325 13824
rect 17359 13852 17371 13855
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 17359 13824 17417 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 17512 13852 17540 13892
rect 17512 13824 17724 13852
rect 17405 13815 17463 13821
rect 17696 13784 17724 13824
rect 17862 13812 17868 13864
rect 17920 13812 17926 13864
rect 18064 13861 18092 13892
rect 18325 13889 18337 13923
rect 18371 13920 18383 13923
rect 18432 13920 18460 14016
rect 18371 13892 18460 13920
rect 19076 13960 19656 13988
rect 18371 13889 18383 13892
rect 18325 13883 18383 13889
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18690 13812 18696 13864
rect 18748 13852 18754 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18748 13824 18889 13852
rect 18748 13812 18754 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 18966 13812 18972 13864
rect 19024 13852 19030 13864
rect 19076 13861 19104 13960
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19628 13929 19656 13960
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19208 13892 19441 13920
rect 19208 13880 19214 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13920 19671 13923
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 19659 13892 20637 13920
rect 19659 13889 19671 13892
rect 19613 13883 19671 13889
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 19024 13824 19073 13852
rect 19024 13812 19030 13824
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19168 13784 19196 13880
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13852 19763 13855
rect 20162 13852 20168 13864
rect 19751 13824 20168 13852
rect 19751 13821 19763 13824
rect 19705 13815 19763 13821
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13852 20867 13855
rect 21468 13852 21496 14016
rect 20855 13824 21496 13852
rect 20855 13821 20867 13824
rect 20809 13815 20867 13821
rect 13096 13756 14044 13784
rect 9585 13747 9643 13753
rect 9950 13716 9956 13728
rect 8404 13688 9956 13716
rect 5592 13676 5598 13688
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 11609 13719 11667 13725
rect 11609 13716 11621 13719
rect 11020 13688 11621 13716
rect 11020 13676 11026 13688
rect 11609 13685 11621 13688
rect 11655 13685 11667 13719
rect 14016 13716 14044 13756
rect 16500 13756 17356 13784
rect 17696 13756 19196 13784
rect 16500 13716 16528 13756
rect 17328 13728 17356 13756
rect 14016 13688 16528 13716
rect 16669 13719 16727 13725
rect 11609 13679 11667 13685
rect 16669 13685 16681 13719
rect 16715 13716 16727 13719
rect 16758 13716 16764 13728
rect 16715 13688 16764 13716
rect 16715 13685 16727 13688
rect 16669 13679 16727 13685
rect 16758 13676 16764 13688
rect 16816 13676 16822 13728
rect 16850 13676 16856 13728
rect 16908 13716 16914 13728
rect 17129 13719 17187 13725
rect 17129 13716 17141 13719
rect 16908 13688 17141 13716
rect 16908 13676 16914 13688
rect 17129 13685 17141 13688
rect 17175 13685 17187 13719
rect 17129 13679 17187 13685
rect 17310 13676 17316 13728
rect 17368 13676 17374 13728
rect 18690 13676 18696 13728
rect 18748 13676 18754 13728
rect 552 13626 23368 13648
rect 552 13574 4366 13626
rect 4418 13574 4430 13626
rect 4482 13574 4494 13626
rect 4546 13574 4558 13626
rect 4610 13574 4622 13626
rect 4674 13574 4686 13626
rect 4738 13574 10366 13626
rect 10418 13574 10430 13626
rect 10482 13574 10494 13626
rect 10546 13574 10558 13626
rect 10610 13574 10622 13626
rect 10674 13574 10686 13626
rect 10738 13574 16366 13626
rect 16418 13574 16430 13626
rect 16482 13574 16494 13626
rect 16546 13574 16558 13626
rect 16610 13574 16622 13626
rect 16674 13574 16686 13626
rect 16738 13574 22366 13626
rect 22418 13574 22430 13626
rect 22482 13574 22494 13626
rect 22546 13574 22558 13626
rect 22610 13574 22622 13626
rect 22674 13574 22686 13626
rect 22738 13574 23368 13626
rect 552 13552 23368 13574
rect 3878 13512 3884 13524
rect 2332 13484 3884 13512
rect 1118 13404 1124 13456
rect 1176 13444 1182 13456
rect 1857 13447 1915 13453
rect 1857 13444 1869 13447
rect 1176 13416 1869 13444
rect 1176 13404 1182 13416
rect 1857 13413 1869 13416
rect 1903 13413 1915 13447
rect 1857 13407 1915 13413
rect 2073 13447 2131 13453
rect 2073 13413 2085 13447
rect 2119 13444 2131 13447
rect 2222 13444 2228 13456
rect 2119 13416 2228 13444
rect 2119 13413 2131 13416
rect 2073 13407 2131 13413
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 1026 13336 1032 13388
rect 1084 13376 1090 13388
rect 2332 13385 2360 13484
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 7837 13515 7895 13521
rect 7837 13481 7849 13515
rect 7883 13512 7895 13515
rect 8570 13512 8576 13524
rect 7883 13484 8576 13512
rect 7883 13481 7895 13484
rect 7837 13475 7895 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 8680 13484 12434 13512
rect 2590 13453 2596 13456
rect 2584 13407 2596 13453
rect 2648 13444 2654 13456
rect 6914 13444 6920 13456
rect 2648 13416 2684 13444
rect 3436 13416 6920 13444
rect 2590 13404 2596 13407
rect 2648 13404 2654 13416
rect 2317 13379 2375 13385
rect 2317 13376 2329 13379
rect 1084 13348 2329 13376
rect 1084 13336 1090 13348
rect 2317 13345 2329 13348
rect 2363 13345 2375 13379
rect 2317 13339 2375 13345
rect 3436 13184 3464 13416
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 7742 13444 7748 13456
rect 7668 13416 7748 13444
rect 6086 13336 6092 13388
rect 6144 13376 6150 13388
rect 7668 13385 7696 13416
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 8680 13444 8708 13484
rect 8168 13416 8708 13444
rect 8168 13404 8174 13416
rect 10226 13404 10232 13456
rect 10284 13444 10290 13456
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 10284 13416 10425 13444
rect 10284 13404 10290 13416
rect 6273 13379 6331 13385
rect 6273 13376 6285 13379
rect 6144 13348 6285 13376
rect 6144 13336 6150 13348
rect 6273 13345 6285 13348
rect 6319 13376 6331 13379
rect 6365 13379 6423 13385
rect 6365 13376 6377 13379
rect 6319 13348 6377 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 6365 13345 6377 13348
rect 6411 13345 6423 13379
rect 6365 13339 6423 13345
rect 7653 13379 7711 13385
rect 7653 13345 7665 13379
rect 7699 13345 7711 13379
rect 7653 13339 7711 13345
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13345 7895 13379
rect 7837 13339 7895 13345
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 5810 13308 5816 13320
rect 4212 13280 5816 13308
rect 4212 13268 4218 13280
rect 5810 13268 5816 13280
rect 5868 13308 5874 13320
rect 7668 13308 7696 13339
rect 5868 13280 7696 13308
rect 7852 13308 7880 13339
rect 8754 13336 8760 13388
rect 8812 13336 8818 13388
rect 10336 13385 10364 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 12066 13444 12072 13456
rect 10413 13407 10471 13413
rect 10980 13416 12072 13444
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10597 13379 10655 13385
rect 10367 13348 10401 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10597 13345 10609 13379
rect 10643 13376 10655 13379
rect 10778 13376 10784 13388
rect 10643 13348 10784 13376
rect 10643 13345 10655 13348
rect 10597 13339 10655 13345
rect 8202 13308 8208 13320
rect 7852 13280 8208 13308
rect 5868 13268 5874 13280
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 8772 13308 8800 13336
rect 9306 13308 9312 13320
rect 8772 13280 9312 13308
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 10152 13308 10180 13339
rect 10612 13308 10640 13339
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 9640 13280 10640 13308
rect 9640 13268 9646 13280
rect 5902 13200 5908 13252
rect 5960 13240 5966 13252
rect 10980 13240 11008 13416
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 12406 13444 12434 13484
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 17494 13512 17500 13524
rect 13136 13484 17500 13512
rect 13136 13472 13142 13484
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 17770 13472 17776 13524
rect 17828 13512 17834 13524
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17828 13484 17877 13512
rect 17828 13472 17834 13484
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 17865 13475 17923 13481
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 18414 13512 18420 13524
rect 18104 13484 18420 13512
rect 18104 13472 18110 13484
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 18506 13472 18512 13524
rect 18564 13472 18570 13524
rect 18690 13472 18696 13524
rect 18748 13472 18754 13524
rect 18877 13515 18935 13521
rect 18877 13481 18889 13515
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 16117 13447 16175 13453
rect 12406 13416 16068 13444
rect 11146 13336 11152 13388
rect 11204 13336 11210 13388
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 5960 13212 11008 13240
rect 5960 13200 5966 13212
rect 2038 13132 2044 13184
rect 2096 13132 2102 13184
rect 2225 13175 2283 13181
rect 2225 13141 2237 13175
rect 2271 13172 2283 13175
rect 2682 13172 2688 13184
rect 2271 13144 2688 13172
rect 2271 13141 2283 13144
rect 2225 13135 2283 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 3418 13132 3424 13184
rect 3476 13132 3482 13184
rect 3697 13175 3755 13181
rect 3697 13141 3709 13175
rect 3743 13172 3755 13175
rect 5350 13172 5356 13184
rect 3743 13144 5356 13172
rect 3743 13141 3755 13144
rect 3697 13135 3755 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 6086 13132 6092 13184
rect 6144 13132 6150 13184
rect 6454 13132 6460 13184
rect 6512 13132 6518 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 8018 13172 8024 13184
rect 6972 13144 8024 13172
rect 6972 13132 6978 13144
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8941 13175 8999 13181
rect 8941 13141 8953 13175
rect 8987 13172 8999 13175
rect 9950 13172 9956 13184
rect 8987 13144 9956 13172
rect 8987 13141 8999 13144
rect 8941 13135 8999 13141
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 10686 13172 10692 13184
rect 10275 13144 10692 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 10781 13175 10839 13181
rect 10781 13141 10793 13175
rect 10827 13172 10839 13175
rect 10870 13172 10876 13184
rect 10827 13144 10876 13172
rect 10827 13141 10839 13144
rect 10781 13135 10839 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11072 13172 11100 13271
rect 11146 13200 11152 13252
rect 11204 13240 11210 13252
rect 11425 13243 11483 13249
rect 11425 13240 11437 13243
rect 11204 13212 11437 13240
rect 11204 13200 11210 13212
rect 11425 13209 11437 13212
rect 11471 13209 11483 13243
rect 11425 13203 11483 13209
rect 11514 13200 11520 13252
rect 11572 13240 11578 13252
rect 11716 13240 11744 13271
rect 11790 13268 11796 13320
rect 11848 13308 11854 13320
rect 15930 13308 15936 13320
rect 11848 13280 15936 13308
rect 11848 13268 11854 13280
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16040 13308 16068 13416
rect 16117 13413 16129 13447
rect 16163 13444 16175 13447
rect 17954 13444 17960 13456
rect 16163 13416 17960 13444
rect 16163 13413 16175 13416
rect 16117 13407 16175 13413
rect 17954 13404 17960 13416
rect 18012 13404 18018 13456
rect 18708 13444 18736 13472
rect 18064 13416 18736 13444
rect 18892 13444 18920 13475
rect 19150 13472 19156 13524
rect 19208 13472 19214 13524
rect 21545 13515 21603 13521
rect 21545 13481 21557 13515
rect 21591 13481 21603 13515
rect 21545 13475 21603 13481
rect 21450 13444 21456 13456
rect 18892 13416 20024 13444
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 16850 13376 16856 13388
rect 16347 13348 16856 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 18064 13385 18092 13416
rect 17129 13379 17187 13385
rect 17129 13345 17141 13379
rect 17175 13376 17187 13379
rect 17773 13379 17831 13385
rect 17175 13348 17724 13376
rect 17175 13345 17187 13348
rect 17129 13339 17187 13345
rect 16577 13311 16635 13317
rect 16040 13280 16436 13308
rect 16408 13252 16436 13280
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 16758 13308 16764 13320
rect 16623 13280 16764 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 16758 13268 16764 13280
rect 16816 13308 16822 13320
rect 17696 13308 17724 13348
rect 17773 13345 17785 13379
rect 17819 13376 17831 13379
rect 18049 13379 18107 13385
rect 18049 13376 18061 13379
rect 17819 13348 18061 13376
rect 17819 13345 17831 13348
rect 17773 13339 17831 13345
rect 18049 13345 18061 13348
rect 18095 13345 18107 13379
rect 18506 13376 18512 13388
rect 18049 13339 18107 13345
rect 18156 13348 18512 13376
rect 18156 13308 18184 13348
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 19245 13379 19303 13385
rect 19245 13345 19257 13379
rect 19291 13376 19303 13379
rect 19794 13376 19800 13388
rect 19291 13348 19800 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 19794 13336 19800 13348
rect 19852 13336 19858 13388
rect 19996 13385 20024 13416
rect 20180 13416 21456 13444
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 16816 13280 17172 13308
rect 17696 13280 18184 13308
rect 16816 13268 16822 13280
rect 11572 13212 14504 13240
rect 11572 13200 11578 13212
rect 14476 13184 14504 13212
rect 16390 13200 16396 13252
rect 16448 13200 16454 13252
rect 16485 13243 16543 13249
rect 16485 13209 16497 13243
rect 16531 13240 16543 13243
rect 17144 13240 17172 13280
rect 18322 13268 18328 13320
rect 18380 13268 18386 13320
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 20180 13308 20208 13416
rect 21450 13404 21456 13416
rect 21508 13404 21514 13456
rect 21560 13444 21588 13475
rect 21882 13447 21940 13453
rect 21882 13444 21894 13447
rect 21560 13416 21894 13444
rect 21882 13413 21894 13416
rect 21928 13413 21940 13447
rect 21882 13407 21940 13413
rect 21358 13336 21364 13388
rect 21416 13336 21422 13388
rect 18472 13280 20208 13308
rect 18472 13268 18478 13280
rect 20254 13268 20260 13320
rect 20312 13308 20318 13320
rect 21637 13311 21695 13317
rect 21637 13308 21649 13311
rect 20312 13280 21649 13308
rect 20312 13268 20318 13280
rect 21637 13277 21649 13280
rect 21683 13277 21695 13311
rect 21637 13271 21695 13277
rect 21542 13240 21548 13252
rect 16531 13212 17080 13240
rect 17144 13212 21548 13240
rect 16531 13209 16543 13212
rect 16485 13203 16543 13209
rect 12710 13172 12716 13184
rect 11072 13144 12716 13172
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 17052 13181 17080 13212
rect 21542 13200 21548 13212
rect 21600 13200 21606 13252
rect 16669 13175 16727 13181
rect 16669 13172 16681 13175
rect 14516 13144 16681 13172
rect 14516 13132 14522 13144
rect 16669 13141 16681 13144
rect 16715 13141 16727 13175
rect 16669 13135 16727 13141
rect 17037 13175 17095 13181
rect 17037 13141 17049 13175
rect 17083 13172 17095 13175
rect 17586 13172 17592 13184
rect 17083 13144 17592 13172
rect 17083 13141 17095 13144
rect 17037 13135 17095 13141
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 20165 13175 20223 13181
rect 20165 13141 20177 13175
rect 20211 13172 20223 13175
rect 20438 13172 20444 13184
rect 20211 13144 20444 13172
rect 20211 13141 20223 13144
rect 20165 13135 20223 13141
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 23017 13175 23075 13181
rect 23017 13141 23029 13175
rect 23063 13172 23075 13175
rect 23063 13144 23428 13172
rect 23063 13141 23075 13144
rect 23017 13135 23075 13141
rect 552 13082 23368 13104
rect 552 13030 1366 13082
rect 1418 13030 1430 13082
rect 1482 13030 1494 13082
rect 1546 13030 1558 13082
rect 1610 13030 1622 13082
rect 1674 13030 1686 13082
rect 1738 13030 7366 13082
rect 7418 13030 7430 13082
rect 7482 13030 7494 13082
rect 7546 13030 7558 13082
rect 7610 13030 7622 13082
rect 7674 13030 7686 13082
rect 7738 13030 13366 13082
rect 13418 13030 13430 13082
rect 13482 13030 13494 13082
rect 13546 13030 13558 13082
rect 13610 13030 13622 13082
rect 13674 13030 13686 13082
rect 13738 13030 19366 13082
rect 19418 13030 19430 13082
rect 19482 13030 19494 13082
rect 19546 13030 19558 13082
rect 19610 13030 19622 13082
rect 19674 13030 19686 13082
rect 19738 13030 23368 13082
rect 552 13008 23368 13030
rect 1670 12928 1676 12980
rect 1728 12928 1734 12980
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 1857 12971 1915 12977
rect 1857 12968 1869 12971
rect 1820 12940 1869 12968
rect 1820 12928 1826 12940
rect 1857 12937 1869 12940
rect 1903 12937 1915 12971
rect 1857 12931 1915 12937
rect 2038 12928 2044 12980
rect 2096 12928 2102 12980
rect 2222 12928 2228 12980
rect 2280 12968 2286 12980
rect 2317 12971 2375 12977
rect 2317 12968 2329 12971
rect 2280 12940 2329 12968
rect 2280 12928 2286 12940
rect 2317 12937 2329 12940
rect 2363 12937 2375 12971
rect 3329 12971 3387 12977
rect 3329 12968 3341 12971
rect 2317 12931 2375 12937
rect 2516 12940 3341 12968
rect 1305 12903 1363 12909
rect 1305 12869 1317 12903
rect 1351 12900 1363 12903
rect 2056 12900 2084 12928
rect 2406 12900 2412 12912
rect 1351 12872 2084 12900
rect 2148 12872 2412 12900
rect 1351 12869 1363 12872
rect 1305 12863 1363 12869
rect 1578 12832 1584 12844
rect 1228 12804 1584 12832
rect 1228 12773 1256 12804
rect 1578 12792 1584 12804
rect 1636 12832 1642 12844
rect 1636 12804 1992 12832
rect 1636 12792 1642 12804
rect 1964 12773 1992 12804
rect 2148 12773 2176 12872
rect 2406 12860 2412 12872
rect 2464 12860 2470 12912
rect 1213 12767 1271 12773
rect 1213 12733 1225 12767
rect 1259 12733 1271 12767
rect 1213 12727 1271 12733
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1949 12767 2007 12773
rect 1443 12736 1900 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1118 12656 1124 12708
rect 1176 12696 1182 12708
rect 1489 12699 1547 12705
rect 1489 12696 1501 12699
rect 1176 12668 1501 12696
rect 1176 12656 1182 12668
rect 1489 12665 1501 12668
rect 1535 12665 1547 12699
rect 1872 12696 1900 12736
rect 1949 12733 1961 12767
rect 1995 12733 2007 12767
rect 1949 12727 2007 12733
rect 2133 12767 2191 12773
rect 2133 12733 2145 12767
rect 2179 12733 2191 12767
rect 2409 12767 2467 12773
rect 2409 12764 2421 12767
rect 2133 12727 2191 12733
rect 2332 12736 2421 12764
rect 1872 12668 1992 12696
rect 1489 12659 1547 12665
rect 1964 12640 1992 12668
rect 1670 12588 1676 12640
rect 1728 12637 1734 12640
rect 1728 12631 1747 12637
rect 1735 12597 1747 12631
rect 1728 12591 1747 12597
rect 1728 12588 1734 12591
rect 1946 12588 1952 12640
rect 2004 12588 2010 12640
rect 2332 12628 2360 12736
rect 2409 12733 2421 12736
rect 2455 12733 2467 12767
rect 2516 12764 2544 12940
rect 3329 12937 3341 12940
rect 3375 12937 3387 12971
rect 3878 12968 3884 12980
rect 3329 12931 3387 12937
rect 3528 12940 3884 12968
rect 2958 12900 2964 12912
rect 2619 12872 2964 12900
rect 2619 12832 2647 12872
rect 2958 12860 2964 12872
rect 3016 12860 3022 12912
rect 3528 12841 3556 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 5534 12968 5540 12980
rect 5184 12940 5540 12968
rect 5184 12841 5212 12940
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 5902 12928 5908 12980
rect 5960 12928 5966 12980
rect 6454 12928 6460 12980
rect 6512 12928 6518 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 7064 12940 9229 12968
rect 7064 12928 7070 12940
rect 9217 12937 9229 12940
rect 9263 12937 9275 12971
rect 9217 12931 9275 12937
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10100 12940 10732 12968
rect 10100 12928 10106 12940
rect 6273 12903 6331 12909
rect 6273 12869 6285 12903
rect 6319 12900 6331 12903
rect 6472 12900 6500 12928
rect 6319 12872 6500 12900
rect 6319 12869 6331 12872
rect 6273 12863 6331 12869
rect 3513 12835 3571 12841
rect 2619 12804 2731 12832
rect 2703 12773 2731 12804
rect 3513 12801 3525 12835
rect 3559 12801 3571 12835
rect 3513 12795 3571 12801
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 5350 12792 5356 12844
rect 5408 12792 5414 12844
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2516 12736 2605 12764
rect 2409 12727 2467 12733
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12733 2743 12767
rect 2685 12727 2743 12733
rect 2823 12767 2881 12773
rect 2823 12733 2835 12767
rect 2869 12764 2881 12767
rect 2869 12733 2903 12764
rect 2823 12727 2903 12733
rect 2875 12696 2903 12727
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 3237 12767 3295 12773
rect 3237 12764 3249 12767
rect 3016 12736 3249 12764
rect 3016 12724 3022 12736
rect 3237 12733 3249 12736
rect 3283 12733 3295 12767
rect 3237 12727 3295 12733
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12764 3479 12767
rect 3467 12736 4016 12764
rect 3467 12733 3479 12736
rect 3421 12727 3479 12733
rect 3436 12696 3464 12727
rect 2875 12668 3464 12696
rect 3769 12699 3827 12705
rect 3769 12665 3781 12699
rect 3815 12665 3827 12699
rect 3769 12659 3827 12665
rect 3988 12696 4016 12736
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 4856 12736 5457 12764
rect 4856 12724 4862 12736
rect 5445 12733 5457 12736
rect 5491 12733 5503 12767
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5445 12727 5503 12733
rect 5552 12736 6101 12764
rect 5552 12696 5580 12736
rect 6089 12733 6101 12736
rect 6135 12733 6147 12767
rect 6089 12727 6147 12733
rect 6181 12767 6239 12773
rect 6181 12733 6193 12767
rect 6227 12764 6239 12767
rect 6270 12764 6276 12776
rect 6227 12736 6276 12764
rect 6227 12733 6239 12736
rect 6181 12727 6239 12733
rect 6270 12724 6276 12736
rect 6328 12724 6334 12776
rect 6365 12767 6423 12773
rect 6365 12733 6377 12767
rect 6411 12733 6423 12767
rect 6472 12764 6500 12872
rect 6730 12860 6736 12912
rect 6788 12860 6794 12912
rect 10134 12900 10140 12912
rect 7852 12872 10140 12900
rect 6748 12832 6776 12860
rect 6748 12804 6960 12832
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 6472 12736 6561 12764
rect 6365 12727 6423 12733
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 6733 12767 6791 12773
rect 6733 12733 6745 12767
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 6380 12696 6408 12727
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 3988 12668 5580 12696
rect 5828 12668 6316 12696
rect 6380 12668 6653 12696
rect 2958 12628 2964 12640
rect 2332 12600 2964 12628
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12628 3111 12631
rect 3784 12628 3812 12659
rect 3988 12640 4016 12668
rect 3099 12600 3812 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3970 12588 3976 12640
rect 4028 12588 4034 12640
rect 4890 12588 4896 12640
rect 4948 12588 4954 12640
rect 5828 12637 5856 12668
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12597 5871 12631
rect 6288 12628 6316 12668
rect 6641 12665 6653 12668
rect 6687 12665 6699 12699
rect 6641 12659 6699 12665
rect 6748 12628 6776 12727
rect 6822 12724 6828 12776
rect 6880 12724 6886 12776
rect 6932 12764 6960 12804
rect 7852 12764 7880 12872
rect 10134 12860 10140 12872
rect 10192 12860 10198 12912
rect 10704 12900 10732 12940
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 13044 12940 13645 12968
rect 13044 12928 13050 12940
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 13633 12931 13691 12937
rect 15930 12928 15936 12980
rect 15988 12928 15994 12980
rect 16577 12971 16635 12977
rect 16577 12937 16589 12971
rect 16623 12968 16635 12971
rect 17586 12968 17592 12980
rect 16623 12940 17592 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 17586 12928 17592 12940
rect 17644 12968 17650 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 17644 12940 18429 12968
rect 17644 12928 17650 12940
rect 18417 12937 18429 12940
rect 18463 12937 18475 12971
rect 18417 12931 18475 12937
rect 18524 12940 21220 12968
rect 10704 12872 11284 12900
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 9631 12804 10609 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 10686 12792 10692 12844
rect 10744 12792 10750 12844
rect 10870 12792 10876 12844
rect 10928 12792 10934 12844
rect 11256 12841 11284 12872
rect 12894 12860 12900 12912
rect 12952 12860 12958 12912
rect 13372 12872 14228 12900
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12832 11115 12835
rect 11241 12835 11299 12841
rect 11103 12804 11192 12832
rect 11103 12801 11115 12804
rect 11057 12795 11115 12801
rect 6932 12736 7880 12764
rect 9401 12767 9459 12773
rect 9401 12733 9413 12767
rect 9447 12733 9459 12767
rect 9401 12727 9459 12733
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 9858 12764 9864 12776
rect 9723 12736 9864 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 6288 12600 6776 12628
rect 6840 12628 6868 12724
rect 7092 12699 7150 12705
rect 7092 12665 7104 12699
rect 7138 12696 7150 12699
rect 7466 12696 7472 12708
rect 7138 12668 7472 12696
rect 7138 12665 7150 12668
rect 7092 12659 7150 12665
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 9416 12696 9444 12727
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 10704 12764 10732 12792
rect 10781 12767 10839 12773
rect 10781 12764 10793 12767
rect 10704 12736 10793 12764
rect 10781 12733 10793 12736
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12733 11023 12767
rect 11164 12764 11192 12804
rect 11241 12801 11253 12835
rect 11287 12801 11299 12835
rect 11241 12795 11299 12801
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 13372 12841 13400 12872
rect 13265 12835 13323 12841
rect 13265 12832 13277 12835
rect 11940 12804 13277 12832
rect 11940 12792 11946 12804
rect 13265 12801 13277 12804
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 14200 12841 14228 12872
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 15948 12832 15976 12928
rect 16390 12860 16396 12912
rect 16448 12900 16454 12912
rect 18524 12900 18552 12940
rect 19613 12903 19671 12909
rect 19613 12900 19625 12903
rect 16448 12872 18552 12900
rect 19536 12872 19625 12900
rect 16448 12860 16454 12872
rect 18046 12832 18052 12844
rect 14231 12804 14412 12832
rect 15948 12804 18052 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14384 12776 14412 12804
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 18782 12832 18788 12844
rect 18380 12804 18788 12832
rect 18380 12792 18386 12804
rect 18782 12792 18788 12804
rect 18840 12832 18846 12844
rect 19536 12841 19564 12872
rect 19613 12869 19625 12872
rect 19659 12869 19671 12903
rect 19613 12863 19671 12869
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 18840 12804 19533 12832
rect 18840 12792 18846 12804
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 11330 12764 11336 12776
rect 11164 12736 11336 12764
rect 10965 12727 11023 12733
rect 10980 12696 11008 12727
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 11425 12767 11483 12773
rect 11425 12733 11437 12767
rect 11471 12764 11483 12767
rect 11514 12764 11520 12776
rect 11471 12736 11520 12764
rect 11471 12733 11483 12736
rect 11425 12727 11483 12733
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 11606 12724 11612 12776
rect 11664 12724 11670 12776
rect 11698 12724 11704 12776
rect 11756 12724 11762 12776
rect 13078 12764 13084 12776
rect 12452 12736 13084 12764
rect 11238 12696 11244 12708
rect 9416 12668 9674 12696
rect 10980 12668 11244 12696
rect 7282 12628 7288 12640
rect 6840 12600 7288 12628
rect 5813 12591 5871 12597
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 9490 12628 9496 12640
rect 8260 12600 9496 12628
rect 8260 12588 8266 12600
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9646 12628 9674 12668
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 12452 12696 12480 12736
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 13906 12724 13912 12776
rect 13964 12724 13970 12776
rect 14274 12724 14280 12776
rect 14332 12724 14338 12776
rect 14366 12724 14372 12776
rect 14424 12724 14430 12776
rect 14458 12724 14464 12776
rect 14516 12724 14522 12776
rect 16393 12767 16451 12773
rect 16393 12733 16405 12767
rect 16439 12733 16451 12767
rect 16393 12727 16451 12733
rect 16669 12767 16727 12773
rect 16669 12733 16681 12767
rect 16715 12764 16727 12767
rect 17218 12764 17224 12776
rect 16715 12736 17224 12764
rect 16715 12733 16727 12736
rect 16669 12727 16727 12733
rect 16408 12696 16436 12727
rect 17218 12724 17224 12736
rect 17276 12724 17282 12776
rect 18233 12767 18291 12773
rect 18233 12733 18245 12767
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 19245 12767 19303 12773
rect 18555 12736 19196 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 16850 12696 16856 12708
rect 11348 12668 12480 12696
rect 12820 12668 14688 12696
rect 16408 12668 16856 12696
rect 10226 12628 10232 12640
rect 9646 12600 10232 12628
rect 10226 12588 10232 12600
rect 10284 12628 10290 12640
rect 11348 12628 11376 12668
rect 10284 12600 11376 12628
rect 10284 12588 10290 12600
rect 11974 12588 11980 12640
rect 12032 12628 12038 12640
rect 12820 12628 12848 12668
rect 14660 12640 14688 12668
rect 16850 12656 16856 12668
rect 16908 12696 16914 12708
rect 18248 12696 18276 12727
rect 16908 12668 18276 12696
rect 16908 12656 16914 12668
rect 12032 12600 12848 12628
rect 12032 12588 12038 12600
rect 14642 12588 14648 12640
rect 14700 12588 14706 12640
rect 16209 12631 16267 12637
rect 16209 12597 16221 12631
rect 16255 12628 16267 12631
rect 17310 12628 17316 12640
rect 16255 12600 17316 12628
rect 16255 12597 16267 12600
rect 16209 12591 16267 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12628 18107 12631
rect 18782 12628 18788 12640
rect 18095 12600 18788 12628
rect 18095 12597 18107 12600
rect 18049 12591 18107 12597
rect 18782 12588 18788 12600
rect 18840 12588 18846 12640
rect 19168 12628 19196 12736
rect 19245 12733 19257 12767
rect 19291 12733 19303 12767
rect 19245 12727 19303 12733
rect 19260 12696 19288 12727
rect 19794 12724 19800 12776
rect 19852 12764 19858 12776
rect 20165 12767 20223 12773
rect 19852 12736 20024 12764
rect 19852 12724 19858 12736
rect 19996 12708 20024 12736
rect 20165 12733 20177 12767
rect 20211 12764 20223 12767
rect 20254 12764 20260 12776
rect 20211 12736 20260 12764
rect 20211 12733 20223 12736
rect 20165 12727 20223 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20438 12773 20444 12776
rect 20432 12764 20444 12773
rect 20399 12736 20444 12764
rect 20432 12727 20444 12736
rect 20438 12724 20444 12727
rect 20496 12724 20502 12776
rect 21192 12764 21220 12940
rect 21358 12928 21364 12980
rect 21416 12968 21422 12980
rect 21637 12971 21695 12977
rect 21637 12968 21649 12971
rect 21416 12940 21649 12968
rect 21416 12928 21422 12940
rect 21637 12937 21649 12940
rect 21683 12937 21695 12971
rect 23400 12968 23428 13144
rect 21637 12931 21695 12937
rect 22940 12940 23428 12968
rect 21542 12792 21548 12844
rect 21600 12832 21606 12844
rect 22189 12835 22247 12841
rect 22189 12832 22201 12835
rect 21600 12804 22201 12832
rect 21600 12792 21606 12804
rect 22189 12801 22201 12804
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 21192 12736 22109 12764
rect 22097 12733 22109 12736
rect 22143 12764 22155 12767
rect 22940 12764 22968 12940
rect 23290 12832 23296 12844
rect 23032 12804 23296 12832
rect 23032 12773 23060 12804
rect 23290 12792 23296 12804
rect 23348 12792 23354 12844
rect 22143 12736 22968 12764
rect 23017 12767 23075 12773
rect 22143 12733 22155 12736
rect 22097 12727 22155 12733
rect 23017 12733 23029 12767
rect 23063 12733 23075 12767
rect 23017 12727 23075 12733
rect 19886 12696 19892 12708
rect 19260 12668 19892 12696
rect 19886 12656 19892 12668
rect 19944 12656 19950 12708
rect 19978 12656 19984 12708
rect 20036 12656 20042 12708
rect 22005 12699 22063 12705
rect 22005 12665 22017 12699
rect 22051 12696 22063 12699
rect 22186 12696 22192 12708
rect 22051 12668 22192 12696
rect 22051 12665 22063 12668
rect 22005 12659 22063 12665
rect 22186 12656 22192 12668
rect 22244 12656 22250 12708
rect 20162 12628 20168 12640
rect 19168 12600 20168 12628
rect 20162 12588 20168 12600
rect 20220 12588 20226 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 21545 12631 21603 12637
rect 21545 12628 21557 12631
rect 20772 12600 21557 12628
rect 20772 12588 20778 12600
rect 21545 12597 21557 12600
rect 21591 12597 21603 12631
rect 21545 12591 21603 12597
rect 22830 12588 22836 12640
rect 22888 12588 22894 12640
rect 552 12538 23368 12560
rect 552 12486 4366 12538
rect 4418 12486 4430 12538
rect 4482 12486 4494 12538
rect 4546 12486 4558 12538
rect 4610 12486 4622 12538
rect 4674 12486 4686 12538
rect 4738 12486 10366 12538
rect 10418 12486 10430 12538
rect 10482 12486 10494 12538
rect 10546 12486 10558 12538
rect 10610 12486 10622 12538
rect 10674 12486 10686 12538
rect 10738 12486 16366 12538
rect 16418 12486 16430 12538
rect 16482 12486 16494 12538
rect 16546 12486 16558 12538
rect 16610 12486 16622 12538
rect 16674 12486 16686 12538
rect 16738 12486 22366 12538
rect 22418 12486 22430 12538
rect 22482 12486 22494 12538
rect 22546 12486 22558 12538
rect 22610 12486 22622 12538
rect 22674 12486 22686 12538
rect 22738 12486 23368 12538
rect 552 12464 23368 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 1728 12396 2053 12424
rect 1728 12384 1734 12396
rect 2041 12393 2053 12396
rect 2087 12393 2099 12427
rect 2041 12387 2099 12393
rect 2332 12396 3372 12424
rect 1578 12316 1584 12368
rect 1636 12316 1642 12368
rect 1854 12316 1860 12368
rect 1912 12316 1918 12368
rect 1596 12288 1624 12316
rect 1673 12291 1731 12297
rect 1673 12288 1685 12291
rect 1596 12260 1685 12288
rect 1673 12257 1685 12260
rect 1719 12257 1731 12291
rect 1673 12251 1731 12257
rect 1688 12220 1716 12251
rect 1946 12248 1952 12300
rect 2004 12288 2010 12300
rect 2332 12297 2360 12396
rect 2406 12316 2412 12368
rect 2464 12356 2470 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2464 12328 2789 12356
rect 2464 12316 2470 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 2777 12319 2835 12325
rect 3344 12356 3372 12396
rect 4798 12384 4804 12436
rect 4856 12424 4862 12436
rect 5350 12424 5356 12436
rect 4856 12396 5356 12424
rect 4856 12384 4862 12396
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 7466 12384 7472 12436
rect 7524 12384 7530 12436
rect 7576 12396 11100 12424
rect 7576 12356 7604 12396
rect 10870 12356 10876 12368
rect 3344 12328 7604 12356
rect 10520 12328 10876 12356
rect 2317 12291 2375 12297
rect 2317 12288 2329 12291
rect 2004 12260 2329 12288
rect 2004 12248 2010 12260
rect 2317 12257 2329 12260
rect 2363 12257 2375 12291
rect 2317 12251 2375 12257
rect 2498 12248 2504 12300
rect 2556 12248 2562 12300
rect 3344 12297 3372 12328
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12257 3387 12291
rect 3329 12251 3387 12257
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 4304 12260 4445 12288
rect 4304 12248 4310 12260
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 2038 12220 2044 12232
rect 1688 12192 2044 12220
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 1118 12112 1124 12164
rect 1176 12112 1182 12164
rect 1762 12112 1768 12164
rect 1820 12112 1826 12164
rect 2240 12152 2268 12183
rect 2314 12152 2320 12164
rect 2240 12124 2320 12152
rect 2314 12112 2320 12124
rect 2372 12112 2378 12164
rect 2424 12152 2452 12183
rect 2590 12180 2596 12232
rect 2648 12220 2654 12232
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2648 12192 3065 12220
rect 2648 12180 2654 12192
rect 3053 12189 3065 12192
rect 3099 12220 3111 12223
rect 4448 12220 4476 12251
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 4801 12291 4859 12297
rect 4801 12288 4813 12291
rect 4672 12260 4813 12288
rect 4672 12248 4678 12260
rect 4801 12257 4813 12260
rect 4847 12257 4859 12291
rect 4801 12251 4859 12257
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5169 12291 5227 12297
rect 5169 12288 5181 12291
rect 4948 12260 5181 12288
rect 4948 12248 4954 12260
rect 5169 12257 5181 12260
rect 5215 12257 5227 12291
rect 5169 12251 5227 12257
rect 5350 12248 5356 12300
rect 5408 12248 5414 12300
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 5902 12288 5908 12300
rect 5491 12260 5908 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 7834 12288 7840 12300
rect 7699 12260 7840 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 8012 12291 8070 12297
rect 8012 12257 8024 12291
rect 8058 12288 8070 12291
rect 8478 12288 8484 12300
rect 8058 12260 8484 12288
rect 8058 12257 8070 12260
rect 8012 12251 8070 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 10226 12288 10232 12300
rect 9723 12260 10232 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 4706 12220 4712 12232
rect 3099 12192 3812 12220
rect 4448 12192 4712 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3784 12152 3812 12192
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 5368 12220 5396 12248
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5368 12192 5825 12220
rect 5813 12189 5825 12192
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 2424 12124 3556 12152
rect 3784 12124 4936 12152
rect 1136 12084 1164 12112
rect 3528 12096 3556 12124
rect 2406 12084 2412 12096
rect 1136 12056 2412 12084
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 2869 12087 2927 12093
rect 2869 12053 2881 12087
rect 2915 12084 2927 12087
rect 2958 12084 2964 12096
rect 2915 12056 2964 12084
rect 2915 12053 2927 12056
rect 2869 12047 2927 12053
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3510 12044 3516 12096
rect 3568 12044 3574 12096
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4614 12084 4620 12096
rect 4212 12056 4620 12084
rect 4212 12044 4218 12056
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 4908 12084 4936 12124
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 5261 12155 5319 12161
rect 5261 12152 5273 12155
rect 5132 12124 5273 12152
rect 5132 12112 5138 12124
rect 5261 12121 5273 12124
rect 5307 12121 5319 12155
rect 5261 12115 5319 12121
rect 5353 12155 5411 12161
rect 5353 12121 5365 12155
rect 5399 12152 5411 12155
rect 5994 12152 6000 12164
rect 5399 12124 6000 12152
rect 5399 12121 5411 12124
rect 5353 12115 5411 12121
rect 5994 12112 6000 12124
rect 6052 12152 6058 12164
rect 6104 12152 6132 12183
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7340 12192 7757 12220
rect 7340 12180 7346 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 9493 12223 9551 12229
rect 9493 12220 9505 12223
rect 8812 12192 9505 12220
rect 8812 12180 8818 12192
rect 9493 12189 9505 12192
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9953 12223 10011 12229
rect 9953 12220 9965 12223
rect 9824 12192 9965 12220
rect 9824 12180 9830 12192
rect 9953 12189 9965 12192
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10520 12220 10548 12328
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 11072 12356 11100 12396
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 12161 12427 12219 12433
rect 12161 12424 12173 12427
rect 11664 12396 12173 12424
rect 11664 12384 11670 12396
rect 12161 12393 12173 12396
rect 12207 12393 12219 12427
rect 12161 12387 12219 12393
rect 13814 12384 13820 12436
rect 13872 12384 13878 12436
rect 14001 12427 14059 12433
rect 14001 12393 14013 12427
rect 14047 12424 14059 12427
rect 14274 12424 14280 12436
rect 14047 12396 14280 12424
rect 14047 12393 14059 12396
rect 14001 12387 14059 12393
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 15746 12384 15752 12436
rect 15804 12384 15810 12436
rect 17402 12384 17408 12436
rect 17460 12384 17466 12436
rect 13832 12356 13860 12384
rect 11072 12328 12480 12356
rect 10597 12291 10655 12297
rect 10597 12257 10609 12291
rect 10643 12288 10655 12291
rect 10781 12291 10839 12297
rect 10643 12260 10732 12288
rect 10643 12257 10655 12260
rect 10597 12251 10655 12257
rect 10704 12232 10732 12260
rect 10781 12257 10793 12291
rect 10827 12257 10839 12291
rect 10888 12288 10916 12316
rect 12452 12297 12480 12328
rect 13372 12328 13860 12356
rect 10957 12291 11015 12297
rect 10957 12288 10969 12291
rect 10888 12260 10969 12288
rect 10781 12251 10839 12257
rect 10957 12257 10969 12260
rect 11003 12257 11015 12291
rect 10957 12251 11015 12257
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 12345 12291 12403 12297
rect 12345 12288 12357 12291
rect 11471 12260 12357 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 10192 12192 10548 12220
rect 10192 12180 10198 12192
rect 10686 12180 10692 12232
rect 10744 12180 10750 12232
rect 10796 12220 10824 12251
rect 11514 12220 11520 12232
rect 10796 12192 11520 12220
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 6052 12124 6132 12152
rect 6052 12112 6058 12124
rect 4985 12087 5043 12093
rect 4985 12084 4997 12087
rect 4908 12056 4997 12084
rect 4985 12053 4997 12056
rect 5031 12084 5043 12087
rect 5442 12084 5448 12096
rect 5031 12056 5448 12084
rect 5031 12053 5043 12056
rect 4985 12047 5043 12053
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5626 12044 5632 12096
rect 5684 12044 5690 12096
rect 6104 12084 6132 12124
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 9861 12155 9919 12161
rect 9364 12124 9536 12152
rect 9364 12112 9370 12124
rect 6638 12084 6644 12096
rect 6104 12056 6644 12084
rect 6638 12044 6644 12056
rect 6696 12084 6702 12096
rect 7926 12084 7932 12096
rect 6696 12056 7932 12084
rect 6696 12044 6702 12056
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 9125 12087 9183 12093
rect 9125 12053 9137 12087
rect 9171 12084 9183 12087
rect 9398 12084 9404 12096
rect 9171 12056 9404 12084
rect 9171 12053 9183 12056
rect 9125 12047 9183 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9508 12084 9536 12124
rect 9861 12121 9873 12155
rect 9907 12152 9919 12155
rect 10870 12152 10876 12164
rect 9907 12124 10876 12152
rect 9907 12121 9919 12124
rect 9861 12115 9919 12121
rect 10870 12112 10876 12124
rect 10928 12112 10934 12164
rect 11149 12155 11207 12161
rect 11149 12121 11161 12155
rect 11195 12152 11207 12155
rect 11422 12152 11428 12164
rect 11195 12124 11428 12152
rect 11195 12121 11207 12124
rect 11149 12115 11207 12121
rect 11422 12112 11428 12124
rect 11480 12152 11486 12164
rect 11624 12152 11652 12260
rect 12345 12257 12357 12260
rect 12391 12257 12403 12291
rect 12345 12251 12403 12257
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 12529 12291 12587 12297
rect 12529 12257 12541 12291
rect 12575 12288 12587 12291
rect 12575 12260 12848 12288
rect 12575 12257 12587 12260
rect 12529 12251 12587 12257
rect 12820 12232 12848 12260
rect 12986 12248 12992 12300
rect 13044 12248 13050 12300
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 13372 12229 13400 12328
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12257 13691 12291
rect 13633 12251 13691 12257
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 11480 12124 11652 12152
rect 11480 12112 11486 12124
rect 12158 12112 12164 12164
rect 12216 12152 12222 12164
rect 12912 12152 12940 12183
rect 12216 12124 12940 12152
rect 12216 12112 12222 12124
rect 13078 12112 13084 12164
rect 13136 12152 13142 12164
rect 13464 12152 13492 12251
rect 13136 12124 13492 12152
rect 13136 12112 13142 12124
rect 10594 12084 10600 12096
rect 9508 12056 10600 12084
rect 10594 12044 10600 12056
rect 10652 12044 10658 12096
rect 10689 12087 10747 12093
rect 10689 12053 10701 12087
rect 10735 12084 10747 12087
rect 10778 12084 10784 12096
rect 10735 12056 10784 12084
rect 10735 12053 10747 12056
rect 10689 12047 10747 12053
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 11296 12056 11345 12084
rect 11296 12044 11302 12056
rect 11333 12053 11345 12056
rect 11379 12084 11391 12087
rect 12250 12084 12256 12096
rect 11379 12056 12256 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 13648 12084 13676 12251
rect 13722 12248 13728 12300
rect 13780 12248 13786 12300
rect 13832 12297 13860 12328
rect 14090 12316 14096 12368
rect 14148 12356 14154 12368
rect 14734 12356 14740 12368
rect 14148 12328 14740 12356
rect 14148 12316 14154 12328
rect 14734 12316 14740 12328
rect 14792 12356 14798 12368
rect 15764 12356 15792 12384
rect 14792 12328 15792 12356
rect 14792 12316 14798 12328
rect 15930 12316 15936 12368
rect 15988 12356 15994 12368
rect 17230 12359 17288 12365
rect 17230 12356 17242 12359
rect 15988 12328 17242 12356
rect 15988 12316 15994 12328
rect 17230 12325 17242 12328
rect 17276 12325 17288 12359
rect 17230 12319 17288 12325
rect 17420 12356 17448 12384
rect 19058 12356 19064 12368
rect 17420 12328 19064 12356
rect 13832 12291 13899 12297
rect 13832 12260 13853 12291
rect 13841 12257 13853 12260
rect 13887 12257 13899 12291
rect 13841 12251 13899 12257
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16206 12288 16212 12300
rect 15795 12260 16212 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 17420 12288 17448 12328
rect 19058 12316 19064 12328
rect 19116 12356 19122 12368
rect 20254 12356 20260 12368
rect 19116 12328 20260 12356
rect 19116 12316 19122 12328
rect 17497 12291 17555 12297
rect 17497 12288 17509 12291
rect 17420 12260 17509 12288
rect 17497 12257 17509 12260
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 18322 12248 18328 12300
rect 18380 12248 18386 12300
rect 18414 12248 18420 12300
rect 18472 12248 18478 12300
rect 18601 12291 18659 12297
rect 18601 12257 18613 12291
rect 18647 12257 18659 12291
rect 18601 12251 18659 12257
rect 18340 12220 18368 12248
rect 18616 12220 18644 12251
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 20088 12297 20116 12328
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 19806 12291 19864 12297
rect 19806 12288 19818 12291
rect 18748 12260 19818 12288
rect 18748 12248 18754 12260
rect 19806 12257 19818 12260
rect 19852 12257 19864 12291
rect 19806 12251 19864 12257
rect 20073 12291 20131 12297
rect 20073 12257 20085 12291
rect 20119 12257 20131 12291
rect 20073 12251 20131 12257
rect 18782 12220 18788 12232
rect 18340 12192 18788 12220
rect 18782 12180 18788 12192
rect 18840 12180 18846 12232
rect 17586 12112 17592 12164
rect 17644 12152 17650 12164
rect 17644 12124 18828 12152
rect 17644 12112 17650 12124
rect 13320 12056 13676 12084
rect 13320 12044 13326 12056
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 15102 12084 15108 12096
rect 13872 12056 15108 12084
rect 13872 12044 13878 12056
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 15930 12044 15936 12096
rect 15988 12044 15994 12096
rect 16114 12044 16120 12096
rect 16172 12044 16178 12096
rect 18506 12044 18512 12096
rect 18564 12044 18570 12096
rect 18598 12044 18604 12096
rect 18656 12084 18662 12096
rect 18693 12087 18751 12093
rect 18693 12084 18705 12087
rect 18656 12056 18705 12084
rect 18656 12044 18662 12056
rect 18693 12053 18705 12056
rect 18739 12053 18751 12087
rect 18800 12084 18828 12124
rect 22278 12084 22284 12096
rect 18800 12056 22284 12084
rect 18693 12047 18751 12053
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 552 11994 23368 12016
rect 552 11942 1366 11994
rect 1418 11942 1430 11994
rect 1482 11942 1494 11994
rect 1546 11942 1558 11994
rect 1610 11942 1622 11994
rect 1674 11942 1686 11994
rect 1738 11942 7366 11994
rect 7418 11942 7430 11994
rect 7482 11942 7494 11994
rect 7546 11942 7558 11994
rect 7610 11942 7622 11994
rect 7674 11942 7686 11994
rect 7738 11942 13366 11994
rect 13418 11942 13430 11994
rect 13482 11942 13494 11994
rect 13546 11942 13558 11994
rect 13610 11942 13622 11994
rect 13674 11942 13686 11994
rect 13738 11942 19366 11994
rect 19418 11942 19430 11994
rect 19482 11942 19494 11994
rect 19546 11942 19558 11994
rect 19610 11942 19622 11994
rect 19674 11942 19686 11994
rect 19738 11942 23368 11994
rect 552 11920 23368 11942
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 2096 11852 2145 11880
rect 2096 11840 2102 11852
rect 2133 11849 2145 11852
rect 2179 11849 2191 11883
rect 2133 11843 2191 11849
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 2556 11852 4629 11880
rect 2556 11840 2562 11852
rect 4617 11849 4629 11852
rect 4663 11880 4675 11883
rect 5074 11880 5080 11892
rect 4663 11852 5080 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 2056 11744 2084 11840
rect 4246 11772 4252 11824
rect 4304 11812 4310 11824
rect 4525 11815 4583 11821
rect 4525 11812 4537 11815
rect 4304 11784 4537 11812
rect 4304 11772 4310 11784
rect 4525 11781 4537 11784
rect 4571 11781 4583 11815
rect 4525 11775 4583 11781
rect 1596 11716 2084 11744
rect 4632 11744 4660 11843
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 5224 11852 5273 11880
rect 5224 11840 5230 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 11241 11883 11299 11889
rect 11241 11880 11253 11883
rect 10928 11852 11253 11880
rect 10928 11840 10934 11852
rect 11241 11849 11253 11852
rect 11287 11849 11299 11883
rect 11241 11843 11299 11849
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13320 11852 13553 11880
rect 13320 11840 13326 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 14090 11880 14096 11892
rect 13541 11843 13599 11849
rect 13832 11852 14096 11880
rect 4706 11772 4712 11824
rect 4764 11812 4770 11824
rect 10686 11812 10692 11824
rect 4764 11784 10692 11812
rect 4764 11772 4770 11784
rect 10686 11772 10692 11784
rect 10744 11812 10750 11824
rect 10744 11784 11376 11812
rect 10744 11772 10750 11784
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 4632 11716 5549 11744
rect 1596 11685 1624 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5718 11704 5724 11756
rect 5776 11704 5782 11756
rect 6454 11744 6460 11756
rect 6104 11716 6460 11744
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11645 1639 11679
rect 1581 11639 1639 11645
rect 1762 11636 1768 11688
rect 1820 11636 1826 11688
rect 2314 11676 2320 11688
rect 1872 11648 2320 11676
rect 1872 11552 1900 11648
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11676 2559 11679
rect 3234 11676 3240 11688
rect 2547 11648 3240 11676
rect 2547 11645 2559 11648
rect 2501 11639 2559 11645
rect 3234 11636 3240 11648
rect 3292 11636 3298 11688
rect 3510 11636 3516 11688
rect 3568 11636 3574 11688
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 4304 11648 4353 11676
rect 4304 11636 4310 11648
rect 4341 11645 4353 11648
rect 4387 11645 4399 11679
rect 4341 11639 4399 11645
rect 4706 11636 4712 11688
rect 4764 11636 4770 11688
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 4801 11639 4859 11645
rect 5077 11679 5135 11685
rect 5077 11645 5089 11679
rect 5123 11676 5135 11679
rect 5123 11648 5212 11676
rect 5123 11645 5135 11648
rect 5077 11639 5135 11645
rect 3528 11608 3556 11636
rect 4724 11608 4752 11636
rect 3528 11580 4752 11608
rect 4816 11608 4844 11639
rect 4816 11580 5120 11608
rect 5092 11552 5120 11580
rect 5184 11552 5212 11648
rect 5442 11636 5448 11688
rect 5500 11636 5506 11688
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 5902 11676 5908 11688
rect 5675 11648 5908 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 5902 11636 5908 11648
rect 5960 11676 5966 11688
rect 6104 11676 6132 11716
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 10870 11704 10876 11756
rect 10928 11704 10934 11756
rect 10962 11704 10968 11756
rect 11020 11704 11026 11756
rect 5960 11648 6132 11676
rect 6181 11679 6239 11685
rect 5960 11636 5966 11648
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 6227 11648 6868 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 6840 11620 6868 11648
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 10505 11679 10563 11685
rect 7984 11648 10456 11676
rect 7984 11636 7990 11648
rect 6454 11568 6460 11620
rect 6512 11608 6518 11620
rect 6641 11611 6699 11617
rect 6641 11608 6653 11611
rect 6512 11580 6653 11608
rect 6512 11568 6518 11580
rect 6641 11577 6653 11580
rect 6687 11577 6699 11611
rect 6641 11571 6699 11577
rect 6822 11568 6828 11620
rect 6880 11568 6886 11620
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 7248 11580 10149 11608
rect 7248 11568 7254 11580
rect 10137 11577 10149 11580
rect 10183 11577 10195 11611
rect 10137 11571 10195 11577
rect 10226 11568 10232 11620
rect 10284 11608 10290 11620
rect 10321 11611 10379 11617
rect 10321 11608 10333 11611
rect 10284 11580 10333 11608
rect 10284 11568 10290 11580
rect 10321 11577 10333 11580
rect 10367 11577 10379 11611
rect 10428 11608 10456 11648
rect 10505 11645 10517 11679
rect 10551 11676 10563 11679
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10551 11648 10793 11676
rect 10551 11645 10563 11648
rect 10505 11639 10563 11645
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 11054 11636 11060 11688
rect 11112 11636 11118 11688
rect 11348 11676 11376 11784
rect 11514 11772 11520 11824
rect 11572 11812 11578 11824
rect 11572 11784 11652 11812
rect 11572 11772 11578 11784
rect 11422 11704 11428 11756
rect 11480 11704 11486 11756
rect 11624 11753 11652 11784
rect 12158 11772 12164 11824
rect 12216 11772 12222 11824
rect 11609 11747 11667 11753
rect 11609 11713 11621 11747
rect 11655 11713 11667 11747
rect 11609 11707 11667 11713
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11348 11648 11529 11676
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 11698 11636 11704 11688
rect 11756 11636 11762 11688
rect 12176 11676 12204 11772
rect 11808 11648 12204 11676
rect 11808 11608 11836 11648
rect 13722 11636 13728 11688
rect 13780 11636 13786 11688
rect 13832 11685 13860 11852
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11849 14519 11883
rect 14461 11843 14519 11849
rect 14277 11815 14335 11821
rect 14277 11781 14289 11815
rect 14323 11781 14335 11815
rect 14277 11775 14335 11781
rect 13817 11679 13875 11685
rect 13817 11645 13829 11679
rect 13863 11645 13875 11679
rect 13817 11639 13875 11645
rect 14090 11636 14096 11688
rect 14148 11636 14154 11688
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14292 11676 14320 11775
rect 14231 11648 14320 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 10428 11580 11836 11608
rect 10321 11571 10379 11577
rect 12894 11568 12900 11620
rect 12952 11608 12958 11620
rect 13630 11608 13636 11620
rect 12952 11580 13636 11608
rect 12952 11568 12958 11580
rect 13630 11568 13636 11580
rect 13688 11608 13694 11620
rect 13909 11611 13967 11617
rect 13909 11608 13921 11611
rect 13688 11580 13921 11608
rect 13688 11568 13694 11580
rect 13909 11577 13921 11580
rect 13955 11577 13967 11611
rect 13909 11571 13967 11577
rect 14274 11568 14280 11620
rect 14332 11608 14338 11620
rect 14476 11608 14504 11843
rect 16206 11840 16212 11892
rect 16264 11840 16270 11892
rect 17402 11840 17408 11892
rect 17460 11840 17466 11892
rect 18322 11840 18328 11892
rect 18380 11840 18386 11892
rect 18506 11840 18512 11892
rect 18564 11840 18570 11892
rect 18690 11840 18696 11892
rect 18748 11840 18754 11892
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 14936 11716 15301 11744
rect 14936 11688 14964 11716
rect 15289 11713 15301 11716
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 16114 11704 16120 11756
rect 16172 11704 16178 11756
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11744 16911 11747
rect 17126 11744 17132 11756
rect 16899 11716 17132 11744
rect 16899 11713 16911 11716
rect 16853 11707 16911 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 18524 11744 18552 11840
rect 18524 11716 19104 11744
rect 14918 11636 14924 11688
rect 14976 11636 14982 11688
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11645 15163 11679
rect 15105 11639 15163 11645
rect 14332 11580 14504 11608
rect 14332 11568 14338 11580
rect 14642 11568 14648 11620
rect 14700 11568 14706 11620
rect 15120 11608 15148 11639
rect 15378 11636 15384 11688
rect 15436 11636 15442 11688
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11676 15991 11679
rect 16132 11676 16160 11704
rect 15979 11648 16160 11676
rect 16577 11679 16635 11685
rect 15979 11645 15991 11648
rect 15933 11639 15991 11645
rect 16577 11645 16589 11679
rect 16623 11676 16635 11679
rect 17218 11676 17224 11688
rect 16623 11648 17224 11676
rect 16623 11645 16635 11648
rect 16577 11639 16635 11645
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18141 11679 18199 11685
rect 18141 11676 18153 11679
rect 18012 11648 18153 11676
rect 18012 11636 18018 11648
rect 18141 11645 18153 11648
rect 18187 11645 18199 11679
rect 18141 11639 18199 11645
rect 18598 11636 18604 11688
rect 18656 11636 18662 11688
rect 19076 11685 19104 11716
rect 20254 11704 20260 11756
rect 20312 11744 20318 11756
rect 20622 11744 20628 11756
rect 20312 11716 20628 11744
rect 20312 11704 20318 11716
rect 20622 11704 20628 11716
rect 20680 11744 20686 11756
rect 21177 11747 21235 11753
rect 21177 11744 21189 11747
rect 20680 11716 21189 11744
rect 20680 11704 20686 11716
rect 21177 11713 21189 11716
rect 21223 11713 21235 11747
rect 21177 11707 21235 11713
rect 18969 11679 19027 11685
rect 18969 11645 18981 11679
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19061 11679 19119 11685
rect 19061 11645 19073 11679
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 17313 11611 17371 11617
rect 14936 11580 16160 11608
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 1673 11543 1731 11549
rect 1673 11540 1685 11543
rect 1544 11512 1685 11540
rect 1544 11500 1550 11512
rect 1673 11509 1685 11512
rect 1719 11509 1731 11543
rect 1673 11503 1731 11509
rect 1854 11500 1860 11552
rect 1912 11500 1918 11552
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 4893 11543 4951 11549
rect 4893 11540 4905 11543
rect 4028 11512 4905 11540
rect 4028 11500 4034 11512
rect 4893 11509 4905 11512
rect 4939 11509 4951 11543
rect 4893 11503 4951 11509
rect 5074 11500 5080 11552
rect 5132 11500 5138 11552
rect 5166 11500 5172 11552
rect 5224 11500 5230 11552
rect 6089 11543 6147 11549
rect 6089 11509 6101 11543
rect 6135 11540 6147 11543
rect 6362 11540 6368 11552
rect 6135 11512 6368 11540
rect 6135 11509 6147 11512
rect 6089 11503 6147 11509
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 6730 11500 6736 11552
rect 6788 11500 6794 11552
rect 10597 11543 10655 11549
rect 10597 11509 10609 11543
rect 10643 11540 10655 11543
rect 11882 11540 11888 11552
rect 10643 11512 11888 11540
rect 10643 11509 10655 11512
rect 10597 11503 10655 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 13998 11540 14004 11552
rect 12124 11512 14004 11540
rect 12124 11500 12130 11512
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 14445 11543 14503 11549
rect 14445 11509 14457 11543
rect 14491 11540 14503 11543
rect 14550 11540 14556 11552
rect 14491 11512 14556 11540
rect 14491 11509 14503 11512
rect 14445 11503 14503 11509
rect 14550 11500 14556 11512
rect 14608 11540 14614 11552
rect 14936 11540 14964 11580
rect 14608 11512 14964 11540
rect 14608 11500 14614 11512
rect 15010 11500 15016 11552
rect 15068 11500 15074 11552
rect 16132 11549 16160 11580
rect 17313 11577 17325 11611
rect 17359 11608 17371 11611
rect 18616 11608 18644 11636
rect 17359 11580 18644 11608
rect 18984 11608 19012 11639
rect 19150 11636 19156 11688
rect 19208 11636 19214 11688
rect 19337 11679 19395 11685
rect 19337 11645 19349 11679
rect 19383 11676 19395 11679
rect 19886 11676 19892 11688
rect 19383 11648 19892 11676
rect 19383 11645 19395 11648
rect 19337 11639 19395 11645
rect 19886 11636 19892 11648
rect 19944 11676 19950 11688
rect 20346 11676 20352 11688
rect 19944 11648 20352 11676
rect 19944 11636 19950 11648
rect 20346 11636 20352 11648
rect 20404 11636 20410 11688
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11676 20867 11679
rect 21082 11676 21088 11688
rect 20855 11648 21088 11676
rect 20855 11645 20867 11648
rect 20809 11639 20867 11645
rect 21082 11636 21088 11648
rect 21140 11636 21146 11688
rect 20438 11608 20444 11620
rect 18984 11580 20444 11608
rect 17359 11577 17371 11580
rect 17313 11571 17371 11577
rect 20438 11568 20444 11580
rect 20496 11568 20502 11620
rect 20898 11568 20904 11620
rect 20956 11608 20962 11620
rect 21422 11611 21480 11617
rect 21422 11608 21434 11611
rect 20956 11580 21434 11608
rect 20956 11568 20962 11580
rect 21422 11577 21434 11580
rect 21468 11577 21480 11611
rect 21422 11571 21480 11577
rect 16117 11543 16175 11549
rect 16117 11509 16129 11543
rect 16163 11540 16175 11543
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 16163 11512 16681 11540
rect 16163 11509 16175 11512
rect 16117 11503 16175 11509
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 16669 11503 16727 11509
rect 20990 11500 20996 11552
rect 21048 11500 21054 11552
rect 22094 11500 22100 11552
rect 22152 11540 22158 11552
rect 22557 11543 22615 11549
rect 22557 11540 22569 11543
rect 22152 11512 22569 11540
rect 22152 11500 22158 11512
rect 22557 11509 22569 11512
rect 22603 11509 22615 11543
rect 22557 11503 22615 11509
rect 552 11450 23368 11472
rect 552 11398 4366 11450
rect 4418 11398 4430 11450
rect 4482 11398 4494 11450
rect 4546 11398 4558 11450
rect 4610 11398 4622 11450
rect 4674 11398 4686 11450
rect 4738 11398 10366 11450
rect 10418 11398 10430 11450
rect 10482 11398 10494 11450
rect 10546 11398 10558 11450
rect 10610 11398 10622 11450
rect 10674 11398 10686 11450
rect 10738 11398 16366 11450
rect 16418 11398 16430 11450
rect 16482 11398 16494 11450
rect 16546 11398 16558 11450
rect 16610 11398 16622 11450
rect 16674 11398 16686 11450
rect 16738 11398 22366 11450
rect 22418 11398 22430 11450
rect 22482 11398 22494 11450
rect 22546 11398 22558 11450
rect 22610 11398 22622 11450
rect 22674 11398 22686 11450
rect 22738 11398 23368 11450
rect 552 11376 23368 11398
rect 4890 11296 4896 11348
rect 4948 11296 4954 11348
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 5132 11308 5549 11336
rect 5132 11296 5138 11308
rect 5537 11305 5549 11308
rect 5583 11336 5595 11339
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5583 11308 6009 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 5997 11305 6009 11308
rect 6043 11336 6055 11339
rect 6178 11336 6184 11348
rect 6043 11308 6184 11336
rect 6043 11305 6055 11308
rect 5997 11299 6055 11305
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 7101 11339 7159 11345
rect 7101 11305 7113 11339
rect 7147 11336 7159 11339
rect 7190 11336 7196 11348
rect 7147 11308 7196 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 7834 11296 7840 11348
rect 7892 11336 7898 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 7892 11308 7941 11336
rect 7892 11296 7898 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 8750 11339 8808 11345
rect 8750 11336 8762 11339
rect 8536 11308 8762 11336
rect 8536 11296 8542 11308
rect 8750 11305 8762 11308
rect 8796 11305 8808 11339
rect 8750 11299 8808 11305
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 10284 11308 10609 11336
rect 10284 11296 10290 11308
rect 10597 11305 10609 11308
rect 10643 11305 10655 11339
rect 10597 11299 10655 11305
rect 1026 11160 1032 11212
rect 1084 11160 1090 11212
rect 1486 11209 1492 11212
rect 1480 11200 1492 11209
rect 1447 11172 1492 11200
rect 1480 11163 1492 11172
rect 1486 11160 1492 11163
rect 1544 11160 1550 11212
rect 3326 11160 3332 11212
rect 3384 11200 3390 11212
rect 3421 11203 3479 11209
rect 3421 11200 3433 11203
rect 3384 11172 3433 11200
rect 3384 11160 3390 11172
rect 3421 11169 3433 11172
rect 3467 11169 3479 11203
rect 3421 11163 3479 11169
rect 3973 11203 4031 11209
rect 3973 11169 3985 11203
rect 4019 11200 4031 11203
rect 4154 11200 4160 11212
rect 4019 11172 4160 11200
rect 4019 11169 4031 11172
rect 3973 11163 4031 11169
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 4706 11200 4712 11212
rect 4387 11172 4712 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11169 4859 11203
rect 4908 11200 4936 11296
rect 6273 11271 6331 11277
rect 6273 11268 6285 11271
rect 5184 11240 6285 11268
rect 5184 11200 5212 11240
rect 6273 11237 6285 11240
rect 6319 11237 6331 11271
rect 6273 11231 6331 11237
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 6733 11271 6791 11277
rect 6733 11268 6745 11271
rect 6696 11240 6745 11268
rect 6696 11228 6702 11240
rect 6733 11237 6745 11240
rect 6779 11237 6791 11271
rect 6733 11231 6791 11237
rect 8113 11271 8171 11277
rect 8113 11237 8125 11271
rect 8159 11268 8171 11271
rect 8386 11268 8392 11280
rect 8159 11240 8392 11268
rect 8159 11237 8171 11240
rect 8113 11231 8171 11237
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 8665 11271 8723 11277
rect 8665 11237 8677 11271
rect 8711 11268 8723 11271
rect 8711 11240 9260 11268
rect 8711 11237 8723 11240
rect 8665 11231 8723 11237
rect 9232 11212 9260 11240
rect 9950 11228 9956 11280
rect 10008 11268 10014 11280
rect 10612 11268 10640 11299
rect 11054 11296 11060 11348
rect 11112 11296 11118 11348
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 12526 11336 12532 11348
rect 11296 11308 12532 11336
rect 11296 11296 11302 11308
rect 12526 11296 12532 11308
rect 12584 11336 12590 11348
rect 12584 11308 14044 11336
rect 12584 11296 12590 11308
rect 13814 11268 13820 11280
rect 10008 11240 10456 11268
rect 10612 11240 13820 11268
rect 10008 11228 10014 11240
rect 5261 11203 5319 11209
rect 5261 11200 5273 11203
rect 4908 11172 5273 11200
rect 4801 11163 4859 11169
rect 5261 11169 5273 11172
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 1044 11132 1072 11160
rect 1213 11135 1271 11141
rect 1213 11132 1225 11135
rect 1044 11104 1225 11132
rect 1213 11101 1225 11104
rect 1259 11101 1271 11135
rect 4246 11132 4252 11144
rect 1213 11095 1271 11101
rect 2608 11104 4252 11132
rect 2608 11073 2636 11104
rect 4246 11092 4252 11104
rect 4304 11132 4310 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4304 11104 4629 11132
rect 4304 11092 4310 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4816 11132 4844 11163
rect 5350 11160 5356 11212
rect 5408 11160 5414 11212
rect 6365 11203 6423 11209
rect 6365 11169 6377 11203
rect 6411 11200 6423 11203
rect 6546 11200 6552 11212
rect 6411 11172 6552 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 8573 11203 8631 11209
rect 8573 11200 8585 11203
rect 8496 11172 8585 11200
rect 4982 11132 4988 11144
rect 4816 11104 4988 11132
rect 4617 11095 4675 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 6638 11092 6644 11144
rect 6696 11092 6702 11144
rect 8110 11092 8116 11144
rect 8168 11132 8174 11144
rect 8496 11141 8524 11172
rect 8573 11169 8585 11172
rect 8619 11169 8631 11203
rect 8573 11163 8631 11169
rect 8846 11160 8852 11212
rect 8904 11160 8910 11212
rect 9214 11160 9220 11212
rect 9272 11160 9278 11212
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 10428 11209 10456 11240
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 9456 11172 9505 11200
rect 9456 11160 9462 11172
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 8481 11135 8539 11141
rect 8481 11132 8493 11135
rect 8168 11104 8493 11132
rect 8168 11092 8174 11104
rect 8481 11101 8493 11104
rect 8527 11101 8539 11135
rect 9508 11132 9536 11163
rect 10870 11160 10876 11212
rect 10928 11200 10934 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 10928 11172 11253 11200
rect 10928 11160 10934 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 11655 11172 11744 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 11146 11132 11152 11144
rect 9508 11104 11152 11132
rect 8481 11095 8539 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11716 11132 11744 11172
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 13081 11203 13139 11209
rect 13081 11200 13093 11203
rect 12860 11172 13093 11200
rect 12860 11160 12866 11172
rect 13081 11169 13093 11172
rect 13127 11200 13139 11203
rect 13170 11200 13176 11212
rect 13127 11172 13176 11200
rect 13127 11169 13139 11172
rect 13081 11163 13139 11169
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 13906 11200 13912 11212
rect 13372 11172 13912 11200
rect 11517 11095 11575 11101
rect 11624 11104 11744 11132
rect 2593 11067 2651 11073
rect 2593 11033 2605 11067
rect 2639 11033 2651 11067
rect 2593 11027 2651 11033
rect 3878 11024 3884 11076
rect 3936 11024 3942 11076
rect 4338 11064 4344 11076
rect 3988 11036 4344 11064
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 3988 10996 4016 11036
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 5166 11064 5172 11076
rect 4448 11036 5172 11064
rect 3292 10968 4016 10996
rect 3292 10956 3298 10968
rect 4062 10956 4068 11008
rect 4120 10956 4126 11008
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 4448 11005 4476 11036
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 7285 11067 7343 11073
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 11054 11064 11060 11076
rect 7331 11036 8432 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 4433 10999 4491 11005
rect 4433 10996 4445 10999
rect 4304 10968 4445 10996
rect 4304 10956 4310 10968
rect 4433 10965 4445 10968
rect 4479 10965 4491 10999
rect 4433 10959 4491 10965
rect 4525 10999 4583 11005
rect 4525 10965 4537 10999
rect 4571 10996 4583 10999
rect 4798 10996 4804 11008
rect 4571 10968 4804 10996
rect 4571 10965 4583 10968
rect 4525 10959 4583 10965
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 8113 10999 8171 11005
rect 8113 10965 8125 10999
rect 8159 10996 8171 10999
rect 8202 10996 8208 11008
rect 8159 10968 8208 10996
rect 8159 10965 8171 10968
rect 8113 10959 8171 10965
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8404 10996 8432 11036
rect 8588 11036 11060 11064
rect 8588 10996 8616 11036
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11238 11024 11244 11076
rect 11296 11064 11302 11076
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 11296 11036 11437 11064
rect 11296 11024 11302 11036
rect 11425 11033 11437 11036
rect 11471 11033 11483 11067
rect 11425 11027 11483 11033
rect 8404 10968 8616 10996
rect 9214 10956 9220 11008
rect 9272 10996 9278 11008
rect 9309 10999 9367 11005
rect 9309 10996 9321 10999
rect 9272 10968 9321 10996
rect 9272 10956 9278 10968
rect 9309 10965 9321 10968
rect 9355 10965 9367 10999
rect 11072 10996 11100 11024
rect 11532 10996 11560 11095
rect 11624 11076 11652 11104
rect 11882 11092 11888 11144
rect 11940 11092 11946 11144
rect 13372 11141 13400 11172
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 14016 11209 14044 11308
rect 14090 11296 14096 11348
rect 14148 11296 14154 11348
rect 14274 11296 14280 11348
rect 14332 11296 14338 11348
rect 14458 11296 14464 11348
rect 14516 11296 14522 11348
rect 14918 11296 14924 11348
rect 14976 11296 14982 11348
rect 16114 11336 16120 11348
rect 15856 11308 16120 11336
rect 14476 11268 14504 11296
rect 14936 11268 14964 11296
rect 14200 11240 14504 11268
rect 14844 11240 14964 11268
rect 14001 11203 14059 11209
rect 14001 11169 14013 11203
rect 14047 11169 14059 11203
rect 14001 11163 14059 11169
rect 14090 11160 14096 11212
rect 14148 11200 14154 11212
rect 14200 11209 14228 11240
rect 14185 11203 14243 11209
rect 14185 11200 14197 11203
rect 14148 11172 14197 11200
rect 14148 11160 14154 11172
rect 14185 11169 14197 11172
rect 14231 11169 14243 11203
rect 14185 11163 14243 11169
rect 14461 11203 14519 11209
rect 14844 11206 14872 11240
rect 15378 11228 15384 11280
rect 15436 11268 15442 11280
rect 15856 11277 15884 11308
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 19150 11336 19156 11348
rect 18923 11308 19156 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 19886 11336 19892 11348
rect 19720 11308 19892 11336
rect 15657 11271 15715 11277
rect 15657 11268 15669 11271
rect 15436 11240 15669 11268
rect 15436 11228 15442 11240
rect 15657 11237 15669 11240
rect 15703 11237 15715 11271
rect 15657 11231 15715 11237
rect 15841 11271 15899 11277
rect 15841 11237 15853 11271
rect 15887 11237 15899 11271
rect 16390 11268 16396 11280
rect 15841 11231 15899 11237
rect 16040 11240 16396 11268
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 14660 11200 14872 11206
rect 16040 11200 16068 11240
rect 16390 11228 16396 11240
rect 16448 11268 16454 11280
rect 18230 11268 18236 11280
rect 16448 11240 17908 11268
rect 16448 11228 16454 11240
rect 14507 11178 14872 11200
rect 14507 11172 14688 11178
rect 15028 11172 16068 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13630 11092 13636 11144
rect 13688 11132 13694 11144
rect 15028 11132 15056 11172
rect 16114 11160 16120 11212
rect 16172 11160 16178 11212
rect 16758 11160 16764 11212
rect 16816 11160 16822 11212
rect 17586 11160 17592 11212
rect 17644 11160 17650 11212
rect 17880 11209 17908 11240
rect 18064 11240 18236 11268
rect 18064 11209 18092 11240
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 18509 11271 18567 11277
rect 18509 11237 18521 11271
rect 18555 11268 18567 11271
rect 19720 11268 19748 11308
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 20257 11339 20315 11345
rect 20257 11305 20269 11339
rect 20303 11336 20315 11339
rect 20530 11336 20536 11348
rect 20303 11308 20536 11336
rect 20303 11305 20315 11308
rect 20257 11299 20315 11305
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 20622 11296 20628 11348
rect 20680 11296 20686 11348
rect 20990 11296 20996 11348
rect 21048 11336 21054 11348
rect 21048 11308 21404 11336
rect 21048 11296 21054 11308
rect 18555 11240 19748 11268
rect 18555 11237 18567 11240
rect 18509 11231 18567 11237
rect 19794 11228 19800 11280
rect 19852 11268 19858 11280
rect 20165 11271 20223 11277
rect 20165 11268 20177 11271
rect 19852 11240 20177 11268
rect 19852 11228 19858 11240
rect 20165 11237 20177 11240
rect 20211 11268 20223 11271
rect 20640 11268 20668 11296
rect 21376 11268 21404 11308
rect 21514 11271 21572 11277
rect 21514 11268 21526 11271
rect 20211 11240 20392 11268
rect 20640 11240 21312 11268
rect 21376 11240 21526 11268
rect 20211 11237 20223 11240
rect 20165 11231 20223 11237
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11169 18107 11203
rect 18414 11200 18420 11212
rect 18049 11163 18107 11169
rect 18156 11172 18420 11200
rect 13688 11104 15056 11132
rect 13688 11092 13694 11104
rect 15102 11092 15108 11144
rect 15160 11092 15166 11144
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 15436 11104 16221 11132
rect 15436 11092 15442 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16776 11132 16804 11160
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 16776 11104 17325 11132
rect 16209 11095 16267 11101
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 17954 11092 17960 11144
rect 18012 11092 18018 11144
rect 18156 11141 18184 11172
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11200 18751 11203
rect 18782 11200 18788 11212
rect 18739 11172 18788 11200
rect 18739 11169 18751 11172
rect 18693 11163 18751 11169
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11132 18383 11135
rect 19702 11132 19708 11144
rect 18371 11104 19708 11132
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 19702 11092 19708 11104
rect 19760 11092 19766 11144
rect 19981 11135 20039 11141
rect 19981 11101 19993 11135
rect 20027 11132 20039 11135
rect 20364 11132 20392 11240
rect 20622 11160 20628 11212
rect 20680 11200 20686 11212
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 20680 11172 20913 11200
rect 20680 11160 20686 11172
rect 20901 11169 20913 11172
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 21082 11160 21088 11212
rect 21140 11160 21146 11212
rect 21284 11209 21312 11240
rect 21514 11237 21526 11240
rect 21560 11237 21572 11271
rect 21514 11231 21572 11237
rect 21269 11203 21327 11209
rect 21269 11169 21281 11203
rect 21315 11169 21327 11203
rect 21269 11163 21327 11169
rect 20717 11135 20775 11141
rect 20717 11132 20729 11135
rect 20027 11104 20208 11132
rect 20364 11104 20729 11132
rect 20027 11101 20039 11104
rect 19981 11095 20039 11101
rect 11606 11024 11612 11076
rect 11664 11024 11670 11076
rect 13262 11024 13268 11076
rect 13320 11064 13326 11076
rect 20070 11064 20076 11076
rect 13320 11036 20076 11064
rect 13320 11024 13326 11036
rect 20070 11024 20076 11036
rect 20128 11024 20134 11076
rect 20180 11064 20208 11104
rect 20717 11101 20729 11104
rect 20763 11101 20775 11135
rect 20717 11095 20775 11101
rect 20625 11067 20683 11073
rect 20180 11036 20300 11064
rect 20272 11008 20300 11036
rect 20625 11033 20637 11067
rect 20671 11064 20683 11067
rect 20671 11036 20760 11064
rect 20671 11033 20683 11036
rect 20625 11027 20683 11033
rect 20732 11008 20760 11036
rect 11072 10968 11560 10996
rect 9309 10959 9367 10965
rect 15470 10956 15476 11008
rect 15528 10956 15534 11008
rect 17770 10956 17776 11008
rect 17828 10996 17834 11008
rect 20254 10996 20260 11008
rect 17828 10968 20260 10996
rect 17828 10956 17834 10968
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 20714 10956 20720 11008
rect 20772 10956 20778 11008
rect 22278 10956 22284 11008
rect 22336 10996 22342 11008
rect 22649 10999 22707 11005
rect 22649 10996 22661 10999
rect 22336 10968 22661 10996
rect 22336 10956 22342 10968
rect 22649 10965 22661 10968
rect 22695 10965 22707 10999
rect 22649 10959 22707 10965
rect 552 10906 23368 10928
rect 552 10854 1366 10906
rect 1418 10854 1430 10906
rect 1482 10854 1494 10906
rect 1546 10854 1558 10906
rect 1610 10854 1622 10906
rect 1674 10854 1686 10906
rect 1738 10854 7366 10906
rect 7418 10854 7430 10906
rect 7482 10854 7494 10906
rect 7546 10854 7558 10906
rect 7610 10854 7622 10906
rect 7674 10854 7686 10906
rect 7738 10854 13366 10906
rect 13418 10854 13430 10906
rect 13482 10854 13494 10906
rect 13546 10854 13558 10906
rect 13610 10854 13622 10906
rect 13674 10854 13686 10906
rect 13738 10854 19366 10906
rect 19418 10854 19430 10906
rect 19482 10854 19494 10906
rect 19546 10854 19558 10906
rect 19610 10854 19622 10906
rect 19674 10854 19686 10906
rect 19738 10854 23368 10906
rect 552 10832 23368 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 1857 10795 1915 10801
rect 1857 10792 1869 10795
rect 1820 10764 1869 10792
rect 1820 10752 1826 10764
rect 1857 10761 1869 10764
rect 1903 10761 1915 10795
rect 1857 10755 1915 10761
rect 3694 10752 3700 10804
rect 3752 10792 3758 10804
rect 3973 10795 4031 10801
rect 3973 10792 3985 10795
rect 3752 10764 3985 10792
rect 3752 10752 3758 10764
rect 3973 10761 3985 10764
rect 4019 10761 4031 10795
rect 5258 10792 5264 10804
rect 3973 10755 4031 10761
rect 4356 10764 5264 10792
rect 1762 10616 1768 10668
rect 1820 10616 1826 10668
rect 1854 10548 1860 10600
rect 1912 10588 1918 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1912 10560 1961 10588
rect 1912 10548 1918 10560
rect 1949 10557 1961 10560
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 3510 10588 3516 10600
rect 2087 10560 3516 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4062 10588 4068 10600
rect 4019 10560 4068 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 4356 10597 4384 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 6733 10795 6791 10801
rect 6733 10792 6745 10795
rect 6696 10764 6745 10792
rect 6696 10752 6702 10764
rect 6733 10761 6745 10764
rect 6779 10761 6791 10795
rect 6733 10755 6791 10761
rect 8386 10752 8392 10804
rect 8444 10752 8450 10804
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 9033 10795 9091 10801
rect 9033 10792 9045 10795
rect 8904 10764 9045 10792
rect 8904 10752 8910 10764
rect 9033 10761 9045 10764
rect 9079 10761 9091 10795
rect 9033 10755 9091 10761
rect 9490 10752 9496 10804
rect 9548 10752 9554 10804
rect 10870 10752 10876 10804
rect 10928 10752 10934 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11388 10764 11713 10792
rect 11388 10752 11394 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 11701 10755 11759 10761
rect 12176 10764 12572 10792
rect 4798 10724 4804 10736
rect 4724 10696 4804 10724
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4212 10560 4353 10588
rect 4212 10548 4218 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10588 4491 10591
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 4479 10560 4629 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 4617 10551 4675 10557
rect 4724 10520 4752 10696
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 4908 10696 5948 10724
rect 4908 10665 4936 10696
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5166 10616 5172 10668
rect 5224 10656 5230 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 5224 10628 5273 10656
rect 5224 10616 5230 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5592 10628 5856 10656
rect 5592 10616 5598 10628
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10588 5687 10591
rect 5675 10560 5764 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 5736 10532 5764 10560
rect 5828 10532 5856 10628
rect 5920 10588 5948 10696
rect 8110 10684 8116 10736
rect 8168 10724 8174 10736
rect 9125 10727 9183 10733
rect 9125 10724 9137 10727
rect 8168 10696 9137 10724
rect 8168 10684 8174 10696
rect 9125 10693 9137 10696
rect 9171 10693 9183 10727
rect 9125 10687 9183 10693
rect 6273 10659 6331 10665
rect 6273 10625 6285 10659
rect 6319 10656 6331 10659
rect 6454 10656 6460 10668
rect 6319 10628 6460 10656
rect 6319 10625 6331 10628
rect 6273 10619 6331 10625
rect 6454 10616 6460 10628
rect 6512 10656 6518 10668
rect 6822 10656 6828 10668
rect 6512 10628 6828 10656
rect 6512 10616 6518 10628
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 8496 10628 8800 10656
rect 8496 10600 8524 10628
rect 6362 10588 6368 10600
rect 5920 10560 6368 10588
rect 6362 10548 6368 10560
rect 6420 10588 6426 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6420 10560 6561 10588
rect 6420 10548 6426 10560
rect 6549 10557 6561 10560
rect 6595 10588 6607 10591
rect 6914 10588 6920 10600
rect 6595 10560 6920 10588
rect 6595 10557 6607 10560
rect 6549 10551 6607 10557
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 8478 10548 8484 10600
rect 8536 10548 8542 10600
rect 8772 10597 8800 10628
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 8619 10591 8677 10597
rect 8619 10557 8631 10591
rect 8665 10588 8677 10591
rect 8757 10591 8815 10597
rect 8665 10557 8688 10588
rect 8619 10551 8688 10557
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 5169 10523 5227 10529
rect 5169 10520 5181 10523
rect 4724 10492 5181 10520
rect 5169 10489 5181 10492
rect 5215 10489 5227 10523
rect 5718 10520 5724 10532
rect 5169 10483 5227 10489
rect 5368 10492 5724 10520
rect 3786 10412 3792 10464
rect 3844 10412 3850 10464
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 5368 10452 5396 10492
rect 5718 10480 5724 10492
rect 5776 10480 5782 10532
rect 5810 10480 5816 10532
rect 5868 10520 5874 10532
rect 6825 10523 6883 10529
rect 6825 10520 6837 10523
rect 5868 10492 6837 10520
rect 5868 10480 5874 10492
rect 6825 10489 6837 10492
rect 6871 10489 6883 10523
rect 6825 10483 6883 10489
rect 5123 10424 5396 10452
rect 5445 10455 5503 10461
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 5445 10421 5457 10455
rect 5491 10452 5503 10455
rect 5534 10452 5540 10464
rect 5491 10424 5540 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 8660 10452 8688 10551
rect 8846 10548 8852 10600
rect 8904 10548 8910 10600
rect 9508 10597 9536 10752
rect 11054 10684 11060 10736
rect 11112 10724 11118 10736
rect 12069 10727 12127 10733
rect 12069 10724 12081 10727
rect 11112 10696 12081 10724
rect 11112 10684 11118 10696
rect 12069 10693 12081 10696
rect 12115 10693 12127 10727
rect 12069 10687 12127 10693
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 10008 10628 11345 10656
rect 10008 10616 10014 10628
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 12176 10656 12204 10764
rect 12437 10727 12495 10733
rect 12437 10693 12449 10727
rect 12483 10693 12495 10727
rect 12544 10724 12572 10764
rect 12618 10752 12624 10804
rect 12676 10792 12682 10804
rect 12713 10795 12771 10801
rect 12713 10792 12725 10795
rect 12676 10764 12725 10792
rect 12676 10752 12682 10764
rect 12713 10761 12725 10764
rect 12759 10761 12771 10795
rect 12713 10755 12771 10761
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 13228 10764 14381 10792
rect 13228 10752 13234 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 14369 10755 14427 10761
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 15896 10764 16313 10792
rect 15896 10752 15902 10764
rect 16301 10761 16313 10764
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 17313 10795 17371 10801
rect 17313 10792 17325 10795
rect 16448 10764 17325 10792
rect 16448 10752 16454 10764
rect 17313 10761 17325 10764
rect 17359 10761 17371 10795
rect 17313 10755 17371 10761
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18877 10795 18935 10801
rect 18877 10792 18889 10795
rect 18288 10764 18889 10792
rect 18288 10752 18294 10764
rect 18877 10761 18889 10764
rect 18923 10761 18935 10795
rect 18877 10755 18935 10761
rect 19613 10795 19671 10801
rect 19613 10761 19625 10795
rect 19659 10792 19671 10795
rect 19794 10792 19800 10804
rect 19659 10764 19800 10792
rect 19659 10761 19671 10764
rect 19613 10755 19671 10761
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 19886 10752 19892 10804
rect 19944 10752 19950 10804
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 19996 10764 20269 10792
rect 13541 10727 13599 10733
rect 13541 10724 13553 10727
rect 12544 10696 13553 10724
rect 12437 10687 12495 10693
rect 13541 10693 13553 10696
rect 13587 10693 13599 10727
rect 13906 10724 13912 10736
rect 13541 10687 13599 10693
rect 13648 10696 13912 10724
rect 11333 10619 11391 10625
rect 11538 10628 11836 10656
rect 9493 10591 9551 10597
rect 9216 10569 9274 10575
rect 9216 10535 9228 10569
rect 9262 10535 9274 10569
rect 9493 10557 9505 10591
rect 9539 10588 9551 10591
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 9539 10560 11069 10588
rect 9539 10557 9551 10560
rect 9493 10551 9551 10557
rect 11057 10557 11069 10560
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11241 10591 11299 10597
rect 11241 10588 11253 10591
rect 11204 10560 11253 10588
rect 11204 10548 11210 10560
rect 11241 10557 11253 10560
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 11422 10548 11428 10600
rect 11480 10548 11486 10600
rect 9216 10532 9274 10535
rect 9214 10480 9220 10532
rect 9272 10480 9278 10532
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 11538 10520 11566 10628
rect 11808 10600 11836 10628
rect 11900 10628 12204 10656
rect 11609 10591 11667 10597
rect 11609 10557 11621 10591
rect 11655 10588 11667 10591
rect 11655 10560 11744 10588
rect 11655 10557 11667 10560
rect 11609 10551 11667 10557
rect 9456 10492 11566 10520
rect 11716 10520 11744 10560
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 11900 10597 11928 10628
rect 12452 10600 12480 10687
rect 12802 10616 12808 10668
rect 12860 10616 12866 10668
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 12158 10548 12164 10600
rect 12216 10548 12222 10600
rect 12434 10588 12440 10600
rect 12268 10560 12440 10588
rect 12268 10520 12296 10560
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 12621 10591 12679 10597
rect 12621 10557 12633 10591
rect 12667 10588 12679 10591
rect 12820 10588 12848 10616
rect 12667 10560 12848 10588
rect 12667 10557 12679 10560
rect 12621 10551 12679 10557
rect 12986 10548 12992 10600
rect 13044 10548 13050 10600
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 11716 10492 12296 10520
rect 9456 10480 9462 10492
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 8536 10424 9321 10452
rect 8536 10412 8542 10424
rect 9309 10421 9321 10424
rect 9355 10452 9367 10455
rect 11330 10452 11336 10464
rect 9355 10424 11336 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 11422 10412 11428 10464
rect 11480 10452 11486 10464
rect 13096 10452 13124 10551
rect 13170 10548 13176 10600
rect 13228 10548 13234 10600
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 13372 10520 13400 10551
rect 13648 10520 13676 10696
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 14921 10727 14979 10733
rect 14921 10693 14933 10727
rect 14967 10724 14979 10727
rect 17589 10727 17647 10733
rect 17589 10724 17601 10727
rect 14967 10696 17601 10724
rect 14967 10693 14979 10696
rect 14921 10687 14979 10693
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 15378 10656 15384 10668
rect 13872 10628 14044 10656
rect 13872 10616 13878 10628
rect 13722 10548 13728 10600
rect 13780 10548 13786 10600
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 14016 10597 14044 10628
rect 15120 10628 15384 10656
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10557 14059 10591
rect 14001 10551 14059 10557
rect 14090 10548 14096 10600
rect 14148 10548 14154 10600
rect 14182 10548 14188 10600
rect 14240 10578 14246 10600
rect 14550 10588 14556 10600
rect 14277 10581 14335 10587
rect 14277 10578 14289 10581
rect 14240 10550 14289 10578
rect 14240 10548 14246 10550
rect 14277 10547 14289 10550
rect 14323 10547 14335 10581
rect 14511 10560 14556 10588
rect 14550 10548 14556 10560
rect 14608 10548 14614 10600
rect 14642 10548 14648 10600
rect 14700 10588 14706 10600
rect 15120 10597 15148 10628
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10656 16727 10659
rect 17034 10656 17040 10668
rect 16715 10628 17040 10656
rect 16715 10625 16727 10628
rect 16669 10619 16727 10625
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 17144 10600 17172 10696
rect 17589 10693 17601 10696
rect 17635 10693 17647 10727
rect 17589 10687 17647 10693
rect 19996 10656 20024 10764
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 20257 10755 20315 10761
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 19168 10628 20024 10656
rect 20088 10696 22876 10724
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14700 10560 15025 10588
rect 14700 10548 14706 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15105 10591 15163 10597
rect 15105 10557 15117 10591
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 15286 10548 15292 10600
rect 15344 10548 15350 10600
rect 15657 10591 15715 10597
rect 15657 10557 15669 10591
rect 15703 10588 15715 10591
rect 16114 10588 16120 10600
rect 15703 10560 16120 10588
rect 15703 10557 15715 10560
rect 15657 10551 15715 10557
rect 16114 10548 16120 10560
rect 16172 10548 16178 10600
rect 16206 10548 16212 10600
rect 16264 10588 16270 10600
rect 16485 10591 16543 10597
rect 16485 10588 16497 10591
rect 16264 10560 16497 10588
rect 16264 10548 16270 10560
rect 16485 10557 16497 10560
rect 16531 10557 16543 10591
rect 16485 10551 16543 10557
rect 16577 10591 16635 10597
rect 16577 10557 16589 10591
rect 16623 10557 16635 10591
rect 16577 10551 16635 10557
rect 14277 10541 14335 10547
rect 13814 10520 13820 10532
rect 13372 10492 13820 10520
rect 13814 10480 13820 10492
rect 13872 10480 13878 10532
rect 16592 10520 16620 10551
rect 16758 10548 16764 10600
rect 16816 10548 16822 10600
rect 17126 10548 17132 10600
rect 17184 10548 17190 10600
rect 17405 10591 17463 10597
rect 17405 10557 17417 10591
rect 17451 10588 17463 10591
rect 17586 10588 17592 10600
rect 17451 10560 17592 10588
rect 17451 10557 17463 10560
rect 17405 10551 17463 10557
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 19168 10597 19196 10628
rect 19061 10591 19119 10597
rect 19061 10557 19073 10591
rect 19107 10557 19119 10591
rect 19061 10551 19119 10557
rect 19153 10591 19211 10597
rect 19153 10557 19165 10591
rect 19199 10557 19211 10591
rect 19153 10551 19211 10557
rect 14384 10492 16620 10520
rect 19076 10520 19104 10551
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19392 10560 19441 10588
rect 19392 10548 19398 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 19843 10557 19901 10563
rect 19245 10523 19303 10529
rect 19245 10520 19257 10523
rect 19076 10492 19257 10520
rect 11480 10424 13124 10452
rect 11480 10412 11486 10424
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 14384 10452 14412 10492
rect 19245 10489 19257 10492
rect 19291 10520 19303 10523
rect 19843 10523 19855 10557
rect 19889 10523 19901 10557
rect 20088 10529 20116 10696
rect 22848 10668 22876 10696
rect 20254 10616 20260 10668
rect 20312 10656 20318 10668
rect 21545 10659 21603 10665
rect 21545 10656 21557 10659
rect 20312 10628 21557 10656
rect 20312 10616 20318 10628
rect 21545 10625 21557 10628
rect 21591 10625 21603 10659
rect 21545 10619 21603 10625
rect 22094 10616 22100 10668
rect 22152 10656 22158 10668
rect 22152 10628 22416 10656
rect 22152 10616 22158 10628
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 19843 10520 19901 10523
rect 19291 10492 19748 10520
rect 19291 10489 19303 10492
rect 19245 10483 19303 10489
rect 13228 10424 14412 10452
rect 13228 10412 13234 10424
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 14516 10424 14565 10452
rect 14516 10412 14522 10424
rect 14553 10421 14565 10424
rect 14599 10421 14611 10455
rect 14553 10415 14611 10421
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15378 10452 15384 10464
rect 15335 10424 15384 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 18506 10452 18512 10464
rect 17276 10424 18512 10452
rect 17276 10412 17282 10424
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 19720 10461 19748 10492
rect 19812 10517 19901 10520
rect 20073 10523 20131 10529
rect 19812 10492 19886 10517
rect 19812 10464 19840 10492
rect 20073 10489 20085 10523
rect 20119 10489 20131 10523
rect 20073 10483 20131 10489
rect 19705 10455 19763 10461
rect 19705 10421 19717 10455
rect 19751 10421 19763 10455
rect 19705 10415 19763 10421
rect 19794 10412 19800 10464
rect 19852 10412 19858 10464
rect 19978 10412 19984 10464
rect 20036 10452 20042 10464
rect 20180 10452 20208 10551
rect 20714 10548 20720 10600
rect 20772 10548 20778 10600
rect 20806 10548 20812 10600
rect 20864 10548 20870 10600
rect 22204 10597 22232 10628
rect 21821 10591 21879 10597
rect 21821 10557 21833 10591
rect 21867 10588 21879 10591
rect 22189 10591 22247 10597
rect 22189 10588 22201 10591
rect 21867 10560 22201 10588
rect 21867 10557 21879 10560
rect 21821 10551 21879 10557
rect 22189 10557 22201 10560
rect 22235 10557 22247 10591
rect 22189 10551 22247 10557
rect 22278 10548 22284 10600
rect 22336 10548 22342 10600
rect 22388 10588 22416 10628
rect 22830 10616 22836 10668
rect 22888 10616 22894 10668
rect 22388 10560 22968 10588
rect 20824 10520 20852 10548
rect 21913 10523 21971 10529
rect 21913 10520 21925 10523
rect 20824 10492 21925 10520
rect 21913 10489 21925 10492
rect 21959 10489 21971 10523
rect 21913 10483 21971 10489
rect 22097 10523 22155 10529
rect 22097 10489 22109 10523
rect 22143 10520 22155 10523
rect 22296 10520 22324 10548
rect 22143 10492 22324 10520
rect 22143 10489 22155 10492
rect 22097 10483 22155 10489
rect 22940 10464 22968 10560
rect 20036 10424 20208 10452
rect 20036 10412 20042 10424
rect 21818 10412 21824 10464
rect 21876 10452 21882 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21876 10424 22017 10452
rect 21876 10412 21882 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 22922 10412 22928 10464
rect 22980 10412 22986 10464
rect 552 10362 23368 10384
rect 552 10310 4366 10362
rect 4418 10310 4430 10362
rect 4482 10310 4494 10362
rect 4546 10310 4558 10362
rect 4610 10310 4622 10362
rect 4674 10310 4686 10362
rect 4738 10310 10366 10362
rect 10418 10310 10430 10362
rect 10482 10310 10494 10362
rect 10546 10310 10558 10362
rect 10610 10310 10622 10362
rect 10674 10310 10686 10362
rect 10738 10310 16366 10362
rect 16418 10310 16430 10362
rect 16482 10310 16494 10362
rect 16546 10310 16558 10362
rect 16610 10310 16622 10362
rect 16674 10310 16686 10362
rect 16738 10310 22366 10362
rect 22418 10310 22430 10362
rect 22482 10310 22494 10362
rect 22546 10310 22558 10362
rect 22610 10310 22622 10362
rect 22674 10310 22686 10362
rect 22738 10310 23368 10362
rect 552 10288 23368 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 1857 10251 1915 10257
rect 1857 10248 1869 10251
rect 1820 10220 1869 10248
rect 1820 10208 1826 10220
rect 1857 10217 1869 10220
rect 1903 10217 1915 10251
rect 2130 10248 2136 10260
rect 1857 10211 1915 10217
rect 1964 10220 2136 10248
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 1670 10112 1676 10124
rect 1627 10084 1676 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 1964 10121 1992 10220
rect 2130 10208 2136 10220
rect 2188 10248 2194 10260
rect 2317 10251 2375 10257
rect 2317 10248 2329 10251
rect 2188 10220 2329 10248
rect 2188 10208 2194 10220
rect 2317 10217 2329 10220
rect 2363 10217 2375 10251
rect 6730 10248 6736 10260
rect 2317 10211 2375 10217
rect 3436 10220 6736 10248
rect 2240 10152 2636 10180
rect 2240 10121 2268 10152
rect 2608 10124 2636 10152
rect 2682 10140 2688 10192
rect 2740 10140 2746 10192
rect 3234 10189 3240 10192
rect 3221 10183 3240 10189
rect 3221 10149 3233 10183
rect 3221 10143 3240 10149
rect 3234 10140 3240 10143
rect 3292 10140 3298 10192
rect 3436 10189 3464 10220
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8205 10251 8263 10257
rect 8205 10248 8217 10251
rect 8168 10220 8217 10248
rect 8168 10208 8174 10220
rect 8205 10217 8217 10220
rect 8251 10217 8263 10251
rect 8205 10211 8263 10217
rect 8478 10208 8484 10260
rect 8536 10208 8542 10260
rect 11054 10248 11060 10260
rect 10612 10220 11060 10248
rect 3421 10183 3479 10189
rect 3421 10149 3433 10183
rect 3467 10149 3479 10183
rect 5534 10180 5540 10192
rect 3421 10143 3479 10149
rect 4172 10152 5540 10180
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10081 2007 10115
rect 1949 10075 2007 10081
rect 2133 10115 2191 10121
rect 2133 10081 2145 10115
rect 2179 10081 2191 10115
rect 2133 10075 2191 10081
rect 2225 10115 2283 10121
rect 2225 10081 2237 10115
rect 2271 10081 2283 10115
rect 2225 10075 2283 10081
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10081 2559 10115
rect 2501 10075 2559 10081
rect 1210 10004 1216 10056
rect 1268 10004 1274 10056
rect 1228 9976 1256 10004
rect 1949 9979 2007 9985
rect 1949 9976 1961 9979
rect 1228 9948 1961 9976
rect 1949 9945 1961 9948
rect 1995 9945 2007 9979
rect 1949 9939 2007 9945
rect 1118 9868 1124 9920
rect 1176 9908 1182 9920
rect 1397 9911 1455 9917
rect 1397 9908 1409 9911
rect 1176 9880 1409 9908
rect 1176 9868 1182 9880
rect 1397 9877 1409 9880
rect 1443 9908 1455 9911
rect 2038 9908 2044 9920
rect 1443 9880 2044 9908
rect 1443 9877 1455 9880
rect 1397 9871 1455 9877
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 2148 9908 2176 10075
rect 2516 9976 2544 10075
rect 2590 10072 2596 10124
rect 2648 10072 2654 10124
rect 2823 10115 2881 10121
rect 2823 10081 2835 10115
rect 2869 10081 2881 10115
rect 2823 10075 2881 10081
rect 2838 10044 2866 10075
rect 3326 10072 3332 10124
rect 3384 10112 3390 10124
rect 4172 10112 4200 10152
rect 3384 10084 4200 10112
rect 3384 10072 3390 10084
rect 4246 10072 4252 10124
rect 4304 10112 4310 10124
rect 5368 10121 5396 10152
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 8496 10180 8524 10208
rect 8573 10183 8631 10189
rect 8573 10180 8585 10183
rect 8343 10149 8401 10155
rect 8496 10152 8585 10180
rect 8343 10124 8355 10149
rect 4617 10115 4675 10121
rect 4617 10112 4629 10115
rect 4304 10084 4629 10112
rect 4304 10072 4310 10084
rect 4617 10081 4629 10084
rect 4663 10081 4675 10115
rect 4617 10075 4675 10081
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5353 10075 5411 10081
rect 2961 10047 3019 10053
rect 2838 10016 2912 10044
rect 2884 9988 2912 10016
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 4816 10044 4844 10075
rect 7834 10072 7840 10124
rect 7892 10072 7898 10124
rect 8294 10072 8300 10124
rect 8352 10115 8355 10124
rect 8389 10146 8401 10149
rect 8573 10149 8585 10152
rect 8619 10149 8631 10183
rect 8846 10180 8852 10192
rect 8389 10115 8416 10146
rect 8573 10143 8631 10149
rect 8772 10152 8852 10180
rect 8352 10084 8416 10115
rect 8352 10072 8358 10084
rect 8662 10072 8668 10124
rect 8720 10072 8726 10124
rect 8772 10053 8800 10152
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 9030 10072 9036 10124
rect 9088 10072 9094 10124
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 8757 10047 8815 10053
rect 8757 10044 8769 10047
rect 4816 10016 6040 10044
rect 2961 10007 3019 10013
rect 2774 9976 2780 9988
rect 2516 9948 2780 9976
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 2866 9936 2872 9988
rect 2924 9936 2930 9988
rect 2976 9976 3004 10007
rect 6012 9988 6040 10016
rect 7944 10016 8769 10044
rect 3053 9979 3111 9985
rect 3053 9976 3065 9979
rect 2976 9948 3065 9976
rect 3053 9945 3065 9948
rect 3099 9945 3111 9979
rect 3053 9939 3111 9945
rect 5994 9936 6000 9988
rect 6052 9976 6058 9988
rect 6178 9976 6184 9988
rect 6052 9948 6184 9976
rect 6052 9936 6058 9948
rect 6178 9936 6184 9948
rect 6236 9936 6242 9988
rect 2884 9908 2912 9936
rect 7944 9920 7972 10016
rect 8757 10013 8769 10016
rect 8803 10013 8815 10047
rect 8757 10007 8815 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10044 8999 10047
rect 9048 10044 9076 10072
rect 8987 10016 9076 10044
rect 9232 10044 9260 10075
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10612 10121 10640 10220
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11422 10248 11428 10260
rect 11256 10220 11428 10248
rect 10781 10183 10839 10189
rect 10781 10149 10793 10183
rect 10827 10180 10839 10183
rect 10827 10152 11192 10180
rect 10827 10149 10839 10152
rect 10781 10143 10839 10149
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 10008 10084 10241 10112
rect 10008 10072 10014 10084
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10081 10655 10115
rect 10597 10075 10655 10081
rect 9306 10044 9312 10056
rect 9232 10016 9312 10044
rect 8987 10013 8999 10016
rect 8941 10007 8999 10013
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 10520 10044 10548 10075
rect 10962 10072 10968 10124
rect 11020 10072 11026 10124
rect 11164 10121 11192 10152
rect 11256 10124 11284 10220
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11698 10248 11704 10260
rect 11655 10220 11704 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 13722 10248 13728 10260
rect 11808 10220 13728 10248
rect 11808 10180 11836 10220
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 15286 10248 15292 10260
rect 14148 10220 15292 10248
rect 14148 10208 14154 10220
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 16669 10251 16727 10257
rect 16669 10217 16681 10251
rect 16715 10248 16727 10251
rect 16758 10248 16764 10260
rect 16715 10220 16764 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 16758 10208 16764 10220
rect 16816 10208 16822 10260
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 17221 10251 17279 10257
rect 17221 10248 17233 10251
rect 17184 10220 17233 10248
rect 17184 10208 17190 10220
rect 17221 10217 17233 10220
rect 17267 10248 17279 10251
rect 18690 10248 18696 10260
rect 17267 10220 18696 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 18969 10251 19027 10257
rect 18969 10217 18981 10251
rect 19015 10248 19027 10251
rect 19058 10248 19064 10260
rect 19015 10220 19064 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 19334 10208 19340 10260
rect 19392 10248 19398 10260
rect 20162 10248 20168 10260
rect 19392 10220 20168 10248
rect 19392 10208 19398 10220
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 21542 10208 21548 10260
rect 21600 10208 21606 10260
rect 22186 10208 22192 10260
rect 22244 10208 22250 10260
rect 11440 10152 11836 10180
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10081 11207 10115
rect 11149 10075 11207 10081
rect 11238 10072 11244 10124
rect 11296 10072 11302 10124
rect 11330 10072 11336 10124
rect 11388 10121 11394 10124
rect 11388 10115 11411 10121
rect 11399 10112 11411 10115
rect 11440 10112 11468 10152
rect 12618 10140 12624 10192
rect 12676 10180 12682 10192
rect 13265 10183 13323 10189
rect 12676 10152 13124 10180
rect 12676 10140 12682 10152
rect 12986 10112 12992 10124
rect 11399 10084 11468 10112
rect 11716 10084 12992 10112
rect 11399 10081 11411 10084
rect 11388 10075 11411 10081
rect 11388 10072 11394 10075
rect 11054 10044 11060 10056
rect 10520 10016 11060 10044
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 9033 9979 9091 9985
rect 9033 9976 9045 9979
rect 8680 9948 9045 9976
rect 8680 9920 8708 9948
rect 9033 9945 9045 9948
rect 9079 9945 9091 9979
rect 9033 9939 9091 9945
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 11716 9976 11744 10084
rect 12986 10072 12992 10084
rect 13044 10072 13050 10124
rect 13096 10121 13124 10152
rect 13265 10149 13277 10183
rect 13311 10180 13323 10183
rect 13541 10183 13599 10189
rect 13541 10180 13553 10183
rect 13311 10152 13553 10180
rect 13311 10149 13323 10152
rect 13265 10143 13323 10149
rect 13541 10149 13553 10152
rect 13587 10149 13599 10183
rect 14734 10180 14740 10192
rect 13541 10143 13599 10149
rect 13648 10152 14740 10180
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 13648 10121 13676 10152
rect 14734 10140 14740 10152
rect 14792 10140 14798 10192
rect 21361 10183 21419 10189
rect 21361 10180 21373 10183
rect 16868 10152 21373 10180
rect 16868 10124 16896 10152
rect 21361 10149 21373 10152
rect 21407 10149 21419 10183
rect 21361 10143 21419 10149
rect 21560 10152 22094 10180
rect 13357 10115 13415 10121
rect 13357 10112 13369 10115
rect 13228 10084 13369 10112
rect 13228 10072 13234 10084
rect 13357 10081 13369 10084
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 12710 10004 12716 10056
rect 12768 10004 12774 10056
rect 13464 10044 13492 10075
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14274 10112 14280 10124
rect 14056 10084 14280 10112
rect 14056 10072 14062 10084
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 14458 10072 14464 10124
rect 14516 10072 14522 10124
rect 14829 10115 14887 10121
rect 14829 10081 14841 10115
rect 14875 10112 14887 10115
rect 14875 10084 15608 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 14476 10044 14504 10072
rect 15580 10056 15608 10084
rect 16022 10072 16028 10124
rect 16080 10112 16086 10124
rect 16666 10112 16672 10124
rect 16080 10084 16672 10112
rect 16080 10072 16086 10084
rect 16666 10072 16672 10084
rect 16724 10072 16730 10124
rect 16850 10072 16856 10124
rect 16908 10072 16914 10124
rect 17083 10115 17141 10121
rect 17083 10081 17095 10115
rect 17129 10112 17141 10115
rect 17129 10084 17448 10112
rect 17129 10081 17141 10084
rect 17083 10075 17141 10081
rect 13464 10016 14504 10044
rect 15562 10004 15568 10056
rect 15620 10004 15626 10056
rect 16206 10004 16212 10056
rect 16264 10044 16270 10056
rect 16574 10044 16580 10056
rect 16264 10016 16580 10044
rect 16264 10004 16270 10016
rect 16574 10004 16580 10016
rect 16632 10044 16638 10056
rect 16945 10047 17003 10053
rect 16945 10044 16957 10047
rect 16632 10016 16957 10044
rect 16632 10004 16638 10016
rect 16945 10013 16957 10016
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 17310 10004 17316 10056
rect 17368 10004 17374 10056
rect 17420 10044 17448 10084
rect 17494 10072 17500 10124
rect 17552 10072 17558 10124
rect 17770 10072 17776 10124
rect 17828 10072 17834 10124
rect 18322 10072 18328 10124
rect 18380 10112 18386 10124
rect 19521 10115 19579 10121
rect 19521 10112 19533 10115
rect 18380 10084 19533 10112
rect 18380 10072 18386 10084
rect 19521 10081 19533 10084
rect 19567 10081 19579 10115
rect 19521 10075 19579 10081
rect 17788 10044 17816 10072
rect 17420 10016 17816 10044
rect 19334 10004 19340 10056
rect 19392 10004 19398 10056
rect 19536 10044 19564 10075
rect 19794 10072 19800 10124
rect 19852 10112 19858 10124
rect 20441 10115 20499 10121
rect 20441 10112 20453 10115
rect 19852 10084 20453 10112
rect 19852 10072 19858 10084
rect 20441 10081 20453 10084
rect 20487 10081 20499 10115
rect 20441 10075 20499 10081
rect 21269 10115 21327 10121
rect 21269 10081 21281 10115
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 19886 10044 19892 10056
rect 19536 10016 19892 10044
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 20070 10004 20076 10056
rect 20128 10044 20134 10056
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 20128 10016 20269 10044
rect 20128 10004 20134 10016
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 9272 9948 11744 9976
rect 9272 9936 9278 9948
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 12728 9976 12756 10004
rect 13081 9979 13139 9985
rect 13081 9976 13093 9979
rect 11848 9948 12388 9976
rect 12728 9948 13093 9976
rect 11848 9936 11854 9948
rect 2148 9880 2912 9908
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 3200 9880 3249 9908
rect 3200 9868 3206 9880
rect 3237 9877 3249 9880
rect 3283 9908 3295 9911
rect 4062 9908 4068 9920
rect 3283 9880 4068 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4706 9868 4712 9920
rect 4764 9868 4770 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 6454 9908 6460 9920
rect 5592 9880 6460 9908
rect 5592 9868 5598 9880
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 6549 9911 6607 9917
rect 6549 9877 6561 9911
rect 6595 9908 6607 9911
rect 7282 9908 7288 9920
rect 6595 9880 7288 9908
rect 6595 9877 6607 9880
rect 6549 9871 6607 9877
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 7926 9868 7932 9920
rect 7984 9868 7990 9920
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8389 9911 8447 9917
rect 8389 9908 8401 9911
rect 8352 9880 8401 9908
rect 8352 9868 8358 9880
rect 8389 9877 8401 9880
rect 8435 9908 8447 9911
rect 8662 9908 8668 9920
rect 8435 9880 8668 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 8846 9868 8852 9920
rect 8904 9868 8910 9920
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 9950 9908 9956 9920
rect 9824 9880 9956 9908
rect 9824 9868 9830 9880
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 10321 9911 10379 9917
rect 10321 9877 10333 9911
rect 10367 9908 10379 9911
rect 10870 9908 10876 9920
rect 10367 9880 10876 9908
rect 10367 9877 10379 9880
rect 10321 9871 10379 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 12360 9908 12388 9948
rect 13081 9945 13093 9948
rect 13127 9945 13139 9979
rect 21174 9976 21180 9988
rect 13081 9939 13139 9945
rect 13280 9948 21180 9976
rect 13280 9908 13308 9948
rect 21174 9936 21180 9948
rect 21232 9976 21238 9988
rect 21284 9976 21312 10075
rect 21232 9948 21312 9976
rect 21232 9936 21238 9948
rect 12360 9880 13308 9908
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14642 9908 14648 9920
rect 13964 9880 14648 9908
rect 13964 9868 13970 9880
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 16114 9908 16120 9920
rect 14792 9880 16120 9908
rect 14792 9868 14798 9880
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 19242 9908 19248 9920
rect 16816 9880 19248 9908
rect 16816 9868 16822 9880
rect 19242 9868 19248 9880
rect 19300 9908 19306 9920
rect 20254 9908 20260 9920
rect 19300 9880 20260 9908
rect 19300 9868 19306 9880
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 20622 9868 20628 9920
rect 20680 9868 20686 9920
rect 21376 9908 21404 10143
rect 21560 10056 21588 10152
rect 21634 10072 21640 10124
rect 21692 10112 21698 10124
rect 21913 10115 21971 10121
rect 21913 10112 21925 10115
rect 21692 10084 21925 10112
rect 21692 10072 21698 10084
rect 21913 10081 21925 10084
rect 21959 10081 21971 10115
rect 22066 10112 22094 10152
rect 22373 10115 22431 10121
rect 22066 10084 22324 10112
rect 21913 10075 21971 10081
rect 21542 10004 21548 10056
rect 21600 10004 21606 10056
rect 21726 10004 21732 10056
rect 21784 10004 21790 10056
rect 21821 10047 21879 10053
rect 21821 10013 21833 10047
rect 21867 10013 21879 10047
rect 21821 10007 21879 10013
rect 22005 10047 22063 10053
rect 22005 10013 22017 10047
rect 22051 10044 22063 10047
rect 22186 10044 22192 10056
rect 22051 10016 22192 10044
rect 22051 10013 22063 10016
rect 22005 10007 22063 10013
rect 21560 9976 21588 10004
rect 21836 9976 21864 10007
rect 22186 10004 22192 10016
rect 22244 10004 22250 10056
rect 22296 10044 22324 10084
rect 22373 10081 22385 10115
rect 22419 10112 22431 10115
rect 22462 10112 22468 10124
rect 22419 10084 22468 10112
rect 22419 10081 22431 10084
rect 22373 10075 22431 10081
rect 22462 10072 22468 10084
rect 22520 10072 22526 10124
rect 22557 10047 22615 10053
rect 22557 10044 22569 10047
rect 22296 10016 22569 10044
rect 22557 10013 22569 10016
rect 22603 10013 22615 10047
rect 22557 10007 22615 10013
rect 21560 9948 21864 9976
rect 22738 9908 22744 9920
rect 21376 9880 22744 9908
rect 22738 9868 22744 9880
rect 22796 9868 22802 9920
rect 552 9818 23368 9840
rect 552 9766 1366 9818
rect 1418 9766 1430 9818
rect 1482 9766 1494 9818
rect 1546 9766 1558 9818
rect 1610 9766 1622 9818
rect 1674 9766 1686 9818
rect 1738 9766 7366 9818
rect 7418 9766 7430 9818
rect 7482 9766 7494 9818
rect 7546 9766 7558 9818
rect 7610 9766 7622 9818
rect 7674 9766 7686 9818
rect 7738 9766 13366 9818
rect 13418 9766 13430 9818
rect 13482 9766 13494 9818
rect 13546 9766 13558 9818
rect 13610 9766 13622 9818
rect 13674 9766 13686 9818
rect 13738 9766 19366 9818
rect 19418 9766 19430 9818
rect 19482 9766 19494 9818
rect 19546 9766 19558 9818
rect 19610 9766 19622 9818
rect 19674 9766 19686 9818
rect 19738 9766 23368 9818
rect 552 9744 23368 9766
rect 2501 9707 2559 9713
rect 2501 9673 2513 9707
rect 2547 9704 2559 9707
rect 2590 9704 2596 9716
rect 2547 9676 2596 9704
rect 2547 9673 2559 9676
rect 2501 9667 2559 9673
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 3234 9664 3240 9716
rect 3292 9664 3298 9716
rect 3421 9707 3479 9713
rect 3421 9673 3433 9707
rect 3467 9673 3479 9707
rect 5534 9704 5540 9716
rect 3421 9667 3479 9673
rect 5368 9676 5540 9704
rect 2777 9639 2835 9645
rect 2777 9636 2789 9639
rect 2332 9608 2789 9636
rect 2332 9512 2360 9608
rect 2777 9605 2789 9608
rect 2823 9636 2835 9639
rect 3436 9636 3464 9667
rect 2823 9608 3464 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 3878 9568 3884 9580
rect 2700 9540 3884 9568
rect 2314 9460 2320 9512
rect 2372 9460 2378 9512
rect 2406 9460 2412 9512
rect 2464 9500 2470 9512
rect 2700 9509 2728 9540
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5368 9568 5396 9676
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 11606 9704 11612 9716
rect 6972 9676 11612 9704
rect 6972 9664 6978 9676
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11974 9664 11980 9716
rect 12032 9704 12038 9716
rect 14734 9704 14740 9716
rect 12032 9676 14740 9704
rect 12032 9664 12038 9676
rect 14734 9664 14740 9676
rect 14792 9664 14798 9716
rect 14936 9676 15148 9704
rect 5442 9596 5448 9648
rect 5500 9596 5506 9648
rect 8205 9639 8263 9645
rect 8205 9605 8217 9639
rect 8251 9636 8263 9639
rect 13771 9639 13829 9645
rect 13771 9636 13783 9639
rect 8251 9608 8421 9636
rect 8251 9605 8263 9608
rect 8205 9599 8263 9605
rect 5215 9540 5396 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2464 9472 2697 9500
rect 2464 9460 2470 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 2869 9503 2927 9509
rect 2869 9469 2881 9503
rect 2915 9469 2927 9503
rect 2869 9463 2927 9469
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9500 3019 9503
rect 3142 9500 3148 9512
rect 3007 9472 3148 9500
rect 3007 9469 3019 9472
rect 2961 9463 3019 9469
rect 2884 9432 2912 9463
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3234 9460 3240 9512
rect 3292 9460 3298 9512
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 3252 9432 3280 9460
rect 2884 9404 3280 9432
rect 3436 9432 3464 9463
rect 3510 9460 3516 9512
rect 3568 9460 3574 9512
rect 4154 9500 4160 9512
rect 3620 9472 4160 9500
rect 3620 9432 3648 9472
rect 4154 9460 4160 9472
rect 4212 9500 4218 9512
rect 4706 9500 4712 9512
rect 4212 9472 4712 9500
rect 4212 9460 4218 9472
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 4982 9460 4988 9512
rect 5040 9460 5046 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 3436 9404 3648 9432
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 3878 9432 3884 9444
rect 3743 9404 3884 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 3878 9392 3884 9404
rect 3936 9392 3942 9444
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 3142 9364 3148 9376
rect 2280 9336 3148 9364
rect 2280 9324 2286 9336
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 5092 9364 5120 9463
rect 5258 9460 5264 9512
rect 5316 9460 5322 9512
rect 5828 9500 5856 9554
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 8393 9568 8421 9608
rect 12176 9608 13783 9636
rect 12176 9580 12204 9608
rect 13771 9605 13783 9608
rect 13817 9605 13829 9639
rect 13771 9599 13829 9605
rect 7340 9540 8248 9568
rect 8393 9540 8524 9568
rect 7340 9528 7346 9540
rect 5368 9472 5856 9500
rect 5368 9444 5396 9472
rect 5902 9460 5908 9512
rect 5960 9460 5966 9512
rect 6454 9460 6460 9512
rect 6512 9460 6518 9512
rect 8021 9503 8079 9509
rect 7932 9481 7990 9487
rect 5350 9392 5356 9444
rect 5408 9392 5414 9444
rect 5721 9435 5779 9441
rect 5721 9401 5733 9435
rect 5767 9432 5779 9435
rect 5920 9432 5948 9460
rect 7932 9447 7944 9481
rect 7978 9447 7990 9481
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8110 9500 8116 9512
rect 8067 9472 8116 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8220 9500 8248 9540
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 8220 9472 8401 9500
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8496 9500 8524 9540
rect 12158 9528 12164 9580
rect 12216 9528 12222 9580
rect 12434 9568 12440 9580
rect 12268 9540 12440 9568
rect 8645 9503 8703 9509
rect 8645 9500 8657 9503
rect 8496 9472 8657 9500
rect 8389 9463 8447 9469
rect 8645 9469 8657 9472
rect 8691 9469 8703 9503
rect 8645 9463 8703 9469
rect 8938 9460 8944 9512
rect 8996 9500 9002 9512
rect 9674 9500 9680 9512
rect 8996 9472 9680 9500
rect 8996 9460 9002 9472
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 10226 9460 10232 9512
rect 10284 9500 10290 9512
rect 12268 9509 12296 9540
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 12894 9568 12900 9580
rect 12575 9540 12900 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 12894 9528 12900 9540
rect 12952 9568 12958 9580
rect 13078 9568 13084 9580
rect 12952 9540 13084 9568
rect 12952 9528 12958 9540
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 13446 9568 13452 9580
rect 13228 9540 13452 9568
rect 13228 9528 13234 9540
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13998 9568 14004 9580
rect 13587 9540 14004 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 11057 9503 11115 9509
rect 10284 9472 10916 9500
rect 10284 9460 10290 9472
rect 7932 9444 7990 9447
rect 5767 9404 5948 9432
rect 5767 9401 5779 9404
rect 5721 9395 5779 9401
rect 5994 9392 6000 9444
rect 6052 9392 6058 9444
rect 6089 9435 6147 9441
rect 6089 9401 6101 9435
rect 6135 9432 6147 9435
rect 6546 9432 6552 9444
rect 6135 9404 6552 9432
rect 6135 9401 6147 9404
rect 6089 9395 6147 9401
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 7926 9392 7932 9444
rect 7984 9392 7990 9444
rect 8205 9435 8263 9441
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 8846 9432 8852 9444
rect 8251 9404 8852 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 10778 9432 10784 9444
rect 9692 9404 10784 9432
rect 5902 9364 5908 9376
rect 5092 9336 5908 9364
rect 5902 9324 5908 9336
rect 5960 9364 5966 9376
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 5960 9336 6837 9364
rect 5960 9324 5966 9336
rect 6825 9333 6837 9336
rect 6871 9333 6883 9367
rect 6825 9327 6883 9333
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 9692 9364 9720 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 10888 9432 10916 9472
rect 11057 9469 11069 9503
rect 11103 9500 11115 9503
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11103 9472 12265 9500
rect 11103 9469 11115 9472
rect 11057 9463 11115 9469
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 13722 9500 13728 9512
rect 12253 9463 12311 9469
rect 12406 9472 13728 9500
rect 12406 9432 12434 9472
rect 13722 9460 13728 9472
rect 13780 9460 13786 9512
rect 14936 9500 14964 9676
rect 15010 9596 15016 9648
rect 15068 9596 15074 9648
rect 15120 9636 15148 9676
rect 16758 9664 16764 9716
rect 16816 9664 16822 9716
rect 17034 9664 17040 9716
rect 17092 9704 17098 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 17092 9676 17417 9704
rect 17092 9664 17098 9676
rect 17405 9673 17417 9676
rect 17451 9673 17463 9707
rect 17405 9667 17463 9673
rect 17678 9664 17684 9716
rect 17736 9704 17742 9716
rect 18877 9707 18935 9713
rect 18877 9704 18889 9707
rect 17736 9676 18889 9704
rect 17736 9664 17742 9676
rect 18877 9673 18889 9676
rect 18923 9673 18935 9707
rect 18877 9667 18935 9673
rect 19061 9707 19119 9713
rect 19061 9673 19073 9707
rect 19107 9704 19119 9707
rect 19797 9707 19855 9713
rect 19107 9676 19748 9704
rect 19107 9673 19119 9676
rect 19061 9667 19119 9673
rect 15120 9608 15976 9636
rect 15028 9568 15056 9596
rect 15948 9580 15976 9608
rect 16592 9608 18276 9636
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 15028 9540 15301 9568
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 15657 9571 15715 9577
rect 15657 9537 15669 9571
rect 15703 9537 15715 9571
rect 15657 9531 15715 9537
rect 13832 9472 14964 9500
rect 15013 9503 15071 9509
rect 10888 9404 12434 9432
rect 13078 9392 13084 9444
rect 13136 9432 13142 9444
rect 13832 9432 13860 9472
rect 15013 9469 15025 9503
rect 15059 9469 15071 9503
rect 15013 9463 15071 9469
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9500 15439 9503
rect 15562 9500 15568 9512
rect 15427 9472 15568 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 13136 9404 13860 9432
rect 13136 9392 13142 9404
rect 14182 9392 14188 9444
rect 14240 9432 14246 9444
rect 15028 9432 15056 9463
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15672 9444 15700 9531
rect 15930 9528 15936 9580
rect 15988 9528 15994 9580
rect 16592 9509 16620 9608
rect 18248 9568 18276 9608
rect 18322 9596 18328 9648
rect 18380 9636 18386 9648
rect 19720 9636 19748 9676
rect 19797 9673 19809 9707
rect 19843 9704 19855 9707
rect 20622 9704 20628 9716
rect 19843 9676 20628 9704
rect 19843 9673 19855 9676
rect 19797 9667 19855 9673
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 21174 9664 21180 9716
rect 21232 9664 21238 9716
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 21729 9707 21787 9713
rect 21729 9704 21741 9707
rect 21416 9676 21741 9704
rect 21416 9664 21422 9676
rect 21729 9673 21741 9676
rect 21775 9673 21787 9707
rect 21729 9667 21787 9673
rect 22094 9664 22100 9716
rect 22152 9664 22158 9716
rect 22186 9664 22192 9716
rect 22244 9704 22250 9716
rect 22244 9676 22416 9704
rect 22244 9664 22250 9676
rect 19886 9636 19892 9648
rect 18380 9608 19564 9636
rect 19720 9608 19892 9636
rect 18380 9596 18386 9608
rect 18598 9568 18604 9580
rect 18248 9540 18604 9568
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 16577 9503 16635 9509
rect 16577 9469 16589 9503
rect 16623 9469 16635 9503
rect 16577 9463 16635 9469
rect 14240 9404 15056 9432
rect 14240 9392 14246 9404
rect 15654 9392 15660 9444
rect 15712 9392 15718 9444
rect 7055 9336 9720 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 9766 9324 9772 9376
rect 9824 9324 9830 9376
rect 10873 9367 10931 9373
rect 10873 9333 10885 9367
rect 10919 9364 10931 9367
rect 10962 9364 10968 9376
rect 10919 9336 10968 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 15838 9364 15844 9376
rect 11388 9336 15844 9364
rect 11388 9324 11394 9336
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 16408 9364 16436 9463
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 16761 9503 16819 9509
rect 16761 9500 16773 9503
rect 16724 9472 16773 9500
rect 16724 9460 16730 9472
rect 16761 9469 16773 9472
rect 16807 9469 16819 9503
rect 16761 9463 16819 9469
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9497 17187 9503
rect 17862 9500 17868 9512
rect 17236 9497 17868 9500
rect 17175 9472 17868 9497
rect 17175 9469 17264 9472
rect 17129 9463 17187 9469
rect 17862 9460 17868 9472
rect 17920 9500 17926 9512
rect 18248 9509 18276 9540
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 19150 9528 19156 9580
rect 19208 9528 19214 9580
rect 19536 9577 19564 9608
rect 19886 9596 19892 9608
rect 19944 9596 19950 9648
rect 19981 9639 20039 9645
rect 19981 9605 19993 9639
rect 20027 9636 20039 9639
rect 20530 9636 20536 9648
rect 20027 9608 20536 9636
rect 20027 9605 20039 9608
rect 19981 9599 20039 9605
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 22002 9636 22008 9648
rect 21284 9608 22008 9636
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 20070 9528 20076 9580
rect 20128 9528 20134 9580
rect 21284 9577 21312 9608
rect 22002 9596 22008 9608
rect 22060 9596 22066 9648
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9537 21327 9571
rect 22112 9568 22140 9664
rect 22388 9645 22416 9676
rect 22462 9664 22468 9716
rect 22520 9704 22526 9716
rect 22557 9707 22615 9713
rect 22557 9704 22569 9707
rect 22520 9676 22569 9704
rect 22520 9664 22526 9676
rect 22557 9673 22569 9676
rect 22603 9673 22615 9707
rect 22557 9667 22615 9673
rect 22373 9639 22431 9645
rect 22373 9605 22385 9639
rect 22419 9605 22431 9639
rect 22373 9599 22431 9605
rect 21269 9531 21327 9537
rect 21468 9540 22140 9568
rect 22281 9571 22339 9577
rect 18233 9503 18291 9509
rect 17920 9472 18000 9500
rect 17920 9460 17926 9472
rect 16850 9392 16856 9444
rect 16908 9432 16914 9444
rect 17972 9441 18000 9472
rect 18233 9469 18245 9503
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9469 19395 9503
rect 20088 9485 20116 9528
rect 20073 9479 20131 9485
rect 19886 9475 19892 9478
rect 19337 9463 19395 9469
rect 19843 9469 19892 9475
rect 19352 9448 19394 9463
rect 17957 9435 18015 9441
rect 16908 9404 17908 9432
rect 16908 9392 16914 9404
rect 16758 9364 16764 9376
rect 16408 9336 16764 9364
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 17589 9367 17647 9373
rect 17589 9364 17601 9367
rect 17276 9336 17601 9364
rect 17276 9324 17282 9336
rect 17589 9333 17601 9336
rect 17635 9333 17647 9367
rect 17589 9327 17647 9333
rect 17678 9324 17684 9376
rect 17736 9324 17742 9376
rect 17770 9324 17776 9376
rect 17828 9324 17834 9376
rect 17880 9364 17908 9404
rect 17957 9401 17969 9435
rect 18003 9401 18015 9435
rect 17957 9395 18015 9401
rect 18049 9435 18107 9441
rect 18049 9401 18061 9435
rect 18095 9401 18107 9435
rect 18049 9395 18107 9401
rect 18064 9364 18092 9395
rect 18690 9392 18696 9444
rect 18748 9392 18754 9444
rect 17880 9336 18092 9364
rect 18138 9324 18144 9376
rect 18196 9364 18202 9376
rect 18417 9367 18475 9373
rect 18417 9364 18429 9367
rect 18196 9336 18429 9364
rect 18196 9324 18202 9336
rect 18417 9333 18429 9336
rect 18463 9364 18475 9367
rect 18782 9364 18788 9376
rect 18463 9336 18788 9364
rect 18463 9333 18475 9336
rect 18417 9327 18475 9333
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 18874 9324 18880 9376
rect 18932 9373 18938 9376
rect 18932 9367 18951 9373
rect 18939 9333 18951 9367
rect 19366 9364 19394 9448
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 19613 9435 19671 9441
rect 19613 9432 19625 9435
rect 19576 9404 19625 9432
rect 19576 9392 19582 9404
rect 19613 9401 19625 9404
rect 19659 9401 19671 9435
rect 19843 9435 19855 9469
rect 19889 9435 19892 9469
rect 19843 9429 19892 9435
rect 19886 9426 19892 9429
rect 19944 9426 19950 9478
rect 20073 9445 20085 9479
rect 20119 9445 20131 9479
rect 20806 9460 20812 9512
rect 20864 9500 20870 9512
rect 20993 9503 21051 9509
rect 20993 9500 21005 9503
rect 20864 9472 21005 9500
rect 20864 9460 20870 9472
rect 20993 9469 21005 9472
rect 21039 9469 21051 9503
rect 20993 9463 21051 9469
rect 21082 9460 21088 9512
rect 21140 9460 21146 9512
rect 21468 9509 21496 9540
rect 22281 9537 22293 9571
rect 22327 9568 22339 9571
rect 22480 9568 22508 9664
rect 22327 9540 22508 9568
rect 22327 9537 22339 9540
rect 22281 9531 22339 9537
rect 21419 9503 21496 9509
rect 21419 9469 21431 9503
rect 21465 9472 21496 9503
rect 21545 9503 21603 9509
rect 21465 9469 21477 9472
rect 21419 9463 21477 9469
rect 21545 9469 21557 9503
rect 21591 9469 21603 9503
rect 21545 9463 21603 9469
rect 20073 9439 20131 9445
rect 19613 9395 19671 9401
rect 19978 9364 19984 9376
rect 19366 9336 19984 9364
rect 18932 9327 18951 9333
rect 18932 9324 18938 9327
rect 19978 9324 19984 9336
rect 20036 9364 20042 9376
rect 20257 9367 20315 9373
rect 20257 9364 20269 9367
rect 20036 9336 20269 9364
rect 20036 9324 20042 9336
rect 20257 9333 20269 9336
rect 20303 9333 20315 9367
rect 20257 9327 20315 9333
rect 20714 9324 20720 9376
rect 20772 9324 20778 9376
rect 21560 9364 21588 9463
rect 21634 9460 21640 9512
rect 21692 9500 21698 9512
rect 21821 9503 21879 9509
rect 21821 9500 21833 9503
rect 21692 9472 21833 9500
rect 21692 9460 21698 9472
rect 21821 9469 21833 9472
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 21913 9503 21971 9509
rect 21913 9469 21925 9503
rect 21959 9469 21971 9503
rect 21913 9463 21971 9469
rect 22005 9503 22063 9509
rect 22005 9469 22017 9503
rect 22051 9500 22063 9503
rect 22186 9500 22192 9512
rect 22051 9472 22192 9500
rect 22051 9469 22063 9472
rect 22005 9463 22063 9469
rect 21928 9432 21956 9463
rect 22186 9460 22192 9472
rect 22244 9500 22250 9512
rect 22830 9500 22836 9512
rect 22244 9472 22836 9500
rect 22244 9460 22250 9472
rect 22830 9460 22836 9472
rect 22888 9460 22894 9512
rect 22094 9432 22100 9444
rect 21928 9404 22100 9432
rect 22094 9392 22100 9404
rect 22152 9392 22158 9444
rect 22738 9392 22744 9444
rect 22796 9392 22802 9444
rect 21634 9364 21640 9376
rect 21560 9336 21640 9364
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 22002 9324 22008 9376
rect 22060 9364 22066 9376
rect 22531 9367 22589 9373
rect 22531 9364 22543 9367
rect 22060 9336 22543 9364
rect 22060 9324 22066 9336
rect 22531 9333 22543 9336
rect 22577 9333 22589 9367
rect 22531 9327 22589 9333
rect 552 9274 23368 9296
rect 552 9222 4366 9274
rect 4418 9222 4430 9274
rect 4482 9222 4494 9274
rect 4546 9222 4558 9274
rect 4610 9222 4622 9274
rect 4674 9222 4686 9274
rect 4738 9222 10366 9274
rect 10418 9222 10430 9274
rect 10482 9222 10494 9274
rect 10546 9222 10558 9274
rect 10610 9222 10622 9274
rect 10674 9222 10686 9274
rect 10738 9222 16366 9274
rect 16418 9222 16430 9274
rect 16482 9222 16494 9274
rect 16546 9222 16558 9274
rect 16610 9222 16622 9274
rect 16674 9222 16686 9274
rect 16738 9222 22366 9274
rect 22418 9222 22430 9274
rect 22482 9222 22494 9274
rect 22546 9222 22558 9274
rect 22610 9222 22622 9274
rect 22674 9222 22686 9274
rect 22738 9222 23368 9274
rect 552 9200 23368 9222
rect 2225 9163 2283 9169
rect 2225 9129 2237 9163
rect 2271 9129 2283 9163
rect 3510 9160 3516 9172
rect 2225 9123 2283 9129
rect 2746 9132 3516 9160
rect 2240 9092 2268 9123
rect 2746 9092 2774 9132
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9129 3939 9163
rect 3881 9123 3939 9129
rect 3602 9092 3608 9104
rect 2240 9064 2774 9092
rect 3068 9064 3608 9092
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 1964 8956 1992 8987
rect 2130 8984 2136 9036
rect 2188 8984 2194 9036
rect 2222 8984 2228 9036
rect 2280 8984 2286 9036
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 9024 2375 9027
rect 2406 9024 2412 9036
rect 2363 8996 2412 9024
rect 2363 8993 2375 8996
rect 2317 8987 2375 8993
rect 2332 8956 2360 8987
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 8993 2559 9027
rect 2501 8987 2559 8993
rect 1964 8928 2360 8956
rect 2516 8888 2544 8987
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 3068 9033 3096 9064
rect 3602 9052 3608 9064
rect 3660 9052 3666 9104
rect 2961 9027 3019 9033
rect 2961 9024 2973 9027
rect 2648 8996 2973 9024
rect 2648 8984 2654 8996
rect 2961 8993 2973 8996
rect 3007 8993 3019 9027
rect 2961 8987 3019 8993
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 8993 3111 9027
rect 3053 8987 3111 8993
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 3068 8956 3096 8987
rect 3234 8984 3240 9036
rect 3292 9024 3298 9036
rect 3513 9027 3571 9033
rect 3292 8996 3464 9024
rect 3292 8984 3298 8996
rect 2731 8928 3096 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 3326 8888 3332 8900
rect 2516 8860 3332 8888
rect 2700 8832 2728 8860
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 3436 8888 3464 8996
rect 3513 8993 3525 9027
rect 3559 9024 3571 9027
rect 3896 9024 3924 9123
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 5353 9163 5411 9169
rect 5353 9160 5365 9163
rect 5316 9132 5365 9160
rect 5316 9120 5322 9132
rect 5353 9129 5365 9132
rect 5399 9129 5411 9163
rect 8938 9160 8944 9172
rect 5353 9123 5411 9129
rect 5828 9132 8944 9160
rect 5828 9104 5856 9132
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9122 9120 9128 9172
rect 9180 9120 9186 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 9539 9132 10272 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 5810 9052 5816 9104
rect 5868 9052 5874 9104
rect 9416 9064 9628 9092
rect 9416 9036 9444 9064
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 3559 8996 3832 9024
rect 3896 8996 3985 9024
rect 3559 8993 3571 8996
rect 3513 8987 3571 8993
rect 3602 8916 3608 8968
rect 3660 8916 3666 8968
rect 3804 8956 3832 8996
rect 3973 8993 3985 8996
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 4062 8984 4068 9036
rect 4120 8984 4126 9036
rect 4982 8984 4988 9036
rect 5040 8984 5046 9036
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 5132 8996 5181 9024
rect 5132 8984 5138 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 6181 9027 6239 9033
rect 6181 9024 6193 9027
rect 5592 8996 6193 9024
rect 5592 8984 5598 8996
rect 6181 8993 6193 8996
rect 6227 9024 6239 9027
rect 6822 9024 6828 9036
rect 6227 8996 6828 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 8849 9027 8907 9033
rect 8849 9024 8861 9027
rect 8680 8996 8861 9024
rect 4246 8956 4252 8968
rect 3804 8928 4252 8956
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 6638 8956 6644 8968
rect 5316 8928 6644 8956
rect 5316 8916 5322 8928
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 4341 8891 4399 8897
rect 4341 8888 4353 8891
rect 3436 8860 4353 8888
rect 4341 8857 4353 8860
rect 4387 8857 4399 8891
rect 4341 8851 4399 8857
rect 5626 8848 5632 8900
rect 5684 8888 5690 8900
rect 6086 8888 6092 8900
rect 5684 8860 6092 8888
rect 5684 8848 5690 8860
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 8680 8888 8708 8996
rect 8849 8993 8861 8996
rect 8895 8993 8907 9027
rect 8849 8987 8907 8993
rect 9309 9027 9367 9033
rect 9309 8993 9321 9027
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 9324 8956 9352 8987
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 9600 9033 9628 9064
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 9732 9064 9904 9092
rect 9732 9052 9738 9064
rect 9876 9033 9904 9064
rect 9585 9027 9643 9033
rect 9585 8993 9597 9027
rect 9631 8993 9643 9027
rect 9585 8987 9643 8993
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 9324 8928 9689 8956
rect 9677 8925 9689 8928
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 9766 8888 9772 8900
rect 8680 8860 9772 8888
rect 8680 8832 8708 8860
rect 9766 8848 9772 8860
rect 9824 8888 9830 8900
rect 10060 8888 10088 8919
rect 10244 8900 10272 9132
rect 10318 9120 10324 9172
rect 10376 9120 10382 9172
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 13357 9163 13415 9169
rect 10836 9132 11928 9160
rect 10836 9120 10842 9132
rect 10336 9033 10364 9120
rect 11701 9095 11759 9101
rect 11701 9092 11713 9095
rect 11164 9064 11713 9092
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 10962 8984 10968 9036
rect 11020 8984 11026 9036
rect 11164 9033 11192 9064
rect 11701 9061 11713 9064
rect 11747 9061 11759 9095
rect 11701 9055 11759 9061
rect 11149 9027 11207 9033
rect 11149 8993 11161 9027
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 11238 8984 11244 9036
rect 11296 8984 11302 9036
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 9024 11391 9027
rect 11790 9024 11796 9036
rect 11379 8996 11796 9024
rect 11379 8993 11391 8996
rect 11333 8987 11391 8993
rect 11256 8956 11284 8984
rect 11606 8956 11612 8968
rect 11256 8928 11612 8956
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 9824 8860 10088 8888
rect 9824 8848 9830 8860
rect 10226 8848 10232 8900
rect 10284 8848 10290 8900
rect 11716 8888 11744 8996
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 11900 9033 11928 9132
rect 12268 9132 13308 9160
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 11348 8860 11744 8888
rect 11900 8888 11928 8987
rect 11974 8984 11980 9036
rect 12032 8984 12038 9036
rect 12268 9033 12296 9132
rect 12342 9052 12348 9104
rect 12400 9092 12406 9104
rect 12400 9064 12940 9092
rect 12400 9052 12406 9064
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 12492 8996 12541 9024
rect 12492 8984 12498 8996
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 9024 12679 9027
rect 12710 9024 12716 9036
rect 12667 8996 12716 9024
rect 12667 8993 12679 8996
rect 12621 8987 12679 8993
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 12802 8984 12808 9036
rect 12860 8984 12866 9036
rect 12912 9033 12940 9064
rect 12986 9052 12992 9104
rect 13044 9092 13050 9104
rect 13280 9092 13308 9132
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 13446 9160 13452 9172
rect 13403 9132 13452 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 15470 9160 15476 9172
rect 13780 9132 15476 9160
rect 13780 9120 13786 9132
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 15562 9120 15568 9172
rect 15620 9160 15626 9172
rect 15620 9132 16252 9160
rect 15620 9120 15626 9132
rect 16224 9101 16252 9132
rect 17770 9120 17776 9172
rect 17828 9120 17834 9172
rect 18049 9163 18107 9169
rect 18049 9129 18061 9163
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 16209 9095 16267 9101
rect 13044 9064 13216 9092
rect 13280 9064 15792 9092
rect 13044 9052 13050 9064
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 8993 12955 9027
rect 12897 8987 12955 8993
rect 13078 8984 13084 9036
rect 13136 8984 13142 9036
rect 13188 9033 13216 9064
rect 13173 9027 13231 9033
rect 13173 8993 13185 9027
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 13771 9027 13829 9033
rect 13771 8993 13783 9027
rect 13817 8993 13829 9027
rect 13906 9024 13912 9036
rect 13964 9033 13970 9036
rect 13873 8996 13912 9024
rect 13771 8987 13829 8993
rect 12066 8916 12072 8968
rect 12124 8956 12130 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12124 8928 13001 8956
rect 12124 8916 12130 8928
rect 12989 8925 13001 8928
rect 13035 8956 13047 8959
rect 13096 8956 13124 8984
rect 13035 8928 13124 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13786 8888 13814 8987
rect 13906 8984 13912 8996
rect 13964 8987 13973 9033
rect 14013 9029 14071 9035
rect 14013 8995 14025 9029
rect 14059 9026 14071 9029
rect 14185 9027 14243 9033
rect 14059 8998 14127 9026
rect 14059 8995 14071 8998
rect 14013 8989 14071 8995
rect 13964 8984 13970 8987
rect 13906 8888 13912 8900
rect 11900 8860 13676 8888
rect 13786 8860 13912 8888
rect 2682 8780 2688 8832
rect 2740 8780 2746 8832
rect 2774 8780 2780 8832
rect 2832 8780 2838 8832
rect 3142 8780 3148 8832
rect 3200 8780 3206 8832
rect 3697 8823 3755 8829
rect 3697 8789 3709 8823
rect 3743 8820 3755 8823
rect 3786 8820 3792 8832
rect 3743 8792 3792 8820
rect 3743 8789 3755 8792
rect 3697 8783 3755 8789
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 3973 8823 4031 8829
rect 3973 8820 3985 8823
rect 3936 8792 3985 8820
rect 3936 8780 3942 8792
rect 3973 8789 3985 8792
rect 4019 8789 4031 8823
rect 3973 8783 4031 8789
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5960 8792 6009 8820
rect 5960 8780 5966 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 5997 8783 6055 8789
rect 8662 8780 8668 8832
rect 8720 8780 8726 8832
rect 9033 8823 9091 8829
rect 9033 8789 9045 8823
rect 9079 8820 9091 8823
rect 9306 8820 9312 8832
rect 9079 8792 9312 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 9306 8780 9312 8792
rect 9364 8820 9370 8832
rect 11348 8820 11376 8860
rect 9364 8792 11376 8820
rect 9364 8780 9370 8792
rect 11422 8780 11428 8832
rect 11480 8820 11486 8832
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 11480 8792 11621 8820
rect 11480 8780 11486 8792
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11609 8783 11667 8789
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 12161 8823 12219 8829
rect 12161 8820 12173 8823
rect 11848 8792 12173 8820
rect 11848 8780 11854 8792
rect 12161 8789 12173 8792
rect 12207 8820 12219 8823
rect 12250 8820 12256 8832
rect 12207 8792 12256 8820
rect 12207 8789 12219 8792
rect 12161 8783 12219 8789
rect 12250 8780 12256 8792
rect 12308 8780 12314 8832
rect 12342 8780 12348 8832
rect 12400 8780 12406 8832
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 13449 8823 13507 8829
rect 13449 8820 13461 8823
rect 13228 8792 13461 8820
rect 13228 8780 13234 8792
rect 13449 8789 13461 8792
rect 13495 8789 13507 8823
rect 13648 8820 13676 8860
rect 13906 8848 13912 8860
rect 13964 8848 13970 8900
rect 14099 8888 14127 8998
rect 14185 8993 14197 9027
rect 14231 9026 14243 9027
rect 14274 9026 14280 9036
rect 14231 8998 14280 9026
rect 14231 8993 14243 8998
rect 14185 8987 14243 8993
rect 14274 8984 14280 8998
rect 14332 8984 14338 9036
rect 14476 9033 14504 9064
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 8993 14519 9027
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 14461 8987 14519 8993
rect 14660 8996 14749 9024
rect 14660 8968 14688 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 8993 14979 9027
rect 14921 8987 14979 8993
rect 14642 8916 14648 8968
rect 14700 8916 14706 8968
rect 14936 8956 14964 8987
rect 15286 8984 15292 9036
rect 15344 8984 15350 9036
rect 15010 8956 15016 8968
rect 14936 8928 15016 8956
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 14918 8888 14924 8900
rect 14016 8860 14924 8888
rect 14016 8820 14044 8860
rect 14918 8848 14924 8860
rect 14976 8848 14982 8900
rect 13648 8792 14044 8820
rect 14277 8823 14335 8829
rect 13449 8783 13507 8789
rect 14277 8789 14289 8823
rect 14323 8820 14335 8823
rect 14458 8820 14464 8832
rect 14323 8792 14464 8820
rect 14323 8789 14335 8792
rect 14277 8783 14335 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 14826 8780 14832 8832
rect 14884 8780 14890 8832
rect 15304 8820 15332 8984
rect 15764 8888 15792 9064
rect 16209 9061 16221 9095
rect 16255 9061 16267 9095
rect 16209 9055 16267 9061
rect 16758 9052 16764 9104
rect 16816 9092 16822 9104
rect 17586 9092 17592 9104
rect 16816 9064 17592 9092
rect 16816 9052 16822 9064
rect 17586 9052 17592 9064
rect 17644 9092 17650 9104
rect 17681 9095 17739 9101
rect 17681 9092 17693 9095
rect 17644 9064 17693 9092
rect 17644 9052 17650 9064
rect 17681 9061 17693 9064
rect 17727 9061 17739 9095
rect 17681 9055 17739 9061
rect 16776 9017 16804 9052
rect 17037 9027 17095 9033
rect 16761 9011 16819 9017
rect 16761 8977 16773 9011
rect 16807 8977 16819 9011
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 17788 9024 17816 9120
rect 17862 9052 17868 9104
rect 17920 9101 17926 9104
rect 17920 9095 17939 9101
rect 17927 9061 17939 9095
rect 18064 9092 18092 9123
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 20165 9163 20223 9169
rect 18840 9132 20116 9160
rect 18840 9120 18846 9132
rect 20088 9104 20116 9132
rect 20165 9129 20177 9163
rect 20211 9160 20223 9163
rect 20438 9160 20444 9172
rect 20211 9132 20444 9160
rect 20211 9129 20223 9132
rect 20165 9123 20223 9129
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 21726 9120 21732 9172
rect 21784 9160 21790 9172
rect 21821 9163 21879 9169
rect 21821 9160 21833 9163
rect 21784 9132 21833 9160
rect 21784 9120 21790 9132
rect 21821 9129 21833 9132
rect 21867 9129 21879 9163
rect 21821 9123 21879 9129
rect 22186 9120 22192 9172
rect 22244 9120 22250 9172
rect 18874 9092 18880 9104
rect 18064 9064 18880 9092
rect 17920 9055 17939 9061
rect 17920 9052 17926 9055
rect 18874 9052 18880 9064
rect 18932 9092 18938 9104
rect 18932 9064 19288 9092
rect 18932 9052 18938 9064
rect 17083 8996 17816 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 18322 8984 18328 9036
rect 18380 8984 18386 9036
rect 18506 8984 18512 9036
rect 18564 9024 18570 9036
rect 18785 9027 18843 9033
rect 18785 9024 18797 9027
rect 18564 8996 18797 9024
rect 18564 8984 18570 8996
rect 18785 8993 18797 8996
rect 18831 9024 18843 9027
rect 19150 9024 19156 9036
rect 18831 8996 19156 9024
rect 18831 8993 18843 8996
rect 18785 8987 18843 8993
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 19260 9033 19288 9064
rect 20070 9052 20076 9104
rect 20128 9052 20134 9104
rect 21450 9052 21456 9104
rect 21508 9092 21514 9104
rect 21508 9064 21680 9092
rect 21508 9052 21514 9064
rect 19245 9027 19303 9033
rect 19245 8993 19257 9027
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19392 8996 19625 9024
rect 19392 8984 19398 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 19794 8984 19800 9036
rect 19852 8984 19858 9036
rect 19889 9027 19947 9033
rect 19889 8993 19901 9027
rect 19935 9024 19947 9027
rect 19978 9024 19984 9036
rect 19935 8996 19984 9024
rect 19935 8993 19947 8996
rect 19889 8987 19947 8993
rect 19978 8984 19984 8996
rect 20036 9024 20042 9036
rect 20349 9027 20407 9033
rect 20349 9024 20361 9027
rect 20036 8996 20361 9024
rect 20036 8984 20042 8996
rect 20349 8993 20361 8996
rect 20395 8993 20407 9027
rect 20349 8987 20407 8993
rect 20990 8984 20996 9036
rect 21048 9024 21054 9036
rect 21652 9033 21680 9064
rect 21348 9027 21406 9033
rect 21348 9024 21360 9027
rect 21048 8996 21360 9024
rect 21048 8984 21054 8996
rect 21348 8993 21360 8996
rect 21394 9024 21406 9027
rect 21637 9027 21695 9033
rect 21394 8996 21462 9024
rect 21394 8993 21406 8996
rect 21348 8987 21406 8993
rect 16761 8971 16819 8977
rect 17218 8956 17224 8968
rect 16960 8928 17224 8956
rect 16960 8897 16988 8928
rect 17218 8916 17224 8928
rect 17276 8956 17282 8968
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 17276 8928 17325 8956
rect 17276 8916 17282 8928
rect 17313 8925 17325 8928
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 16945 8891 17003 8897
rect 16945 8888 16957 8891
rect 15764 8860 16957 8888
rect 16945 8857 16957 8860
rect 16991 8857 17003 8891
rect 18138 8888 18144 8900
rect 16945 8851 17003 8857
rect 17420 8860 18144 8888
rect 15746 8820 15752 8832
rect 15304 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 15988 8792 16313 8820
rect 15988 8780 15994 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 16301 8783 16359 8789
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17420 8829 17448 8860
rect 18138 8848 18144 8860
rect 18196 8848 18202 8900
rect 18524 8897 18552 8984
rect 19702 8956 19708 8968
rect 19306 8928 19708 8956
rect 18509 8891 18567 8897
rect 18509 8857 18521 8891
rect 18555 8857 18567 8891
rect 18509 8851 18567 8857
rect 18782 8848 18788 8900
rect 18840 8888 18846 8900
rect 18969 8891 19027 8897
rect 18969 8888 18981 8891
rect 18840 8860 18981 8888
rect 18840 8848 18846 8860
rect 18969 8857 18981 8860
rect 19015 8857 19027 8891
rect 18969 8851 19027 8857
rect 19058 8848 19064 8900
rect 19116 8848 19122 8900
rect 19306 8888 19334 8928
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 20162 8956 20168 8968
rect 19996 8928 20168 8956
rect 19996 8897 20024 8928
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 20898 8916 20904 8968
rect 20956 8956 20962 8968
rect 21434 8956 21462 8996
rect 21637 8993 21649 9027
rect 21683 8993 21695 9027
rect 21637 8987 21695 8993
rect 22097 9027 22155 9033
rect 22097 8993 22109 9027
rect 22143 9024 22155 9027
rect 22204 9024 22232 9120
rect 22143 8996 22232 9024
rect 22143 8993 22155 8996
rect 22097 8987 22155 8993
rect 20956 8928 21404 8956
rect 21434 8928 21956 8956
rect 20956 8916 20962 8928
rect 19981 8891 20039 8897
rect 19981 8888 19993 8891
rect 19168 8860 19334 8888
rect 19720 8860 19993 8888
rect 17405 8823 17463 8829
rect 17405 8820 17417 8823
rect 16724 8792 17417 8820
rect 16724 8780 16730 8792
rect 17405 8789 17417 8792
rect 17451 8789 17463 8823
rect 17405 8783 17463 8789
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 17678 8820 17684 8832
rect 17635 8792 17684 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 17678 8780 17684 8792
rect 17736 8780 17742 8832
rect 17770 8780 17776 8832
rect 17828 8820 17834 8832
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 17828 8792 17877 8820
rect 17828 8780 17834 8792
rect 17865 8789 17877 8792
rect 17911 8820 17923 8823
rect 19168 8820 19196 8860
rect 17911 8792 19196 8820
rect 17911 8789 17923 8792
rect 17865 8783 17923 8789
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 19720 8820 19748 8860
rect 19981 8857 19993 8860
rect 20027 8857 20039 8891
rect 21376 8888 21404 8928
rect 21928 8897 21956 8928
rect 21453 8891 21511 8897
rect 21453 8888 21465 8891
rect 21376 8860 21465 8888
rect 19981 8851 20039 8857
rect 21453 8857 21465 8860
rect 21499 8857 21511 8891
rect 21453 8851 21511 8857
rect 21545 8891 21603 8897
rect 21545 8857 21557 8891
rect 21591 8857 21603 8891
rect 21545 8851 21603 8857
rect 21913 8891 21971 8897
rect 21913 8857 21925 8891
rect 21959 8857 21971 8891
rect 21913 8851 21971 8857
rect 19392 8792 19748 8820
rect 19797 8823 19855 8829
rect 19392 8780 19398 8792
rect 19797 8789 19809 8823
rect 19843 8820 19855 8823
rect 19886 8820 19892 8832
rect 19843 8792 19892 8820
rect 19843 8789 19855 8792
rect 19797 8783 19855 8789
rect 19886 8780 19892 8792
rect 19944 8780 19950 8832
rect 20254 8780 20260 8832
rect 20312 8820 20318 8832
rect 20990 8820 20996 8832
rect 20312 8792 20996 8820
rect 20312 8780 20318 8792
rect 20990 8780 20996 8792
rect 21048 8820 21054 8832
rect 21560 8820 21588 8851
rect 21048 8792 21588 8820
rect 21048 8780 21054 8792
rect 552 8730 23368 8752
rect 552 8678 1366 8730
rect 1418 8678 1430 8730
rect 1482 8678 1494 8730
rect 1546 8678 1558 8730
rect 1610 8678 1622 8730
rect 1674 8678 1686 8730
rect 1738 8678 7366 8730
rect 7418 8678 7430 8730
rect 7482 8678 7494 8730
rect 7546 8678 7558 8730
rect 7610 8678 7622 8730
rect 7674 8678 7686 8730
rect 7738 8678 13366 8730
rect 13418 8678 13430 8730
rect 13482 8678 13494 8730
rect 13546 8678 13558 8730
rect 13610 8678 13622 8730
rect 13674 8678 13686 8730
rect 13738 8678 19366 8730
rect 19418 8678 19430 8730
rect 19482 8678 19494 8730
rect 19546 8678 19558 8730
rect 19610 8678 19622 8730
rect 19674 8678 19686 8730
rect 19738 8678 23368 8730
rect 552 8656 23368 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2372 8588 2535 8616
rect 2372 8576 2378 8588
rect 2409 8551 2467 8557
rect 2409 8517 2421 8551
rect 2455 8517 2467 8551
rect 2507 8548 2535 8588
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2648 8588 2697 8616
rect 2648 8576 2654 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 3050 8576 3056 8628
rect 3108 8616 3114 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3108 8588 3249 8616
rect 3108 8576 3114 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3694 8616 3700 8628
rect 3476 8588 3700 8616
rect 3476 8576 3482 8588
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 11425 8619 11483 8625
rect 11425 8616 11437 8619
rect 10928 8588 11437 8616
rect 10928 8576 10934 8588
rect 11425 8585 11437 8588
rect 11471 8616 11483 8619
rect 11790 8616 11796 8628
rect 11471 8588 11796 8616
rect 11471 8585 11483 8588
rect 11425 8579 11483 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12894 8616 12900 8628
rect 12308 8588 12900 8616
rect 12308 8576 12314 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13265 8619 13323 8625
rect 13265 8585 13277 8619
rect 13311 8616 13323 8619
rect 15010 8616 15016 8628
rect 13311 8588 15016 8616
rect 13311 8585 13323 8588
rect 13265 8579 13323 8585
rect 15010 8576 15016 8588
rect 15068 8616 15074 8628
rect 15068 8588 15332 8616
rect 15068 8576 15074 8588
rect 2869 8551 2927 8557
rect 2869 8548 2881 8551
rect 2507 8520 2881 8548
rect 2409 8511 2467 8517
rect 2869 8517 2881 8520
rect 2915 8517 2927 8551
rect 7193 8551 7251 8557
rect 2869 8511 2927 8517
rect 3160 8520 5580 8548
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8381 2283 8415
rect 2424 8412 2452 8511
rect 2501 8415 2559 8421
rect 2501 8412 2513 8415
rect 2424 8384 2513 8412
rect 2225 8375 2283 8381
rect 2501 8381 2513 8384
rect 2547 8412 2559 8415
rect 3053 8415 3111 8421
rect 3053 8412 3065 8415
rect 2547 8384 3065 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 3053 8381 3065 8384
rect 3099 8412 3111 8415
rect 3160 8412 3188 8520
rect 5552 8492 5580 8520
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 9950 8548 9956 8560
rect 7239 8520 9956 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 11054 8508 11060 8560
rect 11112 8508 11118 8560
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 14642 8548 14648 8560
rect 11572 8520 14648 8548
rect 11572 8508 11578 8520
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 4338 8480 4344 8492
rect 3292 8452 4344 8480
rect 3292 8440 3298 8452
rect 3099 8384 3188 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 2240 8288 2268 8375
rect 3326 8372 3332 8424
rect 3384 8412 3390 8424
rect 3528 8421 3556 8452
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5684 8452 5750 8480
rect 5684 8440 5690 8452
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 9674 8480 9680 8492
rect 9646 8440 9680 8480
rect 9732 8440 9738 8492
rect 9128 8424 9180 8430
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3384 8384 3433 8412
rect 3384 8372 3390 8384
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 3513 8415 3571 8421
rect 3513 8381 3525 8415
rect 3559 8381 3571 8415
rect 4709 8415 4767 8421
rect 4709 8412 4721 8415
rect 3513 8375 3571 8381
rect 4264 8384 4721 8412
rect 2682 8304 2688 8356
rect 2740 8344 2746 8356
rect 2777 8347 2835 8353
rect 2777 8344 2789 8347
rect 2740 8316 2789 8344
rect 2740 8304 2746 8316
rect 2777 8313 2789 8316
rect 2823 8313 2835 8347
rect 2777 8307 2835 8313
rect 2961 8347 3019 8353
rect 2961 8313 2973 8347
rect 3007 8344 3019 8347
rect 3237 8347 3295 8353
rect 3007 8316 3188 8344
rect 3007 8313 3019 8316
rect 2961 8307 3019 8313
rect 2222 8236 2228 8288
rect 2280 8236 2286 8288
rect 3160 8276 3188 8316
rect 3237 8313 3249 8347
rect 3283 8344 3295 8347
rect 4154 8344 4160 8356
rect 3283 8316 4160 8344
rect 3283 8313 3295 8316
rect 3237 8307 3295 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 3326 8276 3332 8288
rect 3160 8248 3332 8276
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 3697 8279 3755 8285
rect 3697 8245 3709 8279
rect 3743 8276 3755 8279
rect 3786 8276 3792 8288
rect 3743 8248 3792 8276
rect 3743 8245 3755 8248
rect 3697 8239 3755 8245
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4264 8276 4292 8384
rect 4709 8381 4721 8384
rect 4755 8412 4767 8415
rect 5074 8412 5080 8424
rect 4755 8384 5080 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 5166 8372 5172 8424
rect 5224 8412 5230 8424
rect 6181 8415 6239 8421
rect 6181 8412 6193 8415
rect 5224 8384 6193 8412
rect 5224 8372 5230 8384
rect 6181 8381 6193 8384
rect 6227 8381 6239 8415
rect 6181 8375 6239 8381
rect 6270 8372 6276 8424
rect 6328 8412 6334 8424
rect 6730 8412 6736 8424
rect 6328 8384 6736 8412
rect 6328 8372 6334 8384
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 9646 8412 9674 8440
rect 9180 8384 9674 8412
rect 9968 8412 9996 8508
rect 11072 8480 11100 8508
rect 11974 8480 11980 8492
rect 11072 8452 11980 8480
rect 11256 8421 11284 8452
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 9968 8384 11161 8412
rect 11149 8381 11161 8384
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8381 11299 8415
rect 11241 8375 11299 8381
rect 9128 8366 9180 8372
rect 5902 8304 5908 8356
rect 5960 8304 5966 8356
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 6512 8316 6653 8344
rect 6512 8304 6518 8316
rect 6641 8313 6653 8316
rect 6687 8313 6699 8347
rect 6641 8307 6699 8313
rect 9217 8347 9275 8353
rect 9217 8313 9229 8347
rect 9263 8344 9275 8347
rect 9306 8344 9312 8356
rect 9263 8316 9312 8344
rect 9263 8313 9275 8316
rect 9217 8307 9275 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 11054 8344 11060 8356
rect 11011 8316 11060 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 11164 8344 11192 8375
rect 11330 8372 11336 8424
rect 11388 8412 11394 8424
rect 11514 8412 11520 8424
rect 11388 8384 11520 8412
rect 11388 8372 11394 8384
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 11624 8344 11652 8375
rect 11164 8316 11652 8344
rect 11716 8344 11744 8375
rect 11882 8372 11888 8424
rect 11940 8372 11946 8424
rect 12360 8421 12388 8520
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 14826 8508 14832 8560
rect 14884 8508 14890 8560
rect 14918 8508 14924 8560
rect 14976 8548 14982 8560
rect 15304 8548 15332 8588
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 16301 8619 16359 8625
rect 16301 8616 16313 8619
rect 15896 8588 16313 8616
rect 15896 8576 15902 8588
rect 16301 8585 16313 8588
rect 16347 8585 16359 8619
rect 16301 8579 16359 8585
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 16853 8619 16911 8625
rect 16853 8616 16865 8619
rect 16816 8588 16865 8616
rect 16816 8576 16822 8588
rect 16853 8585 16865 8588
rect 16899 8585 16911 8619
rect 16853 8579 16911 8585
rect 17218 8576 17224 8628
rect 17276 8576 17282 8628
rect 17310 8576 17316 8628
rect 17368 8576 17374 8628
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 18874 8616 18880 8628
rect 18472 8588 18880 8616
rect 18472 8576 18478 8588
rect 18874 8576 18880 8588
rect 18932 8616 18938 8628
rect 19058 8616 19064 8628
rect 18932 8588 19064 8616
rect 18932 8576 18938 8588
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19242 8576 19248 8628
rect 19300 8576 19306 8628
rect 19794 8576 19800 8628
rect 19852 8616 19858 8628
rect 19889 8619 19947 8625
rect 19889 8616 19901 8619
rect 19852 8588 19901 8616
rect 19852 8576 19858 8588
rect 19889 8585 19901 8588
rect 19935 8585 19947 8619
rect 19889 8579 19947 8585
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20349 8619 20407 8625
rect 20349 8616 20361 8619
rect 20128 8588 20361 8616
rect 20128 8576 20134 8588
rect 20349 8585 20361 8588
rect 20395 8616 20407 8619
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 20395 8588 20637 8616
rect 20395 8585 20407 8588
rect 20349 8579 20407 8585
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 20625 8579 20683 8585
rect 20714 8576 20720 8628
rect 20772 8576 20778 8628
rect 21358 8576 21364 8628
rect 21416 8576 21422 8628
rect 21637 8619 21695 8625
rect 21637 8585 21649 8619
rect 21683 8616 21695 8619
rect 22002 8616 22008 8628
rect 21683 8588 22008 8616
rect 21683 8585 21695 8588
rect 21637 8579 21695 8585
rect 22002 8576 22008 8588
rect 22060 8576 22066 8628
rect 15933 8551 15991 8557
rect 15933 8548 15945 8551
rect 14976 8520 15240 8548
rect 15304 8520 15945 8548
rect 14976 8508 14982 8520
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 13170 8480 13176 8492
rect 13096 8452 13176 8480
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12544 8412 12572 8440
rect 13096 8421 13124 8452
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 14090 8480 14096 8492
rect 13412 8452 14096 8480
rect 13412 8440 13418 8452
rect 14090 8440 14096 8452
rect 14148 8480 14154 8492
rect 14458 8480 14464 8492
rect 14148 8452 14464 8480
rect 14148 8440 14154 8452
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14844 8480 14872 8508
rect 15212 8489 15240 8520
rect 15933 8517 15945 8520
rect 15979 8517 15991 8551
rect 17236 8548 17264 8576
rect 17604 8548 17632 8576
rect 15933 8511 15991 8517
rect 16500 8520 17264 8548
rect 17512 8520 17632 8548
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14844 8452 15117 8480
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8449 15255 8483
rect 15197 8443 15255 8449
rect 15378 8440 15384 8492
rect 15436 8480 15442 8492
rect 15436 8452 16252 8480
rect 15436 8440 15442 8452
rect 13081 8415 13139 8421
rect 12544 8384 13032 8412
rect 12544 8344 12572 8384
rect 11716 8316 12572 8344
rect 12894 8304 12900 8356
rect 12952 8304 12958 8356
rect 13004 8344 13032 8384
rect 13081 8381 13093 8415
rect 13127 8381 13139 8415
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 13081 8375 13139 8381
rect 13648 8384 14841 8412
rect 13648 8344 13676 8384
rect 14829 8381 14841 8384
rect 14875 8412 14887 8415
rect 15289 8415 15347 8421
rect 15289 8412 15301 8415
rect 14875 8384 15301 8412
rect 14875 8381 14887 8384
rect 14829 8375 14887 8381
rect 15289 8381 15301 8384
rect 15335 8381 15347 8415
rect 15289 8375 15347 8381
rect 15470 8372 15476 8424
rect 15528 8372 15534 8424
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8412 15807 8415
rect 16022 8412 16028 8424
rect 15795 8384 16028 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 16224 8421 16252 8452
rect 16500 8421 16528 8520
rect 16850 8480 16856 8492
rect 16592 8452 16856 8480
rect 16592 8424 16620 8452
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 17512 8480 17540 8520
rect 19061 8483 19119 8489
rect 17144 8452 17540 8480
rect 17604 8452 19012 8480
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8381 16267 8415
rect 16209 8375 16267 8381
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8381 16543 8415
rect 16485 8375 16543 8381
rect 13004 8316 13676 8344
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 13998 8344 14004 8356
rect 13780 8316 14004 8344
rect 13780 8304 13786 8316
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 14458 8304 14464 8356
rect 14516 8344 14522 8356
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 14516 8316 15669 8344
rect 14516 8304 14522 8316
rect 15657 8313 15669 8316
rect 15703 8313 15715 8347
rect 15657 8307 15715 8313
rect 4120 8248 4292 8276
rect 4120 8236 4126 8248
rect 4338 8236 4344 8288
rect 4396 8276 4402 8288
rect 4893 8279 4951 8285
rect 4893 8276 4905 8279
rect 4396 8248 4905 8276
rect 4396 8236 4402 8248
rect 4893 8245 4905 8248
rect 4939 8245 4951 8279
rect 4893 8239 4951 8245
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 7006 8276 7012 8288
rect 6052 8248 7012 8276
rect 6052 8236 6058 8248
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 11756 8248 12081 8276
rect 11756 8236 11762 8248
rect 12069 8245 12081 8248
rect 12115 8245 12127 8279
rect 12069 8239 12127 8245
rect 12161 8279 12219 8285
rect 12161 8245 12173 8279
rect 12207 8276 12219 8279
rect 12526 8276 12532 8288
rect 12207 8248 12532 8276
rect 12207 8245 12219 8248
rect 12161 8239 12219 8245
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 13078 8276 13084 8288
rect 12860 8248 13084 8276
rect 12860 8236 12866 8248
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 14182 8276 14188 8288
rect 13228 8248 14188 8276
rect 13228 8236 13234 8248
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 16025 8279 16083 8285
rect 16025 8276 16037 8279
rect 15344 8248 16037 8276
rect 15344 8236 15350 8248
rect 16025 8245 16037 8248
rect 16071 8245 16083 8279
rect 16500 8276 16528 8375
rect 16574 8372 16580 8424
rect 16632 8372 16638 8424
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 17144 8421 17172 8452
rect 17037 8415 17095 8421
rect 17037 8412 17049 8415
rect 16724 8384 16896 8412
rect 16724 8372 16730 8384
rect 16868 8353 16896 8384
rect 16960 8384 17049 8412
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8313 16911 8347
rect 16853 8307 16911 8313
rect 16761 8279 16819 8285
rect 16761 8276 16773 8279
rect 16500 8248 16773 8276
rect 16025 8239 16083 8245
rect 16761 8245 16773 8248
rect 16807 8245 16819 8279
rect 16960 8276 16988 8384
rect 17037 8381 17049 8384
rect 17083 8381 17095 8415
rect 17037 8375 17095 8381
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 17310 8372 17316 8424
rect 17368 8412 17374 8424
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 17368 8384 17417 8412
rect 17368 8372 17374 8384
rect 17405 8381 17417 8384
rect 17451 8412 17463 8415
rect 17604 8412 17632 8452
rect 17451 8384 17632 8412
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 17678 8372 17684 8424
rect 17736 8372 17742 8424
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 18877 8415 18935 8421
rect 18877 8412 18889 8415
rect 17920 8384 18889 8412
rect 17920 8372 17926 8384
rect 18877 8381 18889 8384
rect 18923 8381 18935 8415
rect 18984 8412 19012 8452
rect 19061 8449 19073 8483
rect 19107 8480 19119 8483
rect 19260 8480 19288 8576
rect 19978 8548 19984 8560
rect 19107 8452 19288 8480
rect 19444 8520 19984 8548
rect 19107 8449 19119 8452
rect 19061 8443 19119 8449
rect 19334 8412 19340 8424
rect 18984 8384 19340 8412
rect 18877 8375 18935 8381
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 19444 8421 19472 8520
rect 19978 8508 19984 8520
rect 20036 8508 20042 8560
rect 20441 8551 20499 8557
rect 20441 8548 20453 8551
rect 20088 8520 20453 8548
rect 20088 8480 20116 8520
rect 20441 8517 20453 8520
rect 20487 8517 20499 8551
rect 20732 8548 20760 8576
rect 20441 8511 20499 8517
rect 20548 8520 20852 8548
rect 19628 8452 20116 8480
rect 20257 8483 20315 8489
rect 19628 8421 19656 8452
rect 20257 8449 20269 8483
rect 20303 8480 20315 8483
rect 20548 8480 20576 8520
rect 20824 8489 20852 8520
rect 21450 8508 21456 8560
rect 21508 8548 21514 8560
rect 22741 8551 22799 8557
rect 22741 8548 22753 8551
rect 21508 8520 22753 8548
rect 21508 8508 21514 8520
rect 22741 8517 22753 8520
rect 22787 8517 22799 8551
rect 22741 8511 22799 8517
rect 20303 8452 20576 8480
rect 20809 8483 20867 8489
rect 20303 8449 20315 8452
rect 20257 8443 20315 8449
rect 20809 8449 20821 8483
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 21266 8440 21272 8492
rect 21324 8440 21330 8492
rect 21634 8440 21640 8492
rect 21692 8480 21698 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21692 8452 22017 8480
rect 21692 8440 21698 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22922 8480 22928 8492
rect 22005 8443 22063 8449
rect 22664 8452 22928 8480
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8381 19487 8415
rect 19429 8375 19487 8381
rect 19613 8415 19671 8421
rect 19613 8381 19625 8415
rect 19659 8381 19671 8415
rect 19613 8375 19671 8381
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8412 20131 8415
rect 20530 8412 20536 8424
rect 20119 8384 20536 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 20530 8372 20536 8384
rect 20588 8412 20594 8424
rect 20625 8415 20683 8421
rect 20625 8412 20637 8415
rect 20588 8384 20637 8412
rect 20588 8372 20594 8384
rect 20625 8381 20637 8384
rect 20671 8381 20683 8415
rect 20625 8375 20683 8381
rect 20901 8415 20959 8421
rect 20901 8381 20913 8415
rect 20947 8412 20959 8415
rect 20947 8384 21312 8412
rect 20947 8381 20959 8384
rect 20901 8375 20959 8381
rect 17696 8344 17724 8372
rect 21284 8356 21312 8384
rect 21358 8372 21364 8424
rect 21416 8412 21422 8424
rect 22664 8421 22692 8452
rect 22922 8440 22928 8452
rect 22980 8440 22986 8492
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 21416 8384 21465 8412
rect 21416 8372 21422 8384
rect 21453 8381 21465 8384
rect 21499 8412 21511 8415
rect 21729 8415 21787 8421
rect 21729 8412 21741 8415
rect 21499 8384 21741 8412
rect 21499 8381 21511 8384
rect 21453 8375 21511 8381
rect 21729 8381 21741 8384
rect 21775 8381 21787 8415
rect 21729 8375 21787 8381
rect 22649 8415 22707 8421
rect 22649 8381 22661 8415
rect 22695 8381 22707 8415
rect 22649 8375 22707 8381
rect 22833 8415 22891 8421
rect 22833 8381 22845 8415
rect 22879 8381 22891 8415
rect 22833 8375 22891 8381
rect 19978 8344 19984 8356
rect 17696 8316 19984 8344
rect 19978 8304 19984 8316
rect 20036 8304 20042 8356
rect 20254 8304 20260 8356
rect 20312 8344 20318 8356
rect 20349 8347 20407 8353
rect 20349 8344 20361 8347
rect 20312 8316 20361 8344
rect 20312 8304 20318 8316
rect 20349 8313 20361 8316
rect 20395 8313 20407 8347
rect 20349 8307 20407 8313
rect 21174 8304 21180 8356
rect 21232 8304 21238 8356
rect 21266 8304 21272 8356
rect 21324 8304 21330 8356
rect 21744 8344 21772 8375
rect 22848 8344 22876 8375
rect 21744 8316 22876 8344
rect 17586 8276 17592 8288
rect 16960 8248 17592 8276
rect 16761 8239 16819 8245
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 18690 8236 18696 8288
rect 18748 8236 18754 8288
rect 19521 8279 19579 8285
rect 19521 8245 19533 8279
rect 19567 8276 19579 8279
rect 19794 8276 19800 8288
rect 19567 8248 19800 8276
rect 19567 8245 19579 8248
rect 19521 8239 19579 8245
rect 19794 8236 19800 8248
rect 19852 8236 19858 8288
rect 552 8186 23368 8208
rect 552 8134 4366 8186
rect 4418 8134 4430 8186
rect 4482 8134 4494 8186
rect 4546 8134 4558 8186
rect 4610 8134 4622 8186
rect 4674 8134 4686 8186
rect 4738 8134 10366 8186
rect 10418 8134 10430 8186
rect 10482 8134 10494 8186
rect 10546 8134 10558 8186
rect 10610 8134 10622 8186
rect 10674 8134 10686 8186
rect 10738 8134 16366 8186
rect 16418 8134 16430 8186
rect 16482 8134 16494 8186
rect 16546 8134 16558 8186
rect 16610 8134 16622 8186
rect 16674 8134 16686 8186
rect 16738 8134 22366 8186
rect 22418 8134 22430 8186
rect 22482 8134 22494 8186
rect 22546 8134 22558 8186
rect 22610 8134 22622 8186
rect 22674 8134 22686 8186
rect 22738 8134 23368 8186
rect 552 8112 23368 8134
rect 2222 8032 2228 8084
rect 2280 8072 2286 8084
rect 2280 8044 3280 8072
rect 2280 8032 2286 8044
rect 1118 7945 1124 7948
rect 1112 7899 1124 7945
rect 1118 7896 1124 7899
rect 1176 7896 1182 7948
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 3252 7945 3280 8044
rect 3418 8032 3424 8084
rect 3476 8032 3482 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 3568 8044 3893 8072
rect 3568 8032 3574 8044
rect 3881 8041 3893 8044
rect 3927 8072 3939 8075
rect 4062 8072 4068 8084
rect 3927 8044 4068 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4982 8032 4988 8084
rect 5040 8032 5046 8084
rect 5074 8032 5080 8084
rect 5132 8032 5138 8084
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 5994 8072 6000 8084
rect 5224 8044 6000 8072
rect 5224 8032 5230 8044
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 6144 8044 7113 8072
rect 6144 8032 6150 8044
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 7101 8035 7159 8041
rect 11149 8075 11207 8081
rect 11149 8041 11161 8075
rect 11195 8072 11207 8075
rect 11882 8072 11888 8084
rect 11195 8044 11888 8072
rect 11195 8041 11207 8044
rect 11149 8035 11207 8041
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 13722 8072 13728 8084
rect 12492 8044 13728 8072
rect 12492 8032 12498 8044
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 13872 8044 14412 8072
rect 13872 8032 13878 8044
rect 3326 7964 3332 8016
rect 3384 8004 3390 8016
rect 5000 8004 5028 8032
rect 3384 7976 5028 8004
rect 3384 7964 3390 7976
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 2740 7908 2789 7936
rect 2740 7896 2746 7908
rect 2777 7905 2789 7908
rect 2823 7936 2835 7939
rect 3237 7939 3295 7945
rect 2823 7908 3188 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 842 7828 848 7880
rect 900 7828 906 7880
rect 3050 7828 3056 7880
rect 3108 7828 3114 7880
rect 3160 7868 3188 7908
rect 3237 7905 3249 7939
rect 3283 7936 3295 7939
rect 3510 7936 3516 7948
rect 3283 7908 3516 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 5000 7945 5028 7976
rect 3697 7939 3755 7945
rect 3697 7905 3709 7939
rect 3743 7936 3755 7939
rect 4065 7939 4123 7945
rect 3743 7908 4016 7936
rect 3743 7905 3755 7908
rect 3697 7899 3755 7905
rect 3160 7840 3740 7868
rect 3142 7760 3148 7812
rect 3200 7800 3206 7812
rect 3605 7803 3663 7809
rect 3605 7800 3617 7803
rect 3200 7772 3617 7800
rect 3200 7760 3206 7772
rect 3252 7741 3280 7772
rect 3605 7769 3617 7772
rect 3651 7769 3663 7803
rect 3605 7763 3663 7769
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7701 3295 7735
rect 3712 7732 3740 7840
rect 3988 7812 4016 7908
rect 4065 7905 4077 7939
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7905 5043 7939
rect 5092 7936 5120 8032
rect 6178 7964 6184 8016
rect 6236 7970 6242 8016
rect 6236 7964 6316 7970
rect 6638 7964 6644 8016
rect 6696 7964 6702 8016
rect 11514 7964 11520 8016
rect 11572 8004 11578 8016
rect 12526 8004 12532 8016
rect 11572 7976 11652 8004
rect 11572 7964 11578 7976
rect 6196 7945 6316 7964
rect 5261 7939 5319 7945
rect 6196 7942 6324 7945
rect 5261 7936 5273 7939
rect 5092 7908 5273 7936
rect 4985 7899 5043 7905
rect 5261 7905 5273 7908
rect 5307 7905 5319 7939
rect 5261 7899 5319 7905
rect 6266 7939 6324 7942
rect 6266 7905 6278 7939
rect 6312 7905 6324 7939
rect 6266 7899 6324 7905
rect 6353 7939 6411 7945
rect 6353 7905 6365 7939
rect 6399 7938 6411 7939
rect 6399 7936 6500 7938
rect 6656 7936 6684 7964
rect 6399 7910 6684 7936
rect 6399 7905 6411 7910
rect 6472 7908 6684 7910
rect 6733 7939 6791 7945
rect 6353 7899 6411 7905
rect 6733 7905 6745 7939
rect 6779 7936 6791 7939
rect 6822 7936 6828 7948
rect 6779 7908 6828 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 3970 7760 3976 7812
rect 4028 7760 4034 7812
rect 4080 7732 4108 7899
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 9306 7896 9312 7948
rect 9364 7896 9370 7948
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 10226 7936 10232 7948
rect 9631 7908 10232 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11146 7896 11152 7948
rect 11204 7896 11210 7948
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11624 7945 11652 7976
rect 11716 7976 12532 8004
rect 11716 7945 11744 7976
rect 12526 7964 12532 7976
rect 12584 7964 12590 8016
rect 12728 7976 13860 8004
rect 12728 7948 12756 7976
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 11296 7908 11345 7936
rect 11296 7896 11302 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 11701 7939 11759 7945
rect 11701 7905 11713 7939
rect 11747 7905 11759 7939
rect 11701 7899 11759 7905
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 12342 7936 12348 7948
rect 11931 7908 12348 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 12342 7896 12348 7908
rect 12400 7936 12406 7948
rect 12710 7936 12716 7948
rect 12400 7908 12716 7936
rect 12400 7896 12406 7908
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 13832 7945 13860 7976
rect 13725 7939 13783 7945
rect 13725 7936 13737 7939
rect 13320 7908 13737 7936
rect 13320 7896 13326 7908
rect 13725 7905 13737 7908
rect 13771 7905 13783 7939
rect 13725 7899 13783 7905
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7905 13875 7939
rect 13817 7899 13875 7905
rect 13998 7896 14004 7948
rect 14056 7896 14062 7948
rect 14090 7896 14096 7948
rect 14148 7896 14154 7948
rect 14182 7896 14188 7948
rect 14240 7896 14246 7948
rect 14384 7945 14412 8044
rect 14826 8032 14832 8084
rect 14884 8032 14890 8084
rect 14918 8032 14924 8084
rect 14976 8072 14982 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 14976 8044 15577 8072
rect 14976 8032 14982 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 17034 8032 17040 8084
rect 17092 8032 17098 8084
rect 17221 8075 17279 8081
rect 17221 8041 17233 8075
rect 17267 8072 17279 8075
rect 20349 8075 20407 8081
rect 17267 8044 18552 8072
rect 17267 8041 17279 8044
rect 17221 8035 17279 8041
rect 14844 8004 14872 8032
rect 17052 8004 17080 8032
rect 14476 7976 14780 8004
rect 14844 7976 15424 8004
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7905 14427 7939
rect 14369 7899 14427 7905
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 5684 7840 5842 7868
rect 5684 7828 5690 7840
rect 8846 7828 8852 7880
rect 8904 7828 8910 7880
rect 11164 7868 11192 7896
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11164 7840 11529 7868
rect 11517 7837 11529 7840
rect 11563 7868 11575 7871
rect 13170 7868 13176 7880
rect 11563 7840 13176 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 14108 7868 14136 7896
rect 14476 7868 14504 7976
rect 14642 7896 14648 7948
rect 14700 7896 14706 7948
rect 14752 7936 14780 7976
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 14752 7908 14841 7936
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 15286 7896 15292 7948
rect 15344 7896 15350 7948
rect 15396 7945 15424 7976
rect 16960 7976 17080 8004
rect 17313 8007 17371 8013
rect 16960 7945 16988 7976
rect 17313 7973 17325 8007
rect 17359 8004 17371 8007
rect 17494 8004 17500 8016
rect 17359 7976 17500 8004
rect 17359 7973 17371 7976
rect 17313 7967 17371 7973
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 18524 8004 18552 8044
rect 20349 8041 20361 8075
rect 20395 8072 20407 8075
rect 20809 8075 20867 8081
rect 20809 8072 20821 8075
rect 20395 8044 20821 8072
rect 20395 8041 20407 8044
rect 20349 8035 20407 8041
rect 20809 8041 20821 8044
rect 20855 8041 20867 8075
rect 20809 8035 20867 8041
rect 20717 8007 20775 8013
rect 20717 8004 20729 8007
rect 18524 7976 20729 8004
rect 20717 7973 20729 7976
rect 20763 7973 20775 8007
rect 20717 7967 20775 7973
rect 15381 7939 15439 7945
rect 15381 7905 15393 7939
rect 15427 7905 15439 7939
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 15381 7899 15439 7905
rect 16684 7908 16865 7936
rect 14108 7840 14504 7868
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 15470 7868 15476 7880
rect 14599 7840 15476 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 7208 7772 11100 7800
rect 7208 7744 7236 7772
rect 3712 7704 4108 7732
rect 3237 7695 3295 7701
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 5350 7732 5356 7744
rect 4212 7704 5356 7732
rect 4212 7692 4218 7704
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 5445 7735 5503 7741
rect 5445 7701 5457 7735
rect 5491 7732 5503 7735
rect 5994 7732 6000 7744
rect 5491 7704 6000 7732
rect 5491 7701 5503 7704
rect 5445 7695 5503 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 7190 7692 7196 7744
rect 7248 7692 7254 7744
rect 7282 7692 7288 7744
rect 7340 7692 7346 7744
rect 11072 7732 11100 7772
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 11606 7800 11612 7812
rect 11204 7772 11612 7800
rect 11204 7760 11210 7772
rect 11606 7760 11612 7772
rect 11664 7800 11670 7812
rect 15105 7803 15163 7809
rect 15105 7800 15117 7803
rect 11664 7772 12112 7800
rect 11664 7760 11670 7772
rect 11974 7732 11980 7744
rect 11072 7704 11980 7732
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 12084 7732 12112 7772
rect 14200 7772 15117 7800
rect 14200 7732 14228 7772
rect 15105 7769 15117 7772
rect 15151 7769 15163 7803
rect 16684 7800 16712 7908
rect 16853 7905 16865 7908
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 16945 7939 17003 7945
rect 16945 7905 16957 7939
rect 16991 7905 17003 7939
rect 16945 7899 17003 7905
rect 17037 7939 17095 7945
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 18690 7936 18696 7948
rect 17083 7908 18696 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 18690 7896 18696 7908
rect 18748 7936 18754 7948
rect 19705 7939 19763 7945
rect 19705 7936 19717 7939
rect 18748 7908 19717 7936
rect 18748 7896 18754 7908
rect 19705 7905 19717 7908
rect 19751 7905 19763 7939
rect 19705 7899 19763 7905
rect 19794 7896 19800 7948
rect 19852 7936 19858 7948
rect 20165 7939 20223 7945
rect 19852 7908 20116 7936
rect 19852 7896 19858 7908
rect 16758 7828 16764 7880
rect 16816 7868 16822 7880
rect 17770 7868 17776 7880
rect 16816 7840 17776 7868
rect 16816 7828 16822 7840
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 19978 7828 19984 7880
rect 20036 7828 20042 7880
rect 20088 7868 20116 7908
rect 20165 7905 20177 7939
rect 20211 7936 20223 7939
rect 20530 7936 20536 7948
rect 20211 7908 20536 7936
rect 20211 7905 20223 7908
rect 20165 7899 20223 7905
rect 20530 7896 20536 7908
rect 20588 7896 20594 7948
rect 20806 7896 20812 7948
rect 20864 7936 20870 7948
rect 21617 7939 21675 7945
rect 21617 7936 21629 7939
rect 20864 7908 21629 7936
rect 20864 7896 20870 7908
rect 21617 7905 21629 7908
rect 21663 7905 21675 7939
rect 21617 7899 21675 7905
rect 20254 7868 20260 7880
rect 20088 7840 20260 7868
rect 20254 7828 20260 7840
rect 20312 7868 20318 7880
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 20312 7840 20453 7868
rect 20312 7828 20318 7840
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20926 7871 20984 7877
rect 20926 7868 20938 7871
rect 20772 7840 20938 7868
rect 20772 7828 20778 7840
rect 20926 7837 20938 7840
rect 20972 7837 20984 7871
rect 20926 7831 20984 7837
rect 21361 7871 21419 7877
rect 21361 7837 21373 7871
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21376 7800 21404 7831
rect 16684 7772 16804 7800
rect 15105 7763 15163 7769
rect 16776 7744 16804 7772
rect 18800 7772 21404 7800
rect 18800 7744 18828 7772
rect 12084 7704 14228 7732
rect 15013 7735 15071 7741
rect 15013 7701 15025 7735
rect 15059 7732 15071 7735
rect 15470 7732 15476 7744
rect 15059 7704 15476 7732
rect 15059 7701 15071 7704
rect 15013 7695 15071 7701
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 16758 7692 16764 7744
rect 16816 7692 16822 7744
rect 17126 7692 17132 7744
rect 17184 7732 17190 7744
rect 17954 7732 17960 7744
rect 17184 7704 17960 7732
rect 17184 7692 17190 7704
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18782 7692 18788 7744
rect 18840 7692 18846 7744
rect 19429 7735 19487 7741
rect 19429 7701 19441 7735
rect 19475 7732 19487 7735
rect 19978 7732 19984 7744
rect 19475 7704 19984 7732
rect 19475 7701 19487 7704
rect 19429 7695 19487 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 21082 7692 21088 7744
rect 21140 7692 21146 7744
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 22741 7735 22799 7741
rect 22741 7732 22753 7735
rect 21416 7704 22753 7732
rect 21416 7692 21422 7704
rect 22741 7701 22753 7704
rect 22787 7701 22799 7735
rect 22741 7695 22799 7701
rect 552 7642 23368 7664
rect 552 7590 1366 7642
rect 1418 7590 1430 7642
rect 1482 7590 1494 7642
rect 1546 7590 1558 7642
rect 1610 7590 1622 7642
rect 1674 7590 1686 7642
rect 1738 7590 7366 7642
rect 7418 7590 7430 7642
rect 7482 7590 7494 7642
rect 7546 7590 7558 7642
rect 7610 7590 7622 7642
rect 7674 7590 7686 7642
rect 7738 7590 13366 7642
rect 13418 7590 13430 7642
rect 13482 7590 13494 7642
rect 13546 7590 13558 7642
rect 13610 7590 13622 7642
rect 13674 7590 13686 7642
rect 13738 7590 19366 7642
rect 19418 7590 19430 7642
rect 19482 7590 19494 7642
rect 19546 7590 19558 7642
rect 19610 7590 19622 7642
rect 19674 7590 19686 7642
rect 19738 7590 23368 7642
rect 552 7568 23368 7590
rect 1118 7488 1124 7540
rect 1176 7528 1182 7540
rect 1397 7531 1455 7537
rect 1397 7528 1409 7531
rect 1176 7500 1409 7528
rect 1176 7488 1182 7500
rect 1397 7497 1409 7500
rect 1443 7497 1455 7531
rect 1397 7491 1455 7497
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 2924 7500 3249 7528
rect 2924 7488 2930 7500
rect 3237 7497 3249 7500
rect 3283 7497 3295 7531
rect 3237 7491 3295 7497
rect 3326 7488 3332 7540
rect 3384 7488 3390 7540
rect 3697 7531 3755 7537
rect 3697 7497 3709 7531
rect 3743 7497 3755 7531
rect 3697 7491 3755 7497
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 2958 7392 2964 7404
rect 2648 7364 2964 7392
rect 2648 7352 2654 7364
rect 2958 7352 2964 7364
rect 3016 7392 3022 7404
rect 3053 7395 3111 7401
rect 3053 7392 3065 7395
rect 3016 7364 3065 7392
rect 3016 7352 3022 7364
rect 3053 7361 3065 7364
rect 3099 7361 3111 7395
rect 3344 7392 3372 7488
rect 3712 7460 3740 7491
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 7190 7528 7196 7540
rect 5500 7500 7196 7528
rect 5500 7488 5506 7500
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7340 7500 12756 7528
rect 7340 7488 7346 7500
rect 3973 7463 4031 7469
rect 3973 7460 3985 7463
rect 3712 7432 3985 7460
rect 3973 7429 3985 7432
rect 4019 7460 4031 7463
rect 4062 7460 4068 7472
rect 4019 7432 4068 7460
rect 4019 7429 4031 7432
rect 3973 7423 4031 7429
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4154 7420 4160 7472
rect 4212 7420 4218 7472
rect 10870 7420 10876 7472
rect 10928 7460 10934 7472
rect 11882 7460 11888 7472
rect 10928 7432 11888 7460
rect 10928 7420 10934 7432
rect 11882 7420 11888 7432
rect 11940 7420 11946 7472
rect 12728 7460 12756 7500
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 13538 7528 13544 7540
rect 12860 7500 13544 7528
rect 12860 7488 12866 7500
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 15473 7531 15531 7537
rect 13780 7500 15424 7528
rect 13780 7488 13786 7500
rect 14734 7460 14740 7472
rect 12728 7432 14740 7460
rect 5632 7404 5684 7410
rect 3344 7364 3832 7392
rect 3053 7355 3111 7361
rect 3804 7336 3832 7364
rect 7834 7392 7840 7404
rect 5632 7346 5684 7352
rect 7484 7364 7840 7392
rect 1394 7284 1400 7336
rect 1452 7284 1458 7336
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 1854 7324 1860 7336
rect 1627 7296 1860 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 1854 7284 1860 7296
rect 1912 7324 1918 7336
rect 2406 7324 2412 7336
rect 1912 7296 2412 7324
rect 1912 7284 1918 7296
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 3421 7327 3479 7333
rect 2823 7296 3280 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 3252 7268 3280 7296
rect 3421 7293 3433 7327
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3234 7216 3240 7268
rect 3292 7216 3298 7268
rect 3436 7256 3464 7287
rect 3510 7284 3516 7336
rect 3568 7284 3574 7336
rect 3694 7284 3700 7336
rect 3752 7284 3758 7336
rect 3786 7284 3792 7336
rect 3844 7284 3850 7336
rect 4062 7324 4068 7336
rect 3896 7296 4068 7324
rect 3896 7256 3924 7296
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 4304 7296 4721 7324
rect 4304 7284 4310 7296
rect 4709 7293 4721 7296
rect 4755 7324 4767 7327
rect 4982 7324 4988 7336
rect 4755 7296 4988 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5166 7284 5172 7336
rect 5224 7284 5230 7336
rect 7484 7333 7512 7364
rect 7834 7352 7840 7364
rect 7892 7392 7898 7404
rect 12434 7392 12440 7404
rect 7892 7364 12440 7392
rect 7892 7352 7898 7364
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 12526 7352 12532 7404
rect 12584 7392 12590 7404
rect 13170 7392 13176 7404
rect 12584 7364 13176 7392
rect 12584 7352 12590 7364
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 13320 7364 13369 7392
rect 13320 7352 13326 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 9950 7284 9956 7336
rect 10008 7284 10014 7336
rect 10137 7327 10195 7333
rect 10137 7293 10149 7327
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7324 10379 7327
rect 10686 7324 10692 7336
rect 10367 7296 10692 7324
rect 10367 7293 10379 7296
rect 10321 7287 10379 7293
rect 3436 7228 3924 7256
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5258 7256 5264 7268
rect 5123 7228 5264 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 10152 7256 10180 7287
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 10962 7324 10968 7336
rect 10919 7296 10968 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 10226 7256 10232 7268
rect 5592 7228 10088 7256
rect 10152 7228 10232 7256
rect 5592 7216 5598 7228
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 4304 7160 4353 7188
rect 4304 7148 4310 7160
rect 4341 7157 4353 7160
rect 4387 7157 4399 7191
rect 4341 7151 4399 7157
rect 5442 7148 5448 7200
rect 5500 7148 5506 7200
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6454 7188 6460 7200
rect 6227 7160 6460 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 10060 7188 10088 7228
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 10413 7259 10471 7265
rect 10413 7225 10425 7259
rect 10459 7225 10471 7259
rect 10413 7219 10471 7225
rect 10597 7259 10655 7265
rect 10597 7225 10609 7259
rect 10643 7225 10655 7259
rect 10796 7256 10824 7287
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11054 7284 11060 7336
rect 11112 7284 11118 7336
rect 11146 7284 11152 7336
rect 11204 7284 11210 7336
rect 11238 7284 11244 7336
rect 11296 7284 11302 7336
rect 11698 7284 11704 7336
rect 11756 7284 11762 7336
rect 11790 7284 11796 7336
rect 11848 7284 11854 7336
rect 11882 7284 11888 7336
rect 11940 7284 11946 7336
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 11992 7256 12020 7287
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 12986 7324 12992 7336
rect 12860 7296 12992 7324
rect 12860 7284 12866 7296
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7293 13139 7327
rect 13081 7287 13139 7293
rect 10796 7228 12020 7256
rect 12084 7228 12296 7256
rect 10597 7219 10655 7225
rect 10428 7188 10456 7219
rect 10060 7160 10456 7188
rect 10612 7188 10640 7219
rect 11330 7188 11336 7200
rect 10612 7160 11336 7188
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11514 7148 11520 7200
rect 11572 7148 11578 7200
rect 11606 7148 11612 7200
rect 11664 7188 11670 7200
rect 12084 7188 12112 7228
rect 11664 7160 12112 7188
rect 11664 7148 11670 7160
rect 12158 7148 12164 7200
rect 12216 7148 12222 7200
rect 12268 7188 12296 7228
rect 12526 7216 12532 7268
rect 12584 7256 12590 7268
rect 13096 7256 13124 7287
rect 13538 7284 13544 7336
rect 13596 7284 13602 7336
rect 13740 7333 13768 7432
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 14826 7420 14832 7472
rect 14884 7460 14890 7472
rect 15102 7460 15108 7472
rect 14884 7432 15108 7460
rect 14884 7420 14890 7432
rect 15102 7420 15108 7432
rect 15160 7460 15166 7472
rect 15396 7460 15424 7500
rect 15473 7497 15485 7531
rect 15519 7528 15531 7531
rect 15654 7528 15660 7540
rect 15519 7500 15660 7528
rect 15519 7497 15531 7500
rect 15473 7491 15531 7497
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 18690 7528 18696 7540
rect 17635 7500 18696 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 15160 7432 15332 7460
rect 15396 7432 16528 7460
rect 15160 7420 15166 7432
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 13906 7352 13912 7404
rect 13964 7352 13970 7404
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 14752 7392 14780 7420
rect 14752 7364 15240 7392
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 13446 7256 13452 7268
rect 12584 7228 13452 7256
rect 12584 7216 12590 7228
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 13630 7216 13636 7268
rect 13688 7256 13694 7268
rect 14108 7256 14136 7287
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 15212 7333 15240 7364
rect 15304 7333 15332 7432
rect 15470 7352 15476 7404
rect 15528 7352 15534 7404
rect 15838 7352 15844 7404
rect 15896 7392 15902 7404
rect 16500 7401 16528 7432
rect 17402 7420 17408 7472
rect 17460 7420 17466 7472
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 15896 7364 16221 7392
rect 15896 7352 15902 7364
rect 16209 7361 16221 7364
rect 16255 7361 16267 7395
rect 16209 7355 16267 7361
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7392 16543 7395
rect 16758 7392 16764 7404
rect 16531 7364 16764 7392
rect 16531 7361 16543 7364
rect 16485 7355 16543 7361
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 17604 7392 17632 7491
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 18782 7488 18788 7540
rect 18840 7488 18846 7540
rect 19334 7488 19340 7540
rect 19392 7528 19398 7540
rect 20346 7528 20352 7540
rect 19392 7500 20352 7528
rect 19392 7488 19398 7500
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 20806 7488 20812 7540
rect 20864 7488 20870 7540
rect 21082 7488 21088 7540
rect 21140 7488 21146 7540
rect 18800 7460 18828 7488
rect 18800 7432 19012 7460
rect 18984 7401 19012 7432
rect 20530 7420 20536 7472
rect 20588 7460 20594 7472
rect 20993 7463 21051 7469
rect 20993 7460 21005 7463
rect 20588 7432 21005 7460
rect 20588 7420 20594 7432
rect 20993 7429 21005 7432
rect 21039 7429 21051 7463
rect 20993 7423 21051 7429
rect 17773 7395 17831 7401
rect 17773 7392 17785 7395
rect 17144 7364 17632 7392
rect 17696 7364 17785 7392
rect 14553 7327 14611 7333
rect 14553 7324 14565 7327
rect 14240 7296 14565 7324
rect 14240 7284 14246 7296
rect 14553 7293 14565 7296
rect 14599 7293 14611 7327
rect 14553 7287 14611 7293
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7324 14795 7327
rect 15197 7327 15255 7333
rect 14783 7296 15148 7324
rect 14783 7293 14795 7296
rect 14737 7287 14795 7293
rect 13688 7228 14136 7256
rect 13688 7216 13694 7228
rect 14458 7216 14464 7268
rect 14516 7256 14522 7268
rect 14660 7256 14688 7287
rect 15013 7259 15071 7265
rect 15013 7256 15025 7259
rect 14516 7228 14688 7256
rect 14752 7228 15025 7256
rect 14516 7216 14522 7228
rect 13722 7188 13728 7200
rect 12268 7160 13728 7188
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 14277 7191 14335 7197
rect 14277 7188 14289 7191
rect 13872 7160 14289 7188
rect 13872 7148 13878 7160
rect 14277 7157 14289 7160
rect 14323 7157 14335 7191
rect 14277 7151 14335 7157
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 14752 7188 14780 7228
rect 15013 7225 15025 7228
rect 15059 7225 15071 7259
rect 15120 7256 15148 7296
rect 15197 7293 15209 7327
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7293 15347 7327
rect 15289 7287 15347 7293
rect 15488 7256 15516 7352
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7324 15623 7327
rect 16850 7324 16856 7336
rect 15611 7296 16856 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 17144 7333 17172 7364
rect 17696 7336 17724 7364
rect 17773 7361 17785 7364
rect 17819 7361 17831 7395
rect 18969 7395 19027 7401
rect 17773 7355 17831 7361
rect 17972 7364 18828 7392
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7293 17187 7327
rect 17497 7327 17555 7333
rect 17497 7324 17509 7327
rect 17129 7287 17187 7293
rect 17236 7296 17509 7324
rect 15120 7228 15516 7256
rect 15013 7219 15071 7225
rect 17236 7200 17264 7296
rect 17497 7293 17509 7296
rect 17543 7293 17555 7327
rect 17497 7287 17555 7293
rect 17678 7284 17684 7336
rect 17736 7284 17742 7336
rect 17972 7333 18000 7364
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 18138 7284 18144 7336
rect 18196 7284 18202 7336
rect 18322 7284 18328 7336
rect 18380 7284 18386 7336
rect 18690 7284 18696 7336
rect 18748 7284 18754 7336
rect 18800 7333 18828 7364
rect 18969 7361 18981 7395
rect 19015 7361 19027 7395
rect 21100 7392 21128 7488
rect 18969 7355 19027 7361
rect 20640 7364 21128 7392
rect 18785 7327 18843 7333
rect 18785 7293 18797 7327
rect 18831 7293 18843 7327
rect 18785 7287 18843 7293
rect 18874 7284 18880 7336
rect 18932 7284 18938 7336
rect 18984 7324 19012 7355
rect 19794 7324 19800 7336
rect 18984 7296 19800 7324
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 20640 7333 20668 7364
rect 20625 7327 20683 7333
rect 20625 7293 20637 7327
rect 20671 7293 20683 7327
rect 20625 7287 20683 7293
rect 21085 7327 21143 7333
rect 21085 7293 21097 7327
rect 21131 7324 21143 7327
rect 21358 7324 21364 7336
rect 21131 7296 21364 7324
rect 21131 7293 21143 7296
rect 21085 7287 21143 7293
rect 21358 7284 21364 7296
rect 21416 7284 21422 7336
rect 17405 7259 17463 7265
rect 17405 7225 17417 7259
rect 17451 7256 17463 7259
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 17451 7228 17785 7256
rect 17451 7225 17463 7228
rect 17405 7219 17463 7225
rect 17773 7225 17785 7228
rect 17819 7225 17831 7259
rect 18233 7259 18291 7265
rect 18233 7256 18245 7259
rect 17773 7219 17831 7225
rect 17972 7228 18245 7256
rect 17972 7200 18000 7228
rect 18233 7225 18245 7228
rect 18279 7225 18291 7259
rect 19214 7259 19272 7265
rect 19214 7256 19226 7259
rect 18233 7219 18291 7225
rect 18524 7228 19226 7256
rect 14700 7160 14780 7188
rect 14921 7191 14979 7197
rect 14700 7148 14706 7160
rect 14921 7157 14933 7191
rect 14967 7188 14979 7191
rect 17034 7188 17040 7200
rect 14967 7160 17040 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 17218 7148 17224 7200
rect 17276 7148 17282 7200
rect 17954 7148 17960 7200
rect 18012 7148 18018 7200
rect 18524 7197 18552 7228
rect 19214 7225 19226 7228
rect 19260 7225 19272 7259
rect 19214 7219 19272 7225
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7157 18567 7191
rect 18509 7151 18567 7157
rect 552 7098 23368 7120
rect 552 7046 4366 7098
rect 4418 7046 4430 7098
rect 4482 7046 4494 7098
rect 4546 7046 4558 7098
rect 4610 7046 4622 7098
rect 4674 7046 4686 7098
rect 4738 7046 10366 7098
rect 10418 7046 10430 7098
rect 10482 7046 10494 7098
rect 10546 7046 10558 7098
rect 10610 7046 10622 7098
rect 10674 7046 10686 7098
rect 10738 7046 16366 7098
rect 16418 7046 16430 7098
rect 16482 7046 16494 7098
rect 16546 7046 16558 7098
rect 16610 7046 16622 7098
rect 16674 7046 16686 7098
rect 16738 7046 22366 7098
rect 22418 7046 22430 7098
rect 22482 7046 22494 7098
rect 22546 7046 22558 7098
rect 22610 7046 22622 7098
rect 22674 7046 22686 7098
rect 22738 7046 23368 7098
rect 552 7024 23368 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 1765 6987 1823 6993
rect 1765 6984 1777 6987
rect 1452 6956 1777 6984
rect 1452 6944 1458 6956
rect 1765 6953 1777 6956
rect 1811 6953 1823 6987
rect 1765 6947 1823 6953
rect 2130 6944 2136 6996
rect 2188 6944 2194 6996
rect 2406 6944 2412 6996
rect 2464 6944 2470 6996
rect 3329 6987 3387 6993
rect 2516 6956 3280 6984
rect 2148 6916 2176 6944
rect 2516 6916 2544 6956
rect 2590 6925 2596 6928
rect 2148 6888 2544 6916
rect 2577 6919 2596 6925
rect 2577 6885 2589 6919
rect 2577 6879 2596 6885
rect 2590 6876 2596 6879
rect 2648 6876 2654 6928
rect 2777 6919 2835 6925
rect 2777 6885 2789 6919
rect 2823 6916 2835 6919
rect 2958 6916 2964 6928
rect 2823 6888 2964 6916
rect 2823 6885 2835 6888
rect 2777 6879 2835 6885
rect 2958 6876 2964 6888
rect 3016 6916 3022 6928
rect 3252 6916 3280 6956
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 3510 6984 3516 6996
rect 3375 6956 3516 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 3605 6987 3663 6993
rect 3605 6953 3617 6987
rect 3651 6953 3663 6987
rect 3605 6947 3663 6953
rect 3620 6916 3648 6947
rect 3786 6944 3792 6996
rect 3844 6944 3850 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 5258 6984 5264 6996
rect 4120 6956 5264 6984
rect 4120 6944 4126 6956
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 6086 6944 6092 6996
rect 6144 6984 6150 6996
rect 6144 6956 6224 6984
rect 6144 6944 6150 6956
rect 5442 6916 5448 6928
rect 3016 6888 3188 6916
rect 3252 6888 5448 6916
rect 3016 6876 3022 6888
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2087 6820 2774 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 2746 6780 2774 6820
rect 2866 6808 2872 6860
rect 2924 6808 2930 6860
rect 3160 6857 3188 6888
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 6196 6916 6224 6956
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 6420 6956 7389 6984
rect 6420 6944 6426 6956
rect 7377 6953 7389 6956
rect 7423 6984 7435 6987
rect 7423 6956 9076 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 9048 6928 9076 6956
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10226 6984 10232 6996
rect 10008 6956 10232 6984
rect 10008 6944 10014 6956
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 11146 6944 11152 6996
rect 11204 6944 11210 6996
rect 11330 6944 11336 6996
rect 11388 6984 11394 6996
rect 11698 6984 11704 6996
rect 11388 6956 11704 6984
rect 11388 6944 11394 6956
rect 11698 6944 11704 6956
rect 11756 6984 11762 6996
rect 12066 6984 12072 6996
rect 11756 6956 12072 6984
rect 11756 6944 11762 6956
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12400 6956 12664 6984
rect 12400 6944 12406 6956
rect 6273 6919 6331 6925
rect 6273 6916 6285 6919
rect 6196 6888 6285 6916
rect 6273 6885 6285 6888
rect 6319 6885 6331 6919
rect 6273 6879 6331 6885
rect 6454 6876 6460 6928
rect 6512 6916 6518 6928
rect 8294 6916 8300 6928
rect 6512 6888 7135 6916
rect 6512 6876 6518 6888
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6817 3203 6851
rect 3145 6811 3203 6817
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6817 3387 6851
rect 3329 6811 3387 6817
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 3602 6848 3608 6860
rect 3467 6820 3608 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 3234 6780 3240 6792
rect 2746 6752 3240 6780
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3344 6712 3372 6811
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 3694 6808 3700 6860
rect 3752 6848 3758 6860
rect 3970 6848 3976 6860
rect 3752 6820 3976 6848
rect 3752 6808 3758 6820
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6817 4215 6851
rect 4617 6851 4675 6857
rect 4617 6848 4629 6851
rect 4157 6811 4215 6817
rect 4264 6820 4629 6848
rect 3620 6780 3648 6808
rect 4172 6780 4200 6811
rect 4264 6792 4292 6820
rect 4617 6817 4629 6820
rect 4663 6848 4675 6851
rect 4798 6848 4804 6860
rect 4663 6820 4804 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 5902 6808 5908 6860
rect 5960 6848 5966 6860
rect 6012 6848 6224 6854
rect 6549 6851 6607 6857
rect 6549 6848 6561 6851
rect 5960 6826 6561 6848
rect 5960 6820 6040 6826
rect 6196 6820 6561 6826
rect 5960 6808 5966 6820
rect 6549 6817 6561 6820
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6848 6699 6851
rect 6730 6848 6736 6860
rect 6687 6820 6736 6848
rect 6687 6817 6699 6820
rect 6641 6811 6699 6817
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 7006 6808 7012 6860
rect 7064 6808 7070 6860
rect 7107 6848 7135 6888
rect 7852 6888 8300 6916
rect 7852 6857 7880 6888
rect 8294 6876 8300 6888
rect 8352 6916 8358 6928
rect 8570 6916 8576 6928
rect 8352 6888 8576 6916
rect 8352 6876 8358 6888
rect 8570 6876 8576 6888
rect 8628 6876 8634 6928
rect 9030 6876 9036 6928
rect 9088 6876 9094 6928
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 11164 6916 11192 6944
rect 12636 6928 12664 6956
rect 13170 6944 13176 6996
rect 13228 6944 13234 6996
rect 13446 6944 13452 6996
rect 13504 6944 13510 6996
rect 14001 6987 14059 6993
rect 14001 6953 14013 6987
rect 14047 6984 14059 6987
rect 16758 6984 16764 6996
rect 14047 6956 14872 6984
rect 14047 6953 14059 6956
rect 14001 6947 14059 6953
rect 10744 6888 11008 6916
rect 11164 6888 11560 6916
rect 10744 6876 10750 6888
rect 7837 6851 7895 6857
rect 7107 6820 7420 6848
rect 3620 6752 4200 6780
rect 4172 6712 4200 6752
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 7392 6780 7420 6820
rect 7837 6817 7849 6851
rect 7883 6817 7895 6851
rect 7837 6811 7895 6817
rect 8380 6851 8438 6857
rect 8380 6817 8392 6851
rect 8426 6848 8438 6851
rect 9582 6848 9588 6860
rect 8426 6820 9588 6848
rect 8426 6817 8438 6820
rect 8380 6811 8438 6817
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 10980 6857 11008 6888
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 10965 6851 11023 6857
rect 10965 6817 10977 6851
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 5684 6752 6118 6780
rect 7392 6752 8125 6780
rect 5684 6740 5690 6752
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 4433 6715 4491 6721
rect 4433 6712 4445 6715
rect 3344 6684 3924 6712
rect 4172 6684 4445 6712
rect 1946 6604 1952 6656
rect 2004 6604 2010 6656
rect 2593 6647 2651 6653
rect 2593 6613 2605 6647
rect 2639 6644 2651 6647
rect 2866 6644 2872 6656
rect 2639 6616 2872 6644
rect 2639 6613 2651 6616
rect 2593 6607 2651 6613
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3786 6644 3792 6656
rect 3099 6616 3792 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 3896 6644 3924 6684
rect 4433 6681 4445 6684
rect 4479 6681 4491 6715
rect 4433 6675 4491 6681
rect 7561 6715 7619 6721
rect 7561 6681 7573 6715
rect 7607 6712 7619 6715
rect 9416 6712 9444 6740
rect 9493 6715 9551 6721
rect 9493 6712 9505 6715
rect 7607 6684 8156 6712
rect 9416 6684 9505 6712
rect 7607 6681 7619 6684
rect 7561 6675 7619 6681
rect 4154 6644 4160 6656
rect 3896 6616 4160 6644
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 5074 6644 5080 6656
rect 4387 6616 5080 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 5074 6604 5080 6616
rect 5132 6644 5138 6656
rect 6270 6644 6276 6656
rect 5132 6616 6276 6644
rect 5132 6604 5138 6616
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 8018 6604 8024 6656
rect 8076 6604 8082 6656
rect 8128 6644 8156 6684
rect 9493 6681 9505 6684
rect 9539 6681 9551 6715
rect 9493 6675 9551 6681
rect 10612 6656 10640 6811
rect 10796 6780 10824 6811
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11149 6851 11207 6857
rect 11149 6848 11161 6851
rect 11112 6820 11161 6848
rect 11112 6808 11118 6820
rect 11149 6817 11161 6820
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 11256 6780 11284 6811
rect 11330 6808 11336 6860
rect 11388 6808 11394 6860
rect 11532 6857 11560 6888
rect 12618 6876 12624 6928
rect 12676 6876 12682 6928
rect 13188 6916 13216 6944
rect 13464 6916 13492 6944
rect 13188 6888 13400 6916
rect 13464 6888 14320 6916
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 11606 6808 11612 6860
rect 11664 6808 11670 6860
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 11940 6820 12265 6848
rect 11940 6808 11946 6820
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 12253 6811 12311 6817
rect 13265 6851 13323 6857
rect 13265 6817 13277 6851
rect 13311 6817 13323 6851
rect 13372 6848 13400 6888
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13372 6820 13461 6848
rect 13265 6811 13323 6817
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 11624 6780 11652 6808
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 10796 6752 11652 6780
rect 11900 6752 11989 6780
rect 10689 6715 10747 6721
rect 10689 6681 10701 6715
rect 10735 6712 10747 6715
rect 10870 6712 10876 6724
rect 10735 6684 10876 6712
rect 10735 6681 10747 6684
rect 10689 6675 10747 6681
rect 10870 6672 10876 6684
rect 10928 6672 10934 6724
rect 11072 6684 11836 6712
rect 9398 6644 9404 6656
rect 8128 6616 9404 6644
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 10594 6604 10600 6656
rect 10652 6604 10658 6656
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 11072 6644 11100 6684
rect 10836 6616 11100 6644
rect 10836 6604 10842 6616
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11808 6653 11836 6684
rect 11900 6656 11928 6752
rect 11977 6749 11989 6752
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6749 12219 6783
rect 12161 6743 12219 6749
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11296 6616 11713 6644
rect 11296 6604 11302 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 11793 6647 11851 6653
rect 11793 6613 11805 6647
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 11882 6604 11888 6656
rect 11940 6604 11946 6656
rect 12176 6644 12204 6743
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 13280 6780 13308 6811
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13780 6820 13829 6848
rect 13780 6808 13786 6820
rect 13817 6817 13829 6820
rect 13863 6817 13875 6851
rect 13817 6811 13875 6817
rect 13998 6808 14004 6860
rect 14056 6808 14062 6860
rect 14090 6808 14096 6860
rect 14148 6808 14154 6860
rect 14292 6857 14320 6888
rect 14277 6851 14335 6857
rect 14277 6817 14289 6851
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6848 14611 6851
rect 14734 6848 14740 6860
rect 14599 6820 14740 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 12768 6752 13308 6780
rect 13541 6783 13599 6789
rect 12768 6740 12774 6752
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 14016 6780 14044 6808
rect 13679 6752 14044 6780
rect 14292 6780 14320 6811
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 14844 6857 14872 6956
rect 16592 6956 16764 6984
rect 15654 6876 15660 6928
rect 15712 6916 15718 6928
rect 16114 6916 16120 6928
rect 15712 6888 16120 6916
rect 15712 6876 15718 6888
rect 16114 6876 16120 6888
rect 16172 6876 16178 6928
rect 16592 6857 16620 6956
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 17034 6944 17040 6996
rect 17092 6984 17098 6996
rect 17402 6984 17408 6996
rect 17092 6956 17408 6984
rect 17092 6944 17098 6956
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 21266 6944 21272 6996
rect 21324 6944 21330 6996
rect 17954 6916 17960 6928
rect 17328 6888 17960 6916
rect 17328 6857 17356 6888
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 21008 6888 21404 6916
rect 14829 6851 14887 6857
rect 14829 6817 14841 6851
rect 14875 6817 14887 6851
rect 14829 6811 14887 6817
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6817 16635 6851
rect 17313 6851 17371 6857
rect 17313 6848 17325 6851
rect 16577 6811 16635 6817
rect 16684 6820 17325 6848
rect 16684 6780 16712 6820
rect 17313 6817 17325 6820
rect 17359 6817 17371 6851
rect 17313 6811 17371 6817
rect 17497 6851 17555 6857
rect 17497 6817 17509 6851
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6848 17647 6851
rect 17862 6848 17868 6860
rect 17635 6820 17868 6848
rect 17635 6817 17647 6820
rect 17589 6811 17647 6817
rect 17218 6780 17224 6792
rect 14292 6752 16712 6780
rect 16776 6752 17224 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 13078 6672 13084 6724
rect 13136 6712 13142 6724
rect 13446 6712 13452 6724
rect 13136 6684 13452 6712
rect 13136 6672 13142 6684
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 13556 6712 13584 6743
rect 13906 6712 13912 6724
rect 13556 6684 13912 6712
rect 13906 6672 13912 6684
rect 13964 6672 13970 6724
rect 16776 6721 16804 6752
rect 17218 6740 17224 6752
rect 17276 6780 17282 6792
rect 17512 6780 17540 6811
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 20346 6808 20352 6860
rect 20404 6848 20410 6860
rect 21008 6848 21036 6888
rect 20404 6820 21036 6848
rect 21085 6851 21143 6857
rect 20404 6808 20410 6820
rect 21085 6817 21097 6851
rect 21131 6817 21143 6851
rect 21376 6848 21404 6888
rect 21545 6851 21603 6857
rect 21545 6848 21557 6851
rect 21376 6820 21557 6848
rect 21085 6811 21143 6817
rect 21545 6817 21557 6820
rect 21591 6817 21603 6851
rect 21545 6811 21603 6817
rect 21729 6851 21787 6857
rect 21729 6817 21741 6851
rect 21775 6848 21787 6851
rect 21818 6848 21824 6860
rect 21775 6820 21824 6848
rect 21775 6817 21787 6820
rect 21729 6811 21787 6817
rect 17276 6752 17540 6780
rect 17276 6740 17282 6752
rect 18690 6740 18696 6792
rect 18748 6740 18754 6792
rect 21100 6780 21128 6811
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 21910 6808 21916 6860
rect 21968 6848 21974 6860
rect 22005 6851 22063 6857
rect 22005 6848 22017 6851
rect 21968 6820 22017 6848
rect 21968 6808 21974 6820
rect 22005 6817 22017 6820
rect 22051 6817 22063 6851
rect 22005 6811 22063 6817
rect 21100 6752 21772 6780
rect 16761 6715 16819 6721
rect 16761 6712 16773 6715
rect 14108 6684 16773 6712
rect 14108 6644 14136 6684
rect 16761 6681 16773 6684
rect 16807 6681 16819 6715
rect 16761 6675 16819 6681
rect 17313 6715 17371 6721
rect 17313 6681 17325 6715
rect 17359 6712 17371 6715
rect 18708 6712 18736 6740
rect 17359 6684 18736 6712
rect 17359 6681 17371 6684
rect 17313 6675 17371 6681
rect 21744 6656 21772 6752
rect 12176 6616 14136 6644
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 14458 6644 14464 6656
rect 14231 6616 14464 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 14918 6644 14924 6656
rect 14700 6616 14924 6644
rect 14700 6604 14706 6616
rect 14918 6604 14924 6616
rect 14976 6604 14982 6656
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6644 15071 6647
rect 15102 6644 15108 6656
rect 15059 6616 15108 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 20901 6647 20959 6653
rect 20901 6644 20913 6647
rect 20772 6616 20913 6644
rect 20772 6604 20778 6616
rect 20901 6613 20913 6616
rect 20947 6613 20959 6647
rect 20901 6607 20959 6613
rect 21634 6604 21640 6656
rect 21692 6604 21698 6656
rect 21726 6604 21732 6656
rect 21784 6644 21790 6656
rect 21821 6647 21879 6653
rect 21821 6644 21833 6647
rect 21784 6616 21833 6644
rect 21784 6604 21790 6616
rect 21821 6613 21833 6616
rect 21867 6613 21879 6647
rect 21821 6607 21879 6613
rect 552 6554 23368 6576
rect 552 6502 1366 6554
rect 1418 6502 1430 6554
rect 1482 6502 1494 6554
rect 1546 6502 1558 6554
rect 1610 6502 1622 6554
rect 1674 6502 1686 6554
rect 1738 6502 7366 6554
rect 7418 6502 7430 6554
rect 7482 6502 7494 6554
rect 7546 6502 7558 6554
rect 7610 6502 7622 6554
rect 7674 6502 7686 6554
rect 7738 6502 13366 6554
rect 13418 6502 13430 6554
rect 13482 6502 13494 6554
rect 13546 6502 13558 6554
rect 13610 6502 13622 6554
rect 13674 6502 13686 6554
rect 13738 6502 19366 6554
rect 19418 6502 19430 6554
rect 19482 6502 19494 6554
rect 19546 6502 19558 6554
rect 19610 6502 19622 6554
rect 19674 6502 19686 6554
rect 19738 6502 23368 6554
rect 552 6480 23368 6502
rect 1946 6400 1952 6452
rect 2004 6440 2010 6452
rect 2225 6443 2283 6449
rect 2225 6440 2237 6443
rect 2004 6412 2237 6440
rect 2004 6400 2010 6412
rect 2225 6409 2237 6412
rect 2271 6409 2283 6443
rect 2225 6403 2283 6409
rect 1581 6375 1639 6381
rect 1581 6341 1593 6375
rect 1627 6372 1639 6375
rect 1670 6372 1676 6384
rect 1627 6344 1676 6372
rect 1627 6341 1639 6344
rect 1581 6335 1639 6341
rect 1670 6332 1676 6344
rect 1728 6372 1734 6384
rect 1728 6344 2084 6372
rect 1728 6332 1734 6344
rect 1762 6264 1768 6316
rect 1820 6264 1826 6316
rect 1489 6239 1547 6245
rect 1489 6205 1501 6239
rect 1535 6205 1547 6239
rect 1489 6199 1547 6205
rect 1504 6100 1532 6199
rect 1946 6196 1952 6248
rect 2004 6196 2010 6248
rect 2056 6245 2084 6344
rect 2240 6304 2268 6403
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 2590 6440 2596 6452
rect 2464 6412 2596 6440
rect 2464 6400 2470 6412
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 3602 6440 3608 6452
rect 2823 6412 3608 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5994 6440 6000 6452
rect 5592 6412 6000 6440
rect 5592 6400 5598 6412
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 8570 6400 8576 6452
rect 8628 6400 8634 6452
rect 10502 6440 10508 6452
rect 9646 6412 10508 6440
rect 8018 6332 8024 6384
rect 8076 6372 8082 6384
rect 8941 6375 8999 6381
rect 8941 6372 8953 6375
rect 8076 6344 8953 6372
rect 8076 6332 8082 6344
rect 8941 6341 8953 6344
rect 8987 6341 8999 6375
rect 8941 6335 8999 6341
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 9646 6372 9674 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 12066 6440 12072 6452
rect 10652 6412 12072 6440
rect 10652 6400 10658 6412
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12802 6400 12808 6452
rect 12860 6440 12866 6452
rect 12860 6412 13768 6440
rect 12860 6400 12866 6412
rect 13740 6384 13768 6412
rect 17586 6400 17592 6452
rect 17644 6440 17650 6452
rect 20714 6440 20720 6452
rect 17644 6412 20720 6440
rect 17644 6400 17650 6412
rect 20714 6400 20720 6412
rect 20772 6440 20778 6452
rect 20901 6443 20959 6449
rect 20901 6440 20913 6443
rect 20772 6412 20913 6440
rect 20772 6400 20778 6412
rect 20901 6409 20913 6412
rect 20947 6409 20959 6443
rect 20901 6403 20959 6409
rect 21818 6400 21824 6452
rect 21876 6440 21882 6452
rect 22833 6443 22891 6449
rect 22833 6440 22845 6443
rect 21876 6412 22845 6440
rect 21876 6400 21882 6412
rect 22833 6409 22845 6412
rect 22879 6409 22891 6443
rect 22833 6403 22891 6409
rect 11514 6372 11520 6384
rect 9088 6344 9674 6372
rect 10888 6344 11192 6372
rect 9088 6332 9094 6344
rect 10888 6316 10916 6344
rect 2240 6276 2360 6304
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6236 2099 6239
rect 2222 6236 2228 6248
rect 2087 6208 2228 6236
rect 2087 6205 2099 6208
rect 2041 6199 2099 6205
rect 2222 6196 2228 6208
rect 2280 6196 2286 6248
rect 2332 6245 2360 6276
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 3844 6276 5672 6304
rect 3844 6264 3850 6276
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6205 2375 6239
rect 2317 6199 2375 6205
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6205 2559 6239
rect 2501 6199 2559 6205
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 2516 6168 2544 6199
rect 5534 6196 5540 6248
rect 5592 6196 5598 6248
rect 5644 6236 5672 6276
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 5776 6276 5842 6304
rect 5776 6264 5782 6276
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 10870 6304 10876 6316
rect 7156 6276 10876 6304
rect 7156 6264 7162 6276
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 11164 6313 11192 6344
rect 11256 6344 11520 6372
rect 11256 6313 11284 6344
rect 11514 6332 11520 6344
rect 11572 6332 11578 6384
rect 11716 6344 13676 6372
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6273 11299 6307
rect 11241 6267 11299 6273
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11422 6304 11428 6316
rect 11379 6276 11428 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 11716 6313 11744 6344
rect 11700 6307 11758 6313
rect 11700 6273 11712 6307
rect 11746 6273 11758 6307
rect 11700 6267 11758 6273
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 13648 6304 13676 6344
rect 13722 6332 13728 6384
rect 13780 6372 13786 6384
rect 13909 6375 13967 6381
rect 13909 6372 13921 6375
rect 13780 6344 13921 6372
rect 13780 6332 13786 6344
rect 13909 6341 13921 6344
rect 13955 6341 13967 6375
rect 13909 6335 13967 6341
rect 14182 6332 14188 6384
rect 14240 6372 14246 6384
rect 15010 6372 15016 6384
rect 14240 6344 15016 6372
rect 14240 6332 14246 6344
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 13648 6276 15056 6304
rect 15028 6248 15056 6276
rect 15286 6264 15292 6316
rect 15344 6264 15350 6316
rect 18782 6304 18788 6316
rect 17880 6276 18184 6304
rect 17880 6248 17908 6276
rect 5644 6208 6132 6236
rect 1811 6140 2544 6168
rect 2961 6171 3019 6177
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 4982 6168 4988 6180
rect 3007 6140 4988 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 4982 6128 4988 6140
rect 5040 6128 5046 6180
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 5997 6171 6055 6177
rect 5997 6168 6009 6171
rect 5500 6140 6009 6168
rect 5500 6128 5506 6140
rect 5997 6137 6009 6140
rect 6043 6137 6055 6171
rect 6104 6168 6132 6208
rect 6178 6196 6184 6248
rect 6236 6236 6242 6248
rect 6273 6239 6331 6245
rect 6273 6236 6285 6239
rect 6236 6208 6285 6236
rect 6236 6196 6242 6208
rect 6273 6205 6285 6208
rect 6319 6205 6331 6239
rect 6273 6199 6331 6205
rect 6365 6239 6423 6245
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 6546 6236 6552 6248
rect 6411 6208 6552 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 10594 6236 10600 6248
rect 6656 6208 10600 6236
rect 6656 6168 6684 6208
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 11514 6236 11520 6248
rect 11103 6208 11520 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 11606 6196 11612 6248
rect 11664 6196 11670 6248
rect 11803 6239 11861 6245
rect 11803 6205 11815 6239
rect 11849 6205 11861 6239
rect 13725 6239 13783 6245
rect 11803 6199 11861 6205
rect 12084 6208 13676 6236
rect 6104 6140 6684 6168
rect 5997 6131 6055 6137
rect 6730 6128 6736 6180
rect 6788 6128 6794 6180
rect 11330 6168 11336 6180
rect 7024 6140 11336 6168
rect 1946 6100 1952 6112
rect 1504 6072 1952 6100
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2406 6060 2412 6112
rect 2464 6060 2470 6112
rect 2774 6109 2780 6112
rect 2751 6103 2780 6109
rect 2751 6069 2763 6103
rect 2751 6063 2780 6069
rect 2774 6060 2780 6063
rect 2832 6060 2838 6112
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 7024 6100 7052 6140
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 5776 6072 7052 6100
rect 7101 6103 7159 6109
rect 5776 6060 5782 6072
rect 7101 6069 7113 6103
rect 7147 6100 7159 6103
rect 7190 6100 7196 6112
rect 7147 6072 7196 6100
rect 7147 6069 7159 6072
rect 7101 6063 7159 6069
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 7282 6060 7288 6112
rect 7340 6060 7346 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 8352 6072 8401 6100
rect 8352 6060 8358 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10284 6072 10885 6100
rect 10284 6060 10290 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 11808 6100 11836 6199
rect 12084 6168 12112 6208
rect 11992 6140 12112 6168
rect 11992 6112 12020 6140
rect 12158 6128 12164 6180
rect 12216 6128 12222 6180
rect 12345 6171 12403 6177
rect 12345 6137 12357 6171
rect 12391 6168 12403 6171
rect 12802 6168 12808 6180
rect 12391 6140 12808 6168
rect 12391 6137 12403 6140
rect 12345 6131 12403 6137
rect 12802 6128 12808 6140
rect 12860 6128 12866 6180
rect 13648 6168 13676 6208
rect 13725 6205 13737 6239
rect 13771 6236 13783 6239
rect 13814 6236 13820 6248
rect 13771 6208 13820 6236
rect 13771 6205 13783 6208
rect 13725 6199 13783 6205
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 13906 6196 13912 6248
rect 13964 6236 13970 6248
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13964 6208 14013 6236
rect 13964 6196 13970 6208
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 14844 6168 14872 6199
rect 15010 6196 15016 6248
rect 15068 6196 15074 6248
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 15197 6239 15255 6245
rect 15197 6236 15209 6239
rect 15160 6208 15209 6236
rect 15160 6196 15166 6208
rect 15197 6205 15209 6208
rect 15243 6205 15255 6239
rect 15197 6199 15255 6205
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6205 15439 6239
rect 15381 6199 15439 6205
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6236 15531 6239
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 15519 6208 16129 6236
rect 15519 6205 15531 6208
rect 15473 6199 15531 6205
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 16117 6199 16175 6205
rect 16393 6239 16451 6245
rect 16393 6205 16405 6239
rect 16439 6236 16451 6239
rect 16850 6236 16856 6248
rect 16439 6208 16856 6236
rect 16439 6205 16451 6208
rect 16393 6199 16451 6205
rect 13648 6140 14872 6168
rect 11974 6100 11980 6112
rect 11808 6072 11980 6100
rect 10873 6063 10931 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12069 6103 12127 6109
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12250 6100 12256 6112
rect 12115 6072 12256 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12526 6060 12532 6112
rect 12584 6060 12590 6112
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13541 6103 13599 6109
rect 13541 6100 13553 6103
rect 13044 6072 13553 6100
rect 13044 6060 13050 6072
rect 13541 6069 13553 6072
rect 13587 6069 13599 6103
rect 14844 6100 14872 6140
rect 14921 6171 14979 6177
rect 14921 6137 14933 6171
rect 14967 6168 14979 6171
rect 15396 6168 15424 6199
rect 16850 6196 16856 6208
rect 16908 6236 16914 6248
rect 16908 6208 17816 6236
rect 16908 6196 16914 6208
rect 17788 6180 17816 6208
rect 17862 6196 17868 6248
rect 17920 6196 17926 6248
rect 17954 6196 17960 6248
rect 18012 6196 18018 6248
rect 18156 6245 18184 6276
rect 18340 6276 18788 6304
rect 18340 6248 18368 6276
rect 18782 6264 18788 6276
rect 18840 6304 18846 6316
rect 18840 6276 19104 6304
rect 18840 6264 18846 6276
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 18322 6196 18328 6248
rect 18380 6196 18386 6248
rect 19076 6245 19104 6276
rect 20990 6264 20996 6316
rect 21048 6264 21054 6316
rect 21266 6304 21272 6316
rect 21100 6276 21272 6304
rect 18693 6239 18751 6245
rect 18693 6205 18705 6239
rect 18739 6205 18751 6239
rect 18693 6199 18751 6205
rect 19061 6239 19119 6245
rect 19061 6205 19073 6239
rect 19107 6205 19119 6239
rect 19061 6199 19119 6205
rect 15749 6171 15807 6177
rect 15749 6168 15761 6171
rect 14967 6140 15424 6168
rect 15488 6140 15761 6168
rect 14967 6137 14979 6140
rect 14921 6131 14979 6137
rect 15488 6100 15516 6140
rect 15749 6137 15761 6140
rect 15795 6137 15807 6171
rect 15749 6131 15807 6137
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 15988 6140 16252 6168
rect 15988 6128 15994 6140
rect 14844 6072 15516 6100
rect 15657 6103 15715 6109
rect 13541 6063 13599 6069
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 16114 6100 16120 6112
rect 15703 6072 16120 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 16224 6109 16252 6140
rect 17770 6128 17776 6180
rect 17828 6128 17834 6180
rect 18049 6171 18107 6177
rect 18049 6137 18061 6171
rect 18095 6168 18107 6171
rect 18708 6168 18736 6199
rect 19794 6196 19800 6248
rect 19852 6236 19858 6248
rect 21100 6236 21128 6276
rect 21266 6264 21272 6276
rect 21324 6304 21330 6316
rect 21453 6307 21511 6313
rect 21453 6304 21465 6307
rect 21324 6276 21465 6304
rect 21324 6264 21330 6276
rect 21453 6273 21465 6276
rect 21499 6273 21511 6307
rect 21453 6267 21511 6273
rect 19852 6208 21128 6236
rect 21177 6239 21235 6245
rect 19852 6196 19858 6208
rect 21177 6205 21189 6239
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 18095 6140 18736 6168
rect 18877 6171 18935 6177
rect 18095 6137 18107 6140
rect 18049 6131 18107 6137
rect 18877 6137 18889 6171
rect 18923 6137 18935 6171
rect 18877 6131 18935 6137
rect 18969 6171 19027 6177
rect 18969 6137 18981 6171
rect 19015 6137 19027 6171
rect 18969 6131 19027 6137
rect 16209 6103 16267 6109
rect 16209 6069 16221 6103
rect 16255 6069 16267 6103
rect 16209 6063 16267 6069
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 18892 6100 18920 6131
rect 18196 6072 18920 6100
rect 18984 6100 19012 6131
rect 20898 6128 20904 6180
rect 20956 6128 20962 6180
rect 20990 6128 20996 6180
rect 21048 6168 21054 6180
rect 21192 6168 21220 6199
rect 21698 6171 21756 6177
rect 21698 6168 21710 6171
rect 21048 6140 21220 6168
rect 21284 6140 21710 6168
rect 21048 6128 21054 6140
rect 19058 6100 19064 6112
rect 18984 6072 19064 6100
rect 18196 6060 18202 6072
rect 19058 6060 19064 6072
rect 19116 6060 19122 6112
rect 19245 6103 19303 6109
rect 19245 6069 19257 6103
rect 19291 6100 19303 6103
rect 21284 6100 21312 6140
rect 21698 6137 21710 6140
rect 21744 6137 21756 6171
rect 21698 6131 21756 6137
rect 19291 6072 21312 6100
rect 21361 6103 21419 6109
rect 19291 6069 19303 6072
rect 19245 6063 19303 6069
rect 21361 6069 21373 6103
rect 21407 6100 21419 6103
rect 21542 6100 21548 6112
rect 21407 6072 21548 6100
rect 21407 6069 21419 6072
rect 21361 6063 21419 6069
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 552 6010 23368 6032
rect 552 5958 4366 6010
rect 4418 5958 4430 6010
rect 4482 5958 4494 6010
rect 4546 5958 4558 6010
rect 4610 5958 4622 6010
rect 4674 5958 4686 6010
rect 4738 5958 10366 6010
rect 10418 5958 10430 6010
rect 10482 5958 10494 6010
rect 10546 5958 10558 6010
rect 10610 5958 10622 6010
rect 10674 5958 10686 6010
rect 10738 5958 16366 6010
rect 16418 5958 16430 6010
rect 16482 5958 16494 6010
rect 16546 5958 16558 6010
rect 16610 5958 16622 6010
rect 16674 5958 16686 6010
rect 16738 5958 22366 6010
rect 22418 5958 22430 6010
rect 22482 5958 22494 6010
rect 22546 5958 22558 6010
rect 22610 5958 22622 6010
rect 22674 5958 22686 6010
rect 22738 5958 23368 6010
rect 552 5936 23368 5958
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 3786 5896 3792 5908
rect 2004 5868 3792 5896
rect 2004 5856 2010 5868
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 6730 5896 6736 5908
rect 5500 5868 6736 5896
rect 5500 5856 5506 5868
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 7190 5896 7196 5908
rect 7064 5868 7196 5896
rect 7064 5856 7070 5868
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 8113 5899 8171 5905
rect 8113 5865 8125 5899
rect 8159 5896 8171 5899
rect 8202 5896 8208 5908
rect 8159 5868 8208 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8386 5856 8392 5908
rect 8444 5856 8450 5908
rect 8481 5899 8539 5905
rect 8481 5865 8493 5899
rect 8527 5896 8539 5899
rect 8570 5896 8576 5908
rect 8527 5868 8576 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9674 5896 9680 5908
rect 8680 5868 9680 5896
rect 2038 5788 2044 5840
rect 2096 5788 2102 5840
rect 2332 5800 2774 5828
rect 842 5720 848 5772
rect 900 5760 906 5772
rect 2332 5769 2360 5800
rect 2317 5763 2375 5769
rect 2317 5760 2329 5763
rect 900 5732 2329 5760
rect 900 5720 906 5732
rect 2317 5729 2329 5732
rect 2363 5729 2375 5763
rect 2317 5723 2375 5729
rect 2406 5720 2412 5772
rect 2464 5760 2470 5772
rect 2573 5763 2631 5769
rect 2573 5760 2585 5763
rect 2464 5732 2585 5760
rect 2464 5720 2470 5732
rect 2573 5729 2585 5732
rect 2619 5729 2631 5763
rect 2746 5760 2774 5800
rect 5828 5800 6500 5828
rect 4982 5760 4988 5772
rect 2746 5732 4988 5760
rect 2573 5723 2631 5729
rect 4982 5720 4988 5732
rect 5040 5760 5046 5772
rect 5828 5769 5856 5800
rect 6472 5772 6500 5800
rect 6638 5788 6644 5840
rect 6696 5828 6702 5840
rect 8021 5831 8079 5837
rect 8021 5828 8033 5831
rect 6696 5800 8033 5828
rect 6696 5788 6702 5800
rect 8021 5797 8033 5800
rect 8067 5828 8079 5831
rect 8680 5828 8708 5868
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 11606 5856 11612 5908
rect 11664 5856 11670 5908
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12250 5896 12256 5908
rect 12124 5868 12256 5896
rect 12124 5856 12130 5868
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12526 5856 12532 5908
rect 12584 5856 12590 5908
rect 12802 5856 12808 5908
rect 12860 5856 12866 5908
rect 14918 5896 14924 5908
rect 14016 5868 14924 5896
rect 8067 5800 8708 5828
rect 9048 5800 11376 5828
rect 8067 5797 8079 5800
rect 8021 5791 8079 5797
rect 9048 5772 9076 5800
rect 5813 5763 5871 5769
rect 5813 5760 5825 5763
rect 5040 5732 5825 5760
rect 5040 5720 5046 5732
rect 5813 5729 5825 5732
rect 5859 5729 5871 5763
rect 5813 5723 5871 5729
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 6069 5763 6127 5769
rect 6069 5760 6081 5763
rect 5960 5732 6081 5760
rect 5960 5720 5966 5732
rect 6069 5729 6081 5732
rect 6115 5729 6127 5763
rect 6069 5723 6127 5729
rect 6454 5720 6460 5772
rect 6512 5720 6518 5772
rect 7098 5720 7104 5772
rect 7156 5720 7162 5772
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5760 7619 5763
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 7607 5732 7849 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 7837 5729 7849 5732
rect 7883 5729 7895 5763
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 7837 5723 7895 5729
rect 7944 5732 8217 5760
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 3384 5664 5028 5692
rect 3384 5652 3390 5664
rect 2056 5596 2360 5624
rect 2056 5565 2084 5596
rect 2041 5559 2099 5565
rect 2041 5525 2053 5559
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 2222 5516 2228 5568
rect 2280 5516 2286 5568
rect 2332 5556 2360 5596
rect 3620 5596 4936 5624
rect 3620 5556 3648 5596
rect 2332 5528 3648 5556
rect 3694 5516 3700 5568
rect 3752 5516 3758 5568
rect 4908 5565 4936 5596
rect 4893 5559 4951 5565
rect 4893 5525 4905 5559
rect 4939 5525 4951 5559
rect 5000 5556 5028 5664
rect 5074 5652 5080 5704
rect 5132 5652 5138 5704
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 5184 5624 5212 5655
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5692 5411 5695
rect 5718 5692 5724 5704
rect 5399 5664 5724 5692
rect 5399 5661 5411 5664
rect 5353 5655 5411 5661
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 5626 5624 5632 5636
rect 5184 5596 5632 5624
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 7116 5624 7144 5720
rect 7576 5692 7604 5723
rect 7944 5704 7972 5732
rect 8205 5729 8217 5732
rect 8251 5760 8263 5763
rect 8665 5763 8723 5769
rect 8665 5760 8677 5763
rect 8251 5732 8677 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8665 5729 8677 5732
rect 8711 5729 8723 5763
rect 9030 5758 9036 5772
rect 8665 5723 8723 5729
rect 8864 5730 9036 5758
rect 6748 5596 7144 5624
rect 7208 5664 7604 5692
rect 6748 5556 6776 5596
rect 7208 5568 7236 5664
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8864 5701 8892 5730
rect 9030 5720 9036 5730
rect 9088 5720 9094 5772
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5760 9183 5763
rect 9306 5760 9312 5772
rect 9171 5732 9312 5760
rect 9171 5729 9183 5732
rect 9125 5723 9183 5729
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 9582 5720 9588 5772
rect 9640 5720 9646 5772
rect 10134 5720 10140 5772
rect 10192 5760 10198 5772
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 10192 5732 10793 5760
rect 10192 5720 10198 5732
rect 10781 5729 10793 5732
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 10870 5720 10876 5772
rect 10928 5720 10934 5772
rect 10962 5720 10968 5772
rect 11020 5720 11026 5772
rect 11348 5769 11376 5800
rect 11514 5788 11520 5840
rect 11572 5828 11578 5840
rect 11974 5828 11980 5840
rect 11572 5800 11980 5828
rect 11572 5788 11578 5800
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5729 11207 5763
rect 11149 5723 11207 5729
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11241 5723 11299 5729
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 8757 5695 8815 5701
rect 8757 5692 8769 5695
rect 8444 5664 8769 5692
rect 8444 5652 8450 5664
rect 8757 5661 8769 5664
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 8849 5695 8907 5701
rect 8849 5661 8861 5695
rect 8895 5661 8907 5695
rect 8849 5655 8907 5661
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 7745 5627 7803 5633
rect 7745 5593 7757 5627
rect 7791 5624 7803 5627
rect 8956 5624 8984 5655
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 9600 5692 9628 5720
rect 9272 5664 9628 5692
rect 10888 5692 10916 5720
rect 11164 5692 11192 5723
rect 10888 5664 11192 5692
rect 9272 5652 9278 5664
rect 11146 5624 11152 5636
rect 7791 5596 11152 5624
rect 7791 5593 7803 5596
rect 7745 5587 7803 5593
rect 11146 5584 11152 5596
rect 11204 5584 11210 5636
rect 5000 5528 6776 5556
rect 4893 5519 4951 5525
rect 7190 5516 7196 5568
rect 7248 5516 7254 5568
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 9030 5556 9036 5568
rect 7984 5528 9036 5556
rect 7984 5516 7990 5528
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 10597 5559 10655 5565
rect 10597 5525 10609 5559
rect 10643 5556 10655 5559
rect 10778 5556 10784 5568
rect 10643 5528 10784 5556
rect 10643 5525 10655 5528
rect 10597 5519 10655 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 11256 5556 11284 5723
rect 11790 5720 11796 5772
rect 11848 5760 11854 5772
rect 12253 5763 12311 5769
rect 12253 5760 12265 5763
rect 11848 5732 12265 5760
rect 11848 5720 11854 5732
rect 12253 5729 12265 5732
rect 12299 5729 12311 5763
rect 12253 5723 12311 5729
rect 12437 5763 12495 5769
rect 12437 5729 12449 5763
rect 12483 5760 12495 5763
rect 12544 5760 12572 5856
rect 12820 5828 12848 5856
rect 14016 5840 14044 5868
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15010 5856 15016 5908
rect 15068 5896 15074 5908
rect 15473 5899 15531 5905
rect 15473 5896 15485 5899
rect 15068 5868 15485 5896
rect 15068 5856 15074 5868
rect 15473 5865 15485 5868
rect 15519 5865 15531 5899
rect 15473 5859 15531 5865
rect 15930 5856 15936 5908
rect 15988 5856 15994 5908
rect 17034 5856 17040 5908
rect 17092 5896 17098 5908
rect 17586 5896 17592 5908
rect 17092 5868 17592 5896
rect 17092 5856 17098 5868
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 17681 5899 17739 5905
rect 17681 5865 17693 5899
rect 17727 5896 17739 5899
rect 17954 5896 17960 5908
rect 17727 5868 17960 5896
rect 17727 5865 17739 5868
rect 17681 5859 17739 5865
rect 17954 5856 17960 5868
rect 18012 5856 18018 5908
rect 18877 5899 18935 5905
rect 18877 5865 18889 5899
rect 18923 5896 18935 5899
rect 21085 5899 21143 5905
rect 18923 5868 19472 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 13998 5828 14004 5840
rect 12820 5800 14004 5828
rect 12483 5732 12572 5760
rect 12483 5729 12495 5732
rect 12437 5723 12495 5729
rect 12710 5720 12716 5772
rect 12768 5720 12774 5772
rect 12175 5695 12233 5701
rect 12175 5661 12187 5695
rect 12221 5661 12233 5695
rect 12175 5655 12233 5661
rect 12176 5624 12204 5655
rect 12342 5652 12348 5704
rect 12400 5652 12406 5704
rect 12820 5692 12848 5800
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 15746 5828 15752 5840
rect 14936 5800 15752 5828
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 13170 5760 13176 5772
rect 12943 5732 13176 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13170 5720 13176 5732
rect 13228 5720 13234 5772
rect 13262 5720 13268 5772
rect 13320 5720 13326 5772
rect 13449 5763 13507 5769
rect 13449 5729 13461 5763
rect 13495 5760 13507 5763
rect 13725 5763 13783 5769
rect 13725 5760 13737 5763
rect 13495 5732 13737 5760
rect 13495 5729 13507 5732
rect 13449 5723 13507 5729
rect 13725 5729 13737 5732
rect 13771 5729 13783 5763
rect 14936 5760 14964 5800
rect 15746 5788 15752 5800
rect 15804 5788 15810 5840
rect 13725 5723 13783 5729
rect 13832 5732 14964 5760
rect 12989 5695 13047 5701
rect 12989 5692 13001 5695
rect 12820 5664 13001 5692
rect 12989 5661 13001 5664
rect 13035 5661 13047 5695
rect 12989 5655 13047 5661
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13832 5692 13860 5732
rect 15010 5720 15016 5772
rect 15068 5720 15074 5772
rect 15381 5763 15439 5769
rect 15381 5729 15393 5763
rect 15427 5760 15439 5763
rect 15562 5760 15568 5772
rect 15427 5732 15568 5760
rect 15427 5729 15439 5732
rect 15381 5723 15439 5729
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 15948 5760 15976 5856
rect 16868 5800 17172 5828
rect 16868 5772 16896 5800
rect 15703 5732 15976 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 16850 5720 16856 5772
rect 16908 5720 16914 5772
rect 17034 5720 17040 5772
rect 17092 5720 17098 5772
rect 17144 5769 17172 5800
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 18509 5831 18567 5837
rect 17276 5800 18460 5828
rect 17276 5788 17282 5800
rect 17129 5763 17187 5769
rect 17129 5729 17141 5763
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17773 5763 17831 5769
rect 17773 5729 17785 5763
rect 17819 5760 17831 5763
rect 18049 5763 18107 5769
rect 18049 5760 18061 5763
rect 17819 5732 18061 5760
rect 17819 5729 17831 5732
rect 17773 5723 17831 5729
rect 18049 5729 18061 5732
rect 18095 5729 18107 5763
rect 18049 5723 18107 5729
rect 13127 5664 13860 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14001 5695 14059 5701
rect 14001 5692 14013 5695
rect 13964 5664 14013 5692
rect 13964 5652 13970 5664
rect 14001 5661 14013 5664
rect 14047 5661 14059 5695
rect 14001 5655 14059 5661
rect 14642 5652 14648 5704
rect 14700 5652 14706 5704
rect 14918 5652 14924 5704
rect 14976 5652 14982 5704
rect 15028 5692 15056 5720
rect 17604 5692 17632 5723
rect 15028 5664 17632 5692
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 12176 5596 13553 5624
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 13541 5587 13599 5593
rect 12526 5556 12532 5568
rect 11256 5528 12532 5556
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 12621 5559 12679 5565
rect 12621 5525 12633 5559
rect 12667 5556 12679 5559
rect 13170 5556 13176 5568
rect 12667 5528 13176 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 14458 5556 14464 5568
rect 13955 5528 14464 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 14458 5516 14464 5528
rect 14516 5556 14522 5568
rect 14660 5556 14688 5652
rect 14936 5624 14964 5652
rect 14936 5596 15332 5624
rect 14516 5528 14688 5556
rect 14516 5516 14522 5528
rect 15194 5516 15200 5568
rect 15252 5516 15258 5568
rect 15304 5556 15332 5596
rect 17218 5584 17224 5636
rect 17276 5584 17282 5636
rect 16850 5556 16856 5568
rect 15304 5528 16856 5556
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 17236 5556 17264 5584
rect 17313 5559 17371 5565
rect 17313 5556 17325 5559
rect 17236 5528 17325 5556
rect 17313 5525 17325 5528
rect 17359 5525 17371 5559
rect 17604 5556 17632 5664
rect 17862 5652 17868 5704
rect 17920 5652 17926 5704
rect 18064 5624 18092 5723
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 18196 5732 18337 5760
rect 18196 5720 18202 5732
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18432 5760 18460 5800
rect 18509 5797 18521 5831
rect 18555 5828 18567 5831
rect 19061 5831 19119 5837
rect 19061 5828 19073 5831
rect 18555 5800 19073 5828
rect 18555 5797 18567 5800
rect 18509 5791 18567 5797
rect 19061 5797 19073 5800
rect 19107 5797 19119 5831
rect 19444 5828 19472 5868
rect 21085 5865 21097 5899
rect 21131 5896 21143 5899
rect 21131 5868 21588 5896
rect 21131 5865 21143 5868
rect 21085 5859 21143 5865
rect 19950 5831 20008 5837
rect 19950 5828 19962 5831
rect 19444 5800 19962 5828
rect 19061 5791 19119 5797
rect 19950 5797 19962 5800
rect 19996 5797 20008 5831
rect 19950 5791 20008 5797
rect 21560 5828 21588 5868
rect 22094 5856 22100 5908
rect 22152 5856 22158 5908
rect 21560 5800 22232 5828
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 18432 5732 18613 5760
rect 18325 5723 18383 5729
rect 18601 5729 18613 5732
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5760 18751 5763
rect 18782 5760 18788 5772
rect 18739 5732 18788 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 18782 5720 18788 5732
rect 18840 5720 18846 5772
rect 18874 5720 18880 5772
rect 18932 5760 18938 5772
rect 18969 5763 19027 5769
rect 18969 5760 18981 5763
rect 18932 5732 18981 5760
rect 18932 5720 18938 5732
rect 18969 5729 18981 5732
rect 19015 5729 19027 5763
rect 18969 5723 19027 5729
rect 19150 5720 19156 5772
rect 19208 5720 19214 5772
rect 19705 5763 19763 5769
rect 19705 5729 19717 5763
rect 19751 5760 19763 5763
rect 19794 5760 19800 5772
rect 19751 5732 19800 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 21560 5769 21588 5800
rect 21545 5763 21603 5769
rect 21545 5729 21557 5763
rect 21591 5729 21603 5763
rect 21545 5723 21603 5729
rect 21818 5720 21824 5772
rect 21876 5720 21882 5772
rect 21910 5720 21916 5772
rect 21968 5720 21974 5772
rect 22204 5769 22232 5800
rect 22189 5763 22247 5769
rect 22189 5729 22201 5763
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 18892 5624 18920 5720
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5692 21511 5695
rect 21836 5692 21864 5720
rect 21499 5664 21864 5692
rect 21499 5661 21511 5664
rect 21453 5655 21511 5661
rect 18064 5596 18920 5624
rect 21358 5584 21364 5636
rect 21416 5624 21422 5636
rect 21726 5624 21732 5636
rect 21416 5596 21732 5624
rect 21416 5584 21422 5596
rect 21726 5584 21732 5596
rect 21784 5624 21790 5636
rect 22373 5627 22431 5633
rect 22373 5624 22385 5627
rect 21784 5596 22385 5624
rect 21784 5584 21790 5596
rect 22373 5593 22385 5596
rect 22419 5593 22431 5627
rect 22373 5587 22431 5593
rect 19058 5556 19064 5568
rect 17604 5528 19064 5556
rect 17313 5519 17371 5525
rect 19058 5516 19064 5528
rect 19116 5516 19122 5568
rect 21913 5559 21971 5565
rect 21913 5525 21925 5559
rect 21959 5556 21971 5559
rect 22094 5556 22100 5568
rect 21959 5528 22100 5556
rect 21959 5525 21971 5528
rect 21913 5519 21971 5525
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 552 5466 23368 5488
rect 552 5414 1366 5466
rect 1418 5414 1430 5466
rect 1482 5414 1494 5466
rect 1546 5414 1558 5466
rect 1610 5414 1622 5466
rect 1674 5414 1686 5466
rect 1738 5414 7366 5466
rect 7418 5414 7430 5466
rect 7482 5414 7494 5466
rect 7546 5414 7558 5466
rect 7610 5414 7622 5466
rect 7674 5414 7686 5466
rect 7738 5414 13366 5466
rect 13418 5414 13430 5466
rect 13482 5414 13494 5466
rect 13546 5414 13558 5466
rect 13610 5414 13622 5466
rect 13674 5414 13686 5466
rect 13738 5414 19366 5466
rect 19418 5414 19430 5466
rect 19482 5414 19494 5466
rect 19546 5414 19558 5466
rect 19610 5414 19622 5466
rect 19674 5414 19686 5466
rect 19738 5414 23368 5466
rect 552 5392 23368 5414
rect 1762 5312 1768 5364
rect 1820 5312 1826 5364
rect 5353 5355 5411 5361
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 5902 5352 5908 5364
rect 5399 5324 5908 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 6595 5355 6653 5361
rect 6595 5321 6607 5355
rect 6641 5352 6653 5355
rect 6914 5352 6920 5364
rect 6641 5324 6920 5352
rect 6641 5321 6653 5324
rect 6595 5315 6653 5321
rect 6914 5312 6920 5324
rect 6972 5352 6978 5364
rect 7926 5352 7932 5364
rect 6972 5324 7932 5352
rect 6972 5312 6978 5324
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8294 5312 8300 5364
rect 8352 5312 8358 5364
rect 8570 5312 8576 5364
rect 8628 5352 8634 5364
rect 9306 5352 9312 5364
rect 8628 5324 9312 5352
rect 8628 5312 8634 5324
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 11054 5352 11060 5364
rect 10980 5324 11060 5352
rect 1780 5216 1808 5312
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 2774 5284 2780 5296
rect 2179 5256 2780 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 8312 5284 8340 5312
rect 5184 5256 8340 5284
rect 10980 5284 11008 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11698 5352 11704 5364
rect 11204 5324 11704 5352
rect 11204 5312 11210 5324
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 12345 5355 12403 5361
rect 12345 5352 12357 5355
rect 11848 5324 12357 5352
rect 11848 5312 11854 5324
rect 12345 5321 12357 5324
rect 12391 5321 12403 5355
rect 12345 5315 12403 5321
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 14826 5352 14832 5364
rect 13780 5324 14832 5352
rect 13780 5312 13786 5324
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 15746 5352 15752 5364
rect 15620 5324 15752 5352
rect 15620 5312 15626 5324
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16206 5312 16212 5364
rect 16264 5352 16270 5364
rect 17586 5352 17592 5364
rect 16264 5324 17592 5352
rect 16264 5312 16270 5324
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 18509 5355 18567 5361
rect 18509 5321 18521 5355
rect 18555 5352 18567 5355
rect 19150 5352 19156 5364
rect 18555 5324 19156 5352
rect 18555 5321 18567 5324
rect 18509 5315 18567 5321
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 21085 5355 21143 5361
rect 21085 5352 21097 5355
rect 20956 5324 21097 5352
rect 20956 5312 20962 5324
rect 21085 5321 21097 5324
rect 21131 5321 21143 5355
rect 21085 5315 21143 5321
rect 21453 5355 21511 5361
rect 21453 5321 21465 5355
rect 21499 5352 21511 5355
rect 21542 5352 21548 5364
rect 21499 5324 21548 5352
rect 21499 5321 21511 5324
rect 21453 5315 21511 5321
rect 21542 5312 21548 5324
rect 21600 5312 21606 5364
rect 21634 5312 21640 5364
rect 21692 5352 21698 5364
rect 22005 5355 22063 5361
rect 22005 5352 22017 5355
rect 21692 5324 22017 5352
rect 21692 5312 21698 5324
rect 22005 5321 22017 5324
rect 22051 5321 22063 5355
rect 22005 5315 22063 5321
rect 11330 5284 11336 5296
rect 10980 5256 11336 5284
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1780 5188 1961 5216
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 4801 5219 4859 5225
rect 2372 5188 2544 5216
rect 2372 5176 2378 5188
rect 2222 5108 2228 5160
rect 2280 5148 2286 5160
rect 2516 5157 2544 5188
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 5074 5216 5080 5228
rect 4847 5188 5080 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5184 5157 5212 5256
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5684 5188 5733 5216
rect 5684 5176 5690 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5216 6423 5219
rect 6638 5216 6644 5228
rect 6411 5188 6644 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 2501 5151 2559 5157
rect 2280 5120 2452 5148
rect 2280 5108 2286 5120
rect 2424 5080 2452 5120
rect 2501 5117 2513 5151
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5117 4583 5151
rect 4525 5111 4583 5117
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 4540 5080 4568 5111
rect 5442 5108 5448 5160
rect 5500 5108 5506 5160
rect 5736 5148 5764 5179
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 7708 5188 8432 5216
rect 7708 5176 7714 5188
rect 8404 5157 8432 5188
rect 7561 5151 7619 5157
rect 5736 5120 6868 5148
rect 2424 5052 6132 5080
rect 6104 5024 6132 5052
rect 6840 5024 6868 5120
rect 7561 5117 7573 5151
rect 7607 5148 7619 5151
rect 8389 5151 8447 5157
rect 7607 5120 8340 5148
rect 7607 5117 7619 5120
rect 7561 5111 7619 5117
rect 1946 4972 1952 5024
rect 2004 4972 2010 5024
rect 2314 4972 2320 5024
rect 2372 4972 2378 5024
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 5810 5012 5816 5024
rect 3568 4984 5816 5012
rect 3568 4972 3574 4984
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6086 4972 6092 5024
rect 6144 4972 6150 5024
rect 6822 4972 6828 5024
rect 6880 4972 6886 5024
rect 7926 4972 7932 5024
rect 7984 4972 7990 5024
rect 8312 5012 8340 5120
rect 8389 5117 8401 5151
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 8662 5108 8668 5160
rect 8720 5108 8726 5160
rect 9214 5108 9220 5160
rect 9272 5108 9278 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 10980 5157 11008 5256
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 11882 5284 11888 5296
rect 11532 5256 11888 5284
rect 11057 5219 11115 5225
rect 11057 5185 11069 5219
rect 11103 5216 11115 5219
rect 11532 5216 11560 5256
rect 11882 5244 11888 5256
rect 11940 5284 11946 5296
rect 11940 5256 17264 5284
rect 11940 5244 11946 5256
rect 17236 5228 17264 5256
rect 18064 5256 18552 5284
rect 11103 5188 11560 5216
rect 11103 5185 11115 5188
rect 11057 5179 11115 5185
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 9456 5120 10333 5148
rect 9456 5108 9462 5120
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 10735 5120 10793 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 10781 5117 10793 5120
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 10965 5151 11023 5157
rect 10965 5117 10977 5151
rect 11011 5117 11023 5151
rect 10965 5111 11023 5117
rect 11146 5108 11152 5160
rect 11204 5108 11210 5160
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 11422 5148 11428 5160
rect 11379 5120 11428 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 11532 5148 11560 5188
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 15378 5216 15384 5228
rect 12544 5188 14780 5216
rect 12544 5160 12572 5188
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 11532 5120 11805 5148
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 11885 5151 11943 5157
rect 11885 5117 11897 5151
rect 11931 5117 11943 5151
rect 11885 5111 11943 5117
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 9232 5080 9260 5108
rect 8527 5052 9260 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 10008 5052 10517 5080
rect 10008 5040 10014 5052
rect 10505 5049 10517 5052
rect 10551 5080 10563 5083
rect 11606 5080 11612 5092
rect 10551 5052 11612 5080
rect 10551 5049 10563 5052
rect 10505 5043 10563 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 11900 5080 11928 5111
rect 11974 5108 11980 5160
rect 12032 5108 12038 5160
rect 12158 5108 12164 5160
rect 12216 5108 12222 5160
rect 12434 5108 12440 5160
rect 12492 5108 12498 5160
rect 12526 5108 12532 5160
rect 12584 5108 12590 5160
rect 12618 5108 12624 5160
rect 12676 5108 12682 5160
rect 12728 5157 12756 5188
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5117 12771 5151
rect 12713 5111 12771 5117
rect 12802 5108 12808 5160
rect 12860 5108 12866 5160
rect 12989 5151 13047 5157
rect 12989 5117 13001 5151
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 11716 5052 11928 5080
rect 12176 5080 12204 5108
rect 12452 5080 12480 5108
rect 13004 5080 13032 5111
rect 12176 5052 12388 5080
rect 12452 5052 13032 5080
rect 13556 5080 13584 5111
rect 13630 5108 13636 5160
rect 13688 5148 13694 5160
rect 13814 5148 13820 5160
rect 13688 5120 13820 5148
rect 13688 5108 13694 5120
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14182 5108 14188 5160
rect 14240 5108 14246 5160
rect 14200 5080 14228 5108
rect 14550 5080 14556 5092
rect 13556 5052 14556 5080
rect 11716 5024 11744 5052
rect 8570 5012 8576 5024
rect 8312 4984 8576 5012
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 8849 5015 8907 5021
rect 8849 4981 8861 5015
rect 8895 5012 8907 5015
rect 9030 5012 9036 5024
rect 8895 4984 9036 5012
rect 8895 4981 8907 4984
rect 8849 4975 8907 4981
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 11698 4972 11704 5024
rect 11756 4972 11762 5024
rect 12158 4972 12164 5024
rect 12216 4972 12222 5024
rect 12360 5012 12388 5052
rect 14550 5040 14556 5052
rect 14608 5040 14614 5092
rect 13170 5012 13176 5024
rect 12360 4984 13176 5012
rect 13170 4972 13176 4984
rect 13228 4972 13234 5024
rect 14752 5021 14780 5188
rect 14936 5188 15384 5216
rect 14936 5157 14964 5188
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15528 5188 15853 5216
rect 15528 5176 15534 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15930 5176 15936 5228
rect 15988 5176 15994 5228
rect 16022 5176 16028 5228
rect 16080 5216 16086 5228
rect 16206 5216 16212 5228
rect 16080 5188 16212 5216
rect 16080 5176 16086 5188
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 17218 5176 17224 5228
rect 17276 5176 17282 5228
rect 14921 5151 14979 5157
rect 14921 5117 14933 5151
rect 14967 5117 14979 5151
rect 14921 5111 14979 5117
rect 15194 5108 15200 5160
rect 15252 5108 15258 5160
rect 15289 5151 15347 5157
rect 15289 5117 15301 5151
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 15565 5151 15623 5157
rect 15565 5117 15577 5151
rect 15611 5148 15623 5151
rect 15654 5148 15660 5160
rect 15611 5120 15660 5148
rect 15611 5117 15623 5120
rect 15565 5111 15623 5117
rect 14826 5040 14832 5092
rect 14884 5080 14890 5092
rect 15304 5080 15332 5111
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 17034 5108 17040 5160
rect 17092 5148 17098 5160
rect 17681 5151 17739 5157
rect 17681 5148 17693 5151
rect 17092 5120 17693 5148
rect 17092 5108 17098 5120
rect 17681 5117 17693 5120
rect 17727 5148 17739 5151
rect 18064 5148 18092 5256
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5216 18199 5219
rect 18524 5216 18552 5256
rect 18874 5244 18880 5296
rect 18932 5244 18938 5296
rect 20346 5244 20352 5296
rect 20404 5284 20410 5296
rect 21652 5284 21680 5312
rect 20404 5256 21680 5284
rect 20404 5244 20410 5256
rect 21545 5219 21603 5225
rect 21545 5216 21557 5219
rect 18187 5188 18460 5216
rect 18524 5188 21557 5216
rect 18187 5185 18199 5188
rect 18141 5179 18199 5185
rect 18432 5160 18460 5188
rect 21545 5185 21557 5188
rect 21591 5185 21603 5219
rect 21545 5179 21603 5185
rect 22094 5176 22100 5228
rect 22152 5176 22158 5228
rect 18230 5148 18236 5160
rect 17727 5120 18236 5148
rect 17727 5117 17739 5120
rect 17681 5111 17739 5117
rect 18230 5108 18236 5120
rect 18288 5108 18294 5160
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5117 18383 5151
rect 18325 5111 18383 5117
rect 18340 5080 18368 5111
rect 18414 5108 18420 5160
rect 18472 5148 18478 5160
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18472 5120 18705 5148
rect 18472 5108 18478 5120
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18877 5151 18935 5157
rect 18877 5117 18889 5151
rect 18923 5148 18935 5151
rect 20346 5148 20352 5160
rect 18923 5120 20352 5148
rect 18923 5117 18935 5120
rect 18877 5111 18935 5117
rect 18892 5080 18920 5111
rect 20346 5108 20352 5120
rect 20404 5108 20410 5160
rect 21358 5108 21364 5160
rect 21416 5108 21422 5160
rect 21450 5108 21456 5160
rect 21508 5108 21514 5160
rect 21729 5151 21787 5157
rect 21729 5117 21741 5151
rect 21775 5148 21787 5151
rect 21818 5148 21824 5160
rect 21775 5120 21824 5148
rect 21775 5117 21787 5120
rect 21729 5111 21787 5117
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 21910 5108 21916 5160
rect 21968 5108 21974 5160
rect 22112 5147 22140 5176
rect 22097 5141 22155 5147
rect 22097 5107 22109 5141
rect 22143 5107 22155 5141
rect 22097 5101 22155 5107
rect 14884 5052 18000 5080
rect 18340 5052 18920 5080
rect 14884 5040 14890 5052
rect 14737 5015 14795 5021
rect 14737 4981 14749 5015
rect 14783 5012 14795 5015
rect 14918 5012 14924 5024
rect 14783 4984 14924 5012
rect 14783 4981 14795 4984
rect 14737 4975 14795 4981
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 15013 5015 15071 5021
rect 15013 4981 15025 5015
rect 15059 5012 15071 5015
rect 15194 5012 15200 5024
rect 15059 4984 15200 5012
rect 15059 4981 15071 4984
rect 15013 4975 15071 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15654 4972 15660 5024
rect 15712 4972 15718 5024
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16850 5012 16856 5024
rect 16347 4984 16856 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17862 4972 17868 5024
rect 17920 4972 17926 5024
rect 17972 5012 18000 5052
rect 19978 5040 19984 5092
rect 20036 5080 20042 5092
rect 21082 5080 21088 5092
rect 20036 5052 21088 5080
rect 20036 5040 20042 5052
rect 21082 5040 21088 5052
rect 21140 5040 21146 5092
rect 21542 5012 21548 5024
rect 17972 4984 21548 5012
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 552 4922 23368 4944
rect 552 4870 4366 4922
rect 4418 4870 4430 4922
rect 4482 4870 4494 4922
rect 4546 4870 4558 4922
rect 4610 4870 4622 4922
rect 4674 4870 4686 4922
rect 4738 4870 10366 4922
rect 10418 4870 10430 4922
rect 10482 4870 10494 4922
rect 10546 4870 10558 4922
rect 10610 4870 10622 4922
rect 10674 4870 10686 4922
rect 10738 4870 16366 4922
rect 16418 4870 16430 4922
rect 16482 4870 16494 4922
rect 16546 4870 16558 4922
rect 16610 4870 16622 4922
rect 16674 4870 16686 4922
rect 16738 4870 22366 4922
rect 22418 4870 22430 4922
rect 22482 4870 22494 4922
rect 22546 4870 22558 4922
rect 22610 4870 22622 4922
rect 22674 4870 22686 4922
rect 22738 4870 23368 4922
rect 552 4848 23368 4870
rect 2314 4768 2320 4820
rect 2372 4768 2378 4820
rect 2682 4768 2688 4820
rect 2740 4768 2746 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 4154 4808 4160 4820
rect 3467 4780 4160 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 4154 4768 4160 4780
rect 4212 4808 4218 4820
rect 5442 4808 5448 4820
rect 4212 4780 5448 4808
rect 4212 4768 4218 4780
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5537 4811 5595 4817
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 6638 4808 6644 4820
rect 5583 4780 6644 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 8662 4808 8668 4820
rect 7791 4780 8668 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 11885 4811 11943 4817
rect 9456 4780 11560 4808
rect 9456 4768 9462 4780
rect 1572 4743 1630 4749
rect 1572 4709 1584 4743
rect 1618 4740 1630 4743
rect 2332 4740 2360 4768
rect 1618 4712 2360 4740
rect 1618 4709 1630 4712
rect 1572 4703 1630 4709
rect 3694 4700 3700 4752
rect 3752 4740 3758 4752
rect 3752 4712 6040 4740
rect 3752 4700 3758 4712
rect 842 4632 848 4684
rect 900 4672 906 4684
rect 1305 4675 1363 4681
rect 1305 4672 1317 4675
rect 900 4644 1317 4672
rect 900 4632 906 4644
rect 1305 4641 1317 4644
rect 1351 4641 1363 4675
rect 1305 4635 1363 4641
rect 3602 4632 3608 4684
rect 3660 4632 3666 4684
rect 4338 4632 4344 4684
rect 4396 4672 4402 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4396 4644 4813 4672
rect 4396 4632 4402 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 5353 4675 5411 4681
rect 5353 4641 5365 4675
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 3697 4607 3755 4613
rect 3697 4573 3709 4607
rect 3743 4604 3755 4607
rect 3786 4604 3792 4616
rect 3743 4576 3792 4604
rect 3743 4573 3755 4576
rect 3697 4567 3755 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 3988 4536 4016 4567
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 4212 4576 4629 4604
rect 4212 4564 4218 4576
rect 4617 4573 4629 4576
rect 4663 4604 4675 4607
rect 5368 4604 5396 4635
rect 4663 4576 5396 4604
rect 4663 4573 4675 4576
rect 4617 4567 4675 4573
rect 5828 4536 5856 4635
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 6012 4604 6040 4712
rect 6086 4700 6092 4752
rect 6144 4740 6150 4752
rect 11532 4740 11560 4780
rect 11885 4777 11897 4811
rect 11931 4808 11943 4811
rect 12342 4808 12348 4820
rect 11931 4780 12348 4808
rect 11931 4777 11943 4780
rect 11885 4771 11943 4777
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 13541 4811 13599 4817
rect 13541 4808 13553 4811
rect 12860 4780 13553 4808
rect 12860 4768 12866 4780
rect 13541 4777 13553 4780
rect 13587 4777 13599 4811
rect 13541 4771 13599 4777
rect 14734 4768 14740 4820
rect 14792 4768 14798 4820
rect 16850 4768 16856 4820
rect 16908 4768 16914 4820
rect 18509 4811 18567 4817
rect 18509 4777 18521 4811
rect 18555 4808 18567 4811
rect 20806 4808 20812 4820
rect 18555 4780 20812 4808
rect 18555 4777 18567 4780
rect 18509 4771 18567 4777
rect 20806 4768 20812 4780
rect 20864 4768 20870 4820
rect 21085 4811 21143 4817
rect 21085 4777 21097 4811
rect 21131 4808 21143 4811
rect 21174 4808 21180 4820
rect 21131 4780 21180 4808
rect 21131 4777 21143 4780
rect 21085 4771 21143 4777
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 21910 4768 21916 4820
rect 21968 4808 21974 4820
rect 22278 4808 22284 4820
rect 21968 4780 22284 4808
rect 21968 4768 21974 4780
rect 22278 4768 22284 4780
rect 22336 4808 22342 4820
rect 22649 4811 22707 4817
rect 22649 4808 22661 4811
rect 22336 4780 22661 4808
rect 22336 4768 22342 4780
rect 22649 4777 22661 4780
rect 22695 4777 22707 4811
rect 22649 4771 22707 4777
rect 13906 4740 13912 4752
rect 6144 4712 11100 4740
rect 11532 4712 13912 4740
rect 6144 4700 6150 4712
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7190 4672 7196 4684
rect 6963 4644 7196 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7190 4632 7196 4644
rect 7248 4674 7254 4684
rect 7377 4675 7435 4681
rect 7377 4674 7389 4675
rect 7248 4646 7389 4674
rect 7248 4632 7254 4646
rect 7377 4641 7389 4646
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 7466 4632 7472 4684
rect 7524 4672 7530 4684
rect 7561 4675 7619 4681
rect 7561 4672 7573 4675
rect 7524 4644 7573 4672
rect 7524 4632 7530 4644
rect 7561 4641 7573 4644
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4674 10655 4675
rect 10643 4672 10732 4674
rect 10778 4672 10784 4684
rect 10643 4646 10784 4672
rect 10643 4641 10655 4646
rect 10704 4644 10784 4646
rect 10597 4635 10655 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 11072 4672 11100 4712
rect 11698 4672 11704 4684
rect 11072 4644 11704 4672
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 11882 4632 11888 4684
rect 11940 4632 11946 4684
rect 13078 4632 13084 4684
rect 13136 4632 13142 4684
rect 13740 4681 13768 4712
rect 13906 4700 13912 4712
rect 13964 4700 13970 4752
rect 13998 4700 14004 4752
rect 14056 4700 14062 4752
rect 14752 4740 14780 4768
rect 15930 4740 15936 4752
rect 14752 4712 15936 4740
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4641 13783 4675
rect 13725 4635 13783 4641
rect 13814 4632 13820 4684
rect 13872 4632 13878 4684
rect 14016 4672 14044 4700
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 14016 4644 14105 4672
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 14369 4675 14427 4681
rect 14369 4672 14381 4675
rect 14240 4644 14381 4672
rect 14240 4632 14246 4644
rect 14369 4641 14381 4644
rect 14415 4672 14427 4675
rect 15102 4672 15108 4684
rect 14415 4644 15108 4672
rect 14415 4641 14427 4644
rect 14369 4635 14427 4641
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 15212 4681 15240 4712
rect 15930 4700 15936 4712
rect 15988 4740 15994 4752
rect 15988 4712 16160 4740
rect 15988 4700 15994 4712
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 15378 4632 15384 4684
rect 15436 4632 15442 4684
rect 15562 4632 15568 4684
rect 15620 4632 15626 4684
rect 15746 4632 15752 4684
rect 15804 4632 15810 4684
rect 16132 4681 16160 4712
rect 16206 4700 16212 4752
rect 16264 4740 16270 4752
rect 18049 4743 18107 4749
rect 18049 4740 18061 4743
rect 16264 4712 16528 4740
rect 16264 4700 16270 4712
rect 16500 4681 16528 4712
rect 17788 4712 18061 4740
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 16301 4675 16359 4681
rect 16301 4641 16313 4675
rect 16347 4641 16359 4675
rect 16301 4635 16359 4641
rect 16393 4675 16451 4681
rect 16393 4641 16405 4675
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 16485 4675 16543 4681
rect 16485 4641 16497 4675
rect 16531 4641 16543 4675
rect 16485 4635 16543 4641
rect 16669 4675 16727 4681
rect 16669 4641 16681 4675
rect 16715 4672 16727 4675
rect 17218 4672 17224 4684
rect 16715 4644 17224 4672
rect 16715 4641 16727 4644
rect 16669 4635 16727 4641
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6012 4576 7021 4604
rect 7009 4573 7021 4576
rect 7055 4604 7067 4607
rect 7055 4576 7236 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7208 4548 7236 4576
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 10502 4604 10508 4616
rect 7800 4576 10508 4604
rect 7800 4564 7806 4576
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 11790 4564 11796 4616
rect 11848 4604 11854 4616
rect 11848 4576 12112 4604
rect 11848 4564 11854 4576
rect 6086 4536 6092 4548
rect 3988 4508 5304 4536
rect 5828 4508 6092 4536
rect 5276 4480 5304 4508
rect 6086 4496 6092 4508
rect 6144 4496 6150 4548
rect 7190 4496 7196 4548
rect 7248 4496 7254 4548
rect 7285 4539 7343 4545
rect 7285 4505 7297 4539
rect 7331 4536 7343 4539
rect 7650 4536 7656 4548
rect 7331 4508 7656 4536
rect 7331 4505 7343 4508
rect 7285 4499 7343 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 10781 4539 10839 4545
rect 10781 4505 10793 4539
rect 10827 4536 10839 4539
rect 11974 4536 11980 4548
rect 10827 4508 11980 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 12084 4536 12112 4576
rect 12802 4564 12808 4616
rect 12860 4564 12866 4616
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4604 12955 4607
rect 14001 4607 14059 4613
rect 14001 4604 14013 4607
rect 12943 4576 14013 4604
rect 12943 4573 12955 4576
rect 12897 4567 12955 4573
rect 13096 4548 13124 4576
rect 14001 4573 14013 4576
rect 14047 4604 14059 4607
rect 15286 4604 15292 4616
rect 14047 4576 15292 4604
rect 14047 4573 14059 4576
rect 14001 4567 14059 4573
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4573 15531 4607
rect 16316 4604 16344 4635
rect 15473 4567 15531 4573
rect 15764 4576 16344 4604
rect 16408 4604 16436 4635
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 17788 4604 17816 4712
rect 18049 4709 18061 4712
rect 18095 4740 18107 4743
rect 18230 4740 18236 4752
rect 18095 4712 18236 4740
rect 18095 4709 18107 4712
rect 18049 4703 18107 4709
rect 18230 4700 18236 4712
rect 18288 4740 18294 4752
rect 19794 4740 19800 4752
rect 18288 4712 19800 4740
rect 18288 4700 18294 4712
rect 17862 4632 17868 4684
rect 17920 4672 17926 4684
rect 19536 4681 19564 4712
rect 19794 4700 19800 4712
rect 19852 4700 19858 4752
rect 20438 4740 20444 4752
rect 19904 4712 20444 4740
rect 18325 4675 18383 4681
rect 18325 4672 18337 4675
rect 17920 4644 18337 4672
rect 17920 4632 17926 4644
rect 18325 4641 18337 4644
rect 18371 4641 18383 4675
rect 18325 4635 18383 4641
rect 19061 4675 19119 4681
rect 19061 4641 19073 4675
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 19521 4675 19579 4681
rect 19521 4641 19533 4675
rect 19567 4641 19579 4675
rect 19521 4635 19579 4641
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4672 19671 4675
rect 19904 4672 19932 4712
rect 20438 4700 20444 4712
rect 20496 4700 20502 4752
rect 20625 4743 20683 4749
rect 20625 4709 20637 4743
rect 20671 4740 20683 4743
rect 21634 4740 21640 4752
rect 20671 4712 21640 4740
rect 20671 4709 20683 4712
rect 20625 4703 20683 4709
rect 21634 4700 21640 4712
rect 21692 4700 21698 4752
rect 19659 4644 19932 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 16408 4576 17816 4604
rect 18233 4607 18291 4613
rect 12084 4508 12940 4536
rect 12912 4480 12940 4508
rect 13078 4496 13084 4548
rect 13136 4496 13142 4548
rect 14826 4496 14832 4548
rect 14884 4536 14890 4548
rect 15488 4536 15516 4567
rect 14884 4508 15516 4536
rect 14884 4496 14890 4508
rect 4985 4471 5043 4477
rect 4985 4437 4997 4471
rect 5031 4468 5043 4471
rect 5166 4468 5172 4480
rect 5031 4440 5172 4468
rect 5031 4437 5043 4440
rect 4985 4431 5043 4437
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 12342 4468 12348 4480
rect 5316 4440 12348 4468
rect 5316 4428 5322 4440
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12894 4428 12900 4480
rect 12952 4428 12958 4480
rect 13262 4428 13268 4480
rect 13320 4428 13326 4480
rect 14182 4428 14188 4480
rect 14240 4428 14246 4480
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 15764 4468 15792 4576
rect 18233 4573 18245 4607
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 16390 4496 16396 4548
rect 16448 4536 16454 4548
rect 18248 4536 18276 4567
rect 18690 4564 18696 4616
rect 18748 4604 18754 4616
rect 19076 4604 19104 4635
rect 19978 4632 19984 4684
rect 20036 4632 20042 4684
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 20990 4672 20996 4684
rect 20947 4644 20996 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 21266 4632 21272 4684
rect 21324 4632 21330 4684
rect 21525 4675 21583 4681
rect 21525 4672 21537 4675
rect 21376 4644 21537 4672
rect 18748 4576 19104 4604
rect 19797 4607 19855 4613
rect 18748 4564 18754 4576
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 19996 4604 20024 4632
rect 19843 4576 20024 4604
rect 20809 4607 20867 4613
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 20809 4573 20821 4607
rect 20855 4604 20867 4607
rect 21082 4604 21088 4616
rect 20855 4576 21088 4604
rect 20855 4573 20867 4576
rect 20809 4567 20867 4573
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 21376 4604 21404 4644
rect 21525 4641 21537 4644
rect 21571 4641 21583 4675
rect 21525 4635 21583 4641
rect 21192 4576 21404 4604
rect 19610 4536 19616 4548
rect 16448 4508 19616 4536
rect 16448 4496 16454 4508
rect 19610 4496 19616 4508
rect 19668 4496 19674 4548
rect 20162 4496 20168 4548
rect 20220 4536 20226 4548
rect 20257 4539 20315 4545
rect 20257 4536 20269 4539
rect 20220 4508 20269 4536
rect 20220 4496 20226 4508
rect 20257 4505 20269 4508
rect 20303 4536 20315 4539
rect 20990 4536 20996 4548
rect 20303 4508 20996 4536
rect 20303 4505 20315 4508
rect 20257 4499 20315 4505
rect 20990 4496 20996 4508
rect 21048 4496 21054 4548
rect 14608 4440 15792 4468
rect 15933 4471 15991 4477
rect 14608 4428 14614 4440
rect 15933 4437 15945 4471
rect 15979 4468 15991 4471
rect 16206 4468 16212 4480
rect 15979 4440 16212 4468
rect 15979 4437 15991 4440
rect 15933 4431 15991 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 18325 4471 18383 4477
rect 18325 4437 18337 4471
rect 18371 4468 18383 4471
rect 18414 4468 18420 4480
rect 18371 4440 18420 4468
rect 18371 4437 18383 4440
rect 18325 4431 18383 4437
rect 18414 4428 18420 4440
rect 18472 4428 18478 4480
rect 18874 4428 18880 4480
rect 18932 4428 18938 4480
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4468 19763 4471
rect 19978 4468 19984 4480
rect 19751 4440 19984 4468
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 20714 4428 20720 4480
rect 20772 4428 20778 4480
rect 20806 4428 20812 4480
rect 20864 4468 20870 4480
rect 21192 4468 21220 4576
rect 20864 4440 21220 4468
rect 20864 4428 20870 4440
rect 552 4378 23368 4400
rect 552 4326 1366 4378
rect 1418 4326 1430 4378
rect 1482 4326 1494 4378
rect 1546 4326 1558 4378
rect 1610 4326 1622 4378
rect 1674 4326 1686 4378
rect 1738 4326 7366 4378
rect 7418 4326 7430 4378
rect 7482 4326 7494 4378
rect 7546 4326 7558 4378
rect 7610 4326 7622 4378
rect 7674 4326 7686 4378
rect 7738 4326 13366 4378
rect 13418 4326 13430 4378
rect 13482 4326 13494 4378
rect 13546 4326 13558 4378
rect 13610 4326 13622 4378
rect 13674 4326 13686 4378
rect 13738 4326 19366 4378
rect 19418 4326 19430 4378
rect 19482 4326 19494 4378
rect 19546 4326 19558 4378
rect 19610 4326 19622 4378
rect 19674 4326 19686 4378
rect 19738 4326 23368 4378
rect 552 4304 23368 4326
rect 2685 4267 2743 4273
rect 2685 4233 2697 4267
rect 2731 4264 2743 4267
rect 2774 4264 2780 4276
rect 2731 4236 2780 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 2700 4128 2728 4227
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 3786 4224 3792 4276
rect 3844 4264 3850 4276
rect 7006 4264 7012 4276
rect 3844 4236 7012 4264
rect 3844 4224 3850 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 11606 4224 11612 4276
rect 11664 4264 11670 4276
rect 11664 4236 13584 4264
rect 11664 4224 11670 4236
rect 5902 4196 5908 4208
rect 5552 4168 5908 4196
rect 2056 4100 2728 4128
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4060 1823 4063
rect 1946 4060 1952 4072
rect 1811 4032 1952 4060
rect 1811 4029 1823 4032
rect 1765 4023 1823 4029
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2056 4069 2084 4100
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 4338 4128 4344 4140
rect 2832 4100 4344 4128
rect 2832 4088 2838 4100
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 5552 4128 5580 4168
rect 5902 4156 5908 4168
rect 5960 4196 5966 4208
rect 13446 4196 13452 4208
rect 5960 4168 13452 4196
rect 5960 4156 5966 4168
rect 13446 4156 13452 4168
rect 13504 4156 13510 4208
rect 4663 4100 5028 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 2222 4020 2228 4072
rect 2280 4020 2286 4072
rect 2314 4020 2320 4072
rect 2372 4020 2378 4072
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 3602 4060 3608 4072
rect 2547 4032 3608 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 5000 4069 5028 4100
rect 5092 4100 5580 4128
rect 7653 4131 7711 4137
rect 5092 4069 5120 4100
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 7926 4128 7932 4140
rect 7699 4100 7932 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 7926 4088 7932 4100
rect 7984 4128 7990 4140
rect 7984 4100 8616 4128
rect 7984 4088 7990 4100
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4212 4032 4261 4060
rect 4212 4020 4218 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4029 5135 4063
rect 5077 4023 5135 4029
rect 1854 3884 1860 3936
rect 1912 3933 1918 3936
rect 1912 3887 1921 3933
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2240 3924 2268 4020
rect 5000 3992 5028 4023
rect 5166 4020 5172 4072
rect 5224 4060 5230 4072
rect 5261 4063 5319 4069
rect 5261 4060 5273 4063
rect 5224 4032 5273 4060
rect 5224 4020 5230 4032
rect 5261 4029 5273 4032
rect 5307 4029 5319 4063
rect 5261 4023 5319 4029
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 7883 4032 8401 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 5445 3995 5503 4001
rect 5000 3964 5396 3992
rect 5368 3936 5396 3964
rect 5445 3961 5457 3995
rect 5491 3992 5503 3995
rect 7852 3992 7880 4023
rect 8478 4020 8484 4072
rect 8536 4020 8542 4072
rect 8588 4069 8616 4100
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 9306 4128 9312 4140
rect 9088 4100 9312 4128
rect 9088 4088 9094 4100
rect 8573 4063 8631 4069
rect 8573 4029 8585 4063
rect 8619 4029 8631 4063
rect 8864 4060 8892 4088
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8864 4032 9137 4060
rect 8573 4023 8631 4029
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9232 4046 9260 4100
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9858 4128 9864 4140
rect 9640 4100 9864 4128
rect 9640 4088 9646 4100
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 12584 4100 13032 4128
rect 12584 4088 12590 4100
rect 9125 4023 9183 4029
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 12713 4063 12771 4069
rect 12713 4060 12725 4063
rect 12492 4032 12725 4060
rect 12492 4020 12498 4032
rect 12713 4029 12725 4032
rect 12759 4029 12771 4063
rect 12713 4023 12771 4029
rect 5491 3964 7880 3992
rect 5491 3961 5503 3964
rect 5445 3955 5503 3961
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 10137 3995 10195 4001
rect 10137 3992 10149 3995
rect 9088 3964 10149 3992
rect 9088 3952 9094 3964
rect 10137 3961 10149 3964
rect 10183 3992 10195 3995
rect 10870 3992 10876 4004
rect 10183 3964 10876 3992
rect 10183 3961 10195 3964
rect 10137 3955 10195 3961
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 1995 3896 2268 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 1912 3884 1918 3887
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 8018 3884 8024 3936
rect 8076 3884 8082 3936
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 11422 3924 11428 3936
rect 8444 3896 11428 3924
rect 8444 3884 8450 3896
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 12728 3924 12756 4023
rect 12802 4020 12808 4072
rect 12860 4020 12866 4072
rect 12894 4020 12900 4072
rect 12952 4020 12958 4072
rect 13004 4069 13032 4100
rect 13354 4088 13360 4140
rect 13412 4088 13418 4140
rect 13556 4128 13584 4236
rect 14550 4224 14556 4276
rect 14608 4224 14614 4276
rect 15102 4224 15108 4276
rect 15160 4264 15166 4276
rect 15160 4236 15700 4264
rect 15160 4224 15166 4236
rect 14568 4196 14596 4224
rect 13924 4168 14596 4196
rect 13924 4137 13952 4168
rect 15378 4156 15384 4208
rect 15436 4156 15442 4208
rect 15672 4196 15700 4236
rect 17678 4224 17684 4276
rect 17736 4224 17742 4276
rect 18230 4224 18236 4276
rect 18288 4264 18294 4276
rect 18325 4267 18383 4273
rect 18325 4264 18337 4267
rect 18288 4236 18337 4264
rect 18288 4224 18294 4236
rect 18325 4233 18337 4236
rect 18371 4233 18383 4267
rect 18325 4227 18383 4233
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 20162 4264 20168 4276
rect 18564 4236 20168 4264
rect 18564 4224 18570 4236
rect 20162 4224 20168 4236
rect 20220 4224 20226 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 22002 4264 22008 4276
rect 21416 4236 22008 4264
rect 21416 4224 21422 4236
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 22094 4224 22100 4276
rect 22152 4264 22158 4276
rect 22152 4236 22784 4264
rect 22152 4224 22158 4236
rect 17696 4196 17724 4224
rect 15672 4168 16436 4196
rect 17696 4168 19012 4196
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13556 4100 13829 4128
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4097 13967 4131
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 13909 4091 13967 4097
rect 14016 4100 14381 4128
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 12820 3992 12848 4020
rect 13096 3992 13124 4023
rect 13170 4020 13176 4072
rect 13228 4020 13234 4072
rect 13262 4020 13268 4072
rect 13320 4060 13326 4072
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 13320 4032 13553 4060
rect 13320 4020 13326 4032
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4060 13783 4063
rect 14016 4060 14044 4100
rect 14369 4097 14381 4100
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 15396 4128 15424 4156
rect 15672 4137 15700 4168
rect 16408 4140 16436 4168
rect 15657 4131 15715 4137
rect 14516 4100 15332 4128
rect 15396 4100 15516 4128
rect 14516 4088 14522 4100
rect 13771 4032 14044 4060
rect 14093 4063 14151 4069
rect 13771 4029 13783 4032
rect 13725 4023 13783 4029
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 14182 4060 14188 4072
rect 14139 4032 14188 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 12820 3964 13124 3992
rect 13188 3992 13216 4020
rect 13740 3992 13768 4023
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 14645 4063 14703 4069
rect 14645 4029 14657 4063
rect 14691 4060 14703 4063
rect 15197 4063 15255 4069
rect 15197 4060 15209 4063
rect 14691 4032 15209 4060
rect 14691 4029 14703 4032
rect 14645 4023 14703 4029
rect 15197 4029 15209 4032
rect 15243 4029 15255 4063
rect 15197 4023 15255 4029
rect 13188 3964 13768 3992
rect 14277 3995 14335 4001
rect 14277 3961 14289 3995
rect 14323 3992 14335 3995
rect 15102 3992 15108 4004
rect 14323 3964 15108 3992
rect 14323 3961 14335 3964
rect 14277 3955 14335 3961
rect 15102 3952 15108 3964
rect 15160 3952 15166 4004
rect 14458 3924 14464 3936
rect 12728 3896 14464 3924
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14826 3884 14832 3936
rect 14884 3884 14890 3936
rect 15304 3924 15332 4100
rect 15378 4020 15384 4072
rect 15436 4020 15442 4072
rect 15488 3992 15516 4100
rect 15657 4097 15669 4131
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 15930 4088 15936 4140
rect 15988 4088 15994 4140
rect 16022 4088 16028 4140
rect 16080 4088 16086 4140
rect 16390 4088 16396 4140
rect 16448 4088 16454 4140
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 15562 4020 15568 4072
rect 15620 4020 15626 4072
rect 15749 4063 15807 4069
rect 15749 4029 15761 4063
rect 15795 4029 15807 4063
rect 15948 4059 15976 4088
rect 16117 4063 16175 4069
rect 15749 4023 15807 4029
rect 15933 4053 15991 4059
rect 15764 3992 15792 4023
rect 15933 4019 15945 4053
rect 15979 4019 15991 4053
rect 16117 4029 16129 4063
rect 16163 4029 16175 4063
rect 16117 4023 16175 4029
rect 15933 4013 15991 4019
rect 15488 3964 15792 3992
rect 16132 3924 16160 4023
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 18984 4069 19012 4168
rect 20070 4156 20076 4208
rect 20128 4196 20134 4208
rect 20128 4168 20475 4196
rect 20128 4156 20134 4168
rect 20088 4128 20116 4156
rect 20346 4128 20352 4140
rect 19904 4100 20116 4128
rect 20180 4100 20352 4128
rect 19904 4069 19932 4100
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 16264 4032 16313 4060
rect 16264 4020 16270 4032
rect 16301 4029 16313 4032
rect 16347 4029 16359 4063
rect 16301 4023 16359 4029
rect 18509 4063 18567 4069
rect 18509 4029 18521 4063
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 18969 4063 19027 4069
rect 18969 4029 18981 4063
rect 19015 4029 19027 4063
rect 18969 4023 19027 4029
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4029 19947 4063
rect 19889 4023 19947 4029
rect 18524 3992 18552 4023
rect 19978 4020 19984 4072
rect 20036 4060 20042 4072
rect 20180 4069 20208 4100
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 20447 4128 20475 4168
rect 20622 4156 20628 4208
rect 20680 4196 20686 4208
rect 20680 4168 20944 4196
rect 20680 4156 20686 4168
rect 20447 4100 20576 4128
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 20036 4032 20085 4060
rect 20036 4020 20042 4032
rect 20073 4029 20085 4032
rect 20119 4029 20131 4063
rect 20073 4023 20131 4029
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4029 20223 4063
rect 20165 4023 20223 4029
rect 20257 4063 20315 4069
rect 20257 4029 20269 4063
rect 20303 4060 20315 4063
rect 20438 4060 20444 4072
rect 20303 4032 20444 4060
rect 20303 4029 20315 4032
rect 20257 4023 20315 4029
rect 18598 3992 18604 4004
rect 18524 3964 18604 3992
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 19610 3952 19616 4004
rect 19668 3992 19674 4004
rect 20272 3992 20300 4023
rect 20438 4020 20444 4032
rect 20496 4020 20502 4072
rect 20548 4060 20576 4100
rect 20622 4060 20628 4072
rect 20548 4032 20628 4060
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 20714 4020 20720 4072
rect 20772 4020 20778 4072
rect 20806 4020 20812 4072
rect 20864 4020 20870 4072
rect 20916 4069 20944 4168
rect 21542 4156 21548 4208
rect 21600 4196 21606 4208
rect 21637 4199 21695 4205
rect 21637 4196 21649 4199
rect 21600 4168 21649 4196
rect 21600 4156 21606 4168
rect 21637 4165 21649 4168
rect 21683 4165 21695 4199
rect 22557 4199 22615 4205
rect 22557 4196 22569 4199
rect 21637 4159 21695 4165
rect 21836 4168 22569 4196
rect 20901 4063 20959 4069
rect 20901 4029 20913 4063
rect 20947 4029 20959 4063
rect 20901 4023 20959 4029
rect 20993 4063 21051 4069
rect 20993 4029 21005 4063
rect 21039 4060 21051 4063
rect 21039 4032 21404 4060
rect 21039 4029 21051 4032
rect 20993 4023 21051 4029
rect 19668 3964 20300 3992
rect 20533 3995 20591 4001
rect 19668 3952 19674 3964
rect 20533 3961 20545 3995
rect 20579 3992 20591 3995
rect 20732 3992 20760 4020
rect 20579 3964 20760 3992
rect 20579 3961 20591 3964
rect 20533 3955 20591 3961
rect 15304 3896 16160 3924
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 16485 3927 16543 3933
rect 16485 3924 16497 3927
rect 16356 3896 16497 3924
rect 16356 3884 16362 3896
rect 16485 3893 16497 3896
rect 16531 3893 16543 3927
rect 16485 3887 16543 3893
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 21008 3924 21036 4023
rect 16816 3896 21036 3924
rect 16816 3884 16822 3896
rect 21174 3884 21180 3936
rect 21232 3924 21238 3936
rect 21376 3933 21404 4032
rect 21450 4020 21456 4072
rect 21508 4020 21514 4072
rect 21560 4069 21588 4156
rect 21545 4063 21603 4069
rect 21545 4029 21557 4063
rect 21591 4029 21603 4063
rect 21545 4023 21603 4029
rect 21634 4020 21640 4072
rect 21692 4060 21698 4072
rect 21836 4069 21864 4168
rect 22557 4165 22569 4168
rect 22603 4165 22615 4199
rect 22557 4159 22615 4165
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 21692 4032 21833 4060
rect 21692 4020 21698 4032
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 22097 4063 22155 4069
rect 22097 4029 22109 4063
rect 22143 4060 22155 4063
rect 22278 4060 22284 4072
rect 22143 4032 22284 4060
rect 22143 4029 22155 4032
rect 22097 4023 22155 4029
rect 22278 4020 22284 4032
rect 22336 4020 22342 4072
rect 22756 4069 22784 4236
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 22741 4063 22799 4069
rect 22741 4029 22753 4063
rect 22787 4060 22799 4063
rect 22830 4060 22836 4072
rect 22787 4032 22836 4060
rect 22787 4029 22799 4032
rect 22741 4023 22799 4029
rect 21269 3927 21327 3933
rect 21269 3924 21281 3927
rect 21232 3896 21281 3924
rect 21232 3884 21238 3896
rect 21269 3893 21281 3896
rect 21315 3893 21327 3927
rect 21269 3887 21327 3893
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3893 21419 3927
rect 21468 3924 21496 4020
rect 22002 3952 22008 4004
rect 22060 3992 22066 4004
rect 22186 3992 22192 4004
rect 22060 3964 22192 3992
rect 22060 3952 22066 3964
rect 22186 3952 22192 3964
rect 22244 3992 22250 4004
rect 22480 3992 22508 4023
rect 22830 4020 22836 4032
rect 22888 4020 22894 4072
rect 22244 3964 22508 3992
rect 22244 3952 22250 3964
rect 22281 3927 22339 3933
rect 22281 3924 22293 3927
rect 21468 3896 22293 3924
rect 21361 3887 21419 3893
rect 22281 3893 22293 3896
rect 22327 3893 22339 3927
rect 22281 3887 22339 3893
rect 552 3834 23368 3856
rect 552 3782 4366 3834
rect 4418 3782 4430 3834
rect 4482 3782 4494 3834
rect 4546 3782 4558 3834
rect 4610 3782 4622 3834
rect 4674 3782 4686 3834
rect 4738 3782 10366 3834
rect 10418 3782 10430 3834
rect 10482 3782 10494 3834
rect 10546 3782 10558 3834
rect 10610 3782 10622 3834
rect 10674 3782 10686 3834
rect 10738 3782 16366 3834
rect 16418 3782 16430 3834
rect 16482 3782 16494 3834
rect 16546 3782 16558 3834
rect 16610 3782 16622 3834
rect 16674 3782 16686 3834
rect 16738 3782 22366 3834
rect 22418 3782 22430 3834
rect 22482 3782 22494 3834
rect 22546 3782 22558 3834
rect 22610 3782 22622 3834
rect 22674 3782 22686 3834
rect 22738 3782 23368 3834
rect 552 3760 23368 3782
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 3605 3723 3663 3729
rect 2372 3692 2820 3720
rect 2372 3680 2378 3692
rect 2792 3661 2820 3692
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 4154 3720 4160 3732
rect 3651 3692 4160 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 6365 3723 6423 3729
rect 6365 3689 6377 3723
rect 6411 3720 6423 3723
rect 6914 3720 6920 3732
rect 6411 3692 6920 3720
rect 6411 3689 6423 3692
rect 6365 3683 6423 3689
rect 6914 3680 6920 3692
rect 6972 3720 6978 3732
rect 6972 3692 7052 3720
rect 6972 3680 6978 3692
rect 2777 3655 2835 3661
rect 2777 3621 2789 3655
rect 2823 3621 2835 3655
rect 2777 3615 2835 3621
rect 2961 3655 3019 3661
rect 2961 3621 2973 3655
rect 3007 3652 3019 3655
rect 3418 3652 3424 3664
rect 3007 3624 3424 3652
rect 3007 3621 3019 3624
rect 2961 3615 3019 3621
rect 3418 3612 3424 3624
rect 3476 3652 3482 3664
rect 3786 3652 3792 3664
rect 3476 3624 3792 3652
rect 3476 3612 3482 3624
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 4740 3655 4798 3661
rect 4740 3621 4752 3655
rect 4786 3652 4798 3655
rect 6549 3655 6607 3661
rect 6549 3652 6561 3655
rect 4786 3624 6561 3652
rect 4786 3621 4798 3624
rect 4740 3615 4798 3621
rect 6549 3621 6561 3624
rect 6595 3621 6607 3655
rect 6549 3615 6607 3621
rect 6656 3624 6960 3652
rect 842 3544 848 3596
rect 900 3584 906 3596
rect 1210 3593 1216 3596
rect 937 3587 995 3593
rect 937 3584 949 3587
rect 900 3556 949 3584
rect 900 3544 906 3556
rect 937 3553 949 3556
rect 983 3553 995 3587
rect 937 3547 995 3553
rect 1204 3547 1216 3593
rect 1210 3544 1216 3547
rect 1268 3544 1274 3596
rect 4982 3544 4988 3596
rect 5040 3544 5046 3596
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 6086 3584 6092 3596
rect 5491 3556 6092 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6656 3584 6684 3624
rect 6503 3556 6684 3584
rect 6733 3587 6791 3593
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6733 3553 6745 3587
rect 6779 3553 6791 3587
rect 6733 3547 6791 3553
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3516 6239 3519
rect 6748 3516 6776 3547
rect 6227 3488 6776 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 5074 3408 5080 3460
rect 5132 3408 5138 3460
rect 6012 3448 6040 3479
rect 6638 3448 6644 3460
rect 6012 3420 6644 3448
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 6932 3389 6960 3624
rect 7024 3593 7052 3692
rect 8478 3680 8484 3732
rect 8536 3680 8542 3732
rect 8588 3692 8800 3720
rect 8018 3612 8024 3664
rect 8076 3612 8082 3664
rect 8496 3652 8524 3680
rect 8128 3624 8524 3652
rect 7009 3587 7067 3593
rect 7009 3553 7021 3587
rect 7055 3553 7067 3587
rect 7009 3547 7067 3553
rect 7653 3587 7711 3593
rect 7653 3553 7665 3587
rect 7699 3553 7711 3587
rect 7653 3547 7711 3553
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3584 7987 3587
rect 8036 3584 8064 3612
rect 8128 3593 8156 3624
rect 8588 3593 8616 3692
rect 7975 3556 8064 3584
rect 8113 3587 8171 3593
rect 7975 3553 7987 3556
rect 7929 3547 7987 3553
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8205 3547 8263 3553
rect 8573 3587 8631 3593
rect 8573 3553 8585 3587
rect 8619 3553 8631 3587
rect 8772 3584 8800 3692
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9033 3723 9091 3729
rect 8904 3692 8984 3720
rect 8904 3680 8910 3692
rect 8956 3652 8984 3692
rect 9033 3689 9045 3723
rect 9079 3720 9091 3723
rect 9490 3720 9496 3732
rect 9079 3692 9496 3720
rect 9079 3689 9091 3692
rect 9033 3683 9091 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 10042 3680 10048 3732
rect 10100 3680 10106 3732
rect 10594 3720 10600 3732
rect 10152 3692 10600 3720
rect 10152 3652 10180 3692
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 11790 3720 11796 3732
rect 10704 3692 11796 3720
rect 10410 3652 10416 3664
rect 8956 3624 9444 3652
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8772 3556 9137 3584
rect 8573 3547 8631 3553
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 7282 3408 7288 3460
rect 7340 3448 7346 3460
rect 7668 3448 7696 3547
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3516 8079 3519
rect 8220 3516 8248 3547
rect 9306 3544 9312 3596
rect 9364 3544 9370 3596
rect 9416 3593 9444 3624
rect 9692 3624 10180 3652
rect 10244 3624 10416 3652
rect 9401 3587 9459 3593
rect 9401 3553 9413 3587
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 8067 3488 8524 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 8110 3448 8116 3460
rect 7340 3420 8116 3448
rect 7340 3408 7346 3420
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 8294 3408 8300 3460
rect 8352 3408 8358 3460
rect 8496 3448 8524 3488
rect 8662 3476 8668 3528
rect 8720 3476 8726 3528
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 8849 3519 8907 3525
rect 8849 3485 8861 3519
rect 8895 3516 8907 3519
rect 9030 3516 9036 3528
rect 8895 3488 9036 3516
rect 8895 3485 8907 3488
rect 8849 3479 8907 3485
rect 8772 3448 8800 3479
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 9692 3516 9720 3624
rect 9769 3587 9827 3593
rect 9769 3553 9781 3587
rect 9815 3584 9827 3587
rect 10244 3584 10272 3624
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 10704 3652 10732 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12084 3692 12434 3720
rect 10520 3624 10732 3652
rect 9815 3556 9904 3584
rect 9815 3553 9827 3556
rect 9769 3547 9827 3553
rect 9876 3525 9904 3556
rect 10152 3556 10272 3584
rect 10321 3587 10379 3593
rect 9140 3488 9720 3516
rect 9861 3519 9919 3525
rect 9140 3460 9168 3488
rect 9861 3485 9873 3519
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10152 3516 10180 3556
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 10520 3584 10548 3624
rect 11422 3612 11428 3664
rect 11480 3612 11486 3664
rect 11961 3655 12019 3661
rect 11961 3621 11973 3655
rect 12007 3652 12019 3655
rect 12084 3652 12112 3692
rect 12007 3624 12112 3652
rect 12161 3655 12219 3661
rect 12007 3621 12019 3624
rect 11961 3615 12019 3621
rect 12161 3621 12173 3655
rect 12207 3621 12219 3655
rect 12406 3652 12434 3692
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 13081 3723 13139 3729
rect 13081 3720 13093 3723
rect 12952 3692 13093 3720
rect 12952 3680 12958 3692
rect 13081 3689 13093 3692
rect 13127 3689 13139 3723
rect 13081 3683 13139 3689
rect 13188 3692 14412 3720
rect 13188 3652 13216 3692
rect 12406 3624 13216 3652
rect 12161 3615 12219 3621
rect 10367 3556 10548 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 10594 3544 10600 3596
rect 10652 3544 10658 3596
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3584 10839 3587
rect 10870 3584 10876 3596
rect 10827 3556 10876 3584
rect 10827 3553 10839 3556
rect 10781 3547 10839 3553
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 11440 3584 11468 3612
rect 12176 3584 12204 3615
rect 13446 3612 13452 3664
rect 13504 3612 13510 3664
rect 14182 3652 14188 3664
rect 13924 3624 14188 3652
rect 11440 3556 12204 3584
rect 12253 3587 12311 3593
rect 12253 3553 12265 3587
rect 12299 3584 12311 3587
rect 12342 3584 12348 3596
rect 12299 3556 12348 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 13170 3544 13176 3596
rect 13228 3584 13234 3596
rect 13265 3587 13323 3593
rect 13265 3584 13277 3587
rect 13228 3556 13277 3584
rect 13228 3544 13234 3556
rect 13265 3553 13277 3556
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3584 13415 3587
rect 13464 3584 13492 3612
rect 13924 3596 13952 3624
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 13630 3593 13636 3596
rect 13403 3556 13492 3584
rect 13615 3587 13636 3593
rect 13403 3553 13415 3556
rect 13357 3547 13415 3553
rect 13615 3553 13627 3587
rect 13615 3547 13636 3553
rect 13630 3544 13636 3547
rect 13688 3544 13694 3596
rect 13725 3587 13783 3593
rect 13725 3553 13737 3587
rect 13771 3584 13783 3587
rect 13771 3556 13860 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 13832 3528 13860 3556
rect 13906 3544 13912 3596
rect 13964 3544 13970 3596
rect 9999 3488 10180 3516
rect 10229 3519 10287 3525
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 10502 3516 10508 3528
rect 10275 3488 10508 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 8496 3420 8800 3448
rect 9122 3408 9128 3460
rect 9180 3408 9186 3460
rect 9766 3448 9772 3460
rect 9416 3420 9772 3448
rect 6917 3383 6975 3389
rect 6917 3349 6929 3383
rect 6963 3380 6975 3383
rect 7006 3380 7012 3392
rect 6963 3352 7012 3380
rect 6963 3349 6975 3352
rect 6917 3343 6975 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7837 3383 7895 3389
rect 7837 3349 7849 3383
rect 7883 3380 7895 3383
rect 7926 3380 7932 3392
rect 7883 3352 7932 3380
rect 7883 3349 7895 3352
rect 7837 3343 7895 3349
rect 7926 3340 7932 3352
rect 7984 3380 7990 3392
rect 8312 3380 8340 3408
rect 7984 3352 8340 3380
rect 8389 3383 8447 3389
rect 7984 3340 7990 3352
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 9416 3380 9444 3420
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 9876 3448 9904 3479
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 10689 3451 10747 3457
rect 10689 3448 10701 3451
rect 9876 3420 10701 3448
rect 10689 3417 10701 3420
rect 10735 3417 10747 3451
rect 10689 3411 10747 3417
rect 11054 3408 11060 3460
rect 11112 3448 11118 3460
rect 11241 3451 11299 3457
rect 11241 3448 11253 3451
rect 11112 3420 11253 3448
rect 11112 3408 11118 3420
rect 11241 3417 11253 3420
rect 11287 3417 11299 3451
rect 11624 3448 11652 3479
rect 13814 3476 13820 3528
rect 13872 3476 13878 3528
rect 14384 3516 14412 3692
rect 14918 3680 14924 3732
rect 14976 3680 14982 3732
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15436 3692 18276 3720
rect 15436 3680 15442 3692
rect 14936 3652 14964 3680
rect 16758 3652 16764 3664
rect 14936 3624 15424 3652
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 15105 3587 15163 3593
rect 15105 3584 15117 3587
rect 14516 3556 15117 3584
rect 14516 3544 14522 3556
rect 15105 3553 15117 3556
rect 15151 3553 15163 3587
rect 15105 3547 15163 3553
rect 15286 3544 15292 3596
rect 15344 3544 15350 3596
rect 15396 3593 15424 3624
rect 16132 3624 16764 3652
rect 15381 3587 15439 3593
rect 15381 3553 15393 3587
rect 15427 3553 15439 3587
rect 15381 3547 15439 3553
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 15194 3516 15200 3528
rect 14384 3488 15200 3516
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 15488 3516 15516 3547
rect 15746 3544 15752 3596
rect 15804 3544 15810 3596
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 16132 3593 16160 3624
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 18049 3655 18107 3661
rect 18049 3652 18061 3655
rect 17328 3624 18061 3652
rect 16117 3587 16175 3593
rect 16117 3584 16129 3587
rect 16080 3556 16129 3584
rect 16080 3544 16086 3556
rect 16117 3553 16129 3556
rect 16163 3553 16175 3587
rect 16117 3547 16175 3553
rect 16301 3587 16359 3593
rect 16301 3553 16313 3587
rect 16347 3584 16359 3587
rect 16390 3584 16396 3596
rect 16347 3556 16396 3584
rect 16347 3553 16359 3556
rect 16301 3547 16359 3553
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17328 3593 17356 3624
rect 18049 3621 18061 3624
rect 18095 3621 18107 3655
rect 18049 3615 18107 3621
rect 18248 3652 18276 3692
rect 18598 3680 18604 3732
rect 18656 3680 18662 3732
rect 19179 3723 19237 3729
rect 19179 3689 19191 3723
rect 19225 3720 19237 3723
rect 19886 3720 19892 3732
rect 19225 3692 19892 3720
rect 19225 3689 19237 3692
rect 19179 3683 19237 3689
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 19981 3723 20039 3729
rect 19981 3689 19993 3723
rect 20027 3720 20039 3723
rect 20806 3720 20812 3732
rect 20027 3692 20812 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 21174 3680 21180 3732
rect 21232 3680 21238 3732
rect 22649 3723 22707 3729
rect 22649 3689 22661 3723
rect 22695 3720 22707 3723
rect 22830 3720 22836 3732
rect 22695 3692 22836 3720
rect 22695 3689 22707 3692
rect 22649 3683 22707 3689
rect 22830 3680 22836 3692
rect 22888 3680 22894 3732
rect 18969 3655 19027 3661
rect 18969 3652 18981 3655
rect 18248 3624 18981 3652
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 17276 3556 17325 3584
rect 17276 3544 17282 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17497 3587 17555 3593
rect 17497 3553 17509 3587
rect 17543 3584 17555 3587
rect 17954 3584 17960 3596
rect 17543 3556 17960 3584
rect 17543 3553 17555 3556
rect 17497 3547 17555 3553
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 18248 3593 18276 3624
rect 18969 3621 18981 3624
rect 19015 3652 19027 3655
rect 20898 3652 20904 3664
rect 19015 3624 20904 3652
rect 19015 3621 19027 3624
rect 18969 3615 19027 3621
rect 20898 3612 20904 3624
rect 20956 3612 20962 3664
rect 21192 3652 21220 3680
rect 21514 3655 21572 3661
rect 21514 3652 21526 3655
rect 21192 3624 21526 3652
rect 21514 3621 21526 3624
rect 21560 3621 21572 3655
rect 21514 3615 21572 3621
rect 18141 3587 18199 3593
rect 18141 3553 18153 3587
rect 18187 3553 18199 3587
rect 18141 3547 18199 3553
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3553 18291 3587
rect 18233 3547 18291 3553
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3553 18751 3587
rect 18693 3547 18751 3553
rect 15764 3516 15792 3544
rect 18156 3516 18184 3547
rect 15488 3488 18092 3516
rect 18156 3488 18644 3516
rect 12437 3451 12495 3457
rect 12437 3448 12449 3451
rect 11624 3420 12449 3448
rect 11241 3411 11299 3417
rect 12437 3417 12449 3420
rect 12483 3448 12495 3451
rect 12483 3420 15332 3448
rect 12483 3417 12495 3420
rect 12437 3411 12495 3417
rect 8435 3352 9444 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 9490 3340 9496 3392
rect 9548 3380 9554 3392
rect 10505 3383 10563 3389
rect 10505 3380 10517 3383
rect 9548 3352 10517 3380
rect 9548 3340 9554 3352
rect 10505 3349 10517 3352
rect 10551 3349 10563 3383
rect 10505 3343 10563 3349
rect 10594 3340 10600 3392
rect 10652 3380 10658 3392
rect 11149 3383 11207 3389
rect 11149 3380 11161 3383
rect 10652 3352 11161 3380
rect 10652 3340 10658 3352
rect 11149 3349 11161 3352
rect 11195 3349 11207 3383
rect 11149 3343 11207 3349
rect 11790 3340 11796 3392
rect 11848 3340 11854 3392
rect 11977 3383 12035 3389
rect 11977 3349 11989 3383
rect 12023 3380 12035 3383
rect 12802 3380 12808 3392
rect 12023 3352 12808 3380
rect 12023 3349 12035 3352
rect 11977 3343 12035 3349
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 13078 3340 13084 3392
rect 13136 3380 13142 3392
rect 13541 3383 13599 3389
rect 13541 3380 13553 3383
rect 13136 3352 13553 3380
rect 13136 3340 13142 3352
rect 13541 3349 13553 3352
rect 13587 3349 13599 3383
rect 13541 3343 13599 3349
rect 13817 3383 13875 3389
rect 13817 3349 13829 3383
rect 13863 3380 13875 3383
rect 14458 3380 14464 3392
rect 13863 3352 14464 3380
rect 13863 3349 13875 3352
rect 13817 3343 13875 3349
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 15304 3380 15332 3420
rect 15470 3408 15476 3460
rect 15528 3448 15534 3460
rect 16850 3448 16856 3460
rect 15528 3420 16856 3448
rect 15528 3408 15534 3420
rect 16850 3408 16856 3420
rect 16908 3408 16914 3460
rect 18064 3448 18092 3488
rect 18322 3448 18328 3460
rect 18064 3420 18328 3448
rect 18322 3408 18328 3420
rect 18380 3408 18386 3460
rect 15562 3380 15568 3392
rect 15304 3352 15568 3380
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 15746 3340 15752 3392
rect 15804 3340 15810 3392
rect 16206 3340 16212 3392
rect 16264 3340 16270 3392
rect 17310 3340 17316 3392
rect 17368 3340 17374 3392
rect 18417 3383 18475 3389
rect 18417 3349 18429 3383
rect 18463 3380 18475 3383
rect 18506 3380 18512 3392
rect 18463 3352 18512 3380
rect 18463 3349 18475 3352
rect 18417 3343 18475 3349
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 18616 3380 18644 3488
rect 18708 3460 18736 3547
rect 19610 3544 19616 3596
rect 19668 3544 19674 3596
rect 19794 3544 19800 3596
rect 19852 3544 19858 3596
rect 20257 3587 20315 3593
rect 20257 3553 20269 3587
rect 20303 3584 20315 3587
rect 20806 3584 20812 3596
rect 20303 3556 20812 3584
rect 20303 3553 20315 3556
rect 20257 3547 20315 3553
rect 19978 3516 19984 3528
rect 19076 3488 19984 3516
rect 18690 3408 18696 3460
rect 18748 3448 18754 3460
rect 19076 3448 19104 3488
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 20272 3448 20300 3547
rect 20806 3544 20812 3556
rect 20864 3544 20870 3596
rect 21266 3544 21272 3596
rect 21324 3544 21330 3596
rect 18748 3420 19104 3448
rect 19168 3420 20300 3448
rect 18748 3408 18754 3420
rect 19058 3380 19064 3392
rect 18616 3352 19064 3380
rect 19058 3340 19064 3352
rect 19116 3380 19122 3392
rect 19168 3389 19196 3420
rect 19153 3383 19211 3389
rect 19153 3380 19165 3383
rect 19116 3352 19165 3380
rect 19116 3340 19122 3352
rect 19153 3349 19165 3352
rect 19199 3349 19211 3383
rect 19153 3343 19211 3349
rect 19337 3383 19395 3389
rect 19337 3349 19349 3383
rect 19383 3380 19395 3383
rect 19886 3380 19892 3392
rect 19383 3352 19892 3380
rect 19383 3349 19395 3352
rect 19337 3343 19395 3349
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 20070 3340 20076 3392
rect 20128 3340 20134 3392
rect 552 3290 23368 3312
rect 552 3238 1366 3290
rect 1418 3238 1430 3290
rect 1482 3238 1494 3290
rect 1546 3238 1558 3290
rect 1610 3238 1622 3290
rect 1674 3238 1686 3290
rect 1738 3238 7366 3290
rect 7418 3238 7430 3290
rect 7482 3238 7494 3290
rect 7546 3238 7558 3290
rect 7610 3238 7622 3290
rect 7674 3238 7686 3290
rect 7738 3238 13366 3290
rect 13418 3238 13430 3290
rect 13482 3238 13494 3290
rect 13546 3238 13558 3290
rect 13610 3238 13622 3290
rect 13674 3238 13686 3290
rect 13738 3238 19366 3290
rect 19418 3238 19430 3290
rect 19482 3238 19494 3290
rect 19546 3238 19558 3290
rect 19610 3238 19622 3290
rect 19674 3238 19686 3290
rect 19738 3238 23368 3290
rect 552 3216 23368 3238
rect 1210 3136 1216 3188
rect 1268 3176 1274 3188
rect 1397 3179 1455 3185
rect 1397 3176 1409 3179
rect 1268 3148 1409 3176
rect 1268 3136 1274 3148
rect 1397 3145 1409 3148
rect 1443 3145 1455 3179
rect 1397 3139 1455 3145
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 3237 3179 3295 3185
rect 3237 3176 3249 3179
rect 2823 3148 3249 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 3237 3145 3249 3148
rect 3283 3176 3295 3179
rect 3878 3176 3884 3188
rect 3283 3148 3884 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6638 3176 6644 3188
rect 6595 3148 6644 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 2409 3111 2467 3117
rect 2409 3077 2421 3111
rect 2455 3108 2467 3111
rect 3050 3108 3056 3120
rect 2455 3080 3056 3108
rect 2455 3077 2467 3080
rect 2409 3071 2467 3077
rect 3050 3068 3056 3080
rect 3108 3068 3114 3120
rect 1578 2932 1584 2984
rect 1636 2932 1642 2984
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2941 2007 2975
rect 1949 2935 2007 2941
rect 1964 2904 1992 2935
rect 2314 2932 2320 2984
rect 2372 2932 2378 2984
rect 2498 2932 2504 2984
rect 2556 2932 2562 2984
rect 3050 2972 3056 2984
rect 2746 2947 3056 2972
rect 2731 2944 3056 2947
rect 2731 2941 2789 2944
rect 2731 2907 2743 2941
rect 2777 2907 2789 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 3418 2932 3424 2984
rect 3476 2932 3482 2984
rect 3602 2932 3608 2984
rect 3660 2932 3666 2984
rect 1964 2876 2636 2904
rect 2731 2901 2789 2907
rect 2961 2907 3019 2913
rect 1762 2796 1768 2848
rect 1820 2796 1826 2848
rect 2608 2845 2636 2876
rect 2961 2873 2973 2907
rect 3007 2904 3019 2907
rect 6564 2904 6592 3139
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 7006 3176 7012 3188
rect 6840 3148 7012 3176
rect 6840 3108 6868 3148
rect 7006 3136 7012 3148
rect 7064 3176 7070 3188
rect 12713 3179 12771 3185
rect 7064 3148 9444 3176
rect 7064 3136 7070 3148
rect 6748 3080 6868 3108
rect 6748 2972 6776 3080
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 9416 3108 9444 3148
rect 12713 3145 12725 3179
rect 12759 3176 12771 3179
rect 12986 3176 12992 3188
rect 12759 3148 12992 3176
rect 12759 3145 12771 3148
rect 12713 3139 12771 3145
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13357 3179 13415 3185
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 13998 3176 14004 3188
rect 13403 3148 14004 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 14792 3148 15301 3176
rect 14792 3136 14798 3148
rect 15289 3145 15301 3148
rect 15335 3145 15347 3179
rect 15289 3139 15347 3145
rect 15746 3136 15752 3188
rect 15804 3136 15810 3188
rect 16206 3136 16212 3188
rect 16264 3136 16270 3188
rect 16298 3136 16304 3188
rect 16356 3136 16362 3188
rect 17310 3136 17316 3188
rect 17368 3136 17374 3188
rect 18874 3136 18880 3188
rect 18932 3176 18938 3188
rect 19705 3179 19763 3185
rect 19705 3176 19717 3179
rect 18932 3148 19717 3176
rect 18932 3136 18938 3148
rect 19705 3145 19717 3148
rect 19751 3145 19763 3179
rect 19705 3139 19763 3145
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 21726 3176 21732 3188
rect 20956 3148 21732 3176
rect 20956 3136 20962 3148
rect 21726 3136 21732 3148
rect 21784 3136 21790 3188
rect 9490 3108 9496 3120
rect 9088 3080 9352 3108
rect 9416 3080 9496 3108
rect 9088 3068 9094 3080
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 8570 3040 8576 3052
rect 6880 3012 8576 3040
rect 6880 3000 6886 3012
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 9122 3000 9128 3052
rect 9180 3000 9186 3052
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6748 2944 6929 2972
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2972 7711 2975
rect 7926 2972 7932 2984
rect 7699 2944 7932 2972
rect 7699 2941 7711 2944
rect 7653 2935 7711 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8941 2975 8999 2981
rect 8941 2972 8953 2975
rect 8680 2944 8953 2972
rect 3007 2876 6592 2904
rect 3007 2873 3019 2876
rect 2961 2867 3019 2873
rect 7834 2864 7840 2916
rect 7892 2864 7898 2916
rect 8680 2848 8708 2944
rect 8941 2941 8953 2944
rect 8987 2941 8999 2975
rect 9140 2972 9168 3000
rect 9324 2981 9352 3080
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 9766 3108 9772 3120
rect 9586 3080 9772 3108
rect 9586 2981 9614 3080
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 10502 3068 10508 3120
rect 10560 3068 10566 3120
rect 13556 3080 14964 3108
rect 10520 3040 10548 3068
rect 10781 3043 10839 3049
rect 10781 3040 10793 3043
rect 10520 3012 10793 3040
rect 10781 3009 10793 3012
rect 10827 3040 10839 3043
rect 13556 3040 13584 3080
rect 10827 3012 13584 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 13630 3000 13636 3052
rect 13688 3000 13694 3052
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 13924 3049 13952 3080
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 14458 3000 14464 3052
rect 14516 3000 14522 3052
rect 14550 3000 14556 3052
rect 14608 3000 14614 3052
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 14826 3040 14832 3052
rect 14691 3012 14832 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 9140 2944 9229 2972
rect 8941 2935 8999 2941
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2941 9367 2975
rect 9420 2975 9478 2981
rect 9420 2972 9432 2975
rect 9309 2935 9367 2941
rect 9416 2941 9432 2972
rect 9466 2941 9478 2975
rect 9416 2935 9478 2941
rect 9585 2975 9643 2981
rect 9585 2941 9597 2975
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 9416 2904 9444 2935
rect 9674 2932 9680 2984
rect 9732 2932 9738 2984
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 9824 2944 9965 2972
rect 9824 2932 9830 2944
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 9953 2935 10011 2941
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 10137 2975 10195 2981
rect 10137 2972 10149 2975
rect 10100 2944 10149 2972
rect 10100 2932 10106 2944
rect 10137 2941 10149 2944
rect 10183 2941 10195 2975
rect 10137 2935 10195 2941
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10505 2975 10563 2981
rect 10505 2972 10517 2975
rect 10284 2944 10517 2972
rect 10284 2932 10290 2944
rect 10505 2941 10517 2944
rect 10551 2941 10563 2975
rect 10505 2935 10563 2941
rect 12894 2932 12900 2984
rect 12952 2932 12958 2984
rect 13814 2972 13820 2984
rect 13004 2944 13820 2972
rect 9324 2876 9444 2904
rect 9692 2904 9720 2932
rect 10594 2904 10600 2916
rect 9692 2876 10600 2904
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2805 2651 2839
rect 2593 2799 2651 2805
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 5224 2808 6377 2836
rect 5224 2796 5230 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6365 2799 6423 2805
rect 6549 2839 6607 2845
rect 6549 2805 6561 2839
rect 6595 2836 6607 2839
rect 7469 2839 7527 2845
rect 7469 2836 7481 2839
rect 6595 2808 7481 2836
rect 6595 2805 6607 2808
rect 6549 2799 6607 2805
rect 7469 2805 7481 2808
rect 7515 2805 7527 2839
rect 7469 2799 7527 2805
rect 8662 2796 8668 2848
rect 8720 2796 8726 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 9088 2808 9137 2836
rect 9088 2796 9094 2808
rect 9125 2805 9137 2808
rect 9171 2836 9183 2839
rect 9324 2836 9352 2876
rect 10594 2864 10600 2876
rect 10652 2864 10658 2916
rect 13004 2913 13032 2944
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 13998 2932 14004 2984
rect 14056 2972 14062 2984
rect 14369 2975 14427 2981
rect 14369 2972 14381 2975
rect 14056 2944 14381 2972
rect 14056 2932 14062 2944
rect 14369 2941 14381 2944
rect 14415 2941 14427 2975
rect 14369 2935 14427 2941
rect 12989 2907 13047 2913
rect 12989 2904 13001 2907
rect 11808 2876 13001 2904
rect 11808 2848 11836 2876
rect 12989 2873 13001 2876
rect 13035 2873 13047 2907
rect 12989 2867 13047 2873
rect 13173 2907 13231 2913
rect 13173 2873 13185 2907
rect 13219 2873 13231 2907
rect 13173 2867 13231 2873
rect 9171 2808 9352 2836
rect 9171 2805 9183 2808
rect 9125 2799 9183 2805
rect 9766 2796 9772 2848
rect 9824 2796 9830 2848
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 11054 2836 11060 2848
rect 10367 2808 11060 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11790 2796 11796 2848
rect 11848 2796 11854 2848
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 13078 2836 13084 2848
rect 12400 2808 13084 2836
rect 12400 2796 12406 2808
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 13188 2836 13216 2867
rect 14826 2864 14832 2916
rect 14884 2864 14890 2916
rect 14936 2904 14964 3080
rect 15764 3049 15792 3136
rect 15749 3043 15807 3049
rect 15028 3012 15700 3040
rect 15028 2981 15056 3012
rect 15013 2975 15071 2981
rect 15013 2941 15025 2975
rect 15059 2941 15071 2975
rect 15470 2972 15476 2984
rect 15013 2935 15071 2941
rect 15120 2944 15476 2972
rect 15120 2904 15148 2944
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 15562 2932 15568 2984
rect 15620 2932 15626 2984
rect 15672 2981 15700 3012
rect 15749 3009 15761 3043
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 16022 3000 16028 3052
rect 16080 3000 16086 3052
rect 16224 3049 16252 3136
rect 16316 3108 16344 3136
rect 17328 3108 17356 3136
rect 16316 3080 16436 3108
rect 16209 3043 16267 3049
rect 16209 3009 16221 3043
rect 16255 3009 16267 3043
rect 16209 3003 16267 3009
rect 16298 3000 16304 3052
rect 16356 3000 16362 3052
rect 16408 3049 16436 3080
rect 16960 3080 17356 3108
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3009 16451 3043
rect 16393 3003 16451 3009
rect 15657 2975 15715 2981
rect 15657 2941 15669 2975
rect 15703 2972 15715 2975
rect 16040 2972 16068 3000
rect 15703 2944 16068 2972
rect 16117 2975 16175 2981
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 16117 2941 16129 2975
rect 16163 2941 16175 2975
rect 16117 2935 16175 2941
rect 14936 2876 15148 2904
rect 15197 2907 15255 2913
rect 15197 2873 15209 2907
rect 15243 2904 15255 2907
rect 16132 2904 16160 2935
rect 16574 2932 16580 2984
rect 16632 2932 16638 2984
rect 16960 2981 16988 3080
rect 18506 3068 18512 3120
rect 18564 3108 18570 3120
rect 19426 3108 19432 3120
rect 18564 3080 19432 3108
rect 18564 3068 18570 3080
rect 19426 3068 19432 3080
rect 19484 3068 19490 3120
rect 19889 3111 19947 3117
rect 19889 3077 19901 3111
rect 19935 3077 19947 3111
rect 19889 3071 19947 3077
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18380 3012 18920 3040
rect 18380 3000 18386 3012
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 15243 2876 16160 2904
rect 16669 2907 16727 2913
rect 15243 2873 15255 2876
rect 15197 2867 15255 2873
rect 16669 2873 16681 2907
rect 16715 2904 16727 2907
rect 16758 2904 16764 2916
rect 16715 2876 16764 2904
rect 16715 2873 16727 2876
rect 16669 2867 16727 2873
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 13538 2836 13544 2848
rect 13188 2808 13544 2836
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 14090 2796 14096 2848
rect 14148 2796 14154 2848
rect 14185 2839 14243 2845
rect 14185 2805 14197 2839
rect 14231 2836 14243 2839
rect 15562 2836 15568 2848
rect 14231 2808 15568 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 15930 2796 15936 2848
rect 15988 2796 15994 2848
rect 16206 2796 16212 2848
rect 16264 2836 16270 2848
rect 16960 2836 16988 2935
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 17092 2944 17141 2972
rect 17092 2932 17098 2944
rect 17129 2941 17141 2944
rect 17175 2972 17187 2975
rect 17175 2944 18736 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 18708 2848 18736 2944
rect 18782 2932 18788 2984
rect 18840 2932 18846 2984
rect 16264 2808 16988 2836
rect 16264 2796 16270 2808
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 18785 2839 18843 2845
rect 18785 2836 18797 2839
rect 18748 2808 18797 2836
rect 18748 2796 18754 2808
rect 18785 2805 18797 2808
rect 18831 2805 18843 2839
rect 18892 2836 18920 3012
rect 18969 2975 19027 2981
rect 18969 2941 18981 2975
rect 19015 2972 19027 2975
rect 19058 2972 19064 2984
rect 19015 2944 19064 2972
rect 19015 2941 19027 2944
rect 18969 2935 19027 2941
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 19334 2932 19340 2984
rect 19392 2932 19398 2984
rect 19904 2972 19932 3071
rect 21085 2975 21143 2981
rect 21085 2972 21097 2975
rect 19904 2944 21097 2972
rect 21085 2941 21097 2944
rect 21131 2941 21143 2975
rect 21085 2935 21143 2941
rect 19705 2907 19763 2913
rect 19705 2873 19717 2907
rect 19751 2904 19763 2907
rect 19981 2907 20039 2913
rect 19981 2904 19993 2907
rect 19751 2876 19993 2904
rect 19751 2873 19763 2876
rect 19705 2867 19763 2873
rect 19981 2873 19993 2876
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 20070 2864 20076 2916
rect 20128 2904 20134 2916
rect 20165 2907 20223 2913
rect 20165 2904 20177 2907
rect 20128 2876 20177 2904
rect 20128 2864 20134 2876
rect 20165 2873 20177 2876
rect 20211 2873 20223 2907
rect 20165 2867 20223 2873
rect 20180 2836 20208 2867
rect 20254 2864 20260 2916
rect 20312 2904 20318 2916
rect 20349 2907 20407 2913
rect 20349 2904 20361 2907
rect 20312 2876 20361 2904
rect 20312 2864 20318 2876
rect 20349 2873 20361 2876
rect 20395 2873 20407 2907
rect 20349 2867 20407 2873
rect 18892 2808 20208 2836
rect 18785 2799 18843 2805
rect 21266 2796 21272 2848
rect 21324 2796 21330 2848
rect 552 2746 23368 2768
rect 552 2694 4366 2746
rect 4418 2694 4430 2746
rect 4482 2694 4494 2746
rect 4546 2694 4558 2746
rect 4610 2694 4622 2746
rect 4674 2694 4686 2746
rect 4738 2694 10366 2746
rect 10418 2694 10430 2746
rect 10482 2694 10494 2746
rect 10546 2694 10558 2746
rect 10610 2694 10622 2746
rect 10674 2694 10686 2746
rect 10738 2694 16366 2746
rect 16418 2694 16430 2746
rect 16482 2694 16494 2746
rect 16546 2694 16558 2746
rect 16610 2694 16622 2746
rect 16674 2694 16686 2746
rect 16738 2694 22366 2746
rect 22418 2694 22430 2746
rect 22482 2694 22494 2746
rect 22546 2694 22558 2746
rect 22610 2694 22622 2746
rect 22674 2694 22686 2746
rect 22738 2694 23368 2746
rect 552 2672 23368 2694
rect 2498 2592 2504 2644
rect 2556 2632 2562 2644
rect 4062 2632 4068 2644
rect 2556 2604 4068 2632
rect 2556 2592 2562 2604
rect 1388 2567 1446 2573
rect 1388 2533 1400 2567
rect 1434 2564 1446 2567
rect 1762 2564 1768 2576
rect 1434 2536 1768 2564
rect 1434 2533 1446 2536
rect 1388 2527 1446 2533
rect 1762 2524 1768 2536
rect 1820 2524 1826 2576
rect 1121 2499 1179 2505
rect 1121 2465 1133 2499
rect 1167 2496 1179 2499
rect 1210 2496 1216 2508
rect 1167 2468 1216 2496
rect 1167 2465 1179 2468
rect 1121 2459 1179 2465
rect 1210 2456 1216 2468
rect 1268 2456 1274 2508
rect 2884 2505 2912 2604
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 8938 2592 8944 2644
rect 8996 2632 9002 2644
rect 9769 2635 9827 2641
rect 8996 2604 9536 2632
rect 8996 2592 9002 2604
rect 3602 2524 3608 2576
rect 3660 2564 3666 2576
rect 3660 2536 9168 2564
rect 3660 2524 3666 2536
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3620 2496 3648 2524
rect 3191 2468 3648 2496
rect 3973 2499 4031 2505
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3973 2465 3985 2499
rect 4019 2496 4031 2499
rect 5166 2496 5172 2508
rect 4019 2468 5172 2496
rect 4019 2465 4031 2468
rect 3973 2459 4031 2465
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 4433 2431 4491 2437
rect 4433 2428 4445 2431
rect 3936 2400 4445 2428
rect 3936 2388 3942 2400
rect 4433 2397 4445 2400
rect 4479 2397 4491 2431
rect 4433 2391 4491 2397
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 7282 2428 7288 2440
rect 4755 2400 7288 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 9030 2360 9036 2372
rect 3712 2332 9036 2360
rect 3712 2304 3740 2332
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 3694 2252 3700 2304
rect 3752 2252 3758 2304
rect 3786 2252 3792 2304
rect 3844 2252 3850 2304
rect 7282 2252 7288 2304
rect 7340 2292 7346 2304
rect 8754 2292 8760 2304
rect 7340 2264 8760 2292
rect 7340 2252 7346 2264
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 9140 2292 9168 2536
rect 9214 2524 9220 2576
rect 9272 2524 9278 2576
rect 9508 2573 9536 2604
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 9950 2632 9956 2644
rect 9815 2604 9956 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10778 2632 10784 2644
rect 10284 2604 10784 2632
rect 10284 2592 10290 2604
rect 10778 2592 10784 2604
rect 10836 2632 10842 2644
rect 10836 2604 11468 2632
rect 10836 2592 10842 2604
rect 9493 2567 9551 2573
rect 9493 2533 9505 2567
rect 9539 2533 9551 2567
rect 9493 2527 9551 2533
rect 9677 2567 9735 2573
rect 9677 2533 9689 2567
rect 9723 2564 9735 2567
rect 9858 2564 9864 2576
rect 9723 2536 9864 2564
rect 9723 2533 9735 2536
rect 9677 2527 9735 2533
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 10042 2524 10048 2576
rect 10100 2564 10106 2576
rect 10100 2536 10272 2564
rect 10100 2524 10106 2536
rect 9232 2496 9260 2524
rect 9766 2496 9772 2508
rect 9232 2468 9772 2496
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 9876 2496 9904 2524
rect 10244 2505 10272 2536
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 11112 2536 11376 2564
rect 11112 2524 11118 2536
rect 11348 2505 11376 2536
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9876 2468 9965 2496
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2465 10287 2499
rect 11241 2499 11299 2505
rect 11241 2496 11253 2499
rect 10229 2459 10287 2465
rect 10612 2468 11253 2496
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 9784 2428 9812 2456
rect 10152 2428 10180 2459
rect 9548 2400 9674 2428
rect 9784 2400 10180 2428
rect 9548 2388 9554 2400
rect 9646 2360 9674 2400
rect 10318 2388 10324 2440
rect 10376 2388 10382 2440
rect 9766 2360 9772 2372
rect 9646 2332 9772 2360
rect 9766 2320 9772 2332
rect 9824 2320 9830 2372
rect 10045 2363 10103 2369
rect 10045 2329 10057 2363
rect 10091 2360 10103 2363
rect 10612 2360 10640 2468
rect 11241 2465 11253 2468
rect 11287 2465 11299 2499
rect 11241 2459 11299 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2465 11391 2499
rect 11440 2496 11468 2604
rect 11698 2592 11704 2644
rect 11756 2632 11762 2644
rect 12802 2632 12808 2644
rect 11756 2604 12808 2632
rect 11756 2592 11762 2604
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 13814 2632 13820 2644
rect 12952 2604 13820 2632
rect 12952 2592 12958 2604
rect 13814 2592 13820 2604
rect 13872 2632 13878 2644
rect 14274 2632 14280 2644
rect 13872 2604 14280 2632
rect 13872 2592 13878 2604
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 15194 2592 15200 2644
rect 15252 2632 15258 2644
rect 20254 2632 20260 2644
rect 15252 2604 18184 2632
rect 15252 2592 15258 2604
rect 13170 2524 13176 2576
rect 13228 2524 13234 2576
rect 13538 2524 13544 2576
rect 13596 2524 13602 2576
rect 15654 2524 15660 2576
rect 15712 2564 15718 2576
rect 15712 2536 16344 2564
rect 15712 2524 15718 2536
rect 11609 2499 11667 2505
rect 11609 2496 11621 2499
rect 11440 2468 11621 2496
rect 11333 2459 11391 2465
rect 11609 2465 11621 2468
rect 11655 2465 11667 2499
rect 13188 2489 13216 2524
rect 14277 2499 14335 2505
rect 11609 2459 11667 2465
rect 13173 2483 13231 2489
rect 13173 2449 13185 2483
rect 13219 2449 13231 2483
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 13173 2443 13231 2449
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 10091 2332 10640 2360
rect 10091 2329 10103 2332
rect 10045 2323 10103 2329
rect 10778 2320 10784 2372
rect 10836 2360 10842 2372
rect 11072 2360 11100 2391
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11204 2400 11897 2428
rect 11204 2388 11210 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 14001 2431 14059 2437
rect 11885 2391 11943 2397
rect 13740 2400 13952 2428
rect 10836 2332 11652 2360
rect 10836 2320 10842 2332
rect 11146 2292 11152 2304
rect 9140 2264 11152 2292
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 11514 2252 11520 2304
rect 11572 2252 11578 2304
rect 11624 2292 11652 2332
rect 12802 2320 12808 2372
rect 12860 2360 12866 2372
rect 13740 2360 13768 2400
rect 12860 2332 13768 2360
rect 12860 2320 12866 2332
rect 13814 2320 13820 2372
rect 13872 2320 13878 2372
rect 13924 2360 13952 2400
rect 14001 2397 14013 2431
rect 14047 2428 14059 2431
rect 14292 2428 14320 2459
rect 16206 2456 16212 2508
rect 16264 2456 16270 2508
rect 16316 2505 16344 2536
rect 16850 2524 16856 2576
rect 16908 2524 16914 2576
rect 17862 2564 17868 2576
rect 16960 2536 17868 2564
rect 16301 2499 16359 2505
rect 16301 2465 16313 2499
rect 16347 2465 16359 2499
rect 16301 2459 16359 2465
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2496 16635 2499
rect 16666 2496 16672 2508
rect 16623 2468 16672 2496
rect 16623 2465 16635 2468
rect 16577 2459 16635 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2496 16819 2499
rect 16868 2496 16896 2524
rect 16807 2468 16896 2496
rect 16807 2465 16819 2468
rect 16761 2459 16819 2465
rect 14550 2428 14556 2440
rect 14047 2400 14556 2428
rect 14047 2397 14059 2400
rect 14001 2391 14059 2397
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15528 2400 16129 2428
rect 15528 2388 15534 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16224 2428 16252 2456
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16224 2400 16497 2428
rect 16117 2391 16175 2397
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 16684 2428 16712 2456
rect 16960 2428 16988 2536
rect 17862 2524 17868 2536
rect 17920 2524 17926 2576
rect 17034 2456 17040 2508
rect 17092 2456 17098 2508
rect 16684 2400 16988 2428
rect 16485 2391 16543 2397
rect 16393 2363 16451 2369
rect 13924 2332 16344 2360
rect 12989 2295 13047 2301
rect 12989 2292 13001 2295
rect 11624 2264 13001 2292
rect 12989 2261 13001 2264
rect 13035 2292 13047 2295
rect 13078 2292 13084 2304
rect 13035 2264 13084 2292
rect 13035 2261 13047 2264
rect 12989 2255 13047 2261
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 14093 2295 14151 2301
rect 14093 2292 14105 2295
rect 13320 2264 14105 2292
rect 13320 2252 13326 2264
rect 14093 2261 14105 2264
rect 14139 2261 14151 2295
rect 14093 2255 14151 2261
rect 15010 2252 15016 2304
rect 15068 2292 15074 2304
rect 15746 2292 15752 2304
rect 15068 2264 15752 2292
rect 15068 2252 15074 2264
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 16316 2292 16344 2332
rect 16393 2329 16405 2363
rect 16439 2360 16451 2363
rect 17052 2360 17080 2456
rect 18156 2428 18184 2604
rect 19076 2604 20260 2632
rect 18230 2456 18236 2508
rect 18288 2456 18294 2508
rect 18322 2456 18328 2508
rect 18380 2496 18386 2508
rect 19076 2505 19104 2604
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 20806 2592 20812 2644
rect 20864 2632 20870 2644
rect 22833 2635 22891 2641
rect 22833 2632 22845 2635
rect 20864 2604 22845 2632
rect 20864 2592 20870 2604
rect 22833 2601 22845 2604
rect 22879 2601 22891 2635
rect 22833 2595 22891 2601
rect 19613 2567 19671 2573
rect 19613 2533 19625 2567
rect 19659 2564 19671 2567
rect 19659 2536 19932 2564
rect 19659 2533 19671 2536
rect 19613 2527 19671 2533
rect 18877 2499 18935 2505
rect 18877 2496 18889 2499
rect 18380 2468 18889 2496
rect 18380 2456 18386 2468
rect 18877 2465 18889 2468
rect 18923 2465 18935 2499
rect 18877 2459 18935 2465
rect 19061 2499 19119 2505
rect 19061 2465 19073 2499
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 19334 2456 19340 2508
rect 19392 2456 19398 2508
rect 19702 2456 19708 2508
rect 19760 2456 19766 2508
rect 19904 2505 19932 2536
rect 21266 2524 21272 2576
rect 21324 2564 21330 2576
rect 21698 2567 21756 2573
rect 21698 2564 21710 2567
rect 21324 2536 21710 2564
rect 21324 2524 21330 2536
rect 21698 2533 21710 2536
rect 21744 2533 21756 2567
rect 21698 2527 21756 2533
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 21358 2456 21364 2508
rect 21416 2496 21422 2508
rect 21453 2499 21511 2505
rect 21453 2496 21465 2499
rect 21416 2468 21465 2496
rect 21416 2456 21422 2468
rect 21453 2465 21465 2468
rect 21499 2465 21511 2499
rect 21453 2459 21511 2465
rect 19242 2428 19248 2440
rect 18156 2400 19248 2428
rect 19242 2388 19248 2400
rect 19300 2428 19306 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19300 2400 19441 2428
rect 19300 2388 19306 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 20622 2428 20628 2440
rect 19659 2400 20628 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 16439 2332 17080 2360
rect 16439 2329 16451 2332
rect 16393 2323 16451 2329
rect 17034 2292 17040 2304
rect 16316 2264 17040 2292
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 18325 2295 18383 2301
rect 18325 2261 18337 2295
rect 18371 2292 18383 2295
rect 18414 2292 18420 2304
rect 18371 2264 18420 2292
rect 18371 2261 18383 2264
rect 18325 2255 18383 2261
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 19886 2252 19892 2304
rect 19944 2252 19950 2304
rect 552 2202 23368 2224
rect 552 2150 1366 2202
rect 1418 2150 1430 2202
rect 1482 2150 1494 2202
rect 1546 2150 1558 2202
rect 1610 2150 1622 2202
rect 1674 2150 1686 2202
rect 1738 2150 7366 2202
rect 7418 2150 7430 2202
rect 7482 2150 7494 2202
rect 7546 2150 7558 2202
rect 7610 2150 7622 2202
rect 7674 2150 7686 2202
rect 7738 2150 13366 2202
rect 13418 2150 13430 2202
rect 13482 2150 13494 2202
rect 13546 2150 13558 2202
rect 13610 2150 13622 2202
rect 13674 2150 13686 2202
rect 13738 2150 19366 2202
rect 19418 2150 19430 2202
rect 19482 2150 19494 2202
rect 19546 2150 19558 2202
rect 19610 2150 19622 2202
rect 19674 2150 19686 2202
rect 19738 2150 23368 2202
rect 552 2128 23368 2150
rect 3878 2048 3884 2100
rect 3936 2048 3942 2100
rect 4154 2048 4160 2100
rect 4212 2048 4218 2100
rect 6089 2091 6147 2097
rect 6089 2057 6101 2091
rect 6135 2088 6147 2091
rect 6135 2060 8064 2088
rect 6135 2057 6147 2060
rect 6089 2051 6147 2057
rect 1026 1980 1032 2032
rect 1084 2020 1090 2032
rect 1673 2023 1731 2029
rect 1673 2020 1685 2023
rect 1084 1992 1685 2020
rect 1084 1980 1090 1992
rect 1673 1989 1685 1992
rect 1719 1989 1731 2023
rect 1673 1983 1731 1989
rect 3510 1952 3516 1964
rect 1596 1924 3516 1952
rect 1596 1893 1624 1924
rect 3510 1912 3516 1924
rect 3568 1912 3574 1964
rect 3789 1955 3847 1961
rect 3789 1921 3801 1955
rect 3835 1952 3847 1955
rect 3896 1952 3924 2048
rect 4172 2020 4200 2048
rect 3835 1924 3924 1952
rect 3988 1992 4200 2020
rect 6733 2023 6791 2029
rect 3835 1921 3847 1924
rect 3789 1915 3847 1921
rect 1581 1887 1639 1893
rect 1581 1853 1593 1887
rect 1627 1853 1639 1887
rect 1581 1847 1639 1853
rect 1857 1887 1915 1893
rect 1857 1853 1869 1887
rect 1903 1884 1915 1887
rect 2406 1884 2412 1896
rect 1903 1856 2412 1884
rect 1903 1853 1915 1856
rect 1857 1847 1915 1853
rect 2406 1844 2412 1856
rect 2464 1844 2470 1896
rect 3988 1893 4016 1992
rect 6733 1989 6745 2023
rect 6779 2020 6791 2023
rect 7193 2023 7251 2029
rect 6779 1992 7144 2020
rect 6779 1989 6791 1992
rect 6733 1983 6791 1989
rect 4157 1955 4215 1961
rect 4157 1921 4169 1955
rect 4203 1952 4215 1955
rect 4709 1955 4767 1961
rect 4203 1924 4568 1952
rect 4203 1921 4215 1924
rect 4157 1915 4215 1921
rect 4540 1893 4568 1924
rect 4709 1921 4721 1955
rect 4755 1952 4767 1955
rect 4893 1955 4951 1961
rect 4893 1952 4905 1955
rect 4755 1924 4905 1952
rect 4755 1921 4767 1924
rect 4709 1915 4767 1921
rect 4893 1921 4905 1924
rect 4939 1921 4951 1955
rect 4893 1915 4951 1921
rect 5353 1955 5411 1961
rect 5353 1921 5365 1955
rect 5399 1952 5411 1955
rect 7116 1952 7144 1992
rect 7193 1989 7205 2023
rect 7239 2020 7251 2023
rect 7239 1992 7972 2020
rect 7239 1989 7251 1992
rect 7193 1983 7251 1989
rect 7944 1961 7972 1992
rect 7469 1955 7527 1961
rect 5399 1924 5948 1952
rect 5399 1921 5411 1924
rect 5353 1915 5411 1921
rect 3973 1887 4031 1893
rect 3973 1853 3985 1887
rect 4019 1853 4031 1887
rect 3973 1847 4031 1853
rect 4249 1887 4307 1893
rect 4249 1853 4261 1887
rect 4295 1853 4307 1887
rect 4249 1847 4307 1853
rect 4525 1887 4583 1893
rect 4525 1853 4537 1887
rect 4571 1853 4583 1887
rect 4525 1847 4583 1853
rect 4264 1760 4292 1847
rect 4338 1776 4344 1828
rect 4396 1776 4402 1828
rect 4908 1816 4936 1915
rect 4982 1844 4988 1896
rect 5040 1884 5046 1896
rect 5920 1893 5948 1924
rect 7116 1924 7420 1952
rect 5445 1887 5503 1893
rect 5445 1884 5457 1887
rect 5040 1856 5457 1884
rect 5040 1844 5046 1856
rect 5445 1853 5457 1856
rect 5491 1853 5503 1887
rect 5445 1847 5503 1853
rect 5905 1887 5963 1893
rect 5905 1853 5917 1887
rect 5951 1884 5963 1887
rect 6549 1887 6607 1893
rect 6549 1884 6561 1887
rect 5951 1856 6561 1884
rect 5951 1853 5963 1856
rect 5905 1847 5963 1853
rect 6549 1853 6561 1856
rect 6595 1853 6607 1887
rect 7006 1884 7012 1896
rect 6549 1847 6607 1853
rect 6840 1856 7012 1884
rect 5583 1819 5641 1825
rect 5583 1816 5595 1819
rect 4908 1788 5595 1816
rect 5583 1785 5595 1788
rect 5629 1785 5641 1819
rect 5583 1779 5641 1785
rect 5718 1776 5724 1828
rect 5776 1776 5782 1828
rect 5813 1819 5871 1825
rect 5813 1785 5825 1819
rect 5859 1816 5871 1819
rect 6840 1816 6868 1856
rect 7006 1844 7012 1856
rect 7064 1844 7070 1896
rect 7116 1893 7144 1924
rect 7392 1893 7420 1924
rect 7469 1921 7481 1955
rect 7515 1952 7527 1955
rect 7837 1955 7895 1961
rect 7837 1952 7849 1955
rect 7515 1924 7849 1952
rect 7515 1921 7527 1924
rect 7469 1915 7527 1921
rect 7837 1921 7849 1924
rect 7883 1921 7895 1955
rect 7837 1915 7895 1921
rect 7929 1955 7987 1961
rect 7929 1921 7941 1955
rect 7975 1921 7987 1955
rect 8036 1952 8064 2060
rect 8662 2048 8668 2100
rect 8720 2088 8726 2100
rect 8941 2091 8999 2097
rect 8941 2088 8953 2091
rect 8720 2060 8953 2088
rect 8720 2048 8726 2060
rect 8941 2057 8953 2060
rect 8987 2057 8999 2091
rect 8941 2051 8999 2057
rect 9122 2048 9128 2100
rect 9180 2088 9186 2100
rect 9401 2091 9459 2097
rect 9401 2088 9413 2091
rect 9180 2060 9413 2088
rect 9180 2048 9186 2060
rect 9401 2057 9413 2060
rect 9447 2088 9459 2091
rect 10042 2088 10048 2100
rect 9447 2060 10048 2088
rect 9447 2057 9459 2060
rect 9401 2051 9459 2057
rect 10042 2048 10048 2060
rect 10100 2048 10106 2100
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 11204 2060 18184 2088
rect 11204 2048 11210 2060
rect 18049 2023 18107 2029
rect 18049 2020 18061 2023
rect 8588 1992 9076 2020
rect 8588 1961 8616 1992
rect 9048 1961 9076 1992
rect 9646 1992 18061 2020
rect 8481 1955 8539 1961
rect 8481 1952 8493 1955
rect 8036 1924 8493 1952
rect 7929 1915 7987 1921
rect 8481 1921 8493 1924
rect 8527 1921 8539 1955
rect 8481 1915 8539 1921
rect 8573 1955 8631 1961
rect 8573 1921 8585 1955
rect 8619 1921 8631 1955
rect 9033 1955 9091 1961
rect 8573 1915 8631 1921
rect 8680 1924 8892 1952
rect 7101 1887 7159 1893
rect 7101 1853 7113 1887
rect 7147 1853 7159 1887
rect 7101 1847 7159 1853
rect 7285 1887 7343 1893
rect 7285 1853 7297 1887
rect 7331 1853 7343 1887
rect 7285 1847 7343 1853
rect 7377 1887 7435 1893
rect 7377 1853 7389 1887
rect 7423 1853 7435 1887
rect 7377 1847 7435 1853
rect 7300 1816 7328 1847
rect 5859 1788 6868 1816
rect 6932 1788 7328 1816
rect 7392 1816 7420 1847
rect 7558 1844 7564 1896
rect 7616 1844 7622 1896
rect 7742 1844 7748 1896
rect 7800 1844 7806 1896
rect 8021 1887 8079 1893
rect 8021 1853 8033 1887
rect 8067 1853 8079 1887
rect 8021 1847 8079 1853
rect 7392 1788 7696 1816
rect 5859 1785 5871 1788
rect 5813 1779 5871 1785
rect 6932 1760 6960 1788
rect 7668 1760 7696 1788
rect 7834 1776 7840 1828
rect 7892 1816 7898 1828
rect 8035 1816 8063 1847
rect 8294 1844 8300 1896
rect 8352 1884 8358 1896
rect 8680 1893 8708 1924
rect 8665 1887 8723 1893
rect 8665 1884 8677 1887
rect 8352 1856 8677 1884
rect 8352 1844 8358 1856
rect 8665 1853 8677 1856
rect 8711 1853 8723 1887
rect 8665 1847 8723 1853
rect 8757 1887 8815 1893
rect 8757 1853 8769 1887
rect 8803 1853 8815 1887
rect 8864 1884 8892 1924
rect 9033 1921 9045 1955
rect 9079 1952 9091 1955
rect 9646 1952 9674 1992
rect 18049 1989 18061 1992
rect 18095 1989 18107 2023
rect 18156 2020 18184 2060
rect 18690 2048 18696 2100
rect 18748 2088 18754 2100
rect 18874 2088 18880 2100
rect 18748 2060 18880 2088
rect 18748 2048 18754 2060
rect 18874 2048 18880 2060
rect 18932 2048 18938 2100
rect 21726 2048 21732 2100
rect 21784 2048 21790 2100
rect 18156 1992 21496 2020
rect 18049 1983 18107 1989
rect 9079 1924 9812 1952
rect 9079 1921 9091 1924
rect 9033 1915 9091 1921
rect 9784 1893 9812 1924
rect 9858 1912 9864 1964
rect 9916 1952 9922 1964
rect 10226 1952 10232 1964
rect 9916 1924 10232 1952
rect 9916 1912 9922 1924
rect 10226 1912 10232 1924
rect 10284 1912 10290 1964
rect 10318 1912 10324 1964
rect 10376 1952 10382 1964
rect 10413 1955 10471 1961
rect 10413 1952 10425 1955
rect 10376 1924 10425 1952
rect 10376 1912 10382 1924
rect 10413 1921 10425 1924
rect 10459 1921 10471 1955
rect 10413 1915 10471 1921
rect 10597 1955 10655 1961
rect 10597 1921 10609 1955
rect 10643 1952 10655 1955
rect 11054 1952 11060 1964
rect 10643 1924 11060 1952
rect 10643 1921 10655 1924
rect 10597 1915 10655 1921
rect 11054 1912 11060 1924
rect 11112 1912 11118 1964
rect 12345 1955 12403 1961
rect 12345 1952 12357 1955
rect 11164 1924 12357 1952
rect 11164 1896 11192 1924
rect 12345 1921 12357 1924
rect 12391 1921 12403 1955
rect 12986 1952 12992 1964
rect 12345 1915 12403 1921
rect 12452 1924 12992 1952
rect 9217 1887 9275 1893
rect 9217 1884 9229 1887
rect 8864 1856 9229 1884
rect 8757 1847 8815 1853
rect 9217 1853 9229 1856
rect 9263 1884 9275 1887
rect 9585 1887 9643 1893
rect 9585 1884 9597 1887
rect 9263 1856 9597 1884
rect 9263 1853 9275 1856
rect 9217 1847 9275 1853
rect 9585 1853 9597 1856
rect 9631 1853 9643 1887
rect 9585 1847 9643 1853
rect 9769 1887 9827 1893
rect 9769 1853 9781 1887
rect 9815 1853 9827 1887
rect 9769 1847 9827 1853
rect 9953 1887 10011 1893
rect 9953 1853 9965 1887
rect 9999 1884 10011 1887
rect 10505 1887 10563 1893
rect 10505 1884 10517 1887
rect 9999 1856 10517 1884
rect 9999 1853 10011 1856
rect 9953 1847 10011 1853
rect 10505 1853 10517 1856
rect 10551 1853 10563 1887
rect 10505 1847 10563 1853
rect 10689 1887 10747 1893
rect 10689 1853 10701 1887
rect 10735 1884 10747 1887
rect 10778 1884 10784 1896
rect 10735 1856 10784 1884
rect 10735 1853 10747 1856
rect 10689 1847 10747 1853
rect 7892 1788 8063 1816
rect 7892 1776 7898 1788
rect 8386 1776 8392 1828
rect 8444 1816 8450 1828
rect 8772 1816 8800 1847
rect 10778 1844 10784 1856
rect 10836 1844 10842 1896
rect 11146 1844 11152 1896
rect 11204 1844 11210 1896
rect 11238 1844 11244 1896
rect 11296 1844 11302 1896
rect 11330 1844 11336 1896
rect 11388 1844 11394 1896
rect 11514 1844 11520 1896
rect 11572 1844 11578 1896
rect 12452 1893 12480 1924
rect 12986 1912 12992 1924
rect 13044 1912 13050 1964
rect 13814 1912 13820 1964
rect 13872 1952 13878 1964
rect 15010 1952 15016 1964
rect 13872 1924 15016 1952
rect 13872 1912 13878 1924
rect 15010 1912 15016 1924
rect 15068 1912 15074 1964
rect 15470 1912 15476 1964
rect 15528 1952 15534 1964
rect 15528 1924 15792 1952
rect 15528 1912 15534 1924
rect 12253 1887 12311 1893
rect 12253 1853 12265 1887
rect 12299 1853 12311 1887
rect 12253 1847 12311 1853
rect 12437 1887 12495 1893
rect 12437 1853 12449 1887
rect 12483 1853 12495 1887
rect 12437 1847 12495 1853
rect 11606 1816 11612 1828
rect 8444 1788 8800 1816
rect 10244 1788 11612 1816
rect 8444 1776 8450 1788
rect 1118 1708 1124 1760
rect 1176 1748 1182 1760
rect 1397 1751 1455 1757
rect 1397 1748 1409 1751
rect 1176 1720 1409 1748
rect 1176 1708 1182 1720
rect 1397 1717 1409 1720
rect 1443 1717 1455 1751
rect 1397 1711 1455 1717
rect 4246 1708 4252 1760
rect 4304 1708 4310 1760
rect 6914 1708 6920 1760
rect 6972 1708 6978 1760
rect 7650 1708 7656 1760
rect 7708 1708 7714 1760
rect 7742 1708 7748 1760
rect 7800 1748 7806 1760
rect 8110 1748 8116 1760
rect 7800 1720 8116 1748
rect 7800 1708 7806 1720
rect 8110 1708 8116 1720
rect 8168 1708 8174 1760
rect 8205 1751 8263 1757
rect 8205 1717 8217 1751
rect 8251 1748 8263 1751
rect 8754 1748 8760 1760
rect 8251 1720 8760 1748
rect 8251 1717 8263 1720
rect 8205 1711 8263 1717
rect 8754 1708 8760 1720
rect 8812 1708 8818 1760
rect 10244 1757 10272 1788
rect 11606 1776 11612 1788
rect 11664 1776 11670 1828
rect 12268 1816 12296 1847
rect 13078 1844 13084 1896
rect 13136 1884 13142 1896
rect 15764 1893 15792 1924
rect 16114 1912 16120 1964
rect 16172 1952 16178 1964
rect 16301 1955 16359 1961
rect 16301 1952 16313 1955
rect 16172 1924 16313 1952
rect 16172 1912 16178 1924
rect 16301 1921 16313 1924
rect 16347 1921 16359 1955
rect 16301 1915 16359 1921
rect 16393 1955 16451 1961
rect 16393 1921 16405 1955
rect 16439 1952 16451 1955
rect 16945 1955 17003 1961
rect 16945 1952 16957 1955
rect 16439 1924 16957 1952
rect 16439 1921 16451 1924
rect 16393 1915 16451 1921
rect 16945 1921 16957 1924
rect 16991 1921 17003 1955
rect 16945 1915 17003 1921
rect 17034 1912 17040 1964
rect 17092 1952 17098 1964
rect 20717 1955 20775 1961
rect 20717 1952 20729 1955
rect 17092 1924 20729 1952
rect 17092 1912 17098 1924
rect 20717 1921 20729 1924
rect 20763 1921 20775 1955
rect 21269 1955 21327 1961
rect 21269 1952 21281 1955
rect 20717 1915 20775 1921
rect 20916 1924 21281 1952
rect 15657 1887 15715 1893
rect 15657 1884 15669 1887
rect 13136 1856 15669 1884
rect 13136 1844 13142 1856
rect 15657 1853 15669 1856
rect 15703 1853 15715 1887
rect 15657 1847 15715 1853
rect 15749 1887 15807 1893
rect 15749 1853 15761 1887
rect 15795 1853 15807 1887
rect 15749 1847 15807 1853
rect 15838 1844 15844 1896
rect 15896 1844 15902 1896
rect 15930 1844 15936 1896
rect 15988 1884 15994 1896
rect 16025 1887 16083 1893
rect 16025 1884 16037 1887
rect 15988 1856 16037 1884
rect 15988 1844 15994 1856
rect 16025 1853 16037 1856
rect 16071 1853 16083 1887
rect 16025 1847 16083 1853
rect 16209 1887 16267 1893
rect 16209 1853 16221 1887
rect 16255 1853 16267 1887
rect 16209 1847 16267 1853
rect 16485 1887 16543 1893
rect 16485 1853 16497 1887
rect 16531 1853 16543 1887
rect 16485 1847 16543 1853
rect 13096 1816 13124 1844
rect 12268 1788 13124 1816
rect 13262 1776 13268 1828
rect 13320 1816 13326 1828
rect 13725 1819 13783 1825
rect 13725 1816 13737 1819
rect 13320 1788 13737 1816
rect 13320 1776 13326 1788
rect 13725 1785 13737 1788
rect 13771 1816 13783 1819
rect 13998 1816 14004 1828
rect 13771 1788 14004 1816
rect 13771 1785 13783 1788
rect 13725 1779 13783 1785
rect 13998 1776 14004 1788
rect 14056 1776 14062 1828
rect 14550 1776 14556 1828
rect 14608 1816 14614 1828
rect 14608 1788 15240 1816
rect 14608 1776 14614 1788
rect 15212 1760 15240 1788
rect 15286 1776 15292 1828
rect 15344 1816 15350 1828
rect 16224 1816 16252 1847
rect 15344 1788 16252 1816
rect 16500 1816 16528 1847
rect 16758 1844 16764 1896
rect 16816 1884 16822 1896
rect 17129 1887 17187 1893
rect 17129 1884 17141 1887
rect 16816 1856 17141 1884
rect 16816 1844 16822 1856
rect 17129 1853 17141 1856
rect 17175 1884 17187 1887
rect 17397 1889 17455 1895
rect 17397 1886 17409 1889
rect 17328 1884 17409 1886
rect 17175 1858 17409 1884
rect 17175 1856 17356 1858
rect 17175 1853 17187 1856
rect 17129 1847 17187 1853
rect 17397 1855 17409 1858
rect 17443 1855 17455 1889
rect 17397 1849 17455 1855
rect 17589 1887 17647 1893
rect 17589 1853 17601 1887
rect 17635 1884 17647 1887
rect 17635 1856 17724 1884
rect 17635 1853 17647 1856
rect 17589 1847 17647 1853
rect 17313 1819 17371 1825
rect 16500 1788 16804 1816
rect 15344 1776 15350 1788
rect 10229 1751 10287 1757
rect 10229 1717 10241 1751
rect 10275 1717 10287 1751
rect 10229 1711 10287 1717
rect 10318 1708 10324 1760
rect 10376 1748 10382 1760
rect 10873 1751 10931 1757
rect 10873 1748 10885 1751
rect 10376 1720 10885 1748
rect 10376 1708 10382 1720
rect 10873 1717 10885 1720
rect 10919 1717 10931 1751
rect 10873 1711 10931 1717
rect 11054 1708 11060 1760
rect 11112 1748 11118 1760
rect 13173 1751 13231 1757
rect 13173 1748 13185 1751
rect 11112 1720 13185 1748
rect 11112 1708 11118 1720
rect 13173 1717 13185 1720
rect 13219 1717 13231 1751
rect 13173 1711 13231 1717
rect 13446 1708 13452 1760
rect 13504 1748 13510 1760
rect 13633 1751 13691 1757
rect 13633 1748 13645 1751
rect 13504 1720 13645 1748
rect 13504 1708 13510 1720
rect 13633 1717 13645 1720
rect 13679 1717 13691 1751
rect 13633 1711 13691 1717
rect 14642 1708 14648 1760
rect 14700 1748 14706 1760
rect 15010 1748 15016 1760
rect 14700 1720 15016 1748
rect 14700 1708 14706 1720
rect 15010 1708 15016 1720
rect 15068 1708 15074 1760
rect 15194 1708 15200 1760
rect 15252 1708 15258 1760
rect 15378 1708 15384 1760
rect 15436 1708 15442 1760
rect 15470 1708 15476 1760
rect 15528 1748 15534 1760
rect 16669 1751 16727 1757
rect 16669 1748 16681 1751
rect 15528 1720 16681 1748
rect 15528 1708 15534 1720
rect 16669 1717 16681 1720
rect 16715 1717 16727 1751
rect 16776 1748 16804 1788
rect 17313 1785 17325 1819
rect 17359 1816 17371 1819
rect 17696 1816 17724 1856
rect 17862 1844 17868 1896
rect 17920 1844 17926 1896
rect 20916 1893 20944 1924
rect 21269 1921 21281 1924
rect 21315 1921 21327 1955
rect 21269 1915 21327 1921
rect 21468 1893 21496 1992
rect 21637 1955 21695 1961
rect 21637 1921 21649 1955
rect 21683 1952 21695 1955
rect 21744 1952 21772 2048
rect 22186 1980 22192 2032
rect 22244 1980 22250 2032
rect 22094 1952 22100 1964
rect 21683 1924 21772 1952
rect 21836 1924 22100 1952
rect 21683 1921 21695 1924
rect 21637 1915 21695 1921
rect 18049 1887 18107 1893
rect 18049 1853 18061 1887
rect 18095 1853 18107 1887
rect 18049 1847 18107 1853
rect 19153 1887 19211 1893
rect 19153 1853 19165 1887
rect 19199 1884 19211 1887
rect 20901 1887 20959 1893
rect 19199 1856 19380 1884
rect 19199 1853 19211 1856
rect 19153 1847 19211 1853
rect 18064 1816 18092 1847
rect 17359 1788 18092 1816
rect 17359 1785 17371 1788
rect 17313 1779 17371 1785
rect 18064 1760 18092 1788
rect 18417 1819 18475 1825
rect 18417 1785 18429 1819
rect 18463 1816 18475 1819
rect 18463 1788 18736 1816
rect 18463 1785 18475 1788
rect 18417 1779 18475 1785
rect 17405 1751 17463 1757
rect 17405 1748 17417 1751
rect 16776 1720 17417 1748
rect 16669 1711 16727 1717
rect 17405 1717 17417 1720
rect 17451 1717 17463 1751
rect 17405 1711 17463 1717
rect 18046 1708 18052 1760
rect 18104 1708 18110 1760
rect 18708 1757 18736 1788
rect 19352 1760 19380 1856
rect 20901 1853 20913 1887
rect 20947 1853 20959 1887
rect 20901 1847 20959 1853
rect 21177 1887 21235 1893
rect 21177 1853 21189 1887
rect 21223 1853 21235 1887
rect 21177 1847 21235 1853
rect 21453 1887 21511 1893
rect 21453 1853 21465 1887
rect 21499 1853 21511 1887
rect 21453 1847 21511 1853
rect 21192 1816 21220 1847
rect 21836 1816 21864 1924
rect 22094 1912 22100 1924
rect 22152 1912 22158 1964
rect 21910 1844 21916 1896
rect 21968 1844 21974 1896
rect 22204 1887 22232 1980
rect 22197 1881 22255 1887
rect 22197 1847 22209 1881
rect 22243 1847 22255 1881
rect 22197 1841 22255 1847
rect 21192 1788 21864 1816
rect 18693 1751 18751 1757
rect 18693 1717 18705 1751
rect 18739 1717 18751 1751
rect 18693 1711 18751 1717
rect 19334 1708 19340 1760
rect 19392 1708 19398 1760
rect 21082 1708 21088 1760
rect 21140 1748 21146 1760
rect 22097 1751 22155 1757
rect 22097 1748 22109 1751
rect 21140 1720 22109 1748
rect 21140 1708 21146 1720
rect 22097 1717 22109 1720
rect 22143 1717 22155 1751
rect 22097 1711 22155 1717
rect 552 1658 23368 1680
rect 552 1606 4366 1658
rect 4418 1606 4430 1658
rect 4482 1606 4494 1658
rect 4546 1606 4558 1658
rect 4610 1606 4622 1658
rect 4674 1606 4686 1658
rect 4738 1606 10366 1658
rect 10418 1606 10430 1658
rect 10482 1606 10494 1658
rect 10546 1606 10558 1658
rect 10610 1606 10622 1658
rect 10674 1606 10686 1658
rect 10738 1606 16366 1658
rect 16418 1606 16430 1658
rect 16482 1606 16494 1658
rect 16546 1606 16558 1658
rect 16610 1606 16622 1658
rect 16674 1606 16686 1658
rect 16738 1606 22366 1658
rect 22418 1606 22430 1658
rect 22482 1606 22494 1658
rect 22546 1606 22558 1658
rect 22610 1606 22622 1658
rect 22674 1606 22686 1658
rect 22738 1606 23368 1658
rect 552 1584 23368 1606
rect 1118 1504 1124 1556
rect 1176 1504 1182 1556
rect 1210 1504 1216 1556
rect 1268 1504 1274 1556
rect 3694 1544 3700 1556
rect 1964 1516 3700 1544
rect 1136 1408 1164 1504
rect 1228 1476 1256 1504
rect 1964 1485 1992 1516
rect 3694 1504 3700 1516
rect 3752 1504 3758 1556
rect 3786 1504 3792 1556
rect 3844 1504 3850 1556
rect 3878 1504 3884 1556
rect 3936 1504 3942 1556
rect 4154 1504 4160 1556
rect 4212 1544 4218 1556
rect 4525 1547 4583 1553
rect 4525 1544 4537 1547
rect 4212 1516 4537 1544
rect 4212 1504 4218 1516
rect 4525 1513 4537 1516
rect 4571 1513 4583 1547
rect 4525 1507 4583 1513
rect 6914 1504 6920 1556
rect 6972 1544 6978 1556
rect 7745 1547 7803 1553
rect 6972 1516 7512 1544
rect 6972 1504 6978 1516
rect 1949 1479 2007 1485
rect 1228 1448 1348 1476
rect 1213 1411 1271 1417
rect 1213 1408 1225 1411
rect 1136 1380 1225 1408
rect 1213 1377 1225 1380
rect 1259 1377 1271 1411
rect 1213 1371 1271 1377
rect 1320 1340 1348 1448
rect 1949 1445 1961 1479
rect 1995 1445 2007 1479
rect 1949 1439 2007 1445
rect 2492 1479 2550 1485
rect 2492 1445 2504 1479
rect 2538 1476 2550 1479
rect 3804 1476 3832 1504
rect 2538 1448 3832 1476
rect 2538 1445 2550 1448
rect 2492 1439 2550 1445
rect 3896 1417 3924 1504
rect 5718 1436 5724 1488
rect 5776 1476 5782 1488
rect 5776 1448 7236 1476
rect 5776 1436 5782 1448
rect 3881 1411 3939 1417
rect 3881 1408 3893 1411
rect 3620 1380 3893 1408
rect 2225 1343 2283 1349
rect 2225 1340 2237 1343
rect 1320 1312 2237 1340
rect 2225 1309 2237 1312
rect 2271 1309 2283 1343
rect 2225 1303 2283 1309
rect 1762 1232 1768 1284
rect 1820 1232 1826 1284
rect 3620 1281 3648 1380
rect 3881 1377 3893 1380
rect 3927 1377 3939 1411
rect 4341 1411 4399 1417
rect 4341 1408 4353 1411
rect 3881 1371 3939 1377
rect 4172 1380 4353 1408
rect 4172 1352 4200 1380
rect 4341 1377 4353 1380
rect 4387 1377 4399 1411
rect 4341 1371 4399 1377
rect 4985 1411 5043 1417
rect 4985 1377 4997 1411
rect 5031 1408 5043 1411
rect 5442 1408 5448 1420
rect 5031 1380 5448 1408
rect 5031 1377 5043 1380
rect 4985 1371 5043 1377
rect 5442 1368 5448 1380
rect 5500 1368 5506 1420
rect 3973 1343 4031 1349
rect 3973 1309 3985 1343
rect 4019 1340 4031 1343
rect 4154 1340 4160 1352
rect 4019 1312 4160 1340
rect 4019 1309 4031 1312
rect 3973 1303 4031 1309
rect 4154 1300 4160 1312
rect 4212 1300 4218 1352
rect 4246 1300 4252 1352
rect 4304 1340 4310 1352
rect 4893 1343 4951 1349
rect 4893 1340 4905 1343
rect 4304 1312 4905 1340
rect 4304 1300 4310 1312
rect 4893 1309 4905 1312
rect 4939 1309 4951 1343
rect 4893 1303 4951 1309
rect 3605 1275 3663 1281
rect 3605 1241 3617 1275
rect 3651 1241 3663 1275
rect 3605 1235 3663 1241
rect 5353 1275 5411 1281
rect 5353 1241 5365 1275
rect 5399 1272 5411 1275
rect 5736 1272 5764 1436
rect 6380 1417 6408 1448
rect 6365 1411 6423 1417
rect 6365 1377 6377 1411
rect 6411 1377 6423 1411
rect 6365 1371 6423 1377
rect 6457 1411 6515 1417
rect 6457 1377 6469 1411
rect 6503 1408 6515 1411
rect 6641 1411 6699 1417
rect 6503 1380 6592 1408
rect 6503 1377 6515 1380
rect 6457 1371 6515 1377
rect 6564 1340 6592 1380
rect 6641 1377 6653 1411
rect 6687 1408 6699 1411
rect 6914 1408 6920 1420
rect 6687 1380 6920 1408
rect 6687 1377 6699 1380
rect 6641 1371 6699 1377
rect 6914 1368 6920 1380
rect 6972 1368 6978 1420
rect 7006 1368 7012 1420
rect 7064 1368 7070 1420
rect 7208 1417 7236 1448
rect 7282 1436 7288 1488
rect 7340 1436 7346 1488
rect 7101 1411 7159 1417
rect 7101 1377 7113 1411
rect 7147 1377 7159 1411
rect 7101 1371 7159 1377
rect 7193 1411 7251 1417
rect 7193 1377 7205 1411
rect 7239 1377 7251 1411
rect 7300 1408 7328 1436
rect 7377 1411 7435 1417
rect 7377 1408 7389 1411
rect 7300 1380 7389 1408
rect 7193 1371 7251 1377
rect 7377 1377 7389 1380
rect 7423 1377 7435 1411
rect 7484 1408 7512 1516
rect 7745 1513 7757 1547
rect 7791 1544 7803 1547
rect 7834 1544 7840 1556
rect 7791 1516 7840 1544
rect 7791 1513 7803 1516
rect 7745 1507 7803 1513
rect 7834 1504 7840 1516
rect 7892 1504 7898 1556
rect 9030 1504 9036 1556
rect 9088 1504 9094 1556
rect 9858 1544 9864 1556
rect 9140 1516 9864 1544
rect 9140 1476 9168 1516
rect 9858 1504 9864 1516
rect 9916 1504 9922 1556
rect 10870 1544 10876 1556
rect 9968 1516 10876 1544
rect 9968 1476 9996 1516
rect 10870 1504 10876 1516
rect 10928 1504 10934 1556
rect 11146 1504 11152 1556
rect 11204 1504 11210 1556
rect 13262 1544 13268 1556
rect 12406 1516 13268 1544
rect 8220 1448 9168 1476
rect 9232 1448 9996 1476
rect 8220 1417 8248 1448
rect 7929 1411 7987 1417
rect 7929 1408 7941 1411
rect 7484 1380 7941 1408
rect 7377 1371 7435 1377
rect 7929 1377 7941 1380
rect 7975 1377 7987 1411
rect 7929 1371 7987 1377
rect 8205 1411 8263 1417
rect 8205 1377 8217 1411
rect 8251 1377 8263 1411
rect 8205 1371 8263 1377
rect 7024 1340 7052 1368
rect 6564 1312 7052 1340
rect 7116 1340 7144 1371
rect 8386 1368 8392 1420
rect 8444 1368 8450 1420
rect 8570 1368 8576 1420
rect 8628 1368 8634 1420
rect 9232 1417 9260 1448
rect 9217 1411 9275 1417
rect 9217 1377 9229 1411
rect 9263 1377 9275 1411
rect 9217 1371 9275 1377
rect 9398 1368 9404 1420
rect 9456 1368 9462 1420
rect 9490 1368 9496 1420
rect 9548 1368 9554 1420
rect 9968 1417 9996 1448
rect 10428 1448 11008 1476
rect 9953 1411 10011 1417
rect 9953 1377 9965 1411
rect 9999 1377 10011 1411
rect 9953 1371 10011 1377
rect 10134 1368 10140 1420
rect 10192 1368 10198 1420
rect 10428 1417 10456 1448
rect 10980 1420 11008 1448
rect 10413 1411 10471 1417
rect 10413 1377 10425 1411
rect 10459 1377 10471 1411
rect 10413 1371 10471 1377
rect 10597 1411 10655 1417
rect 10597 1377 10609 1411
rect 10643 1377 10655 1411
rect 10597 1371 10655 1377
rect 7285 1343 7343 1349
rect 7285 1340 7297 1343
rect 7116 1312 7297 1340
rect 7285 1309 7297 1312
rect 7331 1309 7343 1343
rect 7285 1303 7343 1309
rect 7558 1300 7564 1352
rect 7616 1300 7622 1352
rect 7650 1300 7656 1352
rect 7708 1340 7714 1352
rect 8113 1343 8171 1349
rect 8113 1340 8125 1343
rect 7708 1312 8125 1340
rect 7708 1300 7714 1312
rect 8113 1309 8125 1312
rect 8159 1340 8171 1343
rect 8404 1340 8432 1368
rect 8159 1312 8432 1340
rect 8849 1343 8907 1349
rect 8159 1309 8171 1312
rect 8113 1303 8171 1309
rect 8849 1309 8861 1343
rect 8895 1340 8907 1343
rect 9508 1340 9536 1368
rect 8895 1312 9536 1340
rect 8895 1309 8907 1312
rect 8849 1303 8907 1309
rect 9766 1300 9772 1352
rect 9824 1340 9830 1352
rect 10229 1343 10287 1349
rect 10229 1340 10241 1343
rect 9824 1312 10241 1340
rect 9824 1300 9830 1312
rect 10229 1309 10241 1312
rect 10275 1340 10287 1343
rect 10321 1343 10379 1349
rect 10321 1340 10333 1343
rect 10275 1312 10333 1340
rect 10275 1309 10287 1312
rect 10229 1303 10287 1309
rect 10321 1309 10333 1312
rect 10367 1340 10379 1343
rect 10502 1340 10508 1352
rect 10367 1312 10508 1340
rect 10367 1309 10379 1312
rect 10321 1303 10379 1309
rect 10502 1300 10508 1312
rect 10560 1300 10566 1352
rect 10612 1340 10640 1371
rect 10962 1368 10968 1420
rect 11020 1368 11026 1420
rect 11164 1408 11192 1504
rect 12406 1476 12434 1516
rect 13262 1504 13268 1516
rect 13320 1504 13326 1556
rect 13538 1504 13544 1556
rect 13596 1544 13602 1556
rect 15470 1544 15476 1556
rect 13596 1516 15476 1544
rect 13596 1504 13602 1516
rect 15470 1504 15476 1516
rect 15528 1504 15534 1556
rect 15654 1504 15660 1556
rect 15712 1544 15718 1556
rect 15712 1516 16896 1544
rect 15712 1504 15718 1516
rect 11532 1448 12480 1476
rect 11333 1411 11391 1417
rect 11333 1408 11345 1411
rect 11164 1380 11345 1408
rect 11333 1377 11345 1380
rect 11379 1377 11391 1411
rect 11333 1371 11391 1377
rect 11422 1368 11428 1420
rect 11480 1368 11486 1420
rect 11532 1417 11560 1448
rect 11517 1411 11575 1417
rect 11517 1377 11529 1411
rect 11563 1377 11575 1411
rect 11517 1371 11575 1377
rect 11606 1368 11612 1420
rect 11664 1408 11670 1420
rect 11701 1411 11759 1417
rect 11701 1408 11713 1411
rect 11664 1380 11713 1408
rect 11664 1368 11670 1380
rect 11701 1377 11713 1380
rect 11747 1377 11759 1411
rect 11701 1371 11759 1377
rect 12250 1368 12256 1420
rect 12308 1368 12314 1420
rect 12452 1417 12480 1448
rect 13998 1436 14004 1488
rect 14056 1476 14062 1488
rect 14056 1448 14320 1476
rect 14056 1436 14062 1448
rect 12437 1411 12495 1417
rect 12437 1377 12449 1411
rect 12483 1377 12495 1411
rect 12437 1371 12495 1377
rect 13173 1411 13231 1417
rect 13173 1377 13185 1411
rect 13219 1408 13231 1411
rect 13725 1411 13783 1417
rect 13725 1408 13737 1411
rect 13219 1380 13737 1408
rect 13219 1377 13231 1380
rect 13173 1371 13231 1377
rect 13725 1377 13737 1380
rect 13771 1408 13783 1411
rect 13814 1408 13820 1420
rect 13771 1380 13820 1408
rect 13771 1377 13783 1380
rect 13725 1371 13783 1377
rect 13814 1368 13820 1380
rect 13872 1368 13878 1420
rect 13909 1411 13967 1417
rect 13909 1377 13921 1411
rect 13955 1408 13967 1411
rect 14090 1408 14096 1420
rect 13955 1380 14096 1408
rect 13955 1377 13967 1380
rect 13909 1371 13967 1377
rect 14090 1368 14096 1380
rect 14148 1368 14154 1420
rect 14292 1417 14320 1448
rect 14568 1448 15976 1476
rect 14568 1417 14596 1448
rect 15948 1420 15976 1448
rect 14277 1411 14335 1417
rect 14277 1377 14289 1411
rect 14323 1377 14335 1411
rect 14277 1371 14335 1377
rect 14553 1411 14611 1417
rect 14553 1377 14565 1411
rect 14599 1377 14611 1411
rect 14553 1371 14611 1377
rect 14734 1368 14740 1420
rect 14792 1368 14798 1420
rect 14918 1368 14924 1420
rect 14976 1368 14982 1420
rect 15194 1368 15200 1420
rect 15252 1368 15258 1420
rect 15562 1368 15568 1420
rect 15620 1368 15626 1420
rect 15746 1368 15752 1420
rect 15804 1368 15810 1420
rect 15930 1368 15936 1420
rect 15988 1368 15994 1420
rect 16206 1368 16212 1420
rect 16264 1368 16270 1420
rect 16390 1368 16396 1420
rect 16448 1368 16454 1420
rect 16758 1368 16764 1420
rect 16816 1368 16822 1420
rect 16868 1408 16896 1516
rect 17126 1504 17132 1556
rect 17184 1544 17190 1556
rect 17184 1516 17816 1544
rect 17184 1504 17190 1516
rect 17052 1448 17724 1476
rect 16945 1411 17003 1417
rect 16945 1408 16957 1411
rect 16868 1380 16957 1408
rect 16945 1377 16957 1380
rect 16991 1408 17003 1411
rect 17052 1408 17080 1448
rect 17696 1420 17724 1448
rect 16991 1380 17080 1408
rect 16991 1377 17003 1380
rect 16945 1371 17003 1377
rect 17218 1368 17224 1420
rect 17276 1368 17282 1420
rect 17402 1368 17408 1420
rect 17460 1408 17466 1420
rect 17589 1411 17647 1417
rect 17589 1408 17601 1411
rect 17460 1380 17601 1408
rect 17460 1368 17466 1380
rect 17589 1377 17601 1380
rect 17635 1377 17647 1411
rect 17589 1371 17647 1377
rect 17678 1368 17684 1420
rect 17736 1368 17742 1420
rect 17788 1417 17816 1516
rect 19886 1504 19892 1556
rect 19944 1504 19950 1556
rect 22370 1504 22376 1556
rect 22428 1544 22434 1556
rect 22649 1547 22707 1553
rect 22649 1544 22661 1547
rect 22428 1516 22661 1544
rect 22428 1504 22434 1516
rect 22649 1513 22661 1516
rect 22695 1513 22707 1547
rect 22649 1507 22707 1513
rect 18046 1436 18052 1488
rect 18104 1436 18110 1488
rect 17773 1411 17831 1417
rect 17773 1377 17785 1411
rect 17819 1377 17831 1411
rect 19334 1408 19340 1420
rect 18998 1380 19340 1408
rect 17773 1371 17831 1377
rect 19334 1368 19340 1380
rect 19392 1408 19398 1420
rect 19794 1408 19800 1420
rect 19392 1380 19800 1408
rect 19392 1368 19398 1380
rect 19794 1368 19800 1380
rect 19852 1368 19858 1420
rect 19904 1408 19932 1504
rect 22094 1436 22100 1488
rect 22152 1436 22158 1488
rect 21456 1420 21508 1426
rect 19961 1411 20019 1417
rect 19961 1408 19973 1411
rect 19904 1380 19973 1408
rect 19961 1377 19973 1380
rect 20007 1377 20019 1411
rect 21358 1408 21364 1420
rect 19961 1371 20019 1377
rect 20732 1380 21364 1408
rect 12161 1343 12219 1349
rect 12161 1340 12173 1343
rect 10612 1312 11376 1340
rect 5399 1244 5764 1272
rect 7576 1272 7604 1300
rect 11348 1284 11376 1312
rect 11624 1312 12173 1340
rect 8021 1275 8079 1281
rect 8021 1272 8033 1275
rect 7576 1244 8033 1272
rect 5399 1241 5411 1244
rect 5353 1235 5411 1241
rect 8021 1241 8033 1244
rect 8067 1241 8079 1275
rect 8021 1235 8079 1241
rect 8202 1232 8208 1284
rect 8260 1272 8266 1284
rect 11057 1275 11115 1281
rect 11057 1272 11069 1275
rect 8260 1244 11069 1272
rect 8260 1232 8266 1244
rect 11057 1241 11069 1244
rect 11103 1241 11115 1275
rect 11057 1235 11115 1241
rect 11330 1232 11336 1284
rect 11388 1232 11394 1284
rect 11624 1216 11652 1312
rect 12161 1309 12173 1312
rect 12207 1340 12219 1343
rect 12207 1312 12434 1340
rect 12207 1309 12219 1312
rect 12161 1303 12219 1309
rect 12406 1272 12434 1312
rect 12710 1300 12716 1352
rect 12768 1340 12774 1352
rect 13446 1340 13452 1352
rect 12768 1312 13452 1340
rect 12768 1300 12774 1312
rect 13446 1300 13452 1312
rect 13504 1300 13510 1352
rect 14001 1343 14059 1349
rect 14001 1309 14013 1343
rect 14047 1340 14059 1343
rect 14829 1343 14887 1349
rect 14829 1340 14841 1343
rect 14047 1312 14841 1340
rect 14047 1309 14059 1312
rect 14001 1303 14059 1309
rect 14829 1309 14841 1312
rect 14875 1309 14887 1343
rect 15473 1343 15531 1349
rect 15473 1340 15485 1343
rect 14829 1303 14887 1309
rect 15396 1312 15485 1340
rect 14016 1272 14044 1303
rect 15396 1281 15424 1312
rect 15473 1309 15485 1312
rect 15519 1340 15531 1343
rect 16114 1340 16120 1352
rect 15519 1312 16120 1340
rect 15519 1309 15531 1312
rect 15473 1303 15531 1309
rect 16114 1300 16120 1312
rect 16172 1340 16178 1352
rect 16669 1343 16727 1349
rect 16669 1340 16681 1343
rect 16172 1312 16681 1340
rect 16172 1300 16178 1312
rect 16669 1309 16681 1312
rect 16715 1309 16727 1343
rect 17497 1343 17555 1349
rect 17497 1340 17509 1343
rect 16669 1303 16727 1309
rect 16776 1312 17509 1340
rect 14093 1275 14151 1281
rect 14093 1272 14105 1275
rect 12406 1244 14105 1272
rect 14093 1241 14105 1244
rect 14139 1241 14151 1275
rect 14093 1235 14151 1241
rect 15381 1275 15439 1281
rect 15381 1241 15393 1275
rect 15427 1241 15439 1275
rect 15381 1235 15439 1241
rect 15746 1232 15752 1284
rect 15804 1272 15810 1284
rect 16776 1272 16804 1312
rect 17497 1309 17509 1312
rect 17543 1340 17555 1343
rect 18690 1340 18696 1352
rect 17543 1312 18696 1340
rect 17543 1309 17555 1312
rect 17497 1303 17555 1309
rect 18690 1300 18696 1312
rect 18748 1300 18754 1352
rect 18874 1300 18880 1352
rect 18932 1300 18938 1352
rect 19705 1343 19763 1349
rect 19705 1309 19717 1343
rect 19751 1309 19763 1343
rect 19705 1303 19763 1309
rect 15804 1244 16804 1272
rect 17129 1275 17187 1281
rect 15804 1232 15810 1244
rect 17129 1241 17141 1275
rect 17175 1272 17187 1275
rect 19058 1272 19064 1284
rect 17175 1244 19064 1272
rect 17175 1241 17187 1244
rect 17129 1235 17187 1241
rect 19058 1232 19064 1244
rect 19116 1232 19122 1284
rect 14 1164 20 1216
rect 72 1204 78 1216
rect 937 1207 995 1213
rect 937 1204 949 1207
rect 72 1176 949 1204
rect 72 1164 78 1176
rect 937 1173 949 1176
rect 983 1173 995 1207
rect 937 1167 995 1173
rect 7101 1207 7159 1213
rect 7101 1173 7113 1207
rect 7147 1204 7159 1207
rect 8294 1204 8300 1216
rect 7147 1176 8300 1204
rect 7147 1173 7159 1176
rect 7101 1167 7159 1173
rect 8294 1164 8300 1176
rect 8352 1164 8358 1216
rect 8386 1164 8392 1216
rect 8444 1164 8450 1216
rect 8754 1164 8760 1216
rect 8812 1164 8818 1216
rect 9766 1164 9772 1216
rect 9824 1164 9830 1216
rect 10778 1164 10784 1216
rect 10836 1164 10842 1216
rect 11606 1164 11612 1216
rect 11664 1164 11670 1216
rect 12618 1164 12624 1216
rect 12676 1164 12682 1216
rect 12986 1164 12992 1216
rect 13044 1164 13050 1216
rect 13357 1207 13415 1213
rect 13357 1173 13369 1207
rect 13403 1204 13415 1207
rect 13446 1204 13452 1216
rect 13403 1176 13452 1204
rect 13403 1173 13415 1176
rect 13357 1167 13415 1173
rect 13446 1164 13452 1176
rect 13504 1164 13510 1216
rect 13541 1207 13599 1213
rect 13541 1173 13553 1207
rect 13587 1204 13599 1207
rect 13814 1204 13820 1216
rect 13587 1176 13820 1204
rect 13587 1173 13599 1176
rect 13541 1167 13599 1173
rect 13814 1164 13820 1176
rect 13872 1164 13878 1216
rect 14366 1164 14372 1216
rect 14424 1164 14430 1216
rect 15102 1164 15108 1216
rect 15160 1164 15166 1216
rect 15930 1164 15936 1216
rect 15988 1164 15994 1216
rect 16574 1164 16580 1216
rect 16632 1164 16638 1216
rect 17402 1164 17408 1216
rect 17460 1164 17466 1216
rect 17954 1164 17960 1216
rect 18012 1164 18018 1216
rect 19720 1204 19748 1303
rect 20732 1204 20760 1380
rect 21358 1368 21364 1380
rect 21416 1368 21422 1420
rect 22465 1411 22523 1417
rect 22465 1408 22477 1411
rect 21456 1362 21508 1368
rect 22112 1380 22477 1408
rect 21545 1343 21603 1349
rect 21545 1309 21557 1343
rect 21591 1340 21603 1343
rect 21910 1340 21916 1352
rect 21591 1312 21916 1340
rect 21591 1309 21603 1312
rect 21545 1303 21603 1309
rect 21085 1275 21143 1281
rect 21085 1241 21097 1275
rect 21131 1272 21143 1275
rect 21560 1272 21588 1303
rect 21910 1300 21916 1312
rect 21968 1300 21974 1352
rect 22112 1340 22140 1380
rect 22465 1377 22477 1380
rect 22511 1377 22523 1411
rect 22465 1371 22523 1377
rect 22066 1312 22140 1340
rect 21131 1244 21588 1272
rect 21131 1241 21143 1244
rect 21085 1235 21143 1241
rect 21634 1232 21640 1284
rect 21692 1272 21698 1284
rect 22066 1272 22094 1312
rect 21692 1244 22094 1272
rect 21692 1232 21698 1244
rect 19720 1176 20760 1204
rect 552 1114 23368 1136
rect 552 1062 1366 1114
rect 1418 1062 1430 1114
rect 1482 1062 1494 1114
rect 1546 1062 1558 1114
rect 1610 1062 1622 1114
rect 1674 1062 1686 1114
rect 1738 1062 7366 1114
rect 7418 1062 7430 1114
rect 7482 1062 7494 1114
rect 7546 1062 7558 1114
rect 7610 1062 7622 1114
rect 7674 1062 7686 1114
rect 7738 1062 13366 1114
rect 13418 1062 13430 1114
rect 13482 1062 13494 1114
rect 13546 1062 13558 1114
rect 13610 1062 13622 1114
rect 13674 1062 13686 1114
rect 13738 1062 19366 1114
rect 19418 1062 19430 1114
rect 19482 1062 19494 1114
rect 19546 1062 19558 1114
rect 19610 1062 19622 1114
rect 19674 1062 19686 1114
rect 19738 1062 23368 1114
rect 552 1040 23368 1062
rect 1210 960 1216 1012
rect 1268 960 1274 1012
rect 2777 1003 2835 1009
rect 2777 969 2789 1003
rect 2823 1000 2835 1003
rect 4154 1000 4160 1012
rect 2823 972 4160 1000
rect 2823 969 2835 972
rect 2777 963 2835 969
rect 4154 960 4160 972
rect 4212 960 4218 1012
rect 8312 972 9720 1000
rect 1228 864 1256 960
rect 8202 932 8208 944
rect 4540 904 8208 932
rect 1397 867 1455 873
rect 1397 864 1409 867
rect 1228 836 1409 864
rect 1397 833 1409 836
rect 1443 833 1455 867
rect 1397 827 1455 833
rect 1026 756 1032 808
rect 1084 796 1090 808
rect 4540 805 4568 904
rect 8202 892 8208 904
rect 8260 892 8266 944
rect 8312 864 8340 972
rect 8386 892 8392 944
rect 8444 892 8450 944
rect 9033 935 9091 941
rect 9033 901 9045 935
rect 9079 901 9091 935
rect 9033 895 9091 901
rect 5368 836 8340 864
rect 5368 805 5396 836
rect 1213 799 1271 805
rect 1213 796 1225 799
rect 1084 768 1225 796
rect 1084 756 1090 768
rect 1213 765 1225 768
rect 1259 765 1271 799
rect 1213 759 1271 765
rect 3513 799 3571 805
rect 3513 765 3525 799
rect 3559 796 3571 799
rect 4525 799 4583 805
rect 3559 768 4476 796
rect 3559 765 3571 768
rect 3513 759 3571 765
rect 1664 731 1722 737
rect 1664 697 1676 731
rect 1710 728 1722 731
rect 1854 728 1860 740
rect 1710 700 1860 728
rect 1710 697 1722 700
rect 1664 691 1722 697
rect 1854 688 1860 700
rect 1912 688 1918 740
rect 2498 688 2504 740
rect 2556 728 2562 740
rect 3605 731 3663 737
rect 3605 728 3617 731
rect 2556 700 3617 728
rect 2556 688 2562 700
rect 3605 697 3617 700
rect 3651 697 3663 731
rect 3605 691 3663 697
rect 3973 731 4031 737
rect 3973 697 3985 731
rect 4019 697 4031 731
rect 4448 728 4476 768
rect 4525 765 4537 799
rect 4571 765 4583 799
rect 4525 759 4583 765
rect 5353 799 5411 805
rect 5353 765 5365 799
rect 5399 765 5411 799
rect 5353 759 5411 765
rect 6178 756 6184 808
rect 6236 756 6242 808
rect 8404 728 8432 892
rect 8665 799 8723 805
rect 8665 765 8677 799
rect 8711 765 8723 799
rect 8665 759 8723 765
rect 4448 700 8432 728
rect 8680 728 8708 759
rect 8846 756 8852 808
rect 8904 756 8910 808
rect 9048 796 9076 895
rect 9217 799 9275 805
rect 9217 796 9229 799
rect 9048 768 9229 796
rect 9217 765 9229 768
rect 9263 765 9275 799
rect 9217 759 9275 765
rect 9692 728 9720 972
rect 9766 960 9772 1012
rect 9824 960 9830 1012
rect 10778 960 10784 1012
rect 10836 960 10842 1012
rect 11701 1003 11759 1009
rect 11701 969 11713 1003
rect 11747 1000 11759 1003
rect 12066 1000 12072 1012
rect 11747 972 12072 1000
rect 11747 969 11759 972
rect 11701 963 11759 969
rect 12066 960 12072 972
rect 12124 960 12130 1012
rect 12618 960 12624 1012
rect 12676 960 12682 1012
rect 12986 960 12992 1012
rect 13044 960 13050 1012
rect 14366 960 14372 1012
rect 14424 960 14430 1012
rect 15010 960 15016 1012
rect 15068 1000 15074 1012
rect 15746 1000 15752 1012
rect 15068 972 15752 1000
rect 15068 960 15074 972
rect 15746 960 15752 972
rect 15804 960 15810 1012
rect 15930 960 15936 1012
rect 15988 960 15994 1012
rect 16022 960 16028 1012
rect 16080 1000 16086 1012
rect 16209 1003 16267 1009
rect 16209 1000 16221 1003
rect 16080 972 16221 1000
rect 16080 960 16086 972
rect 16209 969 16221 972
rect 16255 969 16267 1003
rect 16209 963 16267 969
rect 17586 960 17592 1012
rect 17644 1000 17650 1012
rect 18785 1003 18843 1009
rect 18785 1000 18797 1003
rect 17644 972 18797 1000
rect 17644 960 17650 972
rect 18785 969 18797 972
rect 18831 969 18843 1003
rect 18785 963 18843 969
rect 19794 960 19800 1012
rect 19852 1000 19858 1012
rect 19852 972 21404 1000
rect 19852 960 19858 972
rect 9784 864 9812 960
rect 9784 836 10088 864
rect 9766 756 9772 808
rect 9824 756 9830 808
rect 10060 805 10088 836
rect 10045 799 10103 805
rect 10045 765 10057 799
rect 10091 765 10103 799
rect 10796 796 10824 960
rect 11606 824 11612 876
rect 11664 824 11670 876
rect 11057 799 11115 805
rect 11057 796 11069 799
rect 10796 768 11069 796
rect 10045 759 10103 765
rect 11057 765 11069 768
rect 11103 765 11115 799
rect 11057 759 11115 765
rect 11514 756 11520 808
rect 11572 796 11578 808
rect 11885 799 11943 805
rect 11885 796 11897 799
rect 11572 768 11897 796
rect 11572 756 11578 768
rect 11885 765 11897 768
rect 11931 765 11943 799
rect 11885 759 11943 765
rect 12069 799 12127 805
rect 12069 765 12081 799
rect 12115 796 12127 799
rect 12161 799 12219 805
rect 12161 796 12173 799
rect 12115 768 12173 796
rect 12115 765 12127 768
rect 12069 759 12127 765
rect 12161 765 12173 768
rect 12207 765 12219 799
rect 12636 796 12664 960
rect 12805 799 12863 805
rect 12805 796 12817 799
rect 12636 768 12817 796
rect 12161 759 12219 765
rect 12805 765 12817 768
rect 12851 765 12863 799
rect 12805 759 12863 765
rect 13004 728 13032 960
rect 13541 799 13599 805
rect 13541 765 13553 799
rect 13587 796 13599 799
rect 13814 796 13820 808
rect 13587 768 13820 796
rect 13587 765 13599 768
rect 13541 759 13599 765
rect 13814 756 13820 768
rect 13872 756 13878 808
rect 14384 796 14412 960
rect 15948 932 15976 960
rect 15948 904 20944 932
rect 15120 836 16712 864
rect 15120 808 15148 836
rect 14461 799 14519 805
rect 14461 796 14473 799
rect 14384 768 14473 796
rect 14461 765 14473 768
rect 14507 765 14519 799
rect 14461 759 14519 765
rect 15102 756 15108 808
rect 15160 756 15166 808
rect 15838 756 15844 808
rect 15896 756 15902 808
rect 16114 756 16120 808
rect 16172 756 16178 808
rect 16393 799 16451 805
rect 16393 765 16405 799
rect 16439 765 16451 799
rect 16393 759 16451 765
rect 8680 700 9628 728
rect 9692 700 13032 728
rect 15856 728 15884 756
rect 16408 728 16436 759
rect 16574 756 16580 808
rect 16632 756 16638 808
rect 16684 805 16712 836
rect 17954 824 17960 876
rect 18012 824 18018 876
rect 18690 824 18696 876
rect 18748 824 18754 876
rect 19058 824 19064 876
rect 19116 864 19122 876
rect 19116 836 20852 864
rect 19116 824 19122 836
rect 16669 799 16727 805
rect 16669 765 16681 799
rect 16715 765 16727 799
rect 16669 759 16727 765
rect 17402 756 17408 808
rect 17460 796 17466 808
rect 17497 799 17555 805
rect 17497 796 17509 799
rect 17460 768 17509 796
rect 17460 756 17466 768
rect 17497 765 17509 768
rect 17543 765 17555 799
rect 17972 796 18000 824
rect 18233 799 18291 805
rect 18233 796 18245 799
rect 17972 768 18245 796
rect 17497 759 17555 765
rect 18233 765 18245 768
rect 18279 765 18291 799
rect 18233 759 18291 765
rect 18966 756 18972 808
rect 19024 756 19030 808
rect 20824 805 20852 836
rect 19981 799 20039 805
rect 19981 796 19993 799
rect 19076 768 19993 796
rect 15856 700 16436 728
rect 16592 728 16620 756
rect 19076 728 19104 768
rect 19981 765 19993 768
rect 20027 765 20039 799
rect 19981 759 20039 765
rect 20809 799 20867 805
rect 20809 765 20821 799
rect 20855 765 20867 799
rect 20809 759 20867 765
rect 16592 700 19104 728
rect 19153 731 19211 737
rect 3973 691 4031 697
rect 1026 620 1032 672
rect 1084 620 1090 672
rect 3326 620 3332 672
rect 3384 620 3390 672
rect 3988 660 4016 691
rect 4062 660 4068 672
rect 3988 632 4068 660
rect 4062 620 4068 632
rect 4120 620 4126 672
rect 4338 620 4344 672
rect 4396 620 4402 672
rect 5166 620 5172 672
rect 5224 620 5230 672
rect 5994 620 6000 672
rect 6052 620 6058 672
rect 8478 620 8484 672
rect 8536 620 8542 672
rect 9122 620 9128 672
rect 9180 660 9186 672
rect 9600 669 9628 700
rect 19153 697 19165 731
rect 19199 728 19211 731
rect 19337 731 19395 737
rect 19337 728 19349 731
rect 19199 700 19349 728
rect 19199 697 19211 700
rect 19153 691 19211 697
rect 19337 697 19349 700
rect 19383 697 19395 731
rect 20916 728 20944 904
rect 21376 873 21404 972
rect 21361 867 21419 873
rect 21361 833 21373 867
rect 21407 833 21419 867
rect 21361 827 21419 833
rect 22094 824 22100 876
rect 22152 824 22158 876
rect 22186 756 22192 808
rect 22244 756 22250 808
rect 22557 799 22615 805
rect 22557 765 22569 799
rect 22603 765 22615 799
rect 22557 759 22615 765
rect 22572 728 22600 759
rect 20916 700 22600 728
rect 19337 691 19395 697
rect 9401 663 9459 669
rect 9401 660 9413 663
rect 9180 632 9413 660
rect 9180 620 9186 632
rect 9401 629 9413 632
rect 9447 629 9459 663
rect 9401 623 9459 629
rect 9585 663 9643 669
rect 9585 629 9597 663
rect 9631 629 9643 663
rect 9585 623 9643 629
rect 9950 620 9956 672
rect 10008 660 10014 672
rect 10229 663 10287 669
rect 10229 660 10241 663
rect 10008 632 10241 660
rect 10008 620 10014 632
rect 10229 629 10241 632
rect 10275 629 10287 663
rect 10229 623 10287 629
rect 11146 620 11152 672
rect 11204 620 11210 672
rect 11606 620 11612 672
rect 11664 660 11670 672
rect 12345 663 12403 669
rect 12345 660 12357 663
rect 11664 632 12357 660
rect 11664 620 11670 632
rect 12345 629 12357 632
rect 12391 629 12403 663
rect 12345 623 12403 629
rect 12618 620 12624 672
rect 12676 620 12682 672
rect 13262 620 13268 672
rect 13320 660 13326 672
rect 13725 663 13783 669
rect 13725 660 13737 663
rect 13320 632 13737 660
rect 13320 620 13326 632
rect 13725 629 13737 632
rect 13771 629 13783 663
rect 13725 623 13783 629
rect 14274 620 14280 672
rect 14332 620 14338 672
rect 16577 663 16635 669
rect 16577 629 16589 663
rect 16623 660 16635 663
rect 16758 660 16764 672
rect 16623 632 16764 660
rect 16623 629 16635 632
rect 16577 623 16635 629
rect 16758 620 16764 632
rect 16816 620 16822 672
rect 16850 620 16856 672
rect 16908 620 16914 672
rect 17402 620 17408 672
rect 17460 660 17466 672
rect 17681 663 17739 669
rect 17681 660 17693 663
rect 17460 632 17693 660
rect 17460 620 17466 632
rect 17681 629 17693 632
rect 17727 629 17739 663
rect 17681 623 17739 629
rect 18414 620 18420 672
rect 18472 620 18478 672
rect 19058 620 19064 672
rect 19116 660 19122 672
rect 19429 663 19487 669
rect 19429 660 19441 663
rect 19116 632 19441 660
rect 19116 620 19122 632
rect 19429 629 19441 632
rect 19475 629 19487 663
rect 19429 623 19487 629
rect 19886 620 19892 672
rect 19944 660 19950 672
rect 20165 663 20223 669
rect 20165 660 20177 663
rect 19944 632 20177 660
rect 19944 620 19950 632
rect 20165 629 20177 632
rect 20211 629 20223 663
rect 20165 623 20223 629
rect 20714 620 20720 672
rect 20772 660 20778 672
rect 20993 663 21051 669
rect 20993 660 21005 663
rect 20772 632 21005 660
rect 20772 620 20778 632
rect 20993 629 21005 632
rect 21039 629 21051 663
rect 20993 623 21051 629
rect 21542 620 21548 672
rect 21600 660 21606 672
rect 22741 663 22799 669
rect 22741 660 22753 663
rect 21600 632 22753 660
rect 21600 620 21606 632
rect 22741 629 22753 632
rect 22787 629 22799 663
rect 22741 623 22799 629
rect 552 570 23368 592
rect 552 518 4366 570
rect 4418 518 4430 570
rect 4482 518 4494 570
rect 4546 518 4558 570
rect 4610 518 4622 570
rect 4674 518 4686 570
rect 4738 518 10366 570
rect 10418 518 10430 570
rect 10482 518 10494 570
rect 10546 518 10558 570
rect 10610 518 10622 570
rect 10674 518 10686 570
rect 10738 518 16366 570
rect 16418 518 16430 570
rect 16482 518 16494 570
rect 16546 518 16558 570
rect 16610 518 16622 570
rect 16674 518 16686 570
rect 16738 518 22366 570
rect 22418 518 22430 570
rect 22482 518 22494 570
rect 22546 518 22558 570
rect 22610 518 22622 570
rect 22674 518 22686 570
rect 22738 518 23368 570
rect 552 496 23368 518
rect 21634 456 21640 468
rect 18892 428 21640 456
rect 5442 348 5448 400
rect 5500 388 5506 400
rect 5500 360 16712 388
rect 5500 348 5506 360
rect 6178 280 6184 332
rect 6236 320 6242 332
rect 15378 320 15384 332
rect 6236 292 15384 320
rect 6236 280 6242 292
rect 15378 280 15384 292
rect 15436 280 15442 332
rect 16684 320 16712 360
rect 16758 348 16764 400
rect 16816 388 16822 400
rect 18892 388 18920 428
rect 21634 416 21640 428
rect 21692 416 21698 468
rect 16816 360 18920 388
rect 16816 348 16822 360
rect 18138 320 18144 332
rect 16684 292 18144 320
rect 18138 280 18144 292
rect 18196 280 18202 332
rect 4062 212 4068 264
rect 4120 252 4126 264
rect 10226 252 10232 264
rect 4120 224 10232 252
rect 4120 212 4126 224
rect 10226 212 10232 224
rect 10284 212 10290 264
rect 12710 252 12716 264
rect 11900 224 12716 252
rect 9490 144 9496 196
rect 9548 184 9554 196
rect 11900 184 11928 224
rect 12710 212 12716 224
rect 12768 212 12774 264
rect 9548 156 11928 184
rect 9548 144 9554 156
<< via1 >>
rect 16212 15376 16264 15428
rect 17224 15376 17276 15428
rect 6552 15308 6604 15360
rect 6736 15308 6788 15360
rect 14464 15308 14516 15360
rect 14740 15308 14792 15360
rect 18052 15308 18104 15360
rect 22284 15308 22336 15360
rect 1366 15206 1418 15258
rect 1430 15206 1482 15258
rect 1494 15206 1546 15258
rect 1558 15206 1610 15258
rect 1622 15206 1674 15258
rect 1686 15206 1738 15258
rect 7366 15206 7418 15258
rect 7430 15206 7482 15258
rect 7494 15206 7546 15258
rect 7558 15206 7610 15258
rect 7622 15206 7674 15258
rect 7686 15206 7738 15258
rect 13366 15206 13418 15258
rect 13430 15206 13482 15258
rect 13494 15206 13546 15258
rect 13558 15206 13610 15258
rect 13622 15206 13674 15258
rect 13686 15206 13738 15258
rect 19366 15206 19418 15258
rect 19430 15206 19482 15258
rect 19494 15206 19546 15258
rect 19558 15206 19610 15258
rect 19622 15206 19674 15258
rect 19686 15206 19738 15258
rect 4620 15147 4672 15156
rect 4620 15113 4629 15147
rect 4629 15113 4663 15147
rect 4663 15113 4672 15147
rect 4620 15104 4672 15113
rect 5172 15147 5224 15156
rect 5172 15113 5181 15147
rect 5181 15113 5215 15147
rect 5215 15113 5224 15147
rect 5172 15104 5224 15113
rect 6184 15147 6236 15156
rect 6184 15113 6193 15147
rect 6193 15113 6227 15147
rect 6227 15113 6236 15147
rect 6184 15104 6236 15113
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 7288 15104 7340 15156
rect 8116 15104 8168 15156
rect 9128 15147 9180 15156
rect 9128 15113 9137 15147
rect 9137 15113 9171 15147
rect 9171 15113 9180 15147
rect 9128 15104 9180 15113
rect 9588 15147 9640 15156
rect 9588 15113 9597 15147
rect 9597 15113 9631 15147
rect 9631 15113 9640 15147
rect 9588 15104 9640 15113
rect 10324 15104 10376 15156
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 14464 15104 14516 15156
rect 2228 14900 2280 14952
rect 4896 14900 4948 14952
rect 6736 14832 6788 14884
rect 6920 14875 6972 14884
rect 6920 14841 6929 14875
rect 6929 14841 6963 14875
rect 6963 14841 6972 14875
rect 6920 14832 6972 14841
rect 7656 14968 7708 15020
rect 18604 15104 18656 15156
rect 17040 15036 17092 15088
rect 17316 15036 17368 15088
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 8576 14900 8628 14952
rect 8944 14943 8996 14952
rect 8944 14909 8953 14943
rect 8953 14909 8987 14943
rect 8987 14909 8996 14943
rect 8944 14900 8996 14909
rect 10140 14900 10192 14952
rect 8668 14832 8720 14884
rect 9496 14832 9548 14884
rect 9680 14832 9732 14884
rect 11980 14832 12032 14884
rect 13268 14900 13320 14952
rect 16764 14968 16816 15020
rect 22284 15036 22336 15088
rect 16856 14900 16908 14952
rect 17684 14900 17736 14952
rect 18420 14900 18472 14952
rect 19156 14900 19208 14952
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 20168 14900 20220 14952
rect 20628 14900 20680 14952
rect 21364 14900 21416 14952
rect 21456 14900 21508 14952
rect 18236 14832 18288 14884
rect 22100 14900 22152 14952
rect 22836 14900 22888 14952
rect 2504 14764 2556 14816
rect 5172 14764 5224 14816
rect 7104 14764 7156 14816
rect 7932 14807 7984 14816
rect 7932 14773 7941 14807
rect 7941 14773 7975 14807
rect 7975 14773 7984 14807
rect 7932 14764 7984 14773
rect 11888 14764 11940 14816
rect 13820 14764 13872 14816
rect 18512 14764 18564 14816
rect 18880 14807 18932 14816
rect 18880 14773 18889 14807
rect 18889 14773 18923 14807
rect 18923 14773 18932 14807
rect 18880 14764 18932 14773
rect 19248 14807 19300 14816
rect 19248 14773 19257 14807
rect 19257 14773 19291 14807
rect 19291 14773 19300 14807
rect 19248 14764 19300 14773
rect 19984 14764 20036 14816
rect 20168 14807 20220 14816
rect 20168 14773 20177 14807
rect 20177 14773 20211 14807
rect 20211 14773 20220 14807
rect 20168 14764 20220 14773
rect 21548 14764 21600 14816
rect 4366 14662 4418 14714
rect 4430 14662 4482 14714
rect 4494 14662 4546 14714
rect 4558 14662 4610 14714
rect 4622 14662 4674 14714
rect 4686 14662 4738 14714
rect 10366 14662 10418 14714
rect 10430 14662 10482 14714
rect 10494 14662 10546 14714
rect 10558 14662 10610 14714
rect 10622 14662 10674 14714
rect 10686 14662 10738 14714
rect 16366 14662 16418 14714
rect 16430 14662 16482 14714
rect 16494 14662 16546 14714
rect 16558 14662 16610 14714
rect 16622 14662 16674 14714
rect 16686 14662 16738 14714
rect 22366 14662 22418 14714
rect 22430 14662 22482 14714
rect 22494 14662 22546 14714
rect 22558 14662 22610 14714
rect 22622 14662 22674 14714
rect 22686 14662 22738 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2412 14603 2464 14612
rect 2412 14569 2421 14603
rect 2421 14569 2455 14603
rect 2455 14569 2464 14603
rect 2412 14560 2464 14569
rect 4896 14560 4948 14612
rect 6644 14560 6696 14612
rect 7656 14560 7708 14612
rect 7932 14560 7984 14612
rect 8944 14560 8996 14612
rect 6092 14535 6144 14544
rect 2504 14467 2556 14476
rect 2504 14433 2513 14467
rect 2513 14433 2547 14467
rect 2547 14433 2556 14467
rect 2504 14424 2556 14433
rect 2872 14467 2924 14476
rect 2872 14433 2906 14467
rect 2906 14433 2924 14467
rect 2872 14424 2924 14433
rect 6092 14501 6101 14535
rect 6101 14501 6135 14535
rect 6135 14501 6144 14535
rect 6092 14492 6144 14501
rect 4344 14424 4396 14476
rect 5356 14424 5408 14476
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 6736 14424 6788 14476
rect 7104 14467 7156 14476
rect 7104 14433 7113 14467
rect 7113 14433 7147 14467
rect 7147 14433 7156 14467
rect 7104 14424 7156 14433
rect 8024 14424 8076 14476
rect 8760 14424 8812 14476
rect 10692 14560 10744 14612
rect 10232 14424 10284 14476
rect 14740 14560 14792 14612
rect 15752 14560 15804 14612
rect 16948 14603 17000 14612
rect 16948 14569 16957 14603
rect 16957 14569 16991 14603
rect 16991 14569 17000 14603
rect 16948 14560 17000 14569
rect 18052 14603 18104 14612
rect 18052 14569 18061 14603
rect 18061 14569 18095 14603
rect 18095 14569 18104 14603
rect 18052 14560 18104 14569
rect 18420 14603 18472 14612
rect 18420 14569 18429 14603
rect 18429 14569 18463 14603
rect 18463 14569 18472 14603
rect 18420 14560 18472 14569
rect 19248 14560 19300 14612
rect 21456 14560 21508 14612
rect 1032 14220 1084 14272
rect 1860 14220 1912 14272
rect 4252 14220 4304 14272
rect 6184 14220 6236 14272
rect 9128 14356 9180 14408
rect 9312 14399 9364 14408
rect 9312 14365 9321 14399
rect 9321 14365 9355 14399
rect 9355 14365 9364 14399
rect 9312 14356 9364 14365
rect 10048 14331 10100 14340
rect 10048 14297 10057 14331
rect 10057 14297 10091 14331
rect 10091 14297 10100 14331
rect 10048 14288 10100 14297
rect 8116 14220 8168 14272
rect 9312 14220 9364 14272
rect 10784 14263 10836 14272
rect 10784 14229 10793 14263
rect 10793 14229 10827 14263
rect 10827 14229 10836 14263
rect 10784 14220 10836 14229
rect 10876 14220 10928 14272
rect 11336 14263 11388 14272
rect 11336 14229 11345 14263
rect 11345 14229 11379 14263
rect 11379 14229 11388 14263
rect 11336 14220 11388 14229
rect 13268 14220 13320 14272
rect 14556 14424 14608 14476
rect 17408 14492 17460 14544
rect 15200 14356 15252 14408
rect 16304 14356 16356 14408
rect 16488 14467 16540 14476
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16488 14424 16540 14433
rect 17592 14424 17644 14476
rect 17040 14356 17092 14408
rect 18236 14424 18288 14476
rect 18604 14424 18656 14476
rect 19984 14467 20036 14476
rect 19984 14433 20018 14467
rect 20018 14433 20036 14467
rect 17960 14399 18012 14408
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 15844 14331 15896 14340
rect 15844 14297 15853 14331
rect 15853 14297 15887 14331
rect 15887 14297 15896 14331
rect 15844 14288 15896 14297
rect 17132 14288 17184 14340
rect 17500 14331 17552 14340
rect 17500 14297 17509 14331
rect 17509 14297 17543 14331
rect 17543 14297 17552 14331
rect 17500 14288 17552 14297
rect 15384 14220 15436 14272
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 17868 14263 17920 14272
rect 17868 14229 17877 14263
rect 17877 14229 17911 14263
rect 17911 14229 17920 14263
rect 17868 14220 17920 14229
rect 18788 14356 18840 14408
rect 19984 14424 20036 14433
rect 18880 14288 18932 14340
rect 18604 14220 18656 14272
rect 1366 14118 1418 14170
rect 1430 14118 1482 14170
rect 1494 14118 1546 14170
rect 1558 14118 1610 14170
rect 1622 14118 1674 14170
rect 1686 14118 1738 14170
rect 7366 14118 7418 14170
rect 7430 14118 7482 14170
rect 7494 14118 7546 14170
rect 7558 14118 7610 14170
rect 7622 14118 7674 14170
rect 7686 14118 7738 14170
rect 13366 14118 13418 14170
rect 13430 14118 13482 14170
rect 13494 14118 13546 14170
rect 13558 14118 13610 14170
rect 13622 14118 13674 14170
rect 13686 14118 13738 14170
rect 19366 14118 19418 14170
rect 19430 14118 19482 14170
rect 19494 14118 19546 14170
rect 19558 14118 19610 14170
rect 19622 14118 19674 14170
rect 19686 14118 19738 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 2412 14016 2464 14068
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 7840 14059 7892 14068
rect 7840 14025 7849 14059
rect 7849 14025 7883 14059
rect 7883 14025 7892 14059
rect 7840 14016 7892 14025
rect 8576 14016 8628 14068
rect 10048 14016 10100 14068
rect 10876 14016 10928 14068
rect 11336 14016 11388 14068
rect 6276 13948 6328 14000
rect 10508 13948 10560 14000
rect 1216 13812 1268 13864
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 1768 13744 1820 13796
rect 2688 13855 2740 13864
rect 2688 13821 2697 13855
rect 2697 13821 2731 13855
rect 2731 13821 2740 13855
rect 2688 13812 2740 13821
rect 3884 13812 3936 13864
rect 4344 13812 4396 13864
rect 6828 13812 6880 13864
rect 7748 13812 7800 13864
rect 8208 13812 8260 13864
rect 6184 13744 6236 13796
rect 2596 13676 2648 13728
rect 5540 13676 5592 13728
rect 8576 13812 8628 13864
rect 9128 13812 9180 13864
rect 9312 13812 9364 13864
rect 11152 13948 11204 14000
rect 11888 13948 11940 14000
rect 10784 13812 10836 13864
rect 11428 13812 11480 13864
rect 11612 13812 11664 13864
rect 12992 13812 13044 13864
rect 14556 14059 14608 14068
rect 14556 14025 14565 14059
rect 14565 14025 14599 14059
rect 14599 14025 14608 14059
rect 14556 14016 14608 14025
rect 16212 14016 16264 14068
rect 16856 14016 16908 14068
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 17868 14016 17920 14068
rect 18420 14016 18472 14068
rect 18604 14016 18656 14068
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 21456 14016 21508 14068
rect 14188 13948 14240 14000
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 15752 13880 15804 13932
rect 15844 13880 15896 13932
rect 13176 13855 13228 13864
rect 13176 13821 13185 13855
rect 13185 13821 13219 13855
rect 13219 13821 13228 13855
rect 13176 13812 13228 13821
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14648 13812 14700 13864
rect 16120 13812 16172 13864
rect 17040 13880 17092 13932
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 18696 13812 18748 13864
rect 18972 13812 19024 13864
rect 19156 13880 19208 13932
rect 20168 13812 20220 13864
rect 9956 13676 10008 13728
rect 10968 13676 11020 13728
rect 16764 13676 16816 13728
rect 16856 13676 16908 13728
rect 17316 13676 17368 13728
rect 18696 13719 18748 13728
rect 18696 13685 18705 13719
rect 18705 13685 18739 13719
rect 18739 13685 18748 13719
rect 18696 13676 18748 13685
rect 4366 13574 4418 13626
rect 4430 13574 4482 13626
rect 4494 13574 4546 13626
rect 4558 13574 4610 13626
rect 4622 13574 4674 13626
rect 4686 13574 4738 13626
rect 10366 13574 10418 13626
rect 10430 13574 10482 13626
rect 10494 13574 10546 13626
rect 10558 13574 10610 13626
rect 10622 13574 10674 13626
rect 10686 13574 10738 13626
rect 16366 13574 16418 13626
rect 16430 13574 16482 13626
rect 16494 13574 16546 13626
rect 16558 13574 16610 13626
rect 16622 13574 16674 13626
rect 16686 13574 16738 13626
rect 22366 13574 22418 13626
rect 22430 13574 22482 13626
rect 22494 13574 22546 13626
rect 22558 13574 22610 13626
rect 22622 13574 22674 13626
rect 22686 13574 22738 13626
rect 1124 13404 1176 13456
rect 2228 13404 2280 13456
rect 1032 13336 1084 13388
rect 3884 13472 3936 13524
rect 8576 13472 8628 13524
rect 2596 13447 2648 13456
rect 2596 13413 2630 13447
rect 2630 13413 2648 13447
rect 2596 13404 2648 13413
rect 6920 13404 6972 13456
rect 6092 13336 6144 13388
rect 7748 13404 7800 13456
rect 8116 13404 8168 13456
rect 10232 13404 10284 13456
rect 4160 13268 4212 13320
rect 5816 13268 5868 13320
rect 8760 13379 8812 13388
rect 8760 13345 8769 13379
rect 8769 13345 8803 13379
rect 8803 13345 8812 13379
rect 8760 13336 8812 13345
rect 8208 13268 8260 13320
rect 9312 13268 9364 13320
rect 9588 13268 9640 13320
rect 10784 13336 10836 13388
rect 5908 13200 5960 13252
rect 12072 13404 12124 13456
rect 13084 13472 13136 13524
rect 17500 13472 17552 13524
rect 17776 13472 17828 13524
rect 18052 13472 18104 13524
rect 18420 13515 18472 13524
rect 18420 13481 18429 13515
rect 18429 13481 18463 13515
rect 18463 13481 18472 13515
rect 18420 13472 18472 13481
rect 18512 13515 18564 13524
rect 18512 13481 18521 13515
rect 18521 13481 18555 13515
rect 18555 13481 18564 13515
rect 18512 13472 18564 13481
rect 18696 13472 18748 13524
rect 11152 13379 11204 13388
rect 11152 13345 11161 13379
rect 11161 13345 11195 13379
rect 11195 13345 11204 13379
rect 11152 13336 11204 13345
rect 2044 13175 2096 13184
rect 2044 13141 2053 13175
rect 2053 13141 2087 13175
rect 2087 13141 2096 13175
rect 2044 13132 2096 13141
rect 2688 13132 2740 13184
rect 3424 13132 3476 13184
rect 5356 13132 5408 13184
rect 6092 13175 6144 13184
rect 6092 13141 6101 13175
rect 6101 13141 6135 13175
rect 6135 13141 6144 13175
rect 6092 13132 6144 13141
rect 6460 13175 6512 13184
rect 6460 13141 6469 13175
rect 6469 13141 6503 13175
rect 6503 13141 6512 13175
rect 6460 13132 6512 13141
rect 6920 13132 6972 13184
rect 8024 13132 8076 13184
rect 9956 13132 10008 13184
rect 10692 13132 10744 13184
rect 10876 13132 10928 13184
rect 11152 13200 11204 13252
rect 11520 13200 11572 13252
rect 11796 13268 11848 13320
rect 15936 13268 15988 13320
rect 17960 13404 18012 13456
rect 19156 13515 19208 13524
rect 19156 13481 19165 13515
rect 19165 13481 19199 13515
rect 19199 13481 19208 13515
rect 19156 13472 19208 13481
rect 16856 13379 16908 13388
rect 16856 13345 16865 13379
rect 16865 13345 16899 13379
rect 16899 13345 16908 13379
rect 16856 13336 16908 13345
rect 16764 13268 16816 13320
rect 18512 13336 18564 13388
rect 19800 13336 19852 13388
rect 16396 13200 16448 13252
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 18420 13268 18472 13320
rect 21456 13404 21508 13456
rect 21364 13379 21416 13388
rect 21364 13345 21373 13379
rect 21373 13345 21407 13379
rect 21407 13345 21416 13379
rect 21364 13336 21416 13345
rect 20260 13268 20312 13320
rect 12716 13132 12768 13184
rect 14464 13132 14516 13184
rect 21548 13200 21600 13252
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 20444 13132 20496 13184
rect 1366 13030 1418 13082
rect 1430 13030 1482 13082
rect 1494 13030 1546 13082
rect 1558 13030 1610 13082
rect 1622 13030 1674 13082
rect 1686 13030 1738 13082
rect 7366 13030 7418 13082
rect 7430 13030 7482 13082
rect 7494 13030 7546 13082
rect 7558 13030 7610 13082
rect 7622 13030 7674 13082
rect 7686 13030 7738 13082
rect 13366 13030 13418 13082
rect 13430 13030 13482 13082
rect 13494 13030 13546 13082
rect 13558 13030 13610 13082
rect 13622 13030 13674 13082
rect 13686 13030 13738 13082
rect 19366 13030 19418 13082
rect 19430 13030 19482 13082
rect 19494 13030 19546 13082
rect 19558 13030 19610 13082
rect 19622 13030 19674 13082
rect 19686 13030 19738 13082
rect 1676 12971 1728 12980
rect 1676 12937 1685 12971
rect 1685 12937 1719 12971
rect 1719 12937 1728 12971
rect 1676 12928 1728 12937
rect 1768 12928 1820 12980
rect 2044 12928 2096 12980
rect 2228 12928 2280 12980
rect 1584 12792 1636 12844
rect 2412 12860 2464 12912
rect 1124 12656 1176 12708
rect 1676 12631 1728 12640
rect 1676 12597 1701 12631
rect 1701 12597 1728 12631
rect 1676 12588 1728 12597
rect 1952 12588 2004 12640
rect 2964 12860 3016 12912
rect 3884 12928 3936 12980
rect 5540 12928 5592 12980
rect 5908 12971 5960 12980
rect 5908 12937 5917 12971
rect 5917 12937 5951 12971
rect 5951 12937 5960 12971
rect 5908 12928 5960 12937
rect 6460 12928 6512 12980
rect 7012 12928 7064 12980
rect 10048 12928 10100 12980
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 2964 12724 3016 12776
rect 4804 12724 4856 12776
rect 6276 12724 6328 12776
rect 6736 12860 6788 12912
rect 2964 12588 3016 12640
rect 3976 12588 4028 12640
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 10140 12860 10192 12912
rect 12992 12928 13044 12980
rect 15936 12928 15988 12980
rect 17592 12928 17644 12980
rect 10692 12792 10744 12844
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 12900 12903 12952 12912
rect 12900 12869 12909 12903
rect 12909 12869 12943 12903
rect 12943 12869 12952 12903
rect 12900 12860 12952 12869
rect 7472 12656 7524 12708
rect 9864 12724 9916 12776
rect 11888 12792 11940 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 16396 12860 16448 12912
rect 18052 12792 18104 12844
rect 18328 12792 18380 12844
rect 18788 12792 18840 12844
rect 11336 12724 11388 12776
rect 11520 12724 11572 12776
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 11704 12767 11756 12776
rect 11704 12733 11713 12767
rect 11713 12733 11747 12767
rect 11747 12733 11756 12767
rect 11704 12724 11756 12733
rect 13084 12767 13136 12776
rect 7288 12588 7340 12640
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 9496 12588 9548 12640
rect 11244 12656 11296 12708
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13912 12767 13964 12776
rect 13912 12733 13921 12767
rect 13921 12733 13955 12767
rect 13955 12733 13964 12767
rect 13912 12724 13964 12733
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 14372 12724 14424 12776
rect 14464 12767 14516 12776
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 17224 12724 17276 12776
rect 10232 12588 10284 12640
rect 11980 12588 12032 12640
rect 16856 12656 16908 12708
rect 14648 12631 14700 12640
rect 14648 12597 14657 12631
rect 14657 12597 14691 12631
rect 14691 12597 14700 12631
rect 14648 12588 14700 12597
rect 17316 12588 17368 12640
rect 18788 12588 18840 12640
rect 19800 12767 19852 12776
rect 19800 12733 19809 12767
rect 19809 12733 19843 12767
rect 19843 12733 19852 12767
rect 19800 12724 19852 12733
rect 20260 12724 20312 12776
rect 20444 12767 20496 12776
rect 20444 12733 20478 12767
rect 20478 12733 20496 12767
rect 20444 12724 20496 12733
rect 21364 12928 21416 12980
rect 21548 12792 21600 12844
rect 23296 12792 23348 12844
rect 19892 12656 19944 12708
rect 19984 12656 20036 12708
rect 22192 12656 22244 12708
rect 20168 12588 20220 12640
rect 20720 12588 20772 12640
rect 22836 12631 22888 12640
rect 22836 12597 22845 12631
rect 22845 12597 22879 12631
rect 22879 12597 22888 12631
rect 22836 12588 22888 12597
rect 4366 12486 4418 12538
rect 4430 12486 4482 12538
rect 4494 12486 4546 12538
rect 4558 12486 4610 12538
rect 4622 12486 4674 12538
rect 4686 12486 4738 12538
rect 10366 12486 10418 12538
rect 10430 12486 10482 12538
rect 10494 12486 10546 12538
rect 10558 12486 10610 12538
rect 10622 12486 10674 12538
rect 10686 12486 10738 12538
rect 16366 12486 16418 12538
rect 16430 12486 16482 12538
rect 16494 12486 16546 12538
rect 16558 12486 16610 12538
rect 16622 12486 16674 12538
rect 16686 12486 16738 12538
rect 22366 12486 22418 12538
rect 22430 12486 22482 12538
rect 22494 12486 22546 12538
rect 22558 12486 22610 12538
rect 22622 12486 22674 12538
rect 22686 12486 22738 12538
rect 1676 12384 1728 12436
rect 1584 12316 1636 12368
rect 1860 12359 1912 12368
rect 1860 12325 1869 12359
rect 1869 12325 1903 12359
rect 1903 12325 1912 12359
rect 1860 12316 1912 12325
rect 1952 12291 2004 12300
rect 1952 12257 1961 12291
rect 1961 12257 1995 12291
rect 1995 12257 2004 12291
rect 2412 12316 2464 12368
rect 4804 12384 4856 12436
rect 5356 12384 5408 12436
rect 7472 12427 7524 12436
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 1952 12248 2004 12257
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 2504 12248 2556 12257
rect 4252 12248 4304 12300
rect 2044 12180 2096 12232
rect 1124 12112 1176 12164
rect 1768 12155 1820 12164
rect 1768 12121 1777 12155
rect 1777 12121 1811 12155
rect 1811 12121 1820 12155
rect 1768 12112 1820 12121
rect 2320 12112 2372 12164
rect 2596 12180 2648 12232
rect 4620 12248 4672 12300
rect 4896 12248 4948 12300
rect 5356 12248 5408 12300
rect 5908 12248 5960 12300
rect 7840 12248 7892 12300
rect 8484 12248 8536 12300
rect 10232 12248 10284 12300
rect 4712 12180 4764 12232
rect 2412 12044 2464 12096
rect 2964 12044 3016 12096
rect 3516 12044 3568 12096
rect 4160 12044 4212 12096
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 5080 12112 5132 12164
rect 6000 12112 6052 12164
rect 7288 12180 7340 12232
rect 8760 12180 8812 12232
rect 9772 12180 9824 12232
rect 10140 12180 10192 12232
rect 10876 12316 10928 12368
rect 11612 12384 11664 12436
rect 13820 12384 13872 12436
rect 14280 12384 14332 12436
rect 15752 12384 15804 12436
rect 17408 12384 17460 12436
rect 10692 12180 10744 12232
rect 11520 12180 11572 12232
rect 5448 12044 5500 12096
rect 5632 12087 5684 12096
rect 5632 12053 5641 12087
rect 5641 12053 5675 12087
rect 5675 12053 5684 12087
rect 5632 12044 5684 12053
rect 9312 12112 9364 12164
rect 6644 12044 6696 12096
rect 7932 12044 7984 12096
rect 9404 12044 9456 12096
rect 10876 12112 10928 12164
rect 11428 12112 11480 12164
rect 12992 12291 13044 12300
rect 12992 12257 13001 12291
rect 13001 12257 13035 12291
rect 13035 12257 13044 12291
rect 12992 12248 13044 12257
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 12808 12180 12860 12232
rect 12164 12112 12216 12164
rect 13084 12112 13136 12164
rect 10600 12044 10652 12096
rect 10784 12044 10836 12096
rect 11244 12044 11296 12096
rect 12256 12044 12308 12096
rect 13268 12044 13320 12096
rect 13728 12291 13780 12300
rect 13728 12257 13737 12291
rect 13737 12257 13771 12291
rect 13771 12257 13780 12291
rect 13728 12248 13780 12257
rect 14096 12316 14148 12368
rect 14740 12316 14792 12368
rect 15936 12316 15988 12368
rect 16212 12248 16264 12300
rect 19064 12316 19116 12368
rect 18328 12248 18380 12300
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 18696 12248 18748 12300
rect 20260 12316 20312 12368
rect 18788 12180 18840 12232
rect 17592 12112 17644 12164
rect 13820 12044 13872 12096
rect 15108 12044 15160 12096
rect 15936 12087 15988 12096
rect 15936 12053 15945 12087
rect 15945 12053 15979 12087
rect 15979 12053 15988 12087
rect 15936 12044 15988 12053
rect 16120 12087 16172 12096
rect 16120 12053 16129 12087
rect 16129 12053 16163 12087
rect 16163 12053 16172 12087
rect 16120 12044 16172 12053
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 18604 12044 18656 12096
rect 22284 12044 22336 12096
rect 1366 11942 1418 11994
rect 1430 11942 1482 11994
rect 1494 11942 1546 11994
rect 1558 11942 1610 11994
rect 1622 11942 1674 11994
rect 1686 11942 1738 11994
rect 7366 11942 7418 11994
rect 7430 11942 7482 11994
rect 7494 11942 7546 11994
rect 7558 11942 7610 11994
rect 7622 11942 7674 11994
rect 7686 11942 7738 11994
rect 13366 11942 13418 11994
rect 13430 11942 13482 11994
rect 13494 11942 13546 11994
rect 13558 11942 13610 11994
rect 13622 11942 13674 11994
rect 13686 11942 13738 11994
rect 19366 11942 19418 11994
rect 19430 11942 19482 11994
rect 19494 11942 19546 11994
rect 19558 11942 19610 11994
rect 19622 11942 19674 11994
rect 19686 11942 19738 11994
rect 2044 11840 2096 11892
rect 2504 11840 2556 11892
rect 4252 11772 4304 11824
rect 5080 11840 5132 11892
rect 5172 11840 5224 11892
rect 10876 11840 10928 11892
rect 13268 11840 13320 11892
rect 4712 11772 4764 11824
rect 10692 11772 10744 11824
rect 5724 11747 5776 11756
rect 5724 11713 5733 11747
rect 5733 11713 5767 11747
rect 5767 11713 5776 11747
rect 5724 11704 5776 11713
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 2320 11679 2372 11688
rect 2320 11645 2329 11679
rect 2329 11645 2363 11679
rect 2363 11645 2372 11679
rect 2320 11636 2372 11645
rect 3240 11679 3292 11688
rect 3240 11645 3249 11679
rect 3249 11645 3283 11679
rect 3283 11645 3292 11679
rect 3240 11636 3292 11645
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 4252 11636 4304 11688
rect 4712 11636 4764 11688
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 5448 11636 5500 11645
rect 5908 11636 5960 11688
rect 6460 11704 6512 11756
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 7932 11636 7984 11688
rect 6460 11568 6512 11620
rect 6828 11568 6880 11620
rect 7196 11568 7248 11620
rect 10232 11568 10284 11620
rect 11060 11679 11112 11688
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 11520 11772 11572 11824
rect 11428 11747 11480 11756
rect 11428 11713 11437 11747
rect 11437 11713 11471 11747
rect 11471 11713 11480 11747
rect 11428 11704 11480 11713
rect 12164 11772 12216 11824
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 14096 11840 14148 11892
rect 14096 11679 14148 11688
rect 14096 11645 14105 11679
rect 14105 11645 14139 11679
rect 14139 11645 14148 11679
rect 14096 11636 14148 11645
rect 12900 11568 12952 11620
rect 13636 11568 13688 11620
rect 14280 11568 14332 11620
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 18328 11883 18380 11892
rect 18328 11849 18337 11883
rect 18337 11849 18371 11883
rect 18371 11849 18380 11883
rect 18328 11840 18380 11849
rect 18512 11840 18564 11892
rect 18696 11883 18748 11892
rect 18696 11849 18705 11883
rect 18705 11849 18739 11883
rect 18739 11849 18748 11883
rect 18696 11840 18748 11849
rect 16120 11704 16172 11756
rect 17132 11704 17184 11756
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 14648 11611 14700 11620
rect 14648 11577 14657 11611
rect 14657 11577 14691 11611
rect 14691 11577 14700 11611
rect 14648 11568 14700 11577
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 17224 11636 17276 11688
rect 17960 11636 18012 11688
rect 18604 11636 18656 11688
rect 20260 11704 20312 11756
rect 20628 11704 20680 11756
rect 1492 11500 1544 11552
rect 1860 11500 1912 11552
rect 3976 11500 4028 11552
rect 5080 11500 5132 11552
rect 5172 11500 5224 11552
rect 6368 11500 6420 11552
rect 6736 11543 6788 11552
rect 6736 11509 6745 11543
rect 6745 11509 6779 11543
rect 6779 11509 6788 11543
rect 6736 11500 6788 11509
rect 11888 11500 11940 11552
rect 12072 11500 12124 11552
rect 14004 11500 14056 11552
rect 14556 11500 14608 11552
rect 15016 11543 15068 11552
rect 15016 11509 15025 11543
rect 15025 11509 15059 11543
rect 15059 11509 15068 11543
rect 15016 11500 15068 11509
rect 19156 11679 19208 11688
rect 19156 11645 19165 11679
rect 19165 11645 19199 11679
rect 19199 11645 19208 11679
rect 19156 11636 19208 11645
rect 19892 11636 19944 11688
rect 20352 11636 20404 11688
rect 21088 11636 21140 11688
rect 20444 11568 20496 11620
rect 20904 11568 20956 11620
rect 20996 11543 21048 11552
rect 20996 11509 21005 11543
rect 21005 11509 21039 11543
rect 21039 11509 21048 11543
rect 20996 11500 21048 11509
rect 22100 11500 22152 11552
rect 4366 11398 4418 11450
rect 4430 11398 4482 11450
rect 4494 11398 4546 11450
rect 4558 11398 4610 11450
rect 4622 11398 4674 11450
rect 4686 11398 4738 11450
rect 10366 11398 10418 11450
rect 10430 11398 10482 11450
rect 10494 11398 10546 11450
rect 10558 11398 10610 11450
rect 10622 11398 10674 11450
rect 10686 11398 10738 11450
rect 16366 11398 16418 11450
rect 16430 11398 16482 11450
rect 16494 11398 16546 11450
rect 16558 11398 16610 11450
rect 16622 11398 16674 11450
rect 16686 11398 16738 11450
rect 22366 11398 22418 11450
rect 22430 11398 22482 11450
rect 22494 11398 22546 11450
rect 22558 11398 22610 11450
rect 22622 11398 22674 11450
rect 22686 11398 22738 11450
rect 4896 11296 4948 11348
rect 5080 11296 5132 11348
rect 6184 11296 6236 11348
rect 7196 11296 7248 11348
rect 7840 11296 7892 11348
rect 8484 11296 8536 11348
rect 10232 11296 10284 11348
rect 1032 11160 1084 11212
rect 1492 11203 1544 11212
rect 1492 11169 1526 11203
rect 1526 11169 1544 11203
rect 1492 11160 1544 11169
rect 3332 11160 3384 11212
rect 4160 11160 4212 11212
rect 4712 11160 4764 11212
rect 6644 11228 6696 11280
rect 8392 11228 8444 11280
rect 9956 11228 10008 11280
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 11244 11296 11296 11348
rect 12532 11296 12584 11348
rect 4252 11092 4304 11144
rect 5356 11203 5408 11212
rect 5356 11169 5365 11203
rect 5365 11169 5399 11203
rect 5399 11169 5408 11203
rect 5356 11160 5408 11169
rect 6552 11160 6604 11212
rect 4988 11092 5040 11144
rect 6644 11092 6696 11144
rect 8116 11092 8168 11144
rect 8852 11203 8904 11212
rect 8852 11169 8861 11203
rect 8861 11169 8895 11203
rect 8895 11169 8904 11203
rect 8852 11160 8904 11169
rect 9220 11160 9272 11212
rect 9404 11160 9456 11212
rect 13820 11228 13872 11280
rect 10876 11160 10928 11212
rect 11152 11092 11204 11144
rect 12808 11160 12860 11212
rect 13176 11160 13228 11212
rect 3884 11067 3936 11076
rect 3884 11033 3893 11067
rect 3893 11033 3927 11067
rect 3927 11033 3936 11067
rect 3884 11024 3936 11033
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 4344 11024 4396 11076
rect 5172 11067 5224 11076
rect 3240 10956 3292 10965
rect 4068 10999 4120 11008
rect 4068 10965 4077 10999
rect 4077 10965 4111 10999
rect 4111 10965 4120 10999
rect 4068 10956 4120 10965
rect 4252 10956 4304 11008
rect 5172 11033 5181 11067
rect 5181 11033 5215 11067
rect 5215 11033 5224 11067
rect 5172 11024 5224 11033
rect 4804 10956 4856 11008
rect 8208 10956 8260 11008
rect 11060 11024 11112 11076
rect 11244 11024 11296 11076
rect 9220 10956 9272 11008
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 13912 11160 13964 11212
rect 14096 11339 14148 11348
rect 14096 11305 14105 11339
rect 14105 11305 14139 11339
rect 14139 11305 14148 11339
rect 14096 11296 14148 11305
rect 14280 11339 14332 11348
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 14464 11296 14516 11348
rect 14924 11296 14976 11348
rect 14096 11160 14148 11212
rect 15384 11228 15436 11280
rect 16120 11296 16172 11348
rect 19156 11296 19208 11348
rect 16396 11228 16448 11280
rect 13636 11092 13688 11144
rect 16120 11203 16172 11212
rect 16120 11169 16129 11203
rect 16129 11169 16163 11203
rect 16163 11169 16172 11203
rect 16120 11160 16172 11169
rect 16764 11160 16816 11212
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 18236 11228 18288 11280
rect 19892 11296 19944 11348
rect 20536 11296 20588 11348
rect 20628 11296 20680 11348
rect 20996 11296 21048 11348
rect 19800 11228 19852 11280
rect 18420 11203 18472 11212
rect 15108 11135 15160 11144
rect 15108 11101 15117 11135
rect 15117 11101 15151 11135
rect 15151 11101 15160 11135
rect 15108 11092 15160 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 18788 11160 18840 11212
rect 19708 11092 19760 11144
rect 20628 11160 20680 11212
rect 21088 11203 21140 11212
rect 21088 11169 21097 11203
rect 21097 11169 21131 11203
rect 21131 11169 21140 11203
rect 21088 11160 21140 11169
rect 11612 11024 11664 11076
rect 13268 11024 13320 11076
rect 20076 11024 20128 11076
rect 15476 10999 15528 11008
rect 15476 10965 15485 10999
rect 15485 10965 15519 10999
rect 15519 10965 15528 10999
rect 15476 10956 15528 10965
rect 17776 10956 17828 11008
rect 20260 10956 20312 11008
rect 20720 10956 20772 11008
rect 22284 10956 22336 11008
rect 1366 10854 1418 10906
rect 1430 10854 1482 10906
rect 1494 10854 1546 10906
rect 1558 10854 1610 10906
rect 1622 10854 1674 10906
rect 1686 10854 1738 10906
rect 7366 10854 7418 10906
rect 7430 10854 7482 10906
rect 7494 10854 7546 10906
rect 7558 10854 7610 10906
rect 7622 10854 7674 10906
rect 7686 10854 7738 10906
rect 13366 10854 13418 10906
rect 13430 10854 13482 10906
rect 13494 10854 13546 10906
rect 13558 10854 13610 10906
rect 13622 10854 13674 10906
rect 13686 10854 13738 10906
rect 19366 10854 19418 10906
rect 19430 10854 19482 10906
rect 19494 10854 19546 10906
rect 19558 10854 19610 10906
rect 19622 10854 19674 10906
rect 19686 10854 19738 10906
rect 1768 10752 1820 10804
rect 3700 10752 3752 10804
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 1860 10548 1912 10600
rect 3516 10548 3568 10600
rect 4068 10548 4120 10600
rect 4160 10548 4212 10600
rect 5264 10752 5316 10804
rect 6644 10752 6696 10804
rect 8392 10795 8444 10804
rect 8392 10761 8401 10795
rect 8401 10761 8435 10795
rect 8435 10761 8444 10795
rect 8392 10752 8444 10761
rect 8852 10752 8904 10804
rect 9496 10752 9548 10804
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 11336 10752 11388 10804
rect 4804 10684 4856 10736
rect 5172 10616 5224 10668
rect 5540 10616 5592 10668
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 8116 10684 8168 10736
rect 6460 10616 6512 10668
rect 6828 10616 6880 10668
rect 6368 10548 6420 10600
rect 6920 10548 6972 10600
rect 8484 10548 8536 10600
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 3792 10412 3844 10421
rect 5724 10480 5776 10532
rect 5816 10480 5868 10532
rect 5540 10412 5592 10464
rect 8484 10412 8536 10464
rect 8852 10591 8904 10600
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 11060 10684 11112 10736
rect 9956 10616 10008 10668
rect 12624 10752 12676 10804
rect 13176 10752 13228 10804
rect 15844 10752 15896 10804
rect 16396 10752 16448 10804
rect 18236 10752 18288 10804
rect 19800 10752 19852 10804
rect 19892 10795 19944 10804
rect 19892 10761 19901 10795
rect 19901 10761 19935 10795
rect 19935 10761 19944 10795
rect 19892 10752 19944 10761
rect 11152 10548 11204 10600
rect 11428 10591 11480 10600
rect 11428 10557 11437 10591
rect 11437 10557 11471 10591
rect 11471 10557 11480 10591
rect 11428 10548 11480 10557
rect 9220 10480 9272 10532
rect 9404 10480 9456 10532
rect 11796 10548 11848 10600
rect 12808 10616 12860 10668
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 12440 10548 12492 10600
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 11336 10412 11388 10464
rect 11428 10412 11480 10464
rect 13176 10591 13228 10600
rect 13176 10557 13185 10591
rect 13185 10557 13219 10591
rect 13219 10557 13228 10591
rect 13176 10548 13228 10557
rect 13912 10684 13964 10736
rect 13820 10616 13872 10668
rect 15384 10659 15436 10668
rect 13728 10591 13780 10600
rect 13728 10557 13737 10591
rect 13737 10557 13771 10591
rect 13771 10557 13780 10591
rect 13728 10548 13780 10557
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 14188 10548 14240 10600
rect 14556 10591 14608 10600
rect 14556 10557 14562 10591
rect 14562 10557 14596 10591
rect 14596 10557 14608 10591
rect 14556 10548 14608 10557
rect 14648 10548 14700 10600
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 15384 10616 15436 10625
rect 17040 10616 17092 10668
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 15292 10591 15344 10600
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 16120 10548 16172 10600
rect 16212 10548 16264 10600
rect 13820 10480 13872 10532
rect 16764 10591 16816 10600
rect 16764 10557 16773 10591
rect 16773 10557 16807 10591
rect 16807 10557 16816 10591
rect 16764 10548 16816 10557
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17592 10548 17644 10600
rect 19340 10548 19392 10600
rect 13176 10412 13228 10464
rect 20260 10616 20312 10668
rect 22100 10616 22152 10668
rect 14464 10412 14516 10464
rect 15384 10412 15436 10464
rect 17224 10412 17276 10464
rect 18512 10412 18564 10464
rect 19800 10412 19852 10464
rect 19984 10412 20036 10464
rect 20720 10591 20772 10600
rect 20720 10557 20729 10591
rect 20729 10557 20763 10591
rect 20763 10557 20772 10591
rect 20720 10548 20772 10557
rect 20812 10548 20864 10600
rect 22284 10548 22336 10600
rect 22836 10616 22888 10668
rect 21824 10412 21876 10464
rect 22928 10412 22980 10464
rect 4366 10310 4418 10362
rect 4430 10310 4482 10362
rect 4494 10310 4546 10362
rect 4558 10310 4610 10362
rect 4622 10310 4674 10362
rect 4686 10310 4738 10362
rect 10366 10310 10418 10362
rect 10430 10310 10482 10362
rect 10494 10310 10546 10362
rect 10558 10310 10610 10362
rect 10622 10310 10674 10362
rect 10686 10310 10738 10362
rect 16366 10310 16418 10362
rect 16430 10310 16482 10362
rect 16494 10310 16546 10362
rect 16558 10310 16610 10362
rect 16622 10310 16674 10362
rect 16686 10310 16738 10362
rect 22366 10310 22418 10362
rect 22430 10310 22482 10362
rect 22494 10310 22546 10362
rect 22558 10310 22610 10362
rect 22622 10310 22674 10362
rect 22686 10310 22738 10362
rect 1768 10208 1820 10260
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 2136 10208 2188 10260
rect 2688 10183 2740 10192
rect 2688 10149 2697 10183
rect 2697 10149 2731 10183
rect 2731 10149 2740 10183
rect 2688 10140 2740 10149
rect 3240 10183 3292 10192
rect 3240 10149 3267 10183
rect 3267 10149 3292 10183
rect 3240 10140 3292 10149
rect 6736 10208 6788 10260
rect 8116 10208 8168 10260
rect 8484 10208 8536 10260
rect 1216 10004 1268 10056
rect 1124 9868 1176 9920
rect 2044 9868 2096 9920
rect 2596 10115 2648 10124
rect 2596 10081 2605 10115
rect 2605 10081 2639 10115
rect 2639 10081 2648 10115
rect 2596 10072 2648 10081
rect 3332 10072 3384 10124
rect 4252 10072 4304 10124
rect 5540 10140 5592 10192
rect 7840 10115 7892 10124
rect 7840 10081 7849 10115
rect 7849 10081 7883 10115
rect 7883 10081 7892 10115
rect 7840 10072 7892 10081
rect 8300 10072 8352 10124
rect 8668 10115 8720 10124
rect 8668 10081 8677 10115
rect 8677 10081 8711 10115
rect 8711 10081 8720 10115
rect 8668 10072 8720 10081
rect 8852 10140 8904 10192
rect 9036 10072 9088 10124
rect 2780 9936 2832 9988
rect 2872 9936 2924 9988
rect 6000 9936 6052 9988
rect 6184 9936 6236 9988
rect 9956 10072 10008 10124
rect 11060 10208 11112 10260
rect 9312 10004 9364 10056
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 11428 10208 11480 10260
rect 11704 10208 11756 10260
rect 13728 10208 13780 10260
rect 14096 10208 14148 10260
rect 15292 10208 15344 10260
rect 16764 10208 16816 10260
rect 17132 10208 17184 10260
rect 18696 10208 18748 10260
rect 19064 10208 19116 10260
rect 19340 10208 19392 10260
rect 20168 10208 20220 10260
rect 21548 10251 21600 10260
rect 21548 10217 21557 10251
rect 21557 10217 21591 10251
rect 21591 10217 21600 10251
rect 21548 10208 21600 10217
rect 22192 10251 22244 10260
rect 22192 10217 22201 10251
rect 22201 10217 22235 10251
rect 22235 10217 22244 10251
rect 22192 10208 22244 10217
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 11336 10115 11388 10124
rect 11336 10081 11365 10115
rect 11365 10081 11388 10115
rect 12624 10140 12676 10192
rect 11336 10072 11388 10081
rect 11060 10004 11112 10056
rect 9220 9936 9272 9988
rect 12992 10072 13044 10124
rect 13176 10072 13228 10124
rect 14740 10140 14792 10192
rect 12716 10004 12768 10056
rect 14004 10072 14056 10124
rect 14280 10072 14332 10124
rect 14464 10072 14516 10124
rect 16028 10072 16080 10124
rect 16672 10072 16724 10124
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 15568 10004 15620 10056
rect 16212 10004 16264 10056
rect 16580 10004 16632 10056
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 17500 10115 17552 10124
rect 17500 10081 17509 10115
rect 17509 10081 17543 10115
rect 17543 10081 17552 10115
rect 17500 10072 17552 10081
rect 17776 10072 17828 10124
rect 18328 10072 18380 10124
rect 19340 10047 19392 10056
rect 19340 10013 19349 10047
rect 19349 10013 19383 10047
rect 19383 10013 19392 10047
rect 19340 10004 19392 10013
rect 19800 10072 19852 10124
rect 19892 10004 19944 10056
rect 20076 10004 20128 10056
rect 11796 9936 11848 9988
rect 3148 9868 3200 9920
rect 4068 9868 4120 9920
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 5540 9911 5592 9920
rect 5540 9877 5549 9911
rect 5549 9877 5583 9911
rect 5583 9877 5592 9911
rect 5540 9868 5592 9877
rect 6460 9868 6512 9920
rect 7288 9868 7340 9920
rect 7932 9868 7984 9920
rect 8300 9868 8352 9920
rect 8668 9868 8720 9920
rect 8852 9911 8904 9920
rect 8852 9877 8861 9911
rect 8861 9877 8895 9911
rect 8895 9877 8904 9911
rect 8852 9868 8904 9877
rect 9772 9868 9824 9920
rect 9956 9868 10008 9920
rect 10876 9868 10928 9920
rect 21180 9936 21232 9988
rect 13912 9868 13964 9920
rect 14648 9911 14700 9920
rect 14648 9877 14657 9911
rect 14657 9877 14691 9911
rect 14691 9877 14700 9911
rect 14648 9868 14700 9877
rect 14740 9868 14792 9920
rect 16120 9868 16172 9920
rect 16764 9868 16816 9920
rect 19248 9868 19300 9920
rect 20260 9868 20312 9920
rect 20628 9911 20680 9920
rect 20628 9877 20637 9911
rect 20637 9877 20671 9911
rect 20671 9877 20680 9911
rect 20628 9868 20680 9877
rect 21640 10072 21692 10124
rect 21548 10004 21600 10056
rect 21732 10047 21784 10056
rect 21732 10013 21741 10047
rect 21741 10013 21775 10047
rect 21775 10013 21784 10047
rect 21732 10004 21784 10013
rect 22192 10004 22244 10056
rect 22468 10072 22520 10124
rect 22744 9868 22796 9920
rect 1366 9766 1418 9818
rect 1430 9766 1482 9818
rect 1494 9766 1546 9818
rect 1558 9766 1610 9818
rect 1622 9766 1674 9818
rect 1686 9766 1738 9818
rect 7366 9766 7418 9818
rect 7430 9766 7482 9818
rect 7494 9766 7546 9818
rect 7558 9766 7610 9818
rect 7622 9766 7674 9818
rect 7686 9766 7738 9818
rect 13366 9766 13418 9818
rect 13430 9766 13482 9818
rect 13494 9766 13546 9818
rect 13558 9766 13610 9818
rect 13622 9766 13674 9818
rect 13686 9766 13738 9818
rect 19366 9766 19418 9818
rect 19430 9766 19482 9818
rect 19494 9766 19546 9818
rect 19558 9766 19610 9818
rect 19622 9766 19674 9818
rect 19686 9766 19738 9818
rect 2596 9664 2648 9716
rect 3240 9707 3292 9716
rect 3240 9673 3249 9707
rect 3249 9673 3283 9707
rect 3283 9673 3292 9707
rect 3240 9664 3292 9673
rect 2320 9460 2372 9512
rect 2412 9460 2464 9512
rect 3884 9528 3936 9580
rect 5540 9664 5592 9716
rect 6920 9664 6972 9716
rect 11612 9664 11664 9716
rect 11980 9664 12032 9716
rect 14740 9664 14792 9716
rect 5448 9639 5500 9648
rect 5448 9605 5457 9639
rect 5457 9605 5491 9639
rect 5491 9605 5500 9639
rect 5448 9596 5500 9605
rect 3148 9460 3200 9512
rect 3240 9460 3292 9512
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 4160 9460 4212 9512
rect 4712 9460 4764 9512
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 3884 9392 3936 9444
rect 2228 9324 2280 9376
rect 3148 9324 3200 9376
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 7288 9528 7340 9580
rect 5908 9460 5960 9512
rect 6460 9503 6512 9512
rect 6460 9469 6469 9503
rect 6469 9469 6503 9503
rect 6503 9469 6512 9503
rect 6460 9460 6512 9469
rect 5356 9392 5408 9444
rect 8116 9460 8168 9512
rect 12164 9528 12216 9580
rect 8944 9460 8996 9512
rect 9680 9460 9732 9512
rect 10232 9460 10284 9512
rect 12440 9528 12492 9580
rect 12900 9528 12952 9580
rect 13084 9528 13136 9580
rect 13176 9528 13228 9580
rect 13452 9528 13504 9580
rect 14004 9528 14056 9580
rect 6000 9435 6052 9444
rect 6000 9401 6009 9435
rect 6009 9401 6043 9435
rect 6043 9401 6052 9435
rect 6000 9392 6052 9401
rect 6552 9392 6604 9444
rect 7932 9392 7984 9444
rect 8852 9392 8904 9444
rect 5908 9324 5960 9376
rect 10784 9392 10836 9444
rect 13728 9460 13780 9512
rect 15016 9596 15068 9648
rect 16764 9707 16816 9716
rect 16764 9673 16773 9707
rect 16773 9673 16807 9707
rect 16807 9673 16816 9707
rect 16764 9664 16816 9673
rect 17040 9664 17092 9716
rect 17684 9664 17736 9716
rect 13084 9392 13136 9444
rect 14188 9392 14240 9444
rect 15568 9460 15620 9512
rect 15936 9528 15988 9580
rect 18328 9596 18380 9648
rect 20628 9664 20680 9716
rect 21180 9707 21232 9716
rect 21180 9673 21189 9707
rect 21189 9673 21223 9707
rect 21223 9673 21232 9707
rect 21180 9664 21232 9673
rect 21364 9664 21416 9716
rect 22100 9664 22152 9716
rect 22192 9664 22244 9716
rect 15660 9392 15712 9444
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 10968 9324 11020 9376
rect 11336 9324 11388 9376
rect 15844 9324 15896 9376
rect 16672 9460 16724 9512
rect 17868 9460 17920 9512
rect 18604 9528 18656 9580
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 19892 9596 19944 9648
rect 20536 9596 20588 9648
rect 20076 9528 20128 9580
rect 22008 9596 22060 9648
rect 22468 9664 22520 9716
rect 16856 9392 16908 9444
rect 16764 9324 16816 9376
rect 17224 9324 17276 9376
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 18696 9435 18748 9444
rect 18696 9401 18705 9435
rect 18705 9401 18739 9435
rect 18739 9401 18748 9435
rect 18696 9392 18748 9401
rect 18144 9324 18196 9376
rect 18788 9324 18840 9376
rect 18880 9367 18932 9376
rect 18880 9333 18905 9367
rect 18905 9333 18932 9367
rect 19524 9392 19576 9444
rect 19892 9426 19944 9478
rect 20812 9460 20864 9512
rect 21088 9503 21140 9512
rect 21088 9469 21097 9503
rect 21097 9469 21131 9503
rect 21131 9469 21140 9503
rect 21088 9460 21140 9469
rect 18880 9324 18932 9333
rect 19984 9324 20036 9376
rect 20720 9367 20772 9376
rect 20720 9333 20729 9367
rect 20729 9333 20763 9367
rect 20763 9333 20772 9367
rect 20720 9324 20772 9333
rect 21640 9460 21692 9512
rect 22192 9460 22244 9512
rect 22836 9460 22888 9512
rect 22100 9392 22152 9444
rect 22744 9435 22796 9444
rect 22744 9401 22753 9435
rect 22753 9401 22787 9435
rect 22787 9401 22796 9435
rect 22744 9392 22796 9401
rect 21640 9324 21692 9376
rect 22008 9324 22060 9376
rect 4366 9222 4418 9274
rect 4430 9222 4482 9274
rect 4494 9222 4546 9274
rect 4558 9222 4610 9274
rect 4622 9222 4674 9274
rect 4686 9222 4738 9274
rect 10366 9222 10418 9274
rect 10430 9222 10482 9274
rect 10494 9222 10546 9274
rect 10558 9222 10610 9274
rect 10622 9222 10674 9274
rect 10686 9222 10738 9274
rect 16366 9222 16418 9274
rect 16430 9222 16482 9274
rect 16494 9222 16546 9274
rect 16558 9222 16610 9274
rect 16622 9222 16674 9274
rect 16686 9222 16738 9274
rect 22366 9222 22418 9274
rect 22430 9222 22482 9274
rect 22494 9222 22546 9274
rect 22558 9222 22610 9274
rect 22622 9222 22674 9274
rect 22686 9222 22738 9274
rect 3516 9120 3568 9172
rect 2136 9027 2188 9036
rect 2136 8993 2145 9027
rect 2145 8993 2179 9027
rect 2179 8993 2188 9027
rect 2136 8984 2188 8993
rect 2228 9027 2280 9036
rect 2228 8993 2237 9027
rect 2237 8993 2271 9027
rect 2271 8993 2280 9027
rect 2228 8984 2280 8993
rect 2412 8984 2464 9036
rect 2596 8984 2648 9036
rect 3608 9052 3660 9104
rect 3240 9027 3292 9036
rect 3240 8993 3249 9027
rect 3249 8993 3283 9027
rect 3283 8993 3292 9027
rect 3240 8984 3292 8993
rect 3332 8848 3384 8900
rect 5264 9120 5316 9172
rect 8944 9120 8996 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 5816 9052 5868 9104
rect 3608 8959 3660 8968
rect 3608 8925 3617 8959
rect 3617 8925 3651 8959
rect 3651 8925 3660 8959
rect 3608 8916 3660 8925
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 4068 8984 4120 8993
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 5080 8984 5132 9036
rect 5540 8984 5592 9036
rect 6828 8984 6880 9036
rect 4252 8916 4304 8968
rect 5264 8916 5316 8968
rect 6644 8916 6696 8968
rect 5632 8848 5684 8900
rect 6092 8848 6144 8900
rect 9404 8984 9456 9036
rect 9680 9052 9732 9104
rect 9772 8848 9824 8900
rect 10324 9120 10376 9172
rect 10784 9120 10836 9172
rect 10968 9027 11020 9036
rect 10968 8993 10977 9027
rect 10977 8993 11011 9027
rect 11011 8993 11020 9027
rect 10968 8984 11020 8993
rect 11244 9027 11296 9036
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 11612 8916 11664 8968
rect 10232 8891 10284 8900
rect 10232 8857 10241 8891
rect 10241 8857 10275 8891
rect 10275 8857 10284 8891
rect 10232 8848 10284 8857
rect 11796 8984 11848 9036
rect 11980 9027 12032 9036
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 11980 8984 12032 8993
rect 12348 9052 12400 9104
rect 12440 8984 12492 9036
rect 12716 8984 12768 9036
rect 12808 9027 12860 9036
rect 12808 8993 12817 9027
rect 12817 8993 12851 9027
rect 12851 8993 12860 9027
rect 12808 8984 12860 8993
rect 12992 9052 13044 9104
rect 13452 9120 13504 9172
rect 13728 9120 13780 9172
rect 15476 9120 15528 9172
rect 15568 9120 15620 9172
rect 17776 9120 17828 9172
rect 13084 8984 13136 9036
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 13912 9027 13964 9036
rect 12072 8916 12124 8968
rect 13912 8993 13927 9027
rect 13927 8993 13961 9027
rect 13961 8993 13964 9027
rect 13912 8984 13964 8993
rect 2688 8780 2740 8832
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 2780 8780 2832 8789
rect 3148 8823 3200 8832
rect 3148 8789 3157 8823
rect 3157 8789 3191 8823
rect 3191 8789 3200 8823
rect 3148 8780 3200 8789
rect 3792 8780 3844 8832
rect 3884 8780 3936 8832
rect 5908 8780 5960 8832
rect 8668 8780 8720 8832
rect 9312 8780 9364 8832
rect 11428 8780 11480 8832
rect 11796 8780 11848 8832
rect 12256 8780 12308 8832
rect 12348 8823 12400 8832
rect 12348 8789 12357 8823
rect 12357 8789 12391 8823
rect 12391 8789 12400 8823
rect 12348 8780 12400 8789
rect 13176 8780 13228 8832
rect 13912 8848 13964 8900
rect 14280 8984 14332 9036
rect 14648 8916 14700 8968
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 15016 8959 15068 8968
rect 15016 8925 15025 8959
rect 15025 8925 15059 8959
rect 15059 8925 15068 8959
rect 15016 8916 15068 8925
rect 14924 8848 14976 8900
rect 14464 8780 14516 8832
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 16764 9052 16816 9104
rect 17592 9052 17644 9104
rect 17868 9095 17920 9104
rect 17868 9061 17893 9095
rect 17893 9061 17920 9095
rect 18788 9120 18840 9172
rect 20444 9120 20496 9172
rect 21732 9120 21784 9172
rect 22192 9120 22244 9172
rect 17868 9052 17920 9061
rect 18880 9052 18932 9104
rect 18328 9027 18380 9036
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 18512 8984 18564 9036
rect 19156 8984 19208 9036
rect 20076 9052 20128 9104
rect 21456 9052 21508 9104
rect 19340 8984 19392 9036
rect 19800 9027 19852 9036
rect 19800 8993 19809 9027
rect 19809 8993 19843 9027
rect 19843 8993 19852 9027
rect 19800 8984 19852 8993
rect 19984 8984 20036 9036
rect 20996 8984 21048 9036
rect 17224 8916 17276 8968
rect 15752 8780 15804 8832
rect 15936 8780 15988 8832
rect 16672 8780 16724 8832
rect 18144 8848 18196 8900
rect 18788 8848 18840 8900
rect 19064 8891 19116 8900
rect 19064 8857 19073 8891
rect 19073 8857 19107 8891
rect 19107 8857 19116 8891
rect 19064 8848 19116 8857
rect 19708 8916 19760 8968
rect 20168 8916 20220 8968
rect 20904 8916 20956 8968
rect 17684 8780 17736 8832
rect 17776 8780 17828 8832
rect 19340 8780 19392 8832
rect 19892 8780 19944 8832
rect 20260 8780 20312 8832
rect 20996 8780 21048 8832
rect 1366 8678 1418 8730
rect 1430 8678 1482 8730
rect 1494 8678 1546 8730
rect 1558 8678 1610 8730
rect 1622 8678 1674 8730
rect 1686 8678 1738 8730
rect 7366 8678 7418 8730
rect 7430 8678 7482 8730
rect 7494 8678 7546 8730
rect 7558 8678 7610 8730
rect 7622 8678 7674 8730
rect 7686 8678 7738 8730
rect 13366 8678 13418 8730
rect 13430 8678 13482 8730
rect 13494 8678 13546 8730
rect 13558 8678 13610 8730
rect 13622 8678 13674 8730
rect 13686 8678 13738 8730
rect 19366 8678 19418 8730
rect 19430 8678 19482 8730
rect 19494 8678 19546 8730
rect 19558 8678 19610 8730
rect 19622 8678 19674 8730
rect 19686 8678 19738 8730
rect 2320 8576 2372 8628
rect 2596 8576 2648 8628
rect 3056 8576 3108 8628
rect 3424 8576 3476 8628
rect 3700 8576 3752 8628
rect 10876 8576 10928 8628
rect 11796 8576 11848 8628
rect 12256 8576 12308 8628
rect 12900 8576 12952 8628
rect 15016 8576 15068 8628
rect 9956 8508 10008 8560
rect 11060 8508 11112 8560
rect 11520 8508 11572 8560
rect 3240 8440 3292 8492
rect 3332 8372 3384 8424
rect 4344 8440 4396 8492
rect 5540 8440 5592 8492
rect 5632 8440 5684 8492
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 9680 8440 9732 8492
rect 2688 8304 2740 8356
rect 2228 8236 2280 8288
rect 4160 8304 4212 8356
rect 3332 8236 3384 8288
rect 3792 8236 3844 8288
rect 4068 8236 4120 8288
rect 5080 8372 5132 8424
rect 5172 8372 5224 8424
rect 6276 8415 6328 8424
rect 6276 8381 6285 8415
rect 6285 8381 6319 8415
rect 6319 8381 6328 8415
rect 6276 8372 6328 8381
rect 6736 8372 6788 8424
rect 9128 8372 9180 8424
rect 11980 8440 12032 8492
rect 5908 8347 5960 8356
rect 5908 8313 5917 8347
rect 5917 8313 5951 8347
rect 5951 8313 5960 8347
rect 5908 8304 5960 8313
rect 6460 8304 6512 8356
rect 9312 8304 9364 8356
rect 11060 8304 11112 8356
rect 11336 8372 11388 8424
rect 11520 8415 11572 8424
rect 11520 8381 11529 8415
rect 11529 8381 11563 8415
rect 11563 8381 11572 8415
rect 11520 8372 11572 8381
rect 11888 8415 11940 8424
rect 11888 8381 11897 8415
rect 11897 8381 11931 8415
rect 11931 8381 11940 8415
rect 11888 8372 11940 8381
rect 14648 8508 14700 8560
rect 14832 8508 14884 8560
rect 14924 8508 14976 8560
rect 15844 8576 15896 8628
rect 16764 8576 16816 8628
rect 17224 8576 17276 8628
rect 17316 8619 17368 8628
rect 17316 8585 17325 8619
rect 17325 8585 17359 8619
rect 17359 8585 17368 8619
rect 17316 8576 17368 8585
rect 17592 8619 17644 8628
rect 17592 8585 17601 8619
rect 17601 8585 17635 8619
rect 17635 8585 17644 8619
rect 17592 8576 17644 8585
rect 18420 8576 18472 8628
rect 18880 8576 18932 8628
rect 19064 8576 19116 8628
rect 19248 8576 19300 8628
rect 19800 8576 19852 8628
rect 20076 8576 20128 8628
rect 20720 8576 20772 8628
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 22008 8576 22060 8628
rect 12532 8440 12584 8492
rect 13176 8440 13228 8492
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 14096 8440 14148 8492
rect 14464 8440 14516 8492
rect 15384 8440 15436 8492
rect 12900 8347 12952 8356
rect 12900 8313 12909 8347
rect 12909 8313 12943 8347
rect 12943 8313 12952 8347
rect 12900 8304 12952 8313
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 16028 8372 16080 8424
rect 16856 8440 16908 8492
rect 13728 8304 13780 8356
rect 14004 8304 14056 8356
rect 14464 8304 14516 8356
rect 4344 8236 4396 8288
rect 6000 8236 6052 8288
rect 7012 8279 7064 8288
rect 7012 8245 7021 8279
rect 7021 8245 7055 8279
rect 7055 8245 7064 8279
rect 7012 8236 7064 8245
rect 11704 8236 11756 8288
rect 12532 8236 12584 8288
rect 12808 8236 12860 8288
rect 13084 8236 13136 8288
rect 13176 8236 13228 8288
rect 14188 8236 14240 8288
rect 15292 8236 15344 8288
rect 16580 8415 16632 8424
rect 16580 8381 16589 8415
rect 16589 8381 16623 8415
rect 16623 8381 16632 8415
rect 16580 8372 16632 8381
rect 16672 8372 16724 8424
rect 17316 8372 17368 8424
rect 17684 8372 17736 8424
rect 17868 8372 17920 8424
rect 19340 8372 19392 8424
rect 19984 8508 20036 8560
rect 21456 8508 21508 8560
rect 21272 8483 21324 8492
rect 21272 8449 21281 8483
rect 21281 8449 21315 8483
rect 21315 8449 21324 8483
rect 21272 8440 21324 8449
rect 21640 8440 21692 8492
rect 20536 8372 20588 8424
rect 21364 8372 21416 8424
rect 22928 8440 22980 8492
rect 19984 8304 20036 8356
rect 20260 8304 20312 8356
rect 21180 8347 21232 8356
rect 21180 8313 21189 8347
rect 21189 8313 21223 8347
rect 21223 8313 21232 8347
rect 21180 8304 21232 8313
rect 21272 8304 21324 8356
rect 17592 8236 17644 8288
rect 18696 8279 18748 8288
rect 18696 8245 18705 8279
rect 18705 8245 18739 8279
rect 18739 8245 18748 8279
rect 18696 8236 18748 8245
rect 19800 8236 19852 8288
rect 4366 8134 4418 8186
rect 4430 8134 4482 8186
rect 4494 8134 4546 8186
rect 4558 8134 4610 8186
rect 4622 8134 4674 8186
rect 4686 8134 4738 8186
rect 10366 8134 10418 8186
rect 10430 8134 10482 8186
rect 10494 8134 10546 8186
rect 10558 8134 10610 8186
rect 10622 8134 10674 8186
rect 10686 8134 10738 8186
rect 16366 8134 16418 8186
rect 16430 8134 16482 8186
rect 16494 8134 16546 8186
rect 16558 8134 16610 8186
rect 16622 8134 16674 8186
rect 16686 8134 16738 8186
rect 22366 8134 22418 8186
rect 22430 8134 22482 8186
rect 22494 8134 22546 8186
rect 22558 8134 22610 8186
rect 22622 8134 22674 8186
rect 22686 8134 22738 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 1124 7939 1176 7948
rect 1124 7905 1158 7939
rect 1158 7905 1176 7939
rect 1124 7896 1176 7905
rect 2688 7896 2740 7948
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 3516 8032 3568 8084
rect 4068 8032 4120 8084
rect 4988 8032 5040 8084
rect 5080 8032 5132 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 6000 8075 6052 8084
rect 5172 8032 5224 8041
rect 6000 8041 6009 8075
rect 6009 8041 6043 8075
rect 6043 8041 6052 8075
rect 6000 8032 6052 8041
rect 6092 8032 6144 8084
rect 11888 8032 11940 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 13728 8032 13780 8084
rect 13820 8032 13872 8084
rect 3332 7964 3384 8016
rect 848 7871 900 7880
rect 848 7837 857 7871
rect 857 7837 891 7871
rect 891 7837 900 7871
rect 848 7828 900 7837
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 3516 7896 3568 7948
rect 3148 7760 3200 7812
rect 6184 7964 6236 8016
rect 6644 7964 6696 8016
rect 11520 7964 11572 8016
rect 3976 7760 4028 7812
rect 6828 7896 6880 7948
rect 9312 7939 9364 7948
rect 9312 7905 9321 7939
rect 9321 7905 9355 7939
rect 9355 7905 9364 7939
rect 9312 7896 9364 7905
rect 10232 7896 10284 7948
rect 11152 7896 11204 7948
rect 11244 7896 11296 7948
rect 12532 7964 12584 8016
rect 12348 7896 12400 7948
rect 12716 7896 12768 7948
rect 13268 7896 13320 7948
rect 14004 7939 14056 7948
rect 14004 7905 14013 7939
rect 14013 7905 14047 7939
rect 14047 7905 14056 7939
rect 14004 7896 14056 7905
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 14188 7939 14240 7948
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 14832 8032 14884 8084
rect 14924 8032 14976 8084
rect 17040 8032 17092 8084
rect 5632 7828 5684 7880
rect 8852 7871 8904 7880
rect 8852 7837 8861 7871
rect 8861 7837 8895 7871
rect 8895 7837 8904 7871
rect 8852 7828 8904 7837
rect 13176 7828 13228 7880
rect 14648 7939 14700 7948
rect 14648 7905 14657 7939
rect 14657 7905 14691 7939
rect 14691 7905 14700 7939
rect 14648 7896 14700 7905
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 17500 7964 17552 8016
rect 15476 7828 15528 7880
rect 4160 7692 4212 7744
rect 5356 7692 5408 7744
rect 6000 7692 6052 7744
rect 7196 7692 7248 7744
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 11152 7760 11204 7812
rect 11612 7760 11664 7812
rect 11980 7692 12032 7744
rect 18696 7896 18748 7948
rect 19800 7896 19852 7948
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 17776 7828 17828 7880
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 20536 7896 20588 7948
rect 20812 7896 20864 7948
rect 20260 7828 20312 7880
rect 20720 7828 20772 7880
rect 15476 7692 15528 7744
rect 16764 7692 16816 7744
rect 17132 7692 17184 7744
rect 17960 7692 18012 7744
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 18788 7692 18840 7701
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 21088 7735 21140 7744
rect 21088 7701 21097 7735
rect 21097 7701 21131 7735
rect 21131 7701 21140 7735
rect 21088 7692 21140 7701
rect 21364 7692 21416 7744
rect 1366 7590 1418 7642
rect 1430 7590 1482 7642
rect 1494 7590 1546 7642
rect 1558 7590 1610 7642
rect 1622 7590 1674 7642
rect 1686 7590 1738 7642
rect 7366 7590 7418 7642
rect 7430 7590 7482 7642
rect 7494 7590 7546 7642
rect 7558 7590 7610 7642
rect 7622 7590 7674 7642
rect 7686 7590 7738 7642
rect 13366 7590 13418 7642
rect 13430 7590 13482 7642
rect 13494 7590 13546 7642
rect 13558 7590 13610 7642
rect 13622 7590 13674 7642
rect 13686 7590 13738 7642
rect 19366 7590 19418 7642
rect 19430 7590 19482 7642
rect 19494 7590 19546 7642
rect 19558 7590 19610 7642
rect 19622 7590 19674 7642
rect 19686 7590 19738 7642
rect 1124 7488 1176 7540
rect 2872 7488 2924 7540
rect 3332 7488 3384 7540
rect 2596 7352 2648 7404
rect 2964 7352 3016 7404
rect 5448 7488 5500 7540
rect 7196 7488 7248 7540
rect 7288 7488 7340 7540
rect 4068 7420 4120 7472
rect 4160 7463 4212 7472
rect 4160 7429 4169 7463
rect 4169 7429 4203 7463
rect 4203 7429 4212 7463
rect 4160 7420 4212 7429
rect 10876 7420 10928 7472
rect 11888 7420 11940 7472
rect 12808 7488 12860 7540
rect 13544 7488 13596 7540
rect 13728 7488 13780 7540
rect 5632 7352 5684 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 1860 7284 1912 7336
rect 2412 7284 2464 7336
rect 3240 7216 3292 7268
rect 3516 7327 3568 7336
rect 3516 7293 3525 7327
rect 3525 7293 3559 7327
rect 3559 7293 3568 7327
rect 3516 7284 3568 7293
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 3792 7327 3844 7336
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 3792 7284 3844 7293
rect 4068 7284 4120 7336
rect 4252 7284 4304 7336
rect 4988 7284 5040 7336
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5172 7284 5224 7293
rect 7840 7352 7892 7404
rect 12440 7352 12492 7404
rect 12532 7352 12584 7404
rect 13176 7352 13228 7404
rect 13268 7352 13320 7404
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 5264 7216 5316 7268
rect 5540 7216 5592 7268
rect 10692 7284 10744 7336
rect 4252 7148 4304 7200
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 6460 7148 6512 7200
rect 10232 7216 10284 7268
rect 10968 7284 11020 7336
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 11152 7327 11204 7336
rect 11152 7293 11161 7327
rect 11161 7293 11195 7327
rect 11195 7293 11204 7327
rect 11152 7284 11204 7293
rect 11244 7327 11296 7336
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 11888 7327 11940 7336
rect 11888 7293 11897 7327
rect 11897 7293 11931 7327
rect 11931 7293 11940 7327
rect 11888 7284 11940 7293
rect 12808 7284 12860 7336
rect 12992 7284 13044 7336
rect 11336 7148 11388 7200
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 11612 7148 11664 7200
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 12532 7216 12584 7268
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 14740 7420 14792 7472
rect 14832 7420 14884 7472
rect 15108 7420 15160 7472
rect 15660 7488 15712 7540
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 13912 7395 13964 7404
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 13452 7216 13504 7268
rect 13636 7216 13688 7268
rect 14188 7284 14240 7336
rect 15476 7352 15528 7404
rect 15844 7352 15896 7404
rect 17408 7463 17460 7472
rect 17408 7429 17417 7463
rect 17417 7429 17451 7463
rect 17451 7429 17460 7463
rect 17408 7420 17460 7429
rect 16764 7352 16816 7404
rect 18696 7488 18748 7540
rect 18788 7488 18840 7540
rect 19340 7488 19392 7540
rect 20352 7531 20404 7540
rect 20352 7497 20361 7531
rect 20361 7497 20395 7531
rect 20395 7497 20404 7531
rect 20352 7488 20404 7497
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 21088 7488 21140 7540
rect 20536 7420 20588 7472
rect 14464 7216 14516 7268
rect 13728 7148 13780 7200
rect 13820 7148 13872 7200
rect 14648 7148 14700 7200
rect 16856 7284 16908 7336
rect 17684 7284 17736 7336
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 18696 7327 18748 7336
rect 18696 7293 18705 7327
rect 18705 7293 18739 7327
rect 18739 7293 18748 7327
rect 18696 7284 18748 7293
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 19800 7284 19852 7336
rect 21364 7284 21416 7336
rect 17040 7148 17092 7200
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 17960 7148 18012 7200
rect 4366 7046 4418 7098
rect 4430 7046 4482 7098
rect 4494 7046 4546 7098
rect 4558 7046 4610 7098
rect 4622 7046 4674 7098
rect 4686 7046 4738 7098
rect 10366 7046 10418 7098
rect 10430 7046 10482 7098
rect 10494 7046 10546 7098
rect 10558 7046 10610 7098
rect 10622 7046 10674 7098
rect 10686 7046 10738 7098
rect 16366 7046 16418 7098
rect 16430 7046 16482 7098
rect 16494 7046 16546 7098
rect 16558 7046 16610 7098
rect 16622 7046 16674 7098
rect 16686 7046 16738 7098
rect 22366 7046 22418 7098
rect 22430 7046 22482 7098
rect 22494 7046 22546 7098
rect 22558 7046 22610 7098
rect 22622 7046 22674 7098
rect 22686 7046 22738 7098
rect 1400 6944 1452 6996
rect 2136 6944 2188 6996
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 2596 6919 2648 6928
rect 2596 6885 2623 6919
rect 2623 6885 2648 6919
rect 2596 6876 2648 6885
rect 2964 6876 3016 6928
rect 3516 6944 3568 6996
rect 3792 6987 3844 6996
rect 3792 6953 3801 6987
rect 3801 6953 3835 6987
rect 3835 6953 3844 6987
rect 3792 6944 3844 6953
rect 4068 6944 4120 6996
rect 5264 6944 5316 6996
rect 6092 6944 6144 6996
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 5448 6876 5500 6928
rect 6368 6944 6420 6996
rect 9956 6944 10008 6996
rect 10232 6944 10284 6996
rect 11152 6944 11204 6996
rect 11336 6944 11388 6996
rect 11704 6944 11756 6996
rect 12072 6944 12124 6996
rect 12348 6944 12400 6996
rect 6460 6876 6512 6928
rect 3240 6740 3292 6792
rect 3608 6808 3660 6860
rect 3700 6808 3752 6860
rect 3976 6851 4028 6860
rect 3976 6817 3985 6851
rect 3985 6817 4019 6851
rect 4019 6817 4028 6851
rect 3976 6808 4028 6817
rect 4804 6808 4856 6860
rect 5908 6808 5960 6860
rect 6736 6808 6788 6860
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 8300 6876 8352 6928
rect 8576 6876 8628 6928
rect 9036 6876 9088 6928
rect 10692 6876 10744 6928
rect 13176 6944 13228 6996
rect 13452 6944 13504 6996
rect 4252 6740 4304 6792
rect 5632 6740 5684 6792
rect 9588 6808 9640 6860
rect 9404 6740 9456 6792
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 2872 6604 2924 6656
rect 3792 6604 3844 6656
rect 4160 6604 4212 6656
rect 5080 6604 5132 6656
rect 6276 6604 6328 6656
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 11060 6808 11112 6860
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 12624 6876 12676 6928
rect 11612 6808 11664 6860
rect 11888 6808 11940 6860
rect 10876 6672 10928 6724
rect 9404 6604 9456 6656
rect 10600 6604 10652 6656
rect 10784 6604 10836 6656
rect 11244 6604 11296 6656
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 11888 6604 11940 6656
rect 12716 6740 12768 6792
rect 13728 6808 13780 6860
rect 14004 6808 14056 6860
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 14096 6808 14148 6817
rect 14740 6808 14792 6860
rect 15660 6876 15712 6928
rect 16120 6876 16172 6928
rect 16764 6944 16816 6996
rect 17040 6944 17092 6996
rect 17408 6944 17460 6996
rect 21272 6987 21324 6996
rect 21272 6953 21281 6987
rect 21281 6953 21315 6987
rect 21315 6953 21324 6987
rect 21272 6944 21324 6953
rect 17960 6876 18012 6928
rect 13084 6672 13136 6724
rect 13452 6672 13504 6724
rect 13912 6672 13964 6724
rect 17224 6740 17276 6792
rect 17868 6808 17920 6860
rect 20352 6808 20404 6860
rect 18696 6740 18748 6792
rect 21824 6808 21876 6860
rect 21916 6808 21968 6860
rect 14464 6604 14516 6656
rect 14648 6647 14700 6656
rect 14648 6613 14657 6647
rect 14657 6613 14691 6647
rect 14691 6613 14700 6647
rect 14648 6604 14700 6613
rect 14924 6604 14976 6656
rect 15108 6604 15160 6656
rect 20720 6604 20772 6656
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 21732 6604 21784 6656
rect 1366 6502 1418 6554
rect 1430 6502 1482 6554
rect 1494 6502 1546 6554
rect 1558 6502 1610 6554
rect 1622 6502 1674 6554
rect 1686 6502 1738 6554
rect 7366 6502 7418 6554
rect 7430 6502 7482 6554
rect 7494 6502 7546 6554
rect 7558 6502 7610 6554
rect 7622 6502 7674 6554
rect 7686 6502 7738 6554
rect 13366 6502 13418 6554
rect 13430 6502 13482 6554
rect 13494 6502 13546 6554
rect 13558 6502 13610 6554
rect 13622 6502 13674 6554
rect 13686 6502 13738 6554
rect 19366 6502 19418 6554
rect 19430 6502 19482 6554
rect 19494 6502 19546 6554
rect 19558 6502 19610 6554
rect 19622 6502 19674 6554
rect 19686 6502 19738 6554
rect 1952 6400 2004 6452
rect 1676 6332 1728 6384
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 2412 6400 2464 6452
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 3608 6400 3660 6452
rect 5540 6400 5592 6452
rect 6000 6400 6052 6452
rect 8576 6443 8628 6452
rect 8576 6409 8585 6443
rect 8585 6409 8619 6443
rect 8619 6409 8628 6443
rect 8576 6400 8628 6409
rect 8024 6332 8076 6384
rect 9036 6332 9088 6384
rect 10508 6400 10560 6452
rect 10600 6400 10652 6452
rect 12072 6400 12124 6452
rect 12808 6400 12860 6452
rect 17592 6400 17644 6452
rect 20720 6400 20772 6452
rect 21824 6400 21876 6452
rect 2228 6196 2280 6248
rect 3792 6264 3844 6316
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 5724 6264 5776 6316
rect 7104 6264 7156 6316
rect 10876 6264 10928 6316
rect 11520 6332 11572 6384
rect 11428 6264 11480 6316
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 13728 6332 13780 6384
rect 14188 6332 14240 6384
rect 15016 6332 15068 6384
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 15292 6264 15344 6273
rect 4988 6128 5040 6180
rect 5448 6128 5500 6180
rect 6184 6196 6236 6248
rect 6552 6196 6604 6248
rect 10600 6196 10652 6248
rect 11520 6196 11572 6248
rect 11612 6239 11664 6248
rect 11612 6205 11620 6239
rect 11620 6205 11654 6239
rect 11654 6205 11664 6239
rect 11612 6196 11664 6205
rect 6736 6171 6788 6180
rect 6736 6137 6745 6171
rect 6745 6137 6779 6171
rect 6779 6137 6788 6171
rect 6736 6128 6788 6137
rect 1952 6060 2004 6112
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 2780 6103 2832 6112
rect 2780 6069 2797 6103
rect 2797 6069 2832 6103
rect 2780 6060 2832 6069
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 11336 6128 11388 6180
rect 5724 6060 5776 6069
rect 7196 6060 7248 6112
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 8300 6060 8352 6112
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 10232 6060 10284 6112
rect 12164 6171 12216 6180
rect 12164 6137 12173 6171
rect 12173 6137 12207 6171
rect 12207 6137 12216 6171
rect 12164 6128 12216 6137
rect 12808 6128 12860 6180
rect 13820 6196 13872 6248
rect 13912 6196 13964 6248
rect 15016 6239 15068 6248
rect 15016 6205 15025 6239
rect 15025 6205 15059 6239
rect 15059 6205 15068 6239
rect 15016 6196 15068 6205
rect 15108 6196 15160 6248
rect 11980 6060 12032 6112
rect 12256 6060 12308 6112
rect 12532 6103 12584 6112
rect 12532 6069 12541 6103
rect 12541 6069 12575 6103
rect 12575 6069 12584 6103
rect 12532 6060 12584 6069
rect 12992 6060 13044 6112
rect 16856 6196 16908 6248
rect 17868 6196 17920 6248
rect 17960 6239 18012 6248
rect 17960 6205 17969 6239
rect 17969 6205 18003 6239
rect 18003 6205 18012 6239
rect 17960 6196 18012 6205
rect 18788 6264 18840 6316
rect 18328 6196 18380 6248
rect 20996 6307 21048 6316
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 15936 6171 15988 6180
rect 15936 6137 15945 6171
rect 15945 6137 15979 6171
rect 15979 6137 15988 6171
rect 15936 6128 15988 6137
rect 16120 6060 16172 6112
rect 17776 6128 17828 6180
rect 19800 6196 19852 6248
rect 21272 6264 21324 6316
rect 18144 6060 18196 6112
rect 20904 6171 20956 6180
rect 20904 6137 20913 6171
rect 20913 6137 20947 6171
rect 20947 6137 20956 6171
rect 20904 6128 20956 6137
rect 20996 6128 21048 6180
rect 19064 6060 19116 6112
rect 21548 6060 21600 6112
rect 4366 5958 4418 6010
rect 4430 5958 4482 6010
rect 4494 5958 4546 6010
rect 4558 5958 4610 6010
rect 4622 5958 4674 6010
rect 4686 5958 4738 6010
rect 10366 5958 10418 6010
rect 10430 5958 10482 6010
rect 10494 5958 10546 6010
rect 10558 5958 10610 6010
rect 10622 5958 10674 6010
rect 10686 5958 10738 6010
rect 16366 5958 16418 6010
rect 16430 5958 16482 6010
rect 16494 5958 16546 6010
rect 16558 5958 16610 6010
rect 16622 5958 16674 6010
rect 16686 5958 16738 6010
rect 22366 5958 22418 6010
rect 22430 5958 22482 6010
rect 22494 5958 22546 6010
rect 22558 5958 22610 6010
rect 22622 5958 22674 6010
rect 22686 5958 22738 6010
rect 1952 5856 2004 5908
rect 3792 5856 3844 5908
rect 5448 5856 5500 5908
rect 6736 5856 6788 5908
rect 7012 5856 7064 5908
rect 7196 5856 7248 5908
rect 8208 5856 8260 5908
rect 8392 5899 8444 5908
rect 8392 5865 8401 5899
rect 8401 5865 8435 5899
rect 8435 5865 8444 5899
rect 8392 5856 8444 5865
rect 8576 5856 8628 5908
rect 2044 5831 2096 5840
rect 2044 5797 2053 5831
rect 2053 5797 2087 5831
rect 2087 5797 2096 5831
rect 2044 5788 2096 5797
rect 848 5720 900 5772
rect 2412 5720 2464 5772
rect 4988 5720 5040 5772
rect 6644 5788 6696 5840
rect 9680 5856 9732 5908
rect 11612 5899 11664 5908
rect 11612 5865 11621 5899
rect 11621 5865 11655 5899
rect 11655 5865 11664 5899
rect 11612 5856 11664 5865
rect 12072 5856 12124 5908
rect 12256 5856 12308 5908
rect 12532 5856 12584 5908
rect 12808 5856 12860 5908
rect 5908 5720 5960 5772
rect 6460 5720 6512 5772
rect 7104 5720 7156 5772
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 3332 5652 3384 5704
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 3700 5559 3752 5568
rect 3700 5525 3709 5559
rect 3709 5525 3743 5559
rect 3743 5525 3752 5559
rect 3700 5516 3752 5525
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5724 5652 5776 5704
rect 5632 5584 5684 5636
rect 7932 5652 7984 5704
rect 8392 5652 8444 5704
rect 9036 5720 9088 5772
rect 9312 5720 9364 5772
rect 9588 5720 9640 5772
rect 10140 5720 10192 5772
rect 10876 5720 10928 5772
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 11520 5788 11572 5840
rect 11980 5788 12032 5840
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 11152 5584 11204 5636
rect 7196 5559 7248 5568
rect 7196 5525 7205 5559
rect 7205 5525 7239 5559
rect 7239 5525 7248 5559
rect 7196 5516 7248 5525
rect 7932 5516 7984 5568
rect 9036 5516 9088 5568
rect 10784 5516 10836 5568
rect 11796 5720 11848 5772
rect 14924 5856 14976 5908
rect 15016 5856 15068 5908
rect 15936 5856 15988 5908
rect 17040 5856 17092 5908
rect 17592 5856 17644 5908
rect 17960 5856 18012 5908
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 14004 5788 14056 5840
rect 13176 5720 13228 5772
rect 13268 5763 13320 5772
rect 13268 5729 13277 5763
rect 13277 5729 13311 5763
rect 13311 5729 13320 5763
rect 13268 5720 13320 5729
rect 15752 5788 15804 5840
rect 15016 5720 15068 5772
rect 15568 5720 15620 5772
rect 16856 5720 16908 5772
rect 17040 5763 17092 5772
rect 17040 5729 17049 5763
rect 17049 5729 17083 5763
rect 17083 5729 17092 5763
rect 17040 5720 17092 5729
rect 17224 5788 17276 5840
rect 13912 5652 13964 5704
rect 14648 5652 14700 5704
rect 14924 5652 14976 5704
rect 12532 5516 12584 5568
rect 13176 5516 13228 5568
rect 14464 5516 14516 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 17224 5584 17276 5636
rect 16856 5559 16908 5568
rect 16856 5525 16865 5559
rect 16865 5525 16899 5559
rect 16899 5525 16908 5559
rect 16856 5516 16908 5525
rect 17868 5695 17920 5704
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 18144 5720 18196 5772
rect 22100 5899 22152 5908
rect 22100 5865 22109 5899
rect 22109 5865 22143 5899
rect 22143 5865 22152 5899
rect 22100 5856 22152 5865
rect 18788 5720 18840 5772
rect 18880 5720 18932 5772
rect 19156 5763 19208 5772
rect 19156 5729 19165 5763
rect 19165 5729 19199 5763
rect 19199 5729 19208 5763
rect 19156 5720 19208 5729
rect 19800 5720 19852 5772
rect 21824 5720 21876 5772
rect 21916 5763 21968 5772
rect 21916 5729 21925 5763
rect 21925 5729 21959 5763
rect 21959 5729 21968 5763
rect 21916 5720 21968 5729
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 21364 5584 21416 5636
rect 21732 5584 21784 5636
rect 19064 5516 19116 5568
rect 22100 5516 22152 5568
rect 1366 5414 1418 5466
rect 1430 5414 1482 5466
rect 1494 5414 1546 5466
rect 1558 5414 1610 5466
rect 1622 5414 1674 5466
rect 1686 5414 1738 5466
rect 7366 5414 7418 5466
rect 7430 5414 7482 5466
rect 7494 5414 7546 5466
rect 7558 5414 7610 5466
rect 7622 5414 7674 5466
rect 7686 5414 7738 5466
rect 13366 5414 13418 5466
rect 13430 5414 13482 5466
rect 13494 5414 13546 5466
rect 13558 5414 13610 5466
rect 13622 5414 13674 5466
rect 13686 5414 13738 5466
rect 19366 5414 19418 5466
rect 19430 5414 19482 5466
rect 19494 5414 19546 5466
rect 19558 5414 19610 5466
rect 19622 5414 19674 5466
rect 19686 5414 19738 5466
rect 1768 5312 1820 5364
rect 5908 5312 5960 5364
rect 6920 5312 6972 5364
rect 7932 5312 7984 5364
rect 8300 5312 8352 5364
rect 8576 5312 8628 5364
rect 9312 5312 9364 5364
rect 2780 5244 2832 5296
rect 11060 5312 11112 5364
rect 11152 5312 11204 5364
rect 11704 5312 11756 5364
rect 11796 5312 11848 5364
rect 13728 5312 13780 5364
rect 14832 5312 14884 5364
rect 15568 5312 15620 5364
rect 15752 5312 15804 5364
rect 16212 5312 16264 5364
rect 17592 5312 17644 5364
rect 19156 5312 19208 5364
rect 20904 5312 20956 5364
rect 21548 5312 21600 5364
rect 21640 5312 21692 5364
rect 2320 5176 2372 5228
rect 2228 5151 2280 5160
rect 2228 5117 2237 5151
rect 2237 5117 2271 5151
rect 2271 5117 2280 5151
rect 5080 5176 5132 5228
rect 5632 5176 5684 5228
rect 2228 5108 2280 5117
rect 5448 5151 5500 5160
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 6644 5176 6696 5228
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 3516 4972 3568 5024
rect 5816 4972 5868 5024
rect 6092 4972 6144 5024
rect 6828 4972 6880 5024
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 9220 5108 9272 5160
rect 9404 5108 9456 5160
rect 11336 5244 11388 5296
rect 11888 5244 11940 5296
rect 11152 5151 11204 5160
rect 11152 5117 11161 5151
rect 11161 5117 11195 5151
rect 11195 5117 11204 5151
rect 11152 5108 11204 5117
rect 11428 5108 11480 5160
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 9956 5040 10008 5092
rect 11612 5040 11664 5092
rect 11980 5151 12032 5160
rect 11980 5117 11989 5151
rect 11989 5117 12023 5151
rect 12023 5117 12032 5151
rect 11980 5108 12032 5117
rect 12164 5108 12216 5160
rect 12440 5108 12492 5160
rect 12532 5108 12584 5160
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 13636 5108 13688 5160
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 14188 5108 14240 5160
rect 8576 4972 8628 5024
rect 9036 4972 9088 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 11704 4972 11756 5024
rect 12164 5015 12216 5024
rect 12164 4981 12173 5015
rect 12173 4981 12207 5015
rect 12207 4981 12216 5015
rect 12164 4972 12216 4981
rect 14556 5040 14608 5092
rect 13176 4972 13228 5024
rect 15384 5176 15436 5228
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16028 5176 16080 5228
rect 16212 5176 16264 5228
rect 17224 5176 17276 5228
rect 15200 5151 15252 5160
rect 15200 5117 15209 5151
rect 15209 5117 15243 5151
rect 15243 5117 15252 5151
rect 15200 5108 15252 5117
rect 14832 5040 14884 5092
rect 15660 5108 15712 5160
rect 17040 5108 17092 5160
rect 18880 5287 18932 5296
rect 18880 5253 18889 5287
rect 18889 5253 18923 5287
rect 18923 5253 18932 5287
rect 18880 5244 18932 5253
rect 20352 5244 20404 5296
rect 22100 5176 22152 5228
rect 18236 5108 18288 5160
rect 18420 5108 18472 5160
rect 20352 5108 20404 5160
rect 21364 5151 21416 5160
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 21456 5151 21508 5160
rect 21456 5117 21465 5151
rect 21465 5117 21499 5151
rect 21499 5117 21508 5151
rect 21456 5108 21508 5117
rect 21824 5108 21876 5160
rect 21916 5151 21968 5160
rect 21916 5117 21925 5151
rect 21925 5117 21959 5151
rect 21959 5117 21968 5151
rect 21916 5108 21968 5117
rect 14924 4972 14976 5024
rect 15200 4972 15252 5024
rect 15660 5015 15712 5024
rect 15660 4981 15669 5015
rect 15669 4981 15703 5015
rect 15703 4981 15712 5015
rect 15660 4972 15712 4981
rect 16856 4972 16908 5024
rect 17868 5015 17920 5024
rect 17868 4981 17877 5015
rect 17877 4981 17911 5015
rect 17911 4981 17920 5015
rect 17868 4972 17920 4981
rect 19984 5040 20036 5092
rect 21088 5040 21140 5092
rect 21548 4972 21600 5024
rect 4366 4870 4418 4922
rect 4430 4870 4482 4922
rect 4494 4870 4546 4922
rect 4558 4870 4610 4922
rect 4622 4870 4674 4922
rect 4686 4870 4738 4922
rect 10366 4870 10418 4922
rect 10430 4870 10482 4922
rect 10494 4870 10546 4922
rect 10558 4870 10610 4922
rect 10622 4870 10674 4922
rect 10686 4870 10738 4922
rect 16366 4870 16418 4922
rect 16430 4870 16482 4922
rect 16494 4870 16546 4922
rect 16558 4870 16610 4922
rect 16622 4870 16674 4922
rect 16686 4870 16738 4922
rect 22366 4870 22418 4922
rect 22430 4870 22482 4922
rect 22494 4870 22546 4922
rect 22558 4870 22610 4922
rect 22622 4870 22674 4922
rect 22686 4870 22738 4922
rect 2320 4768 2372 4820
rect 2688 4811 2740 4820
rect 2688 4777 2697 4811
rect 2697 4777 2731 4811
rect 2731 4777 2740 4811
rect 2688 4768 2740 4777
rect 4160 4768 4212 4820
rect 5448 4768 5500 4820
rect 6644 4768 6696 4820
rect 8668 4768 8720 4820
rect 9404 4768 9456 4820
rect 3700 4700 3752 4752
rect 848 4632 900 4684
rect 3608 4675 3660 4684
rect 3608 4641 3617 4675
rect 3617 4641 3651 4675
rect 3651 4641 3660 4675
rect 3608 4632 3660 4641
rect 4344 4632 4396 4684
rect 3792 4564 3844 4616
rect 4160 4564 4212 4616
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6092 4700 6144 4752
rect 12348 4768 12400 4820
rect 12808 4768 12860 4820
rect 14740 4768 14792 4820
rect 16856 4811 16908 4820
rect 16856 4777 16865 4811
rect 16865 4777 16899 4811
rect 16899 4777 16908 4811
rect 16856 4768 16908 4777
rect 20812 4768 20864 4820
rect 21180 4768 21232 4820
rect 21916 4768 21968 4820
rect 22284 4768 22336 4820
rect 7196 4632 7248 4684
rect 7472 4632 7524 4684
rect 10784 4632 10836 4684
rect 11704 4675 11756 4684
rect 11704 4641 11713 4675
rect 11713 4641 11747 4675
rect 11747 4641 11756 4675
rect 11704 4632 11756 4641
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 13912 4700 13964 4752
rect 14004 4700 14056 4752
rect 13820 4675 13872 4684
rect 13820 4641 13829 4675
rect 13829 4641 13863 4675
rect 13863 4641 13872 4675
rect 13820 4632 13872 4641
rect 14188 4632 14240 4684
rect 15108 4632 15160 4684
rect 15936 4700 15988 4752
rect 15384 4675 15436 4684
rect 15384 4641 15393 4675
rect 15393 4641 15427 4675
rect 15427 4641 15436 4675
rect 15384 4632 15436 4641
rect 15568 4675 15620 4684
rect 15568 4641 15577 4675
rect 15577 4641 15611 4675
rect 15611 4641 15620 4675
rect 15568 4632 15620 4641
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 16212 4700 16264 4752
rect 7748 4564 7800 4616
rect 10508 4564 10560 4616
rect 11796 4564 11848 4616
rect 6092 4496 6144 4548
rect 7196 4496 7248 4548
rect 7656 4496 7708 4548
rect 11980 4496 12032 4548
rect 12808 4607 12860 4616
rect 12808 4573 12817 4607
rect 12817 4573 12851 4607
rect 12851 4573 12860 4607
rect 12808 4564 12860 4573
rect 15292 4564 15344 4616
rect 17224 4632 17276 4684
rect 18236 4700 18288 4752
rect 17868 4632 17920 4684
rect 19800 4700 19852 4752
rect 20444 4700 20496 4752
rect 21640 4700 21692 4752
rect 13084 4496 13136 4548
rect 14832 4496 14884 4548
rect 5172 4428 5224 4480
rect 5264 4428 5316 4480
rect 12348 4428 12400 4480
rect 12900 4428 12952 4480
rect 13268 4471 13320 4480
rect 13268 4437 13277 4471
rect 13277 4437 13311 4471
rect 13311 4437 13320 4471
rect 13268 4428 13320 4437
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 14556 4428 14608 4480
rect 16396 4496 16448 4548
rect 18696 4564 18748 4616
rect 19984 4632 20036 4684
rect 20996 4632 21048 4684
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 21088 4564 21140 4616
rect 19616 4496 19668 4548
rect 20168 4496 20220 4548
rect 20996 4496 21048 4548
rect 16212 4428 16264 4480
rect 18420 4428 18472 4480
rect 18880 4471 18932 4480
rect 18880 4437 18889 4471
rect 18889 4437 18923 4471
rect 18923 4437 18932 4471
rect 18880 4428 18932 4437
rect 19984 4428 20036 4480
rect 20720 4471 20772 4480
rect 20720 4437 20729 4471
rect 20729 4437 20763 4471
rect 20763 4437 20772 4471
rect 20720 4428 20772 4437
rect 20812 4428 20864 4480
rect 1366 4326 1418 4378
rect 1430 4326 1482 4378
rect 1494 4326 1546 4378
rect 1558 4326 1610 4378
rect 1622 4326 1674 4378
rect 1686 4326 1738 4378
rect 7366 4326 7418 4378
rect 7430 4326 7482 4378
rect 7494 4326 7546 4378
rect 7558 4326 7610 4378
rect 7622 4326 7674 4378
rect 7686 4326 7738 4378
rect 13366 4326 13418 4378
rect 13430 4326 13482 4378
rect 13494 4326 13546 4378
rect 13558 4326 13610 4378
rect 13622 4326 13674 4378
rect 13686 4326 13738 4378
rect 19366 4326 19418 4378
rect 19430 4326 19482 4378
rect 19494 4326 19546 4378
rect 19558 4326 19610 4378
rect 19622 4326 19674 4378
rect 19686 4326 19738 4378
rect 2780 4224 2832 4276
rect 3792 4224 3844 4276
rect 7012 4224 7064 4276
rect 11612 4224 11664 4276
rect 1952 4020 2004 4072
rect 2780 4088 2832 4140
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 5908 4156 5960 4208
rect 13452 4156 13504 4208
rect 2228 4020 2280 4072
rect 2320 4063 2372 4072
rect 2320 4029 2329 4063
rect 2329 4029 2363 4063
rect 2363 4029 2372 4063
rect 2320 4020 2372 4029
rect 3608 4020 3660 4072
rect 4160 4020 4212 4072
rect 7932 4088 7984 4140
rect 1860 3927 1912 3936
rect 1860 3893 1875 3927
rect 1875 3893 1909 3927
rect 1909 3893 1912 3927
rect 1860 3884 1912 3893
rect 5172 4020 5224 4072
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 8852 4088 8904 4140
rect 9036 4088 9088 4140
rect 9312 4088 9364 4140
rect 9588 4088 9640 4140
rect 9864 4088 9916 4140
rect 12532 4088 12584 4140
rect 12440 4020 12492 4072
rect 9036 3952 9088 4004
rect 10876 3952 10928 4004
rect 5356 3884 5408 3936
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 8392 3884 8444 3936
rect 11428 3884 11480 3936
rect 12808 4020 12860 4072
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 14556 4224 14608 4276
rect 15108 4224 15160 4276
rect 15384 4156 15436 4208
rect 17684 4224 17736 4276
rect 18236 4224 18288 4276
rect 18512 4224 18564 4276
rect 20168 4224 20220 4276
rect 21364 4224 21416 4276
rect 22008 4267 22060 4276
rect 22008 4233 22017 4267
rect 22017 4233 22051 4267
rect 22051 4233 22060 4267
rect 22008 4224 22060 4233
rect 22100 4224 22152 4276
rect 13176 4020 13228 4072
rect 13268 4020 13320 4072
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 14188 4020 14240 4072
rect 15108 3952 15160 4004
rect 14464 3884 14516 3936
rect 14832 3927 14884 3936
rect 14832 3893 14841 3927
rect 14841 3893 14875 3927
rect 14875 3893 14884 3927
rect 14832 3884 14884 3893
rect 15384 4063 15436 4072
rect 15384 4029 15393 4063
rect 15393 4029 15427 4063
rect 15427 4029 15436 4063
rect 15384 4020 15436 4029
rect 15936 4088 15988 4140
rect 16028 4131 16080 4140
rect 16028 4097 16037 4131
rect 16037 4097 16071 4131
rect 16071 4097 16080 4131
rect 16028 4088 16080 4097
rect 16396 4088 16448 4140
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 16212 4020 16264 4072
rect 20076 4156 20128 4208
rect 19984 4020 20036 4072
rect 20352 4088 20404 4140
rect 20628 4156 20680 4208
rect 18604 3952 18656 4004
rect 19616 3952 19668 4004
rect 20444 4020 20496 4072
rect 20628 4063 20680 4072
rect 20628 4029 20637 4063
rect 20637 4029 20671 4063
rect 20671 4029 20680 4063
rect 20628 4020 20680 4029
rect 20720 4020 20772 4072
rect 20812 4063 20864 4072
rect 20812 4029 20821 4063
rect 20821 4029 20855 4063
rect 20855 4029 20864 4063
rect 20812 4020 20864 4029
rect 21548 4156 21600 4208
rect 16304 3884 16356 3936
rect 16764 3884 16816 3936
rect 21180 3884 21232 3936
rect 21456 4020 21508 4072
rect 21640 4020 21692 4072
rect 22284 4020 22336 4072
rect 22008 3952 22060 4004
rect 22192 3952 22244 4004
rect 22836 4020 22888 4072
rect 4366 3782 4418 3834
rect 4430 3782 4482 3834
rect 4494 3782 4546 3834
rect 4558 3782 4610 3834
rect 4622 3782 4674 3834
rect 4686 3782 4738 3834
rect 10366 3782 10418 3834
rect 10430 3782 10482 3834
rect 10494 3782 10546 3834
rect 10558 3782 10610 3834
rect 10622 3782 10674 3834
rect 10686 3782 10738 3834
rect 16366 3782 16418 3834
rect 16430 3782 16482 3834
rect 16494 3782 16546 3834
rect 16558 3782 16610 3834
rect 16622 3782 16674 3834
rect 16686 3782 16738 3834
rect 22366 3782 22418 3834
rect 22430 3782 22482 3834
rect 22494 3782 22546 3834
rect 22558 3782 22610 3834
rect 22622 3782 22674 3834
rect 22686 3782 22738 3834
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 4160 3680 4212 3732
rect 6920 3680 6972 3732
rect 3424 3612 3476 3664
rect 3792 3612 3844 3664
rect 848 3544 900 3596
rect 1216 3587 1268 3596
rect 1216 3553 1250 3587
rect 1250 3553 1268 3587
rect 1216 3544 1268 3553
rect 4988 3587 5040 3596
rect 4988 3553 4997 3587
rect 4997 3553 5031 3587
rect 5031 3553 5040 3587
rect 4988 3544 5040 3553
rect 6092 3544 6144 3596
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 5080 3451 5132 3460
rect 5080 3417 5089 3451
rect 5089 3417 5123 3451
rect 5123 3417 5132 3451
rect 5080 3408 5132 3417
rect 6644 3408 6696 3460
rect 8484 3680 8536 3732
rect 8024 3612 8076 3664
rect 8852 3680 8904 3732
rect 9496 3680 9548 3732
rect 10048 3723 10100 3732
rect 10048 3689 10057 3723
rect 10057 3689 10091 3723
rect 10091 3689 10100 3723
rect 10048 3680 10100 3689
rect 10600 3680 10652 3732
rect 7288 3408 7340 3460
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 8116 3408 8168 3460
rect 8300 3408 8352 3460
rect 8668 3519 8720 3528
rect 8668 3485 8677 3519
rect 8677 3485 8711 3519
rect 8711 3485 8720 3519
rect 8668 3476 8720 3485
rect 9036 3476 9088 3528
rect 10416 3612 10468 3664
rect 11796 3680 11848 3732
rect 11428 3612 11480 3664
rect 12900 3680 12952 3732
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 10876 3544 10928 3596
rect 13452 3612 13504 3664
rect 12348 3544 12400 3596
rect 13176 3544 13228 3596
rect 14188 3612 14240 3664
rect 13636 3587 13688 3596
rect 13636 3553 13661 3587
rect 13661 3553 13688 3587
rect 13636 3544 13688 3553
rect 13912 3587 13964 3596
rect 13912 3553 13921 3587
rect 13921 3553 13955 3587
rect 13955 3553 13964 3587
rect 13912 3544 13964 3553
rect 9128 3408 9180 3460
rect 7012 3340 7064 3392
rect 7932 3340 7984 3392
rect 9772 3408 9824 3460
rect 10508 3476 10560 3528
rect 11060 3408 11112 3460
rect 13820 3476 13872 3528
rect 14924 3680 14976 3732
rect 15384 3680 15436 3732
rect 14464 3544 14516 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 15200 3476 15252 3528
rect 15752 3544 15804 3596
rect 16028 3544 16080 3596
rect 16764 3612 16816 3664
rect 16396 3544 16448 3596
rect 17224 3544 17276 3596
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 19892 3680 19944 3732
rect 20812 3680 20864 3732
rect 21180 3680 21232 3732
rect 22836 3680 22888 3732
rect 17960 3544 18012 3596
rect 20904 3612 20956 3664
rect 9496 3340 9548 3392
rect 10600 3340 10652 3392
rect 11796 3383 11848 3392
rect 11796 3349 11805 3383
rect 11805 3349 11839 3383
rect 11839 3349 11848 3383
rect 11796 3340 11848 3349
rect 12808 3340 12860 3392
rect 13084 3340 13136 3392
rect 14464 3340 14516 3392
rect 15476 3408 15528 3460
rect 16856 3408 16908 3460
rect 18328 3408 18380 3460
rect 15568 3340 15620 3392
rect 15752 3383 15804 3392
rect 15752 3349 15761 3383
rect 15761 3349 15795 3383
rect 15795 3349 15804 3383
rect 15752 3340 15804 3349
rect 16212 3383 16264 3392
rect 16212 3349 16221 3383
rect 16221 3349 16255 3383
rect 16255 3349 16264 3383
rect 16212 3340 16264 3349
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 18512 3340 18564 3392
rect 19616 3587 19668 3596
rect 19616 3553 19625 3587
rect 19625 3553 19659 3587
rect 19659 3553 19668 3587
rect 19616 3544 19668 3553
rect 19800 3587 19852 3596
rect 19800 3553 19809 3587
rect 19809 3553 19843 3587
rect 19843 3553 19852 3587
rect 19800 3544 19852 3553
rect 18696 3408 18748 3460
rect 19984 3476 20036 3528
rect 20812 3544 20864 3596
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 19064 3340 19116 3392
rect 19892 3340 19944 3392
rect 20076 3383 20128 3392
rect 20076 3349 20085 3383
rect 20085 3349 20119 3383
rect 20119 3349 20128 3383
rect 20076 3340 20128 3349
rect 1366 3238 1418 3290
rect 1430 3238 1482 3290
rect 1494 3238 1546 3290
rect 1558 3238 1610 3290
rect 1622 3238 1674 3290
rect 1686 3238 1738 3290
rect 7366 3238 7418 3290
rect 7430 3238 7482 3290
rect 7494 3238 7546 3290
rect 7558 3238 7610 3290
rect 7622 3238 7674 3290
rect 7686 3238 7738 3290
rect 13366 3238 13418 3290
rect 13430 3238 13482 3290
rect 13494 3238 13546 3290
rect 13558 3238 13610 3290
rect 13622 3238 13674 3290
rect 13686 3238 13738 3290
rect 19366 3238 19418 3290
rect 19430 3238 19482 3290
rect 19494 3238 19546 3290
rect 19558 3238 19610 3290
rect 19622 3238 19674 3290
rect 19686 3238 19738 3290
rect 1216 3136 1268 3188
rect 3884 3136 3936 3188
rect 3056 3068 3108 3120
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 2320 2975 2372 2984
rect 2320 2941 2329 2975
rect 2329 2941 2363 2975
rect 2363 2941 2372 2975
rect 2320 2932 2372 2941
rect 2504 2975 2556 2984
rect 2504 2941 2513 2975
rect 2513 2941 2547 2975
rect 2547 2941 2556 2975
rect 2504 2932 2556 2941
rect 3056 2932 3108 2984
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 3608 2975 3660 2984
rect 3608 2941 3617 2975
rect 3617 2941 3651 2975
rect 3651 2941 3660 2975
rect 3608 2932 3660 2941
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 6644 3136 6696 3188
rect 7012 3136 7064 3188
rect 9036 3068 9088 3120
rect 12992 3136 13044 3188
rect 14004 3136 14056 3188
rect 14740 3136 14792 3188
rect 15752 3136 15804 3188
rect 16212 3136 16264 3188
rect 16304 3136 16356 3188
rect 17316 3136 17368 3188
rect 18880 3136 18932 3188
rect 20904 3136 20956 3188
rect 21732 3136 21784 3188
rect 6828 3000 6880 3052
rect 8576 3000 8628 3052
rect 9128 3000 9180 3052
rect 7932 2932 7984 2984
rect 7840 2907 7892 2916
rect 7840 2873 7849 2907
rect 7849 2873 7883 2907
rect 7883 2873 7892 2907
rect 7840 2864 7892 2873
rect 9496 3068 9548 3120
rect 9772 3068 9824 3120
rect 10508 3068 10560 3120
rect 13636 3043 13688 3052
rect 13636 3009 13645 3043
rect 13645 3009 13679 3043
rect 13679 3009 13688 3043
rect 13636 3000 13688 3009
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 14832 3000 14884 3052
rect 9680 2932 9732 2984
rect 9772 2932 9824 2984
rect 10048 2932 10100 2984
rect 10232 2932 10284 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 13820 2975 13872 2984
rect 5172 2796 5224 2848
rect 8668 2796 8720 2848
rect 9036 2796 9088 2848
rect 10600 2864 10652 2916
rect 13820 2941 13829 2975
rect 13829 2941 13863 2975
rect 13863 2941 13872 2975
rect 13820 2932 13872 2941
rect 14004 2932 14056 2984
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 11060 2796 11112 2848
rect 11796 2796 11848 2848
rect 12348 2796 12400 2848
rect 13084 2796 13136 2848
rect 14832 2907 14884 2916
rect 14832 2873 14841 2907
rect 14841 2873 14875 2907
rect 14875 2873 14884 2907
rect 14832 2864 14884 2873
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 15568 2975 15620 2984
rect 15568 2941 15577 2975
rect 15577 2941 15611 2975
rect 15611 2941 15620 2975
rect 15568 2932 15620 2941
rect 16028 3000 16080 3052
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 16580 2975 16632 2984
rect 16580 2941 16589 2975
rect 16589 2941 16623 2975
rect 16623 2941 16632 2975
rect 16580 2932 16632 2941
rect 18512 3068 18564 3120
rect 19432 3068 19484 3120
rect 18328 3000 18380 3052
rect 16764 2864 16816 2916
rect 13544 2796 13596 2848
rect 14096 2839 14148 2848
rect 14096 2805 14105 2839
rect 14105 2805 14139 2839
rect 14139 2805 14148 2839
rect 14096 2796 14148 2805
rect 15568 2796 15620 2848
rect 15936 2839 15988 2848
rect 15936 2805 15945 2839
rect 15945 2805 15979 2839
rect 15979 2805 15988 2839
rect 15936 2796 15988 2805
rect 16212 2796 16264 2848
rect 17040 2932 17092 2984
rect 18788 2975 18840 2984
rect 18788 2941 18797 2975
rect 18797 2941 18831 2975
rect 18831 2941 18840 2975
rect 18788 2932 18840 2941
rect 18696 2796 18748 2848
rect 19064 2932 19116 2984
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 20076 2864 20128 2916
rect 20260 2864 20312 2916
rect 21272 2839 21324 2848
rect 21272 2805 21281 2839
rect 21281 2805 21315 2839
rect 21315 2805 21324 2839
rect 21272 2796 21324 2805
rect 4366 2694 4418 2746
rect 4430 2694 4482 2746
rect 4494 2694 4546 2746
rect 4558 2694 4610 2746
rect 4622 2694 4674 2746
rect 4686 2694 4738 2746
rect 10366 2694 10418 2746
rect 10430 2694 10482 2746
rect 10494 2694 10546 2746
rect 10558 2694 10610 2746
rect 10622 2694 10674 2746
rect 10686 2694 10738 2746
rect 16366 2694 16418 2746
rect 16430 2694 16482 2746
rect 16494 2694 16546 2746
rect 16558 2694 16610 2746
rect 16622 2694 16674 2746
rect 16686 2694 16738 2746
rect 22366 2694 22418 2746
rect 22430 2694 22482 2746
rect 22494 2694 22546 2746
rect 22558 2694 22610 2746
rect 22622 2694 22674 2746
rect 22686 2694 22738 2746
rect 2504 2635 2556 2644
rect 2504 2601 2513 2635
rect 2513 2601 2547 2635
rect 2547 2601 2556 2635
rect 2504 2592 2556 2601
rect 1768 2524 1820 2576
rect 1216 2456 1268 2508
rect 4068 2592 4120 2644
rect 8944 2592 8996 2644
rect 3608 2524 3660 2576
rect 5172 2456 5224 2508
rect 3884 2388 3936 2440
rect 7288 2388 7340 2440
rect 9036 2320 9088 2372
rect 3700 2252 3752 2304
rect 3792 2295 3844 2304
rect 3792 2261 3801 2295
rect 3801 2261 3835 2295
rect 3835 2261 3844 2295
rect 3792 2252 3844 2261
rect 7288 2252 7340 2304
rect 8760 2252 8812 2304
rect 9220 2524 9272 2576
rect 9956 2592 10008 2644
rect 10232 2592 10284 2644
rect 10784 2592 10836 2644
rect 9864 2524 9916 2576
rect 10048 2524 10100 2576
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 11060 2524 11112 2576
rect 9496 2388 9548 2440
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 9772 2320 9824 2372
rect 11704 2592 11756 2644
rect 12808 2592 12860 2644
rect 12900 2592 12952 2644
rect 13820 2592 13872 2644
rect 14280 2592 14332 2644
rect 15200 2592 15252 2644
rect 13176 2524 13228 2576
rect 13544 2567 13596 2576
rect 13544 2533 13553 2567
rect 13553 2533 13587 2567
rect 13587 2533 13596 2567
rect 13544 2524 13596 2533
rect 15660 2524 15712 2576
rect 10784 2320 10836 2372
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 11152 2252 11204 2304
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 12808 2320 12860 2372
rect 13820 2363 13872 2372
rect 13820 2329 13829 2363
rect 13829 2329 13863 2363
rect 13863 2329 13872 2363
rect 13820 2320 13872 2329
rect 16212 2456 16264 2508
rect 16856 2524 16908 2576
rect 16672 2456 16724 2508
rect 14556 2388 14608 2440
rect 15476 2388 15528 2440
rect 17868 2524 17920 2576
rect 17040 2456 17092 2508
rect 13084 2252 13136 2304
rect 13268 2252 13320 2304
rect 15016 2252 15068 2304
rect 15752 2252 15804 2304
rect 18236 2499 18288 2508
rect 18236 2465 18245 2499
rect 18245 2465 18279 2499
rect 18279 2465 18288 2499
rect 18236 2456 18288 2465
rect 18328 2456 18380 2508
rect 20260 2592 20312 2644
rect 20812 2592 20864 2644
rect 19340 2499 19392 2508
rect 19340 2465 19349 2499
rect 19349 2465 19383 2499
rect 19383 2465 19392 2499
rect 19340 2456 19392 2465
rect 19708 2499 19760 2508
rect 19708 2465 19717 2499
rect 19717 2465 19751 2499
rect 19751 2465 19760 2499
rect 19708 2456 19760 2465
rect 21272 2524 21324 2576
rect 21364 2456 21416 2508
rect 19248 2431 19300 2440
rect 19248 2397 19257 2431
rect 19257 2397 19291 2431
rect 19291 2397 19300 2431
rect 19248 2388 19300 2397
rect 20628 2388 20680 2440
rect 17040 2252 17092 2304
rect 18420 2252 18472 2304
rect 19892 2295 19944 2304
rect 19892 2261 19901 2295
rect 19901 2261 19935 2295
rect 19935 2261 19944 2295
rect 19892 2252 19944 2261
rect 1366 2150 1418 2202
rect 1430 2150 1482 2202
rect 1494 2150 1546 2202
rect 1558 2150 1610 2202
rect 1622 2150 1674 2202
rect 1686 2150 1738 2202
rect 7366 2150 7418 2202
rect 7430 2150 7482 2202
rect 7494 2150 7546 2202
rect 7558 2150 7610 2202
rect 7622 2150 7674 2202
rect 7686 2150 7738 2202
rect 13366 2150 13418 2202
rect 13430 2150 13482 2202
rect 13494 2150 13546 2202
rect 13558 2150 13610 2202
rect 13622 2150 13674 2202
rect 13686 2150 13738 2202
rect 19366 2150 19418 2202
rect 19430 2150 19482 2202
rect 19494 2150 19546 2202
rect 19558 2150 19610 2202
rect 19622 2150 19674 2202
rect 19686 2150 19738 2202
rect 3884 2048 3936 2100
rect 4160 2048 4212 2100
rect 1032 1980 1084 2032
rect 3516 1912 3568 1964
rect 2412 1844 2464 1896
rect 4344 1819 4396 1828
rect 4344 1785 4353 1819
rect 4353 1785 4387 1819
rect 4387 1785 4396 1819
rect 4344 1776 4396 1785
rect 4988 1887 5040 1896
rect 4988 1853 4997 1887
rect 4997 1853 5031 1887
rect 5031 1853 5040 1887
rect 4988 1844 5040 1853
rect 5724 1819 5776 1828
rect 5724 1785 5733 1819
rect 5733 1785 5767 1819
rect 5767 1785 5776 1819
rect 5724 1776 5776 1785
rect 7012 1844 7064 1896
rect 8668 2048 8720 2100
rect 9128 2048 9180 2100
rect 10048 2048 10100 2100
rect 11152 2048 11204 2100
rect 7564 1887 7616 1896
rect 7564 1853 7573 1887
rect 7573 1853 7607 1887
rect 7607 1853 7616 1887
rect 7564 1844 7616 1853
rect 7748 1887 7800 1896
rect 7748 1853 7757 1887
rect 7757 1853 7791 1887
rect 7791 1853 7800 1887
rect 7748 1844 7800 1853
rect 7840 1776 7892 1828
rect 8300 1844 8352 1896
rect 18696 2048 18748 2100
rect 18880 2091 18932 2100
rect 18880 2057 18889 2091
rect 18889 2057 18923 2091
rect 18923 2057 18932 2091
rect 18880 2048 18932 2057
rect 21732 2091 21784 2100
rect 21732 2057 21741 2091
rect 21741 2057 21775 2091
rect 21775 2057 21784 2091
rect 21732 2048 21784 2057
rect 9864 1912 9916 1964
rect 10232 1912 10284 1964
rect 10324 1912 10376 1964
rect 11060 1912 11112 1964
rect 8392 1776 8444 1828
rect 10784 1844 10836 1896
rect 11152 1887 11204 1896
rect 11152 1853 11161 1887
rect 11161 1853 11195 1887
rect 11195 1853 11204 1887
rect 11152 1844 11204 1853
rect 11244 1887 11296 1896
rect 11244 1853 11253 1887
rect 11253 1853 11287 1887
rect 11287 1853 11296 1887
rect 11244 1844 11296 1853
rect 11336 1887 11388 1896
rect 11336 1853 11345 1887
rect 11345 1853 11379 1887
rect 11379 1853 11388 1887
rect 11336 1844 11388 1853
rect 11520 1887 11572 1896
rect 11520 1853 11529 1887
rect 11529 1853 11563 1887
rect 11563 1853 11572 1887
rect 11520 1844 11572 1853
rect 12992 1912 13044 1964
rect 13820 1912 13872 1964
rect 15016 1912 15068 1964
rect 15476 1912 15528 1964
rect 1124 1708 1176 1760
rect 4252 1708 4304 1760
rect 6920 1708 6972 1760
rect 7656 1708 7708 1760
rect 7748 1708 7800 1760
rect 8116 1708 8168 1760
rect 8760 1708 8812 1760
rect 11612 1776 11664 1828
rect 13084 1844 13136 1896
rect 16120 1912 16172 1964
rect 17040 1912 17092 1964
rect 15844 1887 15896 1896
rect 15844 1853 15853 1887
rect 15853 1853 15887 1887
rect 15887 1853 15896 1887
rect 15844 1844 15896 1853
rect 15936 1844 15988 1896
rect 13268 1819 13320 1828
rect 13268 1785 13277 1819
rect 13277 1785 13311 1819
rect 13311 1785 13320 1819
rect 13268 1776 13320 1785
rect 14004 1776 14056 1828
rect 14556 1819 14608 1828
rect 14556 1785 14565 1819
rect 14565 1785 14599 1819
rect 14599 1785 14608 1819
rect 14556 1776 14608 1785
rect 15292 1776 15344 1828
rect 16764 1844 16816 1896
rect 10324 1708 10376 1760
rect 11060 1708 11112 1760
rect 13452 1708 13504 1760
rect 14648 1751 14700 1760
rect 14648 1717 14657 1751
rect 14657 1717 14691 1751
rect 14691 1717 14700 1751
rect 14648 1708 14700 1717
rect 15016 1708 15068 1760
rect 15200 1708 15252 1760
rect 15384 1751 15436 1760
rect 15384 1717 15393 1751
rect 15393 1717 15427 1751
rect 15427 1717 15436 1751
rect 15384 1708 15436 1717
rect 15476 1708 15528 1760
rect 17868 1887 17920 1896
rect 17868 1853 17877 1887
rect 17877 1853 17911 1887
rect 17911 1853 17920 1887
rect 17868 1844 17920 1853
rect 22192 1980 22244 2032
rect 18052 1708 18104 1760
rect 22100 1912 22152 1964
rect 21916 1887 21968 1896
rect 21916 1853 21925 1887
rect 21925 1853 21959 1887
rect 21959 1853 21968 1887
rect 21916 1844 21968 1853
rect 19340 1708 19392 1760
rect 21088 1751 21140 1760
rect 21088 1717 21097 1751
rect 21097 1717 21131 1751
rect 21131 1717 21140 1751
rect 21088 1708 21140 1717
rect 4366 1606 4418 1658
rect 4430 1606 4482 1658
rect 4494 1606 4546 1658
rect 4558 1606 4610 1658
rect 4622 1606 4674 1658
rect 4686 1606 4738 1658
rect 10366 1606 10418 1658
rect 10430 1606 10482 1658
rect 10494 1606 10546 1658
rect 10558 1606 10610 1658
rect 10622 1606 10674 1658
rect 10686 1606 10738 1658
rect 16366 1606 16418 1658
rect 16430 1606 16482 1658
rect 16494 1606 16546 1658
rect 16558 1606 16610 1658
rect 16622 1606 16674 1658
rect 16686 1606 16738 1658
rect 22366 1606 22418 1658
rect 22430 1606 22482 1658
rect 22494 1606 22546 1658
rect 22558 1606 22610 1658
rect 22622 1606 22674 1658
rect 22686 1606 22738 1658
rect 1124 1504 1176 1556
rect 1216 1504 1268 1556
rect 3700 1504 3752 1556
rect 3792 1504 3844 1556
rect 3884 1504 3936 1556
rect 4160 1504 4212 1556
rect 6920 1504 6972 1556
rect 5724 1436 5776 1488
rect 1768 1275 1820 1284
rect 1768 1241 1777 1275
rect 1777 1241 1811 1275
rect 1811 1241 1820 1275
rect 1768 1232 1820 1241
rect 5448 1368 5500 1420
rect 4160 1300 4212 1352
rect 4252 1343 4304 1352
rect 4252 1309 4261 1343
rect 4261 1309 4295 1343
rect 4295 1309 4304 1343
rect 4252 1300 4304 1309
rect 6920 1411 6972 1420
rect 6920 1377 6929 1411
rect 6929 1377 6963 1411
rect 6963 1377 6972 1411
rect 6920 1368 6972 1377
rect 7012 1368 7064 1420
rect 7288 1436 7340 1488
rect 7840 1504 7892 1556
rect 9036 1547 9088 1556
rect 9036 1513 9045 1547
rect 9045 1513 9079 1547
rect 9079 1513 9088 1547
rect 9036 1504 9088 1513
rect 9864 1504 9916 1556
rect 10876 1504 10928 1556
rect 11152 1504 11204 1556
rect 8392 1368 8444 1420
rect 8576 1411 8628 1420
rect 8576 1377 8585 1411
rect 8585 1377 8619 1411
rect 8619 1377 8628 1411
rect 8576 1368 8628 1377
rect 9404 1411 9456 1420
rect 9404 1377 9413 1411
rect 9413 1377 9447 1411
rect 9447 1377 9456 1411
rect 9404 1368 9456 1377
rect 9496 1411 9548 1420
rect 9496 1377 9505 1411
rect 9505 1377 9539 1411
rect 9539 1377 9548 1411
rect 9496 1368 9548 1377
rect 10140 1411 10192 1420
rect 10140 1377 10149 1411
rect 10149 1377 10183 1411
rect 10183 1377 10192 1411
rect 10140 1368 10192 1377
rect 7564 1300 7616 1352
rect 7656 1300 7708 1352
rect 9772 1300 9824 1352
rect 10508 1300 10560 1352
rect 10968 1368 11020 1420
rect 13268 1504 13320 1556
rect 13544 1504 13596 1556
rect 15476 1504 15528 1556
rect 15660 1504 15712 1556
rect 11428 1411 11480 1420
rect 11428 1377 11437 1411
rect 11437 1377 11471 1411
rect 11471 1377 11480 1411
rect 11428 1368 11480 1377
rect 11612 1368 11664 1420
rect 12256 1411 12308 1420
rect 12256 1377 12265 1411
rect 12265 1377 12299 1411
rect 12299 1377 12308 1411
rect 12256 1368 12308 1377
rect 14004 1436 14056 1488
rect 13820 1368 13872 1420
rect 14096 1368 14148 1420
rect 14740 1411 14792 1420
rect 14740 1377 14749 1411
rect 14749 1377 14783 1411
rect 14783 1377 14792 1411
rect 14740 1368 14792 1377
rect 14924 1411 14976 1420
rect 14924 1377 14933 1411
rect 14933 1377 14967 1411
rect 14967 1377 14976 1411
rect 14924 1368 14976 1377
rect 15200 1411 15252 1420
rect 15200 1377 15209 1411
rect 15209 1377 15243 1411
rect 15243 1377 15252 1411
rect 15200 1368 15252 1377
rect 15568 1411 15620 1420
rect 15568 1377 15577 1411
rect 15577 1377 15611 1411
rect 15611 1377 15620 1411
rect 15568 1368 15620 1377
rect 15752 1411 15804 1420
rect 15752 1377 15761 1411
rect 15761 1377 15795 1411
rect 15795 1377 15804 1411
rect 15752 1368 15804 1377
rect 15936 1368 15988 1420
rect 16212 1411 16264 1420
rect 16212 1377 16221 1411
rect 16221 1377 16255 1411
rect 16255 1377 16264 1411
rect 16212 1368 16264 1377
rect 16396 1411 16448 1420
rect 16396 1377 16405 1411
rect 16405 1377 16439 1411
rect 16439 1377 16448 1411
rect 16396 1368 16448 1377
rect 16764 1411 16816 1420
rect 16764 1377 16773 1411
rect 16773 1377 16807 1411
rect 16807 1377 16816 1411
rect 16764 1368 16816 1377
rect 17132 1504 17184 1556
rect 17224 1411 17276 1420
rect 17224 1377 17233 1411
rect 17233 1377 17267 1411
rect 17267 1377 17276 1411
rect 17224 1368 17276 1377
rect 17408 1368 17460 1420
rect 17684 1368 17736 1420
rect 19892 1504 19944 1556
rect 22376 1504 22428 1556
rect 18052 1479 18104 1488
rect 18052 1445 18061 1479
rect 18061 1445 18095 1479
rect 18095 1445 18104 1479
rect 18052 1436 18104 1445
rect 19340 1368 19392 1420
rect 19800 1368 19852 1420
rect 22100 1479 22152 1488
rect 22100 1445 22109 1479
rect 22109 1445 22143 1479
rect 22143 1445 22152 1479
rect 22100 1436 22152 1445
rect 8208 1232 8260 1284
rect 11336 1232 11388 1284
rect 12716 1300 12768 1352
rect 13452 1343 13504 1352
rect 13452 1309 13461 1343
rect 13461 1309 13495 1343
rect 13495 1309 13504 1343
rect 13452 1300 13504 1309
rect 16120 1343 16172 1352
rect 16120 1309 16129 1343
rect 16129 1309 16163 1343
rect 16163 1309 16172 1343
rect 16120 1300 16172 1309
rect 15752 1232 15804 1284
rect 18696 1300 18748 1352
rect 18880 1343 18932 1352
rect 18880 1309 18889 1343
rect 18889 1309 18923 1343
rect 18923 1309 18932 1343
rect 18880 1300 18932 1309
rect 19064 1232 19116 1284
rect 20 1164 72 1216
rect 8300 1164 8352 1216
rect 8392 1207 8444 1216
rect 8392 1173 8401 1207
rect 8401 1173 8435 1207
rect 8435 1173 8444 1207
rect 8392 1164 8444 1173
rect 8760 1207 8812 1216
rect 8760 1173 8769 1207
rect 8769 1173 8803 1207
rect 8803 1173 8812 1207
rect 8760 1164 8812 1173
rect 9772 1207 9824 1216
rect 9772 1173 9781 1207
rect 9781 1173 9815 1207
rect 9815 1173 9824 1207
rect 9772 1164 9824 1173
rect 10784 1207 10836 1216
rect 10784 1173 10793 1207
rect 10793 1173 10827 1207
rect 10827 1173 10836 1207
rect 10784 1164 10836 1173
rect 11612 1164 11664 1216
rect 12624 1207 12676 1216
rect 12624 1173 12633 1207
rect 12633 1173 12667 1207
rect 12667 1173 12676 1207
rect 12624 1164 12676 1173
rect 12992 1207 13044 1216
rect 12992 1173 13001 1207
rect 13001 1173 13035 1207
rect 13035 1173 13044 1207
rect 12992 1164 13044 1173
rect 13452 1164 13504 1216
rect 13820 1164 13872 1216
rect 14372 1207 14424 1216
rect 14372 1173 14381 1207
rect 14381 1173 14415 1207
rect 14415 1173 14424 1207
rect 14372 1164 14424 1173
rect 15108 1207 15160 1216
rect 15108 1173 15117 1207
rect 15117 1173 15151 1207
rect 15151 1173 15160 1207
rect 15108 1164 15160 1173
rect 15936 1207 15988 1216
rect 15936 1173 15945 1207
rect 15945 1173 15979 1207
rect 15979 1173 15988 1207
rect 15936 1164 15988 1173
rect 16580 1207 16632 1216
rect 16580 1173 16589 1207
rect 16589 1173 16623 1207
rect 16623 1173 16632 1207
rect 16580 1164 16632 1173
rect 17408 1207 17460 1216
rect 17408 1173 17417 1207
rect 17417 1173 17451 1207
rect 17451 1173 17460 1207
rect 17408 1164 17460 1173
rect 17960 1207 18012 1216
rect 17960 1173 17969 1207
rect 17969 1173 18003 1207
rect 18003 1173 18012 1207
rect 17960 1164 18012 1173
rect 21364 1368 21416 1420
rect 21456 1368 21508 1420
rect 21916 1300 21968 1352
rect 21640 1232 21692 1284
rect 1366 1062 1418 1114
rect 1430 1062 1482 1114
rect 1494 1062 1546 1114
rect 1558 1062 1610 1114
rect 1622 1062 1674 1114
rect 1686 1062 1738 1114
rect 7366 1062 7418 1114
rect 7430 1062 7482 1114
rect 7494 1062 7546 1114
rect 7558 1062 7610 1114
rect 7622 1062 7674 1114
rect 7686 1062 7738 1114
rect 13366 1062 13418 1114
rect 13430 1062 13482 1114
rect 13494 1062 13546 1114
rect 13558 1062 13610 1114
rect 13622 1062 13674 1114
rect 13686 1062 13738 1114
rect 19366 1062 19418 1114
rect 19430 1062 19482 1114
rect 19494 1062 19546 1114
rect 19558 1062 19610 1114
rect 19622 1062 19674 1114
rect 19686 1062 19738 1114
rect 1216 960 1268 1012
rect 4160 960 4212 1012
rect 1032 756 1084 808
rect 8208 892 8260 944
rect 8392 892 8444 944
rect 1860 688 1912 740
rect 2504 688 2556 740
rect 6184 799 6236 808
rect 6184 765 6193 799
rect 6193 765 6227 799
rect 6227 765 6236 799
rect 6184 756 6236 765
rect 8852 799 8904 808
rect 8852 765 8861 799
rect 8861 765 8895 799
rect 8895 765 8904 799
rect 8852 756 8904 765
rect 9772 960 9824 1012
rect 10784 960 10836 1012
rect 12072 960 12124 1012
rect 12624 960 12676 1012
rect 12992 960 13044 1012
rect 14372 960 14424 1012
rect 15016 960 15068 1012
rect 15752 960 15804 1012
rect 15936 960 15988 1012
rect 16028 960 16080 1012
rect 17592 960 17644 1012
rect 19800 960 19852 1012
rect 9772 799 9824 808
rect 9772 765 9781 799
rect 9781 765 9815 799
rect 9815 765 9824 799
rect 9772 756 9824 765
rect 11612 867 11664 876
rect 11612 833 11621 867
rect 11621 833 11655 867
rect 11655 833 11664 867
rect 11612 824 11664 833
rect 11520 756 11572 808
rect 13820 756 13872 808
rect 15108 756 15160 808
rect 15844 756 15896 808
rect 16120 799 16172 808
rect 16120 765 16129 799
rect 16129 765 16163 799
rect 16163 765 16172 799
rect 16120 756 16172 765
rect 16580 756 16632 808
rect 17960 824 18012 876
rect 18696 867 18748 876
rect 18696 833 18705 867
rect 18705 833 18739 867
rect 18739 833 18748 867
rect 18696 824 18748 833
rect 19064 824 19116 876
rect 17408 756 17460 808
rect 18972 799 19024 808
rect 18972 765 18981 799
rect 18981 765 19015 799
rect 19015 765 19024 799
rect 18972 756 19024 765
rect 1032 663 1084 672
rect 1032 629 1041 663
rect 1041 629 1075 663
rect 1075 629 1084 663
rect 1032 620 1084 629
rect 3332 663 3384 672
rect 3332 629 3341 663
rect 3341 629 3375 663
rect 3375 629 3384 663
rect 3332 620 3384 629
rect 4068 620 4120 672
rect 4344 663 4396 672
rect 4344 629 4353 663
rect 4353 629 4387 663
rect 4387 629 4396 663
rect 4344 620 4396 629
rect 5172 663 5224 672
rect 5172 629 5181 663
rect 5181 629 5215 663
rect 5215 629 5224 663
rect 5172 620 5224 629
rect 6000 663 6052 672
rect 6000 629 6009 663
rect 6009 629 6043 663
rect 6043 629 6052 663
rect 6000 620 6052 629
rect 8484 663 8536 672
rect 8484 629 8493 663
rect 8493 629 8527 663
rect 8527 629 8536 663
rect 8484 620 8536 629
rect 9128 620 9180 672
rect 22100 867 22152 876
rect 22100 833 22109 867
rect 22109 833 22143 867
rect 22143 833 22152 867
rect 22100 824 22152 833
rect 22192 799 22244 808
rect 22192 765 22201 799
rect 22201 765 22235 799
rect 22235 765 22244 799
rect 22192 756 22244 765
rect 9956 620 10008 672
rect 11152 663 11204 672
rect 11152 629 11161 663
rect 11161 629 11195 663
rect 11195 629 11204 663
rect 11152 620 11204 629
rect 11612 620 11664 672
rect 12624 663 12676 672
rect 12624 629 12633 663
rect 12633 629 12667 663
rect 12667 629 12676 663
rect 12624 620 12676 629
rect 13268 620 13320 672
rect 14280 663 14332 672
rect 14280 629 14289 663
rect 14289 629 14323 663
rect 14323 629 14332 663
rect 14280 620 14332 629
rect 16764 620 16816 672
rect 16856 663 16908 672
rect 16856 629 16865 663
rect 16865 629 16899 663
rect 16899 629 16908 663
rect 16856 620 16908 629
rect 17408 620 17460 672
rect 18420 663 18472 672
rect 18420 629 18429 663
rect 18429 629 18463 663
rect 18463 629 18472 663
rect 18420 620 18472 629
rect 19064 620 19116 672
rect 19892 620 19944 672
rect 20720 620 20772 672
rect 21548 620 21600 672
rect 4366 518 4418 570
rect 4430 518 4482 570
rect 4494 518 4546 570
rect 4558 518 4610 570
rect 4622 518 4674 570
rect 4686 518 4738 570
rect 10366 518 10418 570
rect 10430 518 10482 570
rect 10494 518 10546 570
rect 10558 518 10610 570
rect 10622 518 10674 570
rect 10686 518 10738 570
rect 16366 518 16418 570
rect 16430 518 16482 570
rect 16494 518 16546 570
rect 16558 518 16610 570
rect 16622 518 16674 570
rect 16686 518 16738 570
rect 22366 518 22418 570
rect 22430 518 22482 570
rect 22494 518 22546 570
rect 22558 518 22610 570
rect 22622 518 22674 570
rect 22686 518 22738 570
rect 5448 348 5500 400
rect 6184 280 6236 332
rect 15384 280 15436 332
rect 16764 348 16816 400
rect 21640 416 21692 468
rect 18144 280 18196 332
rect 4068 212 4120 264
rect 10232 212 10284 264
rect 9496 144 9548 196
rect 12716 212 12768 264
<< metal2 >>
rect 4434 15722 4490 16000
rect 4434 15694 4660 15722
rect 4434 15600 4490 15694
rect 1364 15260 1740 15269
rect 1420 15258 1444 15260
rect 1500 15258 1524 15260
rect 1580 15258 1604 15260
rect 1660 15258 1684 15260
rect 1420 15206 1430 15258
rect 1674 15206 1684 15258
rect 1420 15204 1444 15206
rect 1500 15204 1524 15206
rect 1580 15204 1604 15206
rect 1660 15204 1684 15206
rect 1364 15195 1740 15204
rect 4632 15162 4660 15694
rect 5170 15600 5226 16000
rect 5906 15722 5962 16000
rect 5906 15694 6224 15722
rect 5906 15600 5962 15694
rect 5184 15162 5212 15600
rect 6196 15162 6224 15694
rect 6642 15600 6698 16000
rect 7378 15722 7434 16000
rect 7300 15694 7434 15722
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 2240 14618 2268 14894
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 1032 14272 1084 14278
rect 1032 14214 1084 14220
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1044 13394 1072 14214
rect 1364 14172 1740 14181
rect 1420 14170 1444 14172
rect 1500 14170 1524 14172
rect 1580 14170 1604 14172
rect 1660 14170 1684 14172
rect 1420 14118 1430 14170
rect 1674 14118 1684 14170
rect 1420 14116 1444 14118
rect 1500 14116 1524 14118
rect 1580 14116 1604 14118
rect 1660 14116 1684 14118
rect 1364 14107 1740 14116
rect 1872 14074 1900 14214
rect 2424 14074 2452 14554
rect 2516 14482 2544 14758
rect 4364 14716 4740 14725
rect 4420 14714 4444 14716
rect 4500 14714 4524 14716
rect 4580 14714 4604 14716
rect 4660 14714 4684 14716
rect 4420 14662 4430 14714
rect 4674 14662 4684 14714
rect 4420 14660 4444 14662
rect 4500 14660 4524 14662
rect 4580 14660 4604 14662
rect 4660 14660 4684 14662
rect 4364 14651 4740 14660
rect 4908 14618 4936 14894
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 5184 14464 5212 14758
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 5356 14476 5408 14482
rect 5184 14436 5356 14464
rect 2884 14074 2912 14418
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 1216 13864 1268 13870
rect 1216 13806 1268 13812
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 1124 13456 1176 13462
rect 1124 13398 1176 13404
rect 1032 13388 1084 13394
rect 1032 13330 1084 13336
rect 1044 11218 1072 13330
rect 1136 12714 1164 13398
rect 1124 12708 1176 12714
rect 1124 12650 1176 12656
rect 1136 12170 1164 12650
rect 1124 12164 1176 12170
rect 1124 12106 1176 12112
rect 1032 11212 1084 11218
rect 1032 11154 1084 11160
rect 1136 9926 1164 12106
rect 1228 10062 1256 13806
rect 1768 13796 1820 13802
rect 1768 13738 1820 13744
rect 1364 13084 1740 13093
rect 1420 13082 1444 13084
rect 1500 13082 1524 13084
rect 1580 13082 1604 13084
rect 1660 13082 1684 13084
rect 1420 13030 1430 13082
rect 1674 13030 1684 13082
rect 1420 13028 1444 13030
rect 1500 13028 1524 13030
rect 1580 13028 1604 13030
rect 1660 13028 1684 13030
rect 1364 13019 1740 13028
rect 1780 12986 1808 13738
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 2056 12986 2084 13126
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 12374 1624 12786
rect 1688 12730 1716 12922
rect 1766 12744 1822 12753
rect 1688 12702 1766 12730
rect 1766 12679 1822 12688
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12442 1716 12582
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1584 12368 1636 12374
rect 1584 12310 1636 12316
rect 1780 12170 1808 12679
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1860 12368 1912 12374
rect 1858 12336 1860 12345
rect 1912 12336 1914 12345
rect 1964 12306 1992 12582
rect 1858 12271 1914 12280
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 1768 12164 1820 12170
rect 1768 12106 1820 12112
rect 1364 11996 1740 12005
rect 1420 11994 1444 11996
rect 1500 11994 1524 11996
rect 1580 11994 1604 11996
rect 1660 11994 1684 11996
rect 1420 11942 1430 11994
rect 1674 11942 1684 11994
rect 1420 11940 1444 11942
rect 1500 11940 1524 11942
rect 1580 11940 1604 11942
rect 1660 11940 1684 11942
rect 1364 11931 1740 11940
rect 2056 11898 2084 12174
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1504 11218 1532 11494
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1364 10908 1740 10917
rect 1420 10906 1444 10908
rect 1500 10906 1524 10908
rect 1580 10906 1604 10908
rect 1660 10906 1684 10908
rect 1420 10854 1430 10906
rect 1674 10854 1684 10906
rect 1420 10852 1444 10854
rect 1500 10852 1524 10854
rect 1580 10852 1604 10854
rect 1660 10852 1684 10854
rect 1364 10843 1740 10852
rect 1780 10810 1808 11630
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1780 10266 1808 10610
rect 1872 10606 1900 11494
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1674 10160 1730 10169
rect 1674 10095 1676 10104
rect 1728 10095 1730 10104
rect 1676 10066 1728 10072
rect 1216 10056 1268 10062
rect 1216 9998 1268 10004
rect 1124 9920 1176 9926
rect 1124 9862 1176 9868
rect 1364 9820 1740 9829
rect 1420 9818 1444 9820
rect 1500 9818 1524 9820
rect 1580 9818 1604 9820
rect 1660 9818 1684 9820
rect 1420 9766 1430 9818
rect 1674 9766 1684 9818
rect 1420 9764 1444 9766
rect 1500 9764 1524 9766
rect 1580 9764 1604 9766
rect 1660 9764 1684 9766
rect 1364 9755 1740 9764
rect 1364 8732 1740 8741
rect 1420 8730 1444 8732
rect 1500 8730 1524 8732
rect 1580 8730 1604 8732
rect 1660 8730 1684 8732
rect 1420 8678 1430 8730
rect 1674 8678 1684 8730
rect 1420 8676 1444 8678
rect 1500 8676 1524 8678
rect 1580 8676 1604 8678
rect 1660 8676 1684 8678
rect 1364 8667 1740 8676
rect 1124 7948 1176 7954
rect 1124 7890 1176 7896
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 5778 888 7822
rect 1136 7546 1164 7890
rect 1364 7644 1740 7653
rect 1420 7642 1444 7644
rect 1500 7642 1524 7644
rect 1580 7642 1604 7644
rect 1660 7642 1684 7644
rect 1420 7590 1430 7642
rect 1674 7590 1684 7642
rect 1420 7588 1444 7590
rect 1500 7588 1524 7590
rect 1580 7588 1604 7590
rect 1660 7588 1684 7590
rect 1364 7579 1740 7588
rect 1124 7540 1176 7546
rect 1124 7482 1176 7488
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 7002 1440 7278
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1780 6798 1808 10202
rect 1872 7342 1900 10542
rect 2148 10266 2176 13806
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13462 2636 13670
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2240 12986 2268 13398
rect 2700 13190 2728 13806
rect 3896 13530 3924 13806
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2412 12912 2464 12918
rect 2964 12912 3016 12918
rect 2464 12872 2636 12900
rect 2412 12854 2464 12860
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2502 12336 2558 12345
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2332 11694 2360 12106
rect 2424 12102 2452 12310
rect 2502 12271 2504 12280
rect 2556 12271 2558 12280
rect 2504 12242 2556 12248
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2516 11898 2544 12242
rect 2608 12238 2636 12872
rect 2964 12854 3016 12860
rect 2976 12782 3004 12854
rect 2964 12776 3016 12782
rect 2962 12744 2964 12753
rect 3016 12744 3018 12753
rect 2962 12679 3018 12688
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2976 12102 3004 12582
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2594 11792 2650 11801
rect 2516 11750 2594 11778
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1364 6556 1740 6565
rect 1420 6554 1444 6556
rect 1500 6554 1524 6556
rect 1580 6554 1604 6556
rect 1660 6554 1684 6556
rect 1420 6502 1430 6554
rect 1674 6502 1684 6554
rect 1420 6500 1444 6502
rect 1500 6500 1524 6502
rect 1580 6500 1604 6502
rect 1660 6500 1684 6502
rect 1364 6491 1740 6500
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 848 5772 900 5778
rect 848 5714 900 5720
rect 860 4690 888 5714
rect 1688 5710 1716 6326
rect 1780 6322 1808 6734
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 6458 1992 6598
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1364 5468 1740 5477
rect 1420 5466 1444 5468
rect 1500 5466 1524 5468
rect 1580 5466 1604 5468
rect 1660 5466 1684 5468
rect 1420 5414 1430 5466
rect 1674 5414 1684 5466
rect 1420 5412 1444 5414
rect 1500 5412 1524 5414
rect 1580 5412 1604 5414
rect 1660 5412 1684 5414
rect 1364 5403 1740 5412
rect 1780 5370 1808 6258
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1964 6118 1992 6190
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5914 1992 6054
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2056 5846 2084 9862
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 9042 2268 9318
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2148 8673 2176 8978
rect 2134 8664 2190 8673
rect 2332 8634 2360 9454
rect 2424 9042 2452 9454
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2134 8599 2190 8608
rect 2320 8628 2372 8634
rect 2148 7002 2176 8599
rect 2320 8570 2372 8576
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2240 8090 2268 8230
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2424 7002 2452 7278
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2412 6452 2464 6458
rect 2332 6412 2412 6440
rect 2228 6248 2280 6254
rect 2332 6236 2360 6412
rect 2412 6394 2464 6400
rect 2280 6208 2360 6236
rect 2228 6190 2280 6196
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 2424 5778 2452 6054
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2516 5658 2544 11750
rect 2594 11727 2650 11736
rect 2976 11529 3004 12038
rect 3436 11801 3464 13126
rect 3896 12986 3924 13466
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3422 11792 3478 11801
rect 3422 11727 3478 11736
rect 3528 11694 3556 12038
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 2962 11520 3018 11529
rect 2962 11455 3018 11464
rect 3252 11014 3280 11630
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 2686 10568 2742 10577
rect 2686 10503 2742 10512
rect 2700 10198 2728 10503
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2608 9722 2636 10066
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2608 8634 2636 8978
rect 2792 8838 2820 9930
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2608 7410 2636 8570
rect 2700 8362 2728 8774
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2596 6928 2648 6934
rect 2596 6870 2648 6876
rect 2608 6458 2636 6870
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2424 5630 2544 5658
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 2240 5250 2268 5510
rect 2240 5234 2360 5250
rect 2240 5228 2372 5234
rect 2240 5222 2320 5228
rect 2320 5170 2372 5176
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 848 4684 900 4690
rect 848 4626 900 4632
rect 860 3602 888 4626
rect 1364 4380 1740 4389
rect 1420 4378 1444 4380
rect 1500 4378 1524 4380
rect 1580 4378 1604 4380
rect 1660 4378 1684 4380
rect 1420 4326 1430 4378
rect 1674 4326 1684 4378
rect 1420 4324 1444 4326
rect 1500 4324 1524 4326
rect 1580 4324 1604 4326
rect 1660 4324 1684 4326
rect 1364 4315 1740 4324
rect 1964 4078 1992 4966
rect 2240 4078 2268 5102
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4826 2360 4966
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 848 3596 900 3602
rect 848 3538 900 3544
rect 1216 3596 1268 3602
rect 1216 3538 1268 3544
rect 860 2774 888 3538
rect 1228 3194 1256 3538
rect 1364 3292 1740 3301
rect 1420 3290 1444 3292
rect 1500 3290 1524 3292
rect 1580 3290 1604 3292
rect 1660 3290 1684 3292
rect 1420 3238 1430 3290
rect 1674 3238 1684 3290
rect 1420 3236 1444 3238
rect 1500 3236 1524 3238
rect 1580 3236 1604 3238
rect 1660 3236 1684 3238
rect 1364 3227 1740 3236
rect 1216 3188 1268 3194
rect 1216 3130 1268 3136
rect 1584 2984 1636 2990
rect 1582 2952 1584 2961
rect 1636 2952 1638 2961
rect 1582 2887 1638 2896
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 860 2746 1256 2774
rect 1228 2514 1256 2746
rect 1780 2582 1808 2790
rect 1768 2576 1820 2582
rect 1768 2518 1820 2524
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1032 2032 1084 2038
rect 1032 1974 1084 1980
rect 20 1216 72 1222
rect 20 1158 72 1164
rect 32 400 60 1158
rect 1044 814 1072 1974
rect 1124 1760 1176 1766
rect 1124 1702 1176 1708
rect 1136 1562 1164 1702
rect 1228 1562 1256 2450
rect 1364 2204 1740 2213
rect 1420 2202 1444 2204
rect 1500 2202 1524 2204
rect 1580 2202 1604 2204
rect 1660 2202 1684 2204
rect 1420 2150 1430 2202
rect 1674 2150 1684 2202
rect 1420 2148 1444 2150
rect 1500 2148 1524 2150
rect 1580 2148 1604 2150
rect 1660 2148 1684 2150
rect 1364 2139 1740 2148
rect 1124 1556 1176 1562
rect 1124 1498 1176 1504
rect 1216 1556 1268 1562
rect 1216 1498 1268 1504
rect 1228 1018 1256 1498
rect 1768 1284 1820 1290
rect 1768 1226 1820 1232
rect 1364 1116 1740 1125
rect 1420 1114 1444 1116
rect 1500 1114 1524 1116
rect 1580 1114 1604 1116
rect 1660 1114 1684 1116
rect 1420 1062 1430 1114
rect 1674 1062 1684 1114
rect 1420 1060 1444 1062
rect 1500 1060 1524 1062
rect 1580 1060 1604 1062
rect 1660 1060 1684 1062
rect 1364 1051 1740 1060
rect 1216 1012 1268 1018
rect 1216 954 1268 960
rect 1032 808 1084 814
rect 1032 750 1084 756
rect 1032 672 1084 678
rect 1780 626 1808 1226
rect 1872 746 1900 3878
rect 2332 3738 2360 4014
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2332 2990 2360 3674
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2424 1902 2452 5630
rect 2700 4826 2728 7890
rect 2884 7546 2912 9930
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9518 3188 9862
rect 3252 9722 3280 10134
rect 3344 10130 3372 11154
rect 3528 10606 3556 11630
rect 3988 11558 4016 12582
rect 4172 12186 4200 13262
rect 4264 12306 4292 14214
rect 4356 13870 4384 14418
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4364 13628 4740 13637
rect 4420 13626 4444 13628
rect 4500 13626 4524 13628
rect 4580 13626 4604 13628
rect 4660 13626 4684 13628
rect 4420 13574 4430 13626
rect 4674 13574 4684 13626
rect 4420 13572 4444 13574
rect 4500 13572 4524 13574
rect 4580 13572 4604 13574
rect 4660 13572 4684 13574
rect 4364 13563 4740 13572
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4364 12540 4740 12549
rect 4420 12538 4444 12540
rect 4500 12538 4524 12540
rect 4580 12538 4604 12540
rect 4660 12538 4684 12540
rect 4420 12486 4430 12538
rect 4674 12486 4684 12538
rect 4420 12484 4444 12486
rect 4500 12484 4524 12486
rect 4580 12484 4604 12486
rect 4660 12484 4684 12486
rect 4364 12475 4740 12484
rect 4816 12442 4844 12718
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4804 12436 4856 12442
rect 4632 12406 4804 12434
rect 4632 12306 4660 12406
rect 4804 12378 4856 12384
rect 4908 12306 4936 12582
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4172 12158 4292 12186
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 8922 3188 9318
rect 3252 9042 3280 9454
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3160 8894 3280 8922
rect 3344 8906 3372 10066
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3528 9178 3556 9454
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3608 9104 3660 9110
rect 3528 9052 3608 9058
rect 3528 9046 3660 9052
rect 3528 9030 3648 9046
rect 3528 8922 3556 9030
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3054 8664 3110 8673
rect 3054 8599 3056 8608
rect 3108 8599 3110 8608
rect 3056 8570 3108 8576
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2870 7440 2926 7449
rect 2870 7375 2926 7384
rect 2964 7404 3016 7410
rect 2884 6866 2912 7375
rect 2964 7346 3016 7352
rect 2976 6934 3004 7346
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6662 2912 6802
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5302 2820 6054
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2700 4128 2728 4762
rect 2792 4282 2820 5238
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2780 4140 2832 4146
rect 2700 4100 2780 4128
rect 2780 4082 2832 4088
rect 3068 3126 3096 7822
rect 3160 7818 3188 8774
rect 3252 8498 3280 8894
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3436 8894 3556 8922
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3436 8786 3464 8894
rect 3344 8758 3464 8786
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3344 8430 3372 8758
rect 3424 8628 3476 8634
rect 3620 8616 3648 8910
rect 3712 8634 3740 10746
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 9625 3832 10406
rect 3790 9616 3846 9625
rect 3896 9586 3924 11018
rect 3790 9551 3846 9560
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3896 8838 3924 9386
rect 3988 9024 4016 11494
rect 4172 11218 4200 12038
rect 4264 11830 4292 12158
rect 4632 12102 4660 12242
rect 4712 12232 4764 12238
rect 4764 12192 4844 12220
rect 4712 12174 4764 12180
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4724 11694 4752 11766
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4264 11150 4292 11630
rect 4364 11452 4740 11461
rect 4420 11450 4444 11452
rect 4500 11450 4524 11452
rect 4580 11450 4604 11452
rect 4660 11450 4684 11452
rect 4420 11398 4430 11450
rect 4674 11398 4684 11450
rect 4420 11396 4444 11398
rect 4500 11396 4524 11398
rect 4580 11396 4604 11398
rect 4660 11396 4684 11398
rect 4364 11387 4740 11396
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4342 11112 4398 11121
rect 4342 11047 4344 11056
rect 4396 11047 4398 11056
rect 4344 11018 4396 11024
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4080 10606 4108 10950
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 4080 9926 4108 9959
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4172 9674 4200 10542
rect 4264 10130 4292 10950
rect 4724 10588 4752 11154
rect 4816 11014 4844 12192
rect 4908 11354 4936 12242
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5092 11898 5120 12106
rect 5184 11898 5212 14436
rect 5356 14418 5408 14424
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12850 5396 13126
rect 5552 12986 5580 13670
rect 6104 13394 6132 14486
rect 6564 14482 6592 15302
rect 6656 15162 6684 15600
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6748 15042 6776 15302
rect 7300 15162 7328 15694
rect 7378 15600 7434 15694
rect 8114 15600 8170 16000
rect 8850 15722 8906 16000
rect 8850 15694 9168 15722
rect 8850 15600 8906 15694
rect 7364 15260 7740 15269
rect 7420 15258 7444 15260
rect 7500 15258 7524 15260
rect 7580 15258 7604 15260
rect 7660 15258 7684 15260
rect 7420 15206 7430 15258
rect 7674 15206 7684 15258
rect 7420 15204 7444 15206
rect 7500 15204 7524 15206
rect 7580 15204 7604 15206
rect 7660 15204 7684 15206
rect 7364 15195 7740 15204
rect 8128 15162 8156 15600
rect 9140 15162 9168 15694
rect 9586 15600 9642 16000
rect 10322 15600 10378 16000
rect 11058 15600 11114 16000
rect 17682 15600 17738 16000
rect 18418 15600 18474 16000
rect 19154 15600 19210 16000
rect 19890 15722 19946 16000
rect 19890 15694 20208 15722
rect 19890 15600 19946 15694
rect 9600 15162 9628 15600
rect 10336 15162 10364 15600
rect 11072 15162 11100 15600
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 13364 15260 13740 15269
rect 13420 15258 13444 15260
rect 13500 15258 13524 15260
rect 13580 15258 13604 15260
rect 13660 15258 13684 15260
rect 13420 15206 13430 15258
rect 13674 15206 13684 15258
rect 13420 15204 13444 15206
rect 13500 15204 13524 15206
rect 13580 15204 13604 15206
rect 13660 15204 13684 15206
rect 13364 15195 13740 15204
rect 14476 15162 14504 15302
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 6656 15014 6776 15042
rect 7656 15020 7708 15026
rect 6656 14618 6684 15014
rect 7656 14962 7708 14968
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 13802 6224 14214
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5356 12844 5408 12850
rect 5276 12804 5356 12832
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5170 11656 5226 11665
rect 5000 11614 5170 11642
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4894 11248 4950 11257
rect 4894 11183 4950 11192
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4816 10742 4844 10950
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4804 10600 4856 10606
rect 4724 10560 4804 10588
rect 4804 10542 4856 10548
rect 4364 10364 4740 10373
rect 4420 10362 4444 10364
rect 4500 10362 4524 10364
rect 4580 10362 4604 10364
rect 4660 10362 4684 10364
rect 4420 10310 4430 10362
rect 4674 10310 4684 10362
rect 4420 10308 4444 10310
rect 4500 10308 4524 10310
rect 4580 10308 4604 10310
rect 4660 10308 4684 10310
rect 4364 10299 4740 10308
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4172 9646 4292 9674
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4068 9036 4120 9042
rect 3988 8996 4068 9024
rect 4068 8978 4120 8984
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3424 8570 3476 8576
rect 3528 8588 3648 8616
rect 3700 8628 3752 8634
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 8022 3372 8230
rect 3436 8090 3464 8570
rect 3528 8090 3556 8588
rect 3700 8570 3752 8576
rect 3804 8514 3832 8774
rect 3620 8486 3832 8514
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3514 7984 3570 7993
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3344 7546 3372 7958
rect 3514 7919 3516 7928
rect 3568 7919 3570 7928
rect 3516 7890 3568 7896
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 6798 3280 7210
rect 3528 7002 3556 7278
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3620 6866 3648 8486
rect 3792 8288 3844 8294
rect 3712 8248 3792 8276
rect 3712 7342 3740 8248
rect 3792 8230 3844 8236
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3804 7002 3832 7278
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3240 6792 3292 6798
rect 3292 6752 3372 6780
rect 3240 6734 3292 6740
rect 3344 5710 3372 6752
rect 3620 6458 3648 6802
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3712 5574 3740 6802
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6322 3832 6598
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3804 5914 3832 6258
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 3068 2990 3096 3062
rect 3436 2990 3464 3606
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 2516 2650 2544 2926
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 3528 1970 3556 4966
rect 3712 4758 3740 5510
rect 3700 4752 3752 4758
rect 3700 4694 3752 4700
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3620 4078 3648 4626
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3804 4282 3832 4558
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3620 2990 3648 4014
rect 3804 3670 3832 4218
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3896 3194 3924 8774
rect 4172 8362 4200 9454
rect 4264 8974 4292 9646
rect 4724 9518 4752 9862
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4364 9276 4740 9285
rect 4420 9274 4444 9276
rect 4500 9274 4524 9276
rect 4580 9274 4604 9276
rect 4660 9274 4684 9276
rect 4420 9222 4430 9274
rect 4674 9222 4684 9274
rect 4420 9220 4444 9222
rect 4500 9220 4524 9222
rect 4580 9220 4604 9222
rect 4660 9220 4684 9222
rect 4364 9211 4740 9220
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4356 8294 4384 8434
rect 4068 8288 4120 8294
rect 4344 8288 4396 8294
rect 4068 8230 4120 8236
rect 4264 8248 4344 8276
rect 4080 8090 4108 8230
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 6866 4016 7754
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7478 4200 7686
rect 4068 7472 4120 7478
rect 4066 7440 4068 7449
rect 4160 7472 4212 7478
rect 4120 7440 4122 7449
rect 4160 7414 4212 7420
rect 4066 7375 4122 7384
rect 4264 7342 4292 8248
rect 4344 8230 4396 8236
rect 4364 8188 4740 8197
rect 4420 8186 4444 8188
rect 4500 8186 4524 8188
rect 4580 8186 4604 8188
rect 4660 8186 4684 8188
rect 4420 8134 4430 8186
rect 4674 8134 4684 8186
rect 4420 8132 4444 8134
rect 4500 8132 4524 8134
rect 4580 8132 4604 8134
rect 4660 8132 4684 8134
rect 4364 8123 4740 8132
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4080 7002 4108 7278
rect 4252 7200 4304 7206
rect 4172 7148 4252 7154
rect 4172 7142 4304 7148
rect 4172 7126 4292 7142
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4172 6662 4200 7126
rect 4364 7100 4740 7109
rect 4420 7098 4444 7100
rect 4500 7098 4524 7100
rect 4580 7098 4604 7100
rect 4660 7098 4684 7100
rect 4420 7046 4430 7098
rect 4674 7046 4684 7098
rect 4420 7044 4444 7046
rect 4500 7044 4524 7046
rect 4580 7044 4604 7046
rect 4660 7044 4684 7046
rect 4364 7035 4740 7044
rect 4816 6866 4844 10542
rect 4908 9500 4936 11183
rect 5000 11150 5028 11614
rect 5170 11591 5226 11600
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5092 11354 5120 11494
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5184 11082 5212 11494
rect 5276 11200 5304 12804
rect 5356 12786 5408 12792
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5368 12306 5396 12378
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5448 12096 5500 12102
rect 5368 12056 5448 12084
rect 5368 11393 5396 12056
rect 5448 12038 5500 12044
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5354 11384 5410 11393
rect 5354 11319 5410 11328
rect 5356 11212 5408 11218
rect 5276 11172 5356 11200
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5184 10674 5212 11018
rect 5276 10810 5304 11172
rect 5356 11154 5408 11160
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5460 9654 5488 11630
rect 5552 10674 5580 12922
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5644 11778 5672 12038
rect 5644 11762 5764 11778
rect 5644 11756 5776 11762
rect 5644 11750 5724 11756
rect 5724 11698 5776 11704
rect 5540 10668 5592 10674
rect 5828 10656 5856 13262
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5920 12986 5948 13194
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5920 11694 5948 12242
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5540 10610 5592 10616
rect 5736 10628 5856 10656
rect 5736 10538 5764 10628
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5816 10532 5868 10538
rect 5816 10474 5868 10480
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10198 5580 10406
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9722 5580 9862
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5448 9648 5500 9654
rect 5828 9602 5856 10474
rect 6012 10112 6040 12106
rect 5448 9590 5500 9596
rect 5736 9574 5856 9602
rect 5920 10084 6040 10112
rect 4988 9512 5040 9518
rect 4908 9472 4988 9500
rect 5264 9512 5316 9518
rect 5040 9472 5212 9500
rect 4988 9454 5040 9460
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5000 8090 5028 8978
rect 5092 8430 5120 8978
rect 5184 8430 5212 9472
rect 5264 9454 5316 9460
rect 5276 9178 5304 9454
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5368 9058 5396 9386
rect 5276 9030 5396 9058
rect 5540 9036 5592 9042
rect 5276 8974 5304 9030
rect 5540 8978 5592 8984
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5092 8090 5120 8366
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5184 7342 5212 8026
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 4826 4200 6598
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4172 4078 4200 4558
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4172 3738 4200 4014
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3620 2582 3648 2926
rect 4264 2774 4292 6734
rect 5000 6186 5028 7278
rect 5276 7274 5304 8910
rect 5552 8498 5580 8978
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5644 8498 5672 8842
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 7886 5672 8434
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 7528 5396 7686
rect 5448 7540 5500 7546
rect 5368 7500 5448 7528
rect 5448 7482 5500 7488
rect 5538 7440 5594 7449
rect 5644 7410 5672 7822
rect 5538 7375 5594 7384
rect 5632 7404 5684 7410
rect 5552 7274 5580 7375
rect 5632 7346 5684 7352
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 4364 6012 4740 6021
rect 4420 6010 4444 6012
rect 4500 6010 4524 6012
rect 4580 6010 4604 6012
rect 4660 6010 4684 6012
rect 4420 5958 4430 6010
rect 4674 5958 4684 6010
rect 4420 5956 4444 5958
rect 4500 5956 4524 5958
rect 4580 5956 4604 5958
rect 4660 5956 4684 5958
rect 4364 5947 4740 5956
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 4364 4924 4740 4933
rect 4420 4922 4444 4924
rect 4500 4922 4524 4924
rect 4580 4922 4604 4924
rect 4660 4922 4684 4924
rect 4420 4870 4430 4922
rect 4674 4870 4684 4922
rect 4420 4868 4444 4870
rect 4500 4868 4524 4870
rect 4580 4868 4604 4870
rect 4660 4868 4684 4870
rect 4364 4859 4740 4868
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4356 4146 4384 4626
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4364 3836 4740 3845
rect 4420 3834 4444 3836
rect 4500 3834 4524 3836
rect 4580 3834 4604 3836
rect 4660 3834 4684 3836
rect 4420 3782 4430 3834
rect 4674 3782 4684 3834
rect 4420 3780 4444 3782
rect 4500 3780 4524 3782
rect 4580 3780 4604 3782
rect 4660 3780 4684 3782
rect 4364 3771 4740 3780
rect 5000 3602 5028 5714
rect 5092 5710 5120 6598
rect 5276 5710 5304 6938
rect 5460 6934 5488 7142
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5460 6186 5488 6870
rect 5644 6798 5672 7346
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5552 6254 5580 6394
rect 5736 6322 5764 9574
rect 5920 9518 5948 10084
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 6012 9450 6040 9930
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5092 5234 5120 5646
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5276 4486 5304 5646
rect 5460 5166 5488 5850
rect 5736 5710 5764 6054
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5644 5234 5672 5578
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5460 4826 5488 5102
rect 5828 5030 5856 9046
rect 5920 8838 5948 9318
rect 6104 8906 6132 13126
rect 6288 12782 6316 13942
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6472 12986 6500 13126
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6196 9994 6224 11290
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5920 8362 5948 8774
rect 6288 8430 6316 12718
rect 6656 12434 6684 14554
rect 6748 14482 6776 14826
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6748 12918 6776 14418
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6840 12782 6868 13806
rect 6932 13462 6960 14826
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7116 14482 7144 14758
rect 7668 14618 7696 14962
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7364 14172 7740 14181
rect 7420 14170 7444 14172
rect 7500 14170 7524 14172
rect 7580 14170 7604 14172
rect 7660 14170 7684 14172
rect 7420 14118 7430 14170
rect 7674 14118 7684 14170
rect 7420 14116 7444 14118
rect 7500 14116 7524 14118
rect 7580 14116 7604 14118
rect 7660 14116 7684 14118
rect 7364 14107 7740 14116
rect 7852 14074 7880 14894
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7944 14618 7972 14758
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7760 13462 7788 13806
rect 6920 13456 6972 13462
rect 7748 13456 7800 13462
rect 6972 13416 7052 13444
rect 6920 13398 6972 13404
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6564 12406 6684 12434
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 11626 6500 11698
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 10606 6408 11494
rect 6472 10674 6500 11562
rect 6564 11218 6592 12406
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6656 11286 6684 12038
rect 6932 11778 6960 13126
rect 7024 12986 7052 13416
rect 7748 13398 7800 13404
rect 8036 13274 8064 14418
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 13462 8156 14214
rect 8588 14074 8616 14894
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8220 13326 8248 13806
rect 8588 13530 8616 13806
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8208 13320 8260 13326
rect 8114 13288 8170 13297
rect 8036 13246 8114 13274
rect 8036 13190 8064 13246
rect 8208 13262 8260 13268
rect 8114 13223 8170 13232
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7364 13084 7740 13093
rect 7420 13082 7444 13084
rect 7500 13082 7524 13084
rect 7580 13082 7604 13084
rect 7660 13082 7684 13084
rect 7420 13030 7430 13082
rect 7674 13030 7684 13082
rect 7420 13028 7444 13030
rect 7500 13028 7524 13030
rect 7580 13028 7604 13030
rect 7660 13028 7684 13030
rect 7364 13019 7740 13028
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 12238 7328 12582
rect 7484 12442 7512 12650
rect 8220 12646 8248 13262
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7472 12436 7524 12442
rect 8680 12434 8708 14826
rect 8956 14618 8984 14894
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8772 13394 8800 14418
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9140 13870 9168 14350
rect 9324 14278 9352 14350
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9324 13870 9352 14214
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8680 12406 8800 12434
rect 7472 12378 7524 12384
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 6748 11750 6960 11778
rect 6748 11558 6776 11750
rect 6826 11656 6882 11665
rect 6826 11591 6828 11600
rect 6880 11591 6882 11600
rect 7196 11620 7248 11626
rect 6828 11562 6880 11568
rect 7196 11562 7248 11568
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9518 6500 9862
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6472 8362 6500 9454
rect 6564 9450 6592 11154
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10810 6684 11086
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 5920 6866 5948 8298
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 8090 6040 8230
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6000 7744 6052 7750
rect 6104 7732 6132 8026
rect 6184 8016 6236 8022
rect 6472 8004 6500 8298
rect 6236 7976 6500 8004
rect 6184 7958 6236 7964
rect 6052 7704 6132 7732
rect 6000 7686 6052 7692
rect 6104 7002 6132 7704
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6092 6996 6144 7002
rect 6368 6996 6420 7002
rect 6092 6938 6144 6944
rect 6288 6956 6368 6984
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 6000 6452 6052 6458
rect 6104 6440 6132 6938
rect 6288 6662 6316 6956
rect 6368 6938 6420 6944
rect 6472 6934 6500 7142
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6052 6412 6132 6440
rect 6000 6394 6052 6400
rect 6104 6236 6132 6412
rect 6184 6248 6236 6254
rect 6104 6208 6184 6236
rect 6184 6190 6236 6196
rect 6472 5778 6500 6870
rect 6564 6254 6592 9386
rect 6656 8974 6684 10746
rect 6748 10266 6776 11494
rect 7208 11354 7236 11562
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7208 11121 7236 11290
rect 7194 11112 7250 11121
rect 7194 11047 7250 11056
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6840 9704 6868 10610
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 10441 6960 10542
rect 6918 10432 6974 10441
rect 6918 10367 6974 10376
rect 7300 9926 7328 12174
rect 7364 11996 7740 12005
rect 7420 11994 7444 11996
rect 7500 11994 7524 11996
rect 7580 11994 7604 11996
rect 7660 11994 7684 11996
rect 7420 11942 7430 11994
rect 7674 11942 7684 11994
rect 7420 11940 7444 11942
rect 7500 11940 7524 11942
rect 7580 11940 7604 11942
rect 7660 11940 7684 11942
rect 7364 11931 7740 11940
rect 7852 11354 7880 12242
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11694 7972 12038
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 8496 11354 8524 12242
rect 8772 12238 8800 12406
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7364 10908 7740 10917
rect 7420 10906 7444 10908
rect 7500 10906 7524 10908
rect 7580 10906 7604 10908
rect 7660 10906 7684 10908
rect 7420 10854 7430 10906
rect 7674 10854 7684 10906
rect 7420 10852 7444 10854
rect 7500 10852 7524 10854
rect 7580 10852 7604 10854
rect 7660 10852 7684 10854
rect 7364 10843 7740 10852
rect 8128 10742 8156 11086
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8116 10736 8168 10742
rect 8220 10713 8248 10950
rect 8404 10810 8432 11222
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8116 10678 8168 10684
rect 8206 10704 8262 10713
rect 8128 10266 8156 10678
rect 8206 10639 8262 10648
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 6920 9716 6972 9722
rect 6840 9676 6920 9704
rect 6920 9658 6972 9664
rect 7300 9586 7328 9862
rect 7364 9820 7740 9829
rect 7420 9818 7444 9820
rect 7500 9818 7524 9820
rect 7580 9818 7604 9820
rect 7660 9818 7684 9820
rect 7420 9766 7430 9818
rect 7674 9766 7684 9818
rect 7420 9764 7444 9766
rect 7500 9764 7524 9766
rect 7580 9764 7604 9766
rect 7660 9764 7684 9766
rect 7364 9755 7740 9764
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6656 8022 6684 8910
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6748 6866 6776 8366
rect 6840 7954 6868 8978
rect 7364 8732 7740 8741
rect 7420 8730 7444 8732
rect 7500 8730 7524 8732
rect 7580 8730 7604 8732
rect 7660 8730 7684 8732
rect 7420 8678 7430 8730
rect 7674 8678 7684 8730
rect 7420 8676 7444 8678
rect 7500 8676 7524 8678
rect 7580 8676 7604 8678
rect 7660 8676 7684 8678
rect 7364 8667 7740 8676
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 7024 6866 7052 8230
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7208 7546 7236 7686
rect 7300 7546 7328 7686
rect 7364 7644 7740 7653
rect 7420 7642 7444 7644
rect 7500 7642 7524 7644
rect 7580 7642 7604 7644
rect 7660 7642 7684 7644
rect 7420 7590 7430 7642
rect 7674 7590 7684 7642
rect 7420 7588 7444 7590
rect 7500 7588 7524 7590
rect 7580 7588 7604 7590
rect 7660 7588 7684 7590
rect 7364 7579 7740 7588
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7852 7410 7880 10066
rect 8220 10010 8248 10639
rect 8484 10600 8536 10606
rect 8536 10560 8708 10588
rect 8484 10542 8536 10548
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8496 10266 8524 10406
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8680 10130 8708 10560
rect 8300 10124 8352 10130
rect 8668 10124 8720 10130
rect 8352 10084 8616 10112
rect 8300 10066 8352 10072
rect 8220 9982 8524 10010
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 7944 9450 7972 9862
rect 8116 9512 8168 9518
rect 8312 9500 8340 9862
rect 8168 9472 8340 9500
rect 8116 9454 8168 9460
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7944 8514 7972 9386
rect 7944 8486 8064 8514
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 8036 6662 8064 8486
rect 8300 6928 8352 6934
rect 8352 6888 8432 6916
rect 8300 6870 8352 6876
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7364 6556 7740 6565
rect 7420 6554 7444 6556
rect 7500 6554 7524 6556
rect 7580 6554 7604 6556
rect 7660 6554 7684 6556
rect 7420 6502 7430 6554
rect 7674 6502 7684 6554
rect 7420 6500 7444 6502
rect 7500 6500 7524 6502
rect 7580 6500 7604 6502
rect 7660 6500 7684 6502
rect 7364 6491 7740 6500
rect 8036 6390 8064 6598
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6748 5914 6776 6122
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 5920 5370 5948 5714
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 6656 5234 6684 5782
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 6104 4758 6132 4966
rect 6656 4826 6684 5170
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6090 4584 6146 4593
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5184 4078 5212 4422
rect 5920 4214 5948 4558
rect 6090 4519 6092 4528
rect 6144 4519 6146 4528
rect 6092 4490 6144 4496
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5368 3534 5396 3878
rect 6104 3602 6132 4490
rect 6642 3632 6698 3641
rect 6092 3596 6144 3602
rect 6642 3567 6698 3576
rect 6092 3538 6144 3544
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 6656 3466 6684 3567
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 5092 2774 5120 3402
rect 6656 3194 6684 3402
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6840 3058 6868 4966
rect 6932 3738 6960 5306
rect 7024 4282 7052 5850
rect 7116 5778 7144 6258
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 7208 5914 7236 6054
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 4690 7236 5510
rect 7300 5273 7328 6054
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7932 5704 7984 5710
rect 7852 5664 7932 5692
rect 7364 5468 7740 5477
rect 7420 5466 7444 5468
rect 7500 5466 7524 5468
rect 7580 5466 7604 5468
rect 7660 5466 7684 5468
rect 7420 5414 7430 5466
rect 7674 5414 7684 5466
rect 7420 5412 7444 5414
rect 7500 5412 7524 5414
rect 7580 5412 7604 5414
rect 7660 5412 7684 5414
rect 7364 5403 7740 5412
rect 7286 5264 7342 5273
rect 7286 5199 7342 5208
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7196 4548 7248 4554
rect 7484 4536 7512 4626
rect 7668 4554 7696 5170
rect 7748 4616 7800 4622
rect 7746 4584 7748 4593
rect 7800 4584 7802 4593
rect 7248 4508 7512 4536
rect 7656 4548 7708 4554
rect 7196 4490 7248 4496
rect 7746 4519 7802 4528
rect 7656 4490 7708 4496
rect 7364 4380 7740 4389
rect 7420 4378 7444 4380
rect 7500 4378 7524 4380
rect 7580 4378 7604 4380
rect 7660 4378 7684 4380
rect 7420 4326 7430 4378
rect 7674 4326 7684 4378
rect 7420 4324 7444 4326
rect 7500 4324 7524 4326
rect 7580 4324 7604 4326
rect 7660 4324 7684 4326
rect 7364 4315 7740 4324
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 7024 3505 7052 4218
rect 7010 3496 7066 3505
rect 7010 3431 7066 3440
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3194 7052 3334
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 4172 2746 4292 2774
rect 4364 2748 4740 2757
rect 4420 2746 4444 2748
rect 4500 2746 4524 2748
rect 4580 2746 4604 2748
rect 4660 2746 4684 2748
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 3608 2576 3660 2582
rect 4080 2553 4108 2586
rect 3608 2518 3660 2524
rect 4066 2544 4122 2553
rect 4066 2479 4122 2488
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 3712 1562 3740 2246
rect 3804 1562 3832 2246
rect 3896 2106 3924 2382
rect 4172 2106 4200 2746
rect 4420 2694 4430 2746
rect 4674 2694 4684 2746
rect 4420 2692 4444 2694
rect 4500 2692 4524 2694
rect 4580 2692 4604 2694
rect 4660 2692 4684 2694
rect 4364 2683 4740 2692
rect 5000 2746 5120 2774
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 3896 1562 3924 2042
rect 4172 1562 4200 2042
rect 5000 1902 5028 2746
rect 5184 2514 5212 2790
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 7300 2446 7328 3402
rect 7364 3292 7740 3301
rect 7420 3290 7444 3292
rect 7500 3290 7524 3292
rect 7580 3290 7604 3292
rect 7660 3290 7684 3292
rect 7420 3238 7430 3290
rect 7674 3238 7684 3290
rect 7420 3236 7444 3238
rect 7500 3236 7524 3238
rect 7580 3236 7604 3238
rect 7660 3236 7684 3238
rect 7364 3227 7740 3236
rect 7852 2961 7880 5664
rect 8220 5681 8248 5850
rect 8206 5672 8262 5681
rect 7932 5646 7984 5652
rect 8128 5630 8206 5658
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7944 5370 7972 5510
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4146 7972 4966
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8036 3777 8064 3878
rect 8022 3768 8078 3777
rect 8022 3703 8078 3712
rect 8036 3670 8064 3703
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 8128 3466 8156 5630
rect 8206 5607 8262 5616
rect 8312 5370 8340 6054
rect 8404 5914 8432 6888
rect 8496 6440 8524 9982
rect 8588 6934 8616 10084
rect 8668 10066 8720 10072
rect 8680 9926 8708 10066
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8498 8708 8774
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8576 6452 8628 6458
rect 8496 6412 8576 6440
rect 8576 6394 8628 6400
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5914 8616 6054
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8206 4720 8262 4729
rect 8206 4655 8262 4664
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 2990 7972 3334
rect 7932 2984 7984 2990
rect 7838 2952 7894 2961
rect 7932 2926 7984 2932
rect 7838 2887 7840 2896
rect 7892 2887 7894 2896
rect 7840 2858 7892 2864
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 4988 1896 5040 1902
rect 4342 1864 4398 1873
rect 4988 1838 5040 1844
rect 7012 1896 7064 1902
rect 7012 1838 7064 1844
rect 4342 1799 4344 1808
rect 4396 1799 4398 1808
rect 5724 1828 5776 1834
rect 4344 1770 4396 1776
rect 5724 1770 5776 1776
rect 4252 1760 4304 1766
rect 4252 1702 4304 1708
rect 3700 1556 3752 1562
rect 3700 1498 3752 1504
rect 3792 1556 3844 1562
rect 3792 1498 3844 1504
rect 3884 1556 3936 1562
rect 3884 1498 3936 1504
rect 4160 1556 4212 1562
rect 4160 1498 4212 1504
rect 4264 1358 4292 1702
rect 4364 1660 4740 1669
rect 4420 1658 4444 1660
rect 4500 1658 4524 1660
rect 4580 1658 4604 1660
rect 4660 1658 4684 1660
rect 4420 1606 4430 1658
rect 4674 1606 4684 1658
rect 4420 1604 4444 1606
rect 4500 1604 4524 1606
rect 4580 1604 4604 1606
rect 4660 1604 4684 1606
rect 4364 1595 4740 1604
rect 5736 1494 5764 1770
rect 6920 1760 6972 1766
rect 6920 1702 6972 1708
rect 6932 1562 6960 1702
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 5724 1488 5776 1494
rect 5724 1430 5776 1436
rect 6932 1426 6960 1498
rect 7024 1442 7052 1838
rect 7300 1494 7328 2246
rect 7364 2204 7740 2213
rect 7420 2202 7444 2204
rect 7500 2202 7524 2204
rect 7580 2202 7604 2204
rect 7660 2202 7684 2204
rect 7420 2150 7430 2202
rect 7674 2150 7684 2202
rect 7420 2148 7444 2150
rect 7500 2148 7524 2150
rect 7580 2148 7604 2150
rect 7660 2148 7684 2150
rect 7364 2139 7740 2148
rect 7562 2000 7618 2009
rect 7562 1935 7618 1944
rect 7576 1902 7604 1935
rect 7564 1896 7616 1902
rect 7564 1838 7616 1844
rect 7748 1896 7800 1902
rect 7748 1838 7800 1844
rect 7288 1488 7340 1494
rect 7024 1436 7288 1442
rect 7024 1430 7340 1436
rect 7024 1426 7328 1430
rect 5448 1420 5500 1426
rect 5448 1362 5500 1368
rect 6920 1420 6972 1426
rect 6920 1362 6972 1368
rect 7012 1420 7328 1426
rect 7064 1414 7328 1420
rect 7012 1362 7064 1368
rect 4160 1352 4212 1358
rect 4160 1294 4212 1300
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 4172 1018 4200 1294
rect 4160 1012 4212 1018
rect 4160 954 4212 960
rect 1860 740 1912 746
rect 1860 682 1912 688
rect 2504 740 2556 746
rect 2504 682 2556 688
rect 1032 614 1084 620
rect 1044 490 1072 614
rect 860 462 1072 490
rect 1688 598 1808 626
rect 860 400 888 462
rect 1688 400 1716 598
rect 2516 400 2544 682
rect 3332 672 3384 678
rect 3332 614 3384 620
rect 4068 672 4120 678
rect 4344 672 4396 678
rect 4068 614 4120 620
rect 4172 632 4344 660
rect 3344 400 3372 614
rect 18 0 74 400
rect 846 0 902 400
rect 1674 0 1730 400
rect 2502 0 2558 400
rect 3330 0 3386 400
rect 4080 270 4108 614
rect 4172 400 4200 632
rect 5172 672 5224 678
rect 4344 614 4396 620
rect 5000 632 5172 660
rect 4364 572 4740 581
rect 4420 570 4444 572
rect 4500 570 4524 572
rect 4580 570 4604 572
rect 4660 570 4684 572
rect 4420 518 4430 570
rect 4674 518 4684 570
rect 4420 516 4444 518
rect 4500 516 4524 518
rect 4580 516 4604 518
rect 4660 516 4684 518
rect 4364 507 4740 516
rect 5000 400 5028 632
rect 5172 614 5224 620
rect 5460 406 5488 1362
rect 7576 1358 7604 1838
rect 7760 1766 7788 1838
rect 7840 1828 7892 1834
rect 7840 1770 7892 1776
rect 7656 1760 7708 1766
rect 7656 1702 7708 1708
rect 7748 1760 7800 1766
rect 7748 1702 7800 1708
rect 7668 1358 7696 1702
rect 7852 1562 7880 1770
rect 8116 1760 8168 1766
rect 8220 1748 8248 4655
rect 8404 3942 8432 5646
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8588 5030 8616 5306
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8680 4826 8708 5102
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8404 3652 8432 3878
rect 8496 3738 8524 4014
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8312 3624 8432 3652
rect 8312 3466 8340 3624
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8588 2145 8616 2994
rect 8680 2854 8708 3470
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8574 2136 8630 2145
rect 8680 2106 8708 2790
rect 8772 2774 8800 12174
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8864 10810 8892 11154
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 10198 8892 10542
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8956 10112 8984 10610
rect 9036 10124 9088 10130
rect 8956 10084 9036 10112
rect 9036 10066 9088 10072
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8864 9450 8892 9862
rect 9048 9761 9076 10066
rect 9034 9752 9090 9761
rect 9034 9687 9090 9696
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8956 9178 8984 9454
rect 9140 9178 9168 13806
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 12170 9352 13262
rect 9508 12889 9536 14826
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9494 12880 9550 12889
rect 9494 12815 9550 12824
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11218 9444 12038
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9232 11014 9260 11154
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10538 9260 10950
rect 9508 10810 9536 12582
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9232 9994 9260 10474
rect 9416 10441 9444 10474
rect 9402 10432 9458 10441
rect 9402 10367 9458 10376
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9324 8838 9352 9998
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9140 7993 9168 8366
rect 9312 8356 9364 8362
rect 9416 8344 9444 8978
rect 9364 8316 9444 8344
rect 9494 8392 9550 8401
rect 9494 8327 9550 8336
rect 9312 8298 9364 8304
rect 9126 7984 9182 7993
rect 9324 7954 9352 8298
rect 9126 7919 9182 7928
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 4146 8892 7822
rect 9508 7698 9536 8327
rect 9416 7670 9536 7698
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 9048 6390 9076 6870
rect 9416 6798 9444 7670
rect 9600 7528 9628 13262
rect 9692 12753 9720 14826
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 10060 14074 10088 14282
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10152 13954 10180 14894
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 10364 14716 10740 14725
rect 10420 14714 10444 14716
rect 10500 14714 10524 14716
rect 10580 14714 10604 14716
rect 10660 14714 10684 14716
rect 10420 14662 10430 14714
rect 10674 14662 10684 14714
rect 10420 14660 10444 14662
rect 10500 14660 10524 14662
rect 10580 14660 10604 14662
rect 10660 14660 10684 14662
rect 10364 14651 10740 14660
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10060 13926 10180 13954
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 13190 9996 13670
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9864 12776 9916 12782
rect 9678 12744 9734 12753
rect 9864 12718 9916 12724
rect 9678 12679 9734 12688
rect 9692 9518 9720 12679
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 12073 9812 12174
rect 9770 12064 9826 12073
rect 9770 11999 9826 12008
rect 9784 9926 9812 11999
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9692 8498 9720 9046
rect 9784 8906 9812 9318
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9876 8809 9904 12718
rect 9968 11286 9996 13126
rect 10060 12986 10088 13926
rect 10244 13462 10272 14418
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10520 13841 10548 13942
rect 10506 13832 10562 13841
rect 10506 13767 10562 13776
rect 10704 13716 10732 14554
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 10796 13870 10824 14214
rect 10888 14074 10916 14214
rect 11348 14074 11376 14214
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11900 14006 11928 14758
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10968 13728 11020 13734
rect 10704 13688 10824 13716
rect 10364 13628 10740 13637
rect 10420 13626 10444 13628
rect 10500 13626 10524 13628
rect 10580 13626 10604 13628
rect 10660 13626 10684 13628
rect 10420 13574 10430 13626
rect 10674 13574 10684 13626
rect 10420 13572 10444 13574
rect 10500 13572 10524 13574
rect 10580 13572 10604 13574
rect 10660 13572 10684 13574
rect 10364 13563 10740 13572
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10796 13394 10824 13688
rect 10968 13670 11020 13676
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9968 10674 9996 11222
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9968 10130 9996 10610
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9862 8800 9918 8809
rect 9862 8735 9918 8744
rect 9968 8650 9996 9862
rect 9784 8622 9996 8650
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9508 7500 9628 7528
rect 9404 6792 9456 6798
rect 9324 6752 9404 6780
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 9324 5778 9352 6752
rect 9404 6734 9456 6740
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9048 5574 9076 5714
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9232 5166 9260 5646
rect 9324 5370 9352 5714
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9416 5166 9444 6598
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9048 4146 9076 4966
rect 9416 4826 9444 5102
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 8864 3738 8892 4082
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 9048 3534 9076 3946
rect 9126 3768 9182 3777
rect 9126 3703 9182 3712
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9048 3126 9076 3470
rect 9140 3466 9168 3703
rect 9324 3602 9352 4082
rect 9508 3738 9536 7500
rect 9586 7440 9642 7449
rect 9586 7375 9642 7384
rect 9600 6866 9628 7375
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9678 6760 9734 6769
rect 9678 6695 9734 6704
rect 9586 6216 9642 6225
rect 9586 6151 9642 6160
rect 9600 5778 9628 6151
rect 9692 5914 9720 6695
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 3913 9628 4082
rect 9586 3904 9642 3913
rect 9586 3839 9642 3848
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9784 3618 9812 8622
rect 9956 8560 10008 8566
rect 9862 8528 9918 8537
rect 9956 8502 10008 8508
rect 9862 8463 9918 8472
rect 9876 4146 9904 8463
rect 9968 7342 9996 8502
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9968 5098 9996 6938
rect 10060 5409 10088 12922
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10152 12345 10180 12854
rect 10704 12850 10732 13126
rect 10888 12850 10916 13126
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10138 12336 10194 12345
rect 10244 12306 10272 12582
rect 10364 12540 10740 12549
rect 10420 12538 10444 12540
rect 10500 12538 10524 12540
rect 10580 12538 10604 12540
rect 10660 12538 10684 12540
rect 10420 12486 10430 12538
rect 10674 12486 10684 12538
rect 10420 12484 10444 12486
rect 10500 12484 10524 12486
rect 10580 12484 10604 12486
rect 10660 12484 10684 12486
rect 10364 12475 10740 12484
rect 10876 12368 10928 12374
rect 10980 12356 11008 13670
rect 11164 13394 11192 13942
rect 11428 13864 11480 13870
rect 11612 13864 11664 13870
rect 11480 13824 11612 13852
rect 11428 13806 11480 13812
rect 11612 13806 11664 13812
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11796 13320 11848 13326
rect 11794 13288 11796 13297
rect 11848 13288 11850 13297
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11520 13252 11572 13258
rect 11794 13223 11850 13232
rect 11520 13194 11572 13200
rect 11164 12753 11192 13194
rect 11532 12782 11560 13194
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11336 12776 11388 12782
rect 11150 12744 11206 12753
rect 11336 12718 11388 12724
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11150 12679 11206 12688
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11150 12608 11206 12617
rect 11150 12543 11206 12552
rect 10928 12328 11008 12356
rect 10876 12310 10928 12316
rect 10138 12271 10194 12280
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10140 12232 10192 12238
rect 10692 12232 10744 12238
rect 10140 12174 10192 12180
rect 10598 12200 10654 12209
rect 10152 5778 10180 12174
rect 10692 12174 10744 12180
rect 10598 12135 10654 12144
rect 10612 12102 10640 12135
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10704 11830 10732 12174
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10796 11744 10824 12038
rect 10888 11898 10916 12106
rect 10876 11892 10928 11898
rect 11164 11880 11192 12543
rect 11256 12102 11284 12650
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10876 11834 10928 11840
rect 10980 11852 11192 11880
rect 10980 11762 11008 11852
rect 10876 11756 10928 11762
rect 10796 11716 10876 11744
rect 10876 11698 10928 11704
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10244 11354 10272 11562
rect 10364 11452 10740 11461
rect 10420 11450 10444 11452
rect 10500 11450 10524 11452
rect 10580 11450 10604 11452
rect 10660 11450 10684 11452
rect 10420 11398 10430 11450
rect 10674 11398 10684 11450
rect 10420 11396 10444 11398
rect 10500 11396 10524 11398
rect 10580 11396 10604 11398
rect 10660 11396 10684 11398
rect 10364 11387 10740 11396
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10888 10810 10916 11154
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10364 10364 10740 10373
rect 10420 10362 10444 10364
rect 10500 10362 10524 10364
rect 10580 10362 10604 10364
rect 10660 10362 10684 10364
rect 10420 10310 10430 10362
rect 10674 10310 10684 10362
rect 10420 10308 10444 10310
rect 10500 10308 10524 10310
rect 10580 10308 10604 10310
rect 10660 10308 10684 10310
rect 10364 10299 10740 10308
rect 10980 10248 11008 11698
rect 11060 11688 11112 11694
rect 11112 11648 11192 11676
rect 11060 11630 11112 11636
rect 11164 11506 11192 11648
rect 11072 11478 11192 11506
rect 11072 11354 11100 11478
rect 11150 11384 11206 11393
rect 11060 11348 11112 11354
rect 11150 11319 11206 11328
rect 11244 11348 11296 11354
rect 11060 11290 11112 11296
rect 11164 11150 11192 11319
rect 11244 11290 11296 11296
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11256 11082 11284 11290
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11072 10742 11100 11018
rect 11348 10810 11376 12718
rect 11624 12442 11652 12718
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11518 12336 11574 12345
rect 11518 12271 11574 12280
rect 11532 12238 11560 12271
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11440 11762 11468 12106
rect 11532 11830 11560 12174
rect 11610 12064 11666 12073
rect 11716 12050 11744 12718
rect 11666 12022 11744 12050
rect 11610 11999 11666 12008
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11440 11064 11468 11698
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11612 11076 11664 11082
rect 11440 11036 11612 11064
rect 11612 11018 11664 11024
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11072 10266 11100 10678
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11428 10600 11480 10606
rect 11480 10560 11560 10588
rect 11428 10542 11480 10548
rect 10704 10220 11008 10248
rect 11060 10260 11112 10266
rect 10232 9512 10284 9518
rect 10704 9489 10732 10220
rect 11060 10202 11112 10208
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10232 9454 10284 9460
rect 10690 9480 10746 9489
rect 10244 9160 10272 9454
rect 10690 9415 10746 9424
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10364 9276 10740 9285
rect 10420 9274 10444 9276
rect 10500 9274 10524 9276
rect 10580 9274 10604 9276
rect 10660 9274 10684 9276
rect 10420 9222 10430 9274
rect 10674 9222 10684 9274
rect 10420 9220 10444 9222
rect 10500 9220 10524 9222
rect 10580 9220 10604 9222
rect 10660 9220 10684 9222
rect 10364 9211 10740 9220
rect 10796 9178 10824 9386
rect 10324 9172 10376 9178
rect 10244 9132 10324 9160
rect 10324 9114 10376 9120
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10230 8936 10286 8945
rect 10230 8871 10232 8880
rect 10284 8871 10286 8880
rect 10232 8842 10284 8848
rect 10336 8276 10364 9114
rect 10888 8634 10916 9862
rect 10980 9382 11008 10066
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9042 11008 9318
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10244 8248 10364 8276
rect 10244 7954 10272 8248
rect 10364 8188 10740 8197
rect 10420 8186 10444 8188
rect 10500 8186 10524 8188
rect 10580 8186 10604 8188
rect 10660 8186 10684 8188
rect 10420 8134 10430 8186
rect 10674 8134 10684 8186
rect 10420 8132 10444 8134
rect 10500 8132 10524 8134
rect 10580 8132 10604 8134
rect 10660 8132 10684 8134
rect 10364 8123 10740 8132
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10230 7576 10286 7585
rect 10230 7511 10286 7520
rect 10244 7274 10272 7511
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10692 7336 10744 7342
rect 10744 7296 10824 7324
rect 10692 7278 10744 7284
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10244 7002 10272 7210
rect 10364 7100 10740 7109
rect 10420 7098 10444 7100
rect 10500 7098 10524 7100
rect 10580 7098 10604 7100
rect 10660 7098 10684 7100
rect 10420 7046 10430 7098
rect 10674 7046 10684 7098
rect 10420 7044 10444 7046
rect 10500 7044 10524 7046
rect 10580 7044 10604 7046
rect 10660 7044 10684 7046
rect 10364 7035 10740 7044
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10692 6928 10744 6934
rect 10796 6916 10824 7296
rect 10744 6888 10824 6916
rect 10692 6870 10744 6876
rect 10888 6730 10916 7414
rect 10980 7342 11008 8978
rect 11072 8566 11100 9998
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 7342 11100 8298
rect 11164 7954 11192 10542
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11348 10130 11376 10406
rect 11440 10266 11468 10406
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11256 9042 11284 10066
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11348 8430 11376 9318
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11164 7342 11192 7754
rect 11256 7342 11284 7890
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10600 6656 10652 6662
rect 10506 6624 10562 6633
rect 10600 6598 10652 6604
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10506 6559 10562 6568
rect 10520 6458 10548 6559
rect 10612 6458 10640 6598
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10612 6254 10640 6394
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10046 5400 10102 5409
rect 10046 5335 10102 5344
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 10244 4162 10272 6054
rect 10364 6012 10740 6021
rect 10420 6010 10444 6012
rect 10500 6010 10524 6012
rect 10580 6010 10604 6012
rect 10660 6010 10684 6012
rect 10420 5958 10430 6010
rect 10674 5958 10684 6010
rect 10420 5956 10444 5958
rect 10500 5956 10524 5958
rect 10580 5956 10604 5958
rect 10660 5956 10684 5958
rect 10364 5947 10740 5956
rect 10796 5658 10824 6598
rect 10874 6352 10930 6361
rect 10874 6287 10876 6296
rect 10928 6287 10930 6296
rect 10876 6258 10928 6264
rect 10874 6080 10930 6089
rect 10874 6015 10930 6024
rect 10888 5778 10916 6015
rect 10980 5778 11008 7278
rect 11152 6996 11204 7002
rect 11256 6984 11284 7278
rect 11348 7206 11376 8366
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11204 6956 11284 6984
rect 11336 6996 11388 7002
rect 11152 6938 11204 6944
rect 11336 6938 11388 6944
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10796 5630 11008 5658
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10364 4924 10740 4933
rect 10420 4922 10444 4924
rect 10500 4922 10524 4924
rect 10580 4922 10604 4924
rect 10660 4922 10684 4924
rect 10420 4870 10430 4922
rect 10674 4870 10684 4922
rect 10420 4868 10444 4870
rect 10500 4868 10524 4870
rect 10580 4868 10604 4870
rect 10660 4868 10684 4870
rect 10364 4859 10740 4868
rect 10796 4690 10824 5510
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10508 4616 10560 4622
rect 10506 4584 10508 4593
rect 10560 4584 10562 4593
rect 10506 4519 10562 4528
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10152 4134 10272 4162
rect 10046 3768 10102 3777
rect 10046 3703 10048 3712
rect 10100 3703 10102 3712
rect 10048 3674 10100 3680
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9600 3590 9812 3618
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 9036 3120 9088 3126
rect 8956 3080 9036 3108
rect 8772 2746 8892 2774
rect 8760 2304 8812 2310
rect 8758 2272 8760 2281
rect 8812 2272 8814 2281
rect 8758 2207 8814 2216
rect 8574 2071 8630 2080
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 8300 1896 8352 1902
rect 8300 1838 8352 1844
rect 8168 1720 8248 1748
rect 8116 1702 8168 1708
rect 7840 1556 7892 1562
rect 7840 1498 7892 1504
rect 7564 1352 7616 1358
rect 7564 1294 7616 1300
rect 7656 1352 7708 1358
rect 7656 1294 7708 1300
rect 8208 1284 8260 1290
rect 8208 1226 8260 1232
rect 7364 1116 7740 1125
rect 7420 1114 7444 1116
rect 7500 1114 7524 1116
rect 7580 1114 7604 1116
rect 7660 1114 7684 1116
rect 7420 1062 7430 1114
rect 7674 1062 7684 1114
rect 7420 1060 7444 1062
rect 7500 1060 7524 1062
rect 7580 1060 7604 1062
rect 7660 1060 7684 1062
rect 7364 1051 7740 1060
rect 8220 950 8248 1226
rect 8312 1222 8340 1838
rect 8392 1828 8444 1834
rect 8392 1770 8444 1776
rect 8404 1426 8432 1770
rect 8760 1760 8812 1766
rect 8760 1702 8812 1708
rect 8574 1456 8630 1465
rect 8392 1420 8444 1426
rect 8574 1391 8576 1400
rect 8392 1362 8444 1368
rect 8628 1391 8630 1400
rect 8576 1362 8628 1368
rect 8772 1222 8800 1702
rect 8300 1216 8352 1222
rect 8300 1158 8352 1164
rect 8392 1216 8444 1222
rect 8392 1158 8444 1164
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8404 950 8432 1158
rect 8208 944 8260 950
rect 8208 886 8260 892
rect 8392 944 8444 950
rect 8392 886 8444 892
rect 8864 814 8892 2746
rect 8956 2650 8984 3080
rect 9036 3062 9088 3068
rect 9140 3058 9168 3402
rect 9496 3392 9548 3398
rect 9600 3369 9628 3590
rect 10152 3516 10180 4134
rect 10364 3836 10740 3845
rect 10420 3834 10444 3836
rect 10500 3834 10524 3836
rect 10580 3834 10604 3836
rect 10660 3834 10684 3836
rect 10420 3782 10430 3834
rect 10674 3782 10684 3834
rect 10420 3780 10444 3782
rect 10500 3780 10524 3782
rect 10580 3780 10604 3782
rect 10660 3780 10684 3782
rect 10364 3771 10740 3780
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10152 3488 10364 3516
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9496 3334 9548 3340
rect 9586 3360 9642 3369
rect 9508 3233 9536 3334
rect 9586 3295 9642 3304
rect 9494 3224 9550 3233
rect 9494 3159 9550 3168
rect 9784 3126 9812 3402
rect 9954 3224 10010 3233
rect 10336 3210 10364 3488
rect 10428 3233 10456 3606
rect 10612 3602 10640 3674
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10010 3182 10088 3210
rect 9954 3159 10010 3168
rect 9496 3120 9548 3126
rect 9772 3120 9824 3126
rect 9678 3088 9734 3097
rect 9548 3068 9678 3074
rect 9496 3062 9678 3068
rect 9128 3052 9180 3058
rect 9508 3046 9678 3062
rect 10060 3074 10088 3182
rect 9772 3062 9824 3068
rect 9678 3023 9734 3032
rect 9128 2994 9180 3000
rect 9784 2990 9812 3062
rect 9968 3046 10088 3074
rect 10152 3182 10364 3210
rect 10414 3224 10470 3233
rect 9680 2984 9732 2990
rect 9600 2944 9680 2972
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9310 2816 9366 2825
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 9048 2564 9076 2790
rect 9600 2802 9628 2944
rect 9680 2926 9732 2932
rect 9772 2984 9824 2990
rect 9824 2932 9904 2938
rect 9772 2926 9904 2932
rect 9784 2910 9904 2926
rect 9772 2848 9824 2854
rect 9366 2774 9628 2802
rect 9770 2816 9772 2825
rect 9824 2816 9826 2825
rect 9310 2751 9366 2760
rect 9770 2751 9826 2760
rect 9494 2680 9550 2689
rect 9494 2615 9550 2624
rect 9770 2680 9826 2689
rect 9770 2615 9826 2624
rect 9220 2576 9272 2582
rect 9048 2536 9220 2564
rect 9220 2518 9272 2524
rect 9508 2446 9536 2615
rect 9784 2514 9812 2615
rect 9876 2582 9904 2910
rect 9968 2650 9996 3046
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10060 2689 10088 2926
rect 10046 2680 10102 2689
rect 9956 2644 10008 2650
rect 10046 2615 10102 2624
rect 9956 2586 10008 2592
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9496 2440 9548 2446
rect 9402 2408 9458 2417
rect 9036 2372 9088 2378
rect 9496 2382 9548 2388
rect 9402 2343 9458 2352
rect 9772 2372 9824 2378
rect 9036 2314 9088 2320
rect 9048 1562 9076 2314
rect 9128 2100 9180 2106
rect 9128 2042 9180 2048
rect 9140 2009 9168 2042
rect 9126 2000 9182 2009
rect 9126 1935 9182 1944
rect 9036 1556 9088 1562
rect 9036 1498 9088 1504
rect 9416 1426 9444 2343
rect 9772 2314 9824 2320
rect 9494 1728 9550 1737
rect 9494 1663 9550 1672
rect 9508 1426 9536 1663
rect 9404 1420 9456 1426
rect 9404 1362 9456 1368
rect 9496 1420 9548 1426
rect 9496 1362 9548 1368
rect 6184 808 6236 814
rect 6184 750 6236 756
rect 8852 808 8904 814
rect 8852 750 8904 756
rect 6000 672 6052 678
rect 5828 632 6000 660
rect 5448 400 5500 406
rect 5828 400 5856 632
rect 6000 614 6052 620
rect 4068 264 4120 270
rect 4068 206 4120 212
rect 4158 0 4214 400
rect 4986 0 5042 400
rect 5448 342 5500 348
rect 5814 0 5870 400
rect 6196 338 6224 750
rect 8484 672 8536 678
rect 8312 632 8484 660
rect 8312 400 8340 632
rect 8484 614 8536 620
rect 9128 672 9180 678
rect 9128 614 9180 620
rect 9140 400 9168 614
rect 6184 332 6236 338
rect 6184 274 6236 280
rect 8298 0 8354 400
rect 9126 0 9182 400
rect 9508 202 9536 1362
rect 9784 1358 9812 2314
rect 10060 2106 10088 2518
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 9876 1562 9904 1906
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 10152 1426 10180 3182
rect 10414 3159 10470 3168
rect 10520 3126 10548 3470
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10244 2650 10272 2926
rect 10612 2922 10640 3334
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10364 2748 10740 2757
rect 10420 2746 10444 2748
rect 10500 2746 10524 2748
rect 10580 2746 10604 2748
rect 10660 2746 10684 2748
rect 10420 2694 10430 2746
rect 10674 2694 10684 2746
rect 10420 2692 10444 2694
rect 10500 2692 10524 2694
rect 10580 2692 10604 2694
rect 10660 2692 10684 2694
rect 10364 2683 10740 2692
rect 10796 2650 10824 4626
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10888 3602 10916 3946
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10244 1970 10272 2586
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10336 1970 10364 2382
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 10324 1964 10376 1970
rect 10324 1906 10376 1912
rect 10796 1902 10824 2314
rect 10874 2000 10930 2009
rect 10874 1935 10930 1944
rect 10784 1896 10836 1902
rect 10244 1822 10364 1850
rect 10784 1838 10836 1844
rect 10140 1420 10192 1426
rect 10140 1362 10192 1368
rect 9772 1352 9824 1358
rect 9772 1294 9824 1300
rect 9772 1216 9824 1222
rect 9772 1158 9824 1164
rect 9784 1018 9812 1158
rect 9772 1012 9824 1018
rect 9772 954 9824 960
rect 9770 912 9826 921
rect 9770 847 9826 856
rect 9784 814 9812 847
rect 9772 808 9824 814
rect 9772 750 9824 756
rect 9956 672 10008 678
rect 9956 614 10008 620
rect 9968 400 9996 614
rect 9496 196 9548 202
rect 9496 138 9548 144
rect 9954 0 10010 400
rect 10244 270 10272 1822
rect 10336 1766 10364 1822
rect 10324 1760 10376 1766
rect 10324 1702 10376 1708
rect 10364 1660 10740 1669
rect 10420 1658 10444 1660
rect 10500 1658 10524 1660
rect 10580 1658 10604 1660
rect 10660 1658 10684 1660
rect 10420 1606 10430 1658
rect 10674 1606 10684 1658
rect 10420 1604 10444 1606
rect 10500 1604 10524 1606
rect 10580 1604 10604 1606
rect 10660 1604 10684 1606
rect 10364 1595 10740 1604
rect 10888 1562 10916 1935
rect 10876 1556 10928 1562
rect 10876 1498 10928 1504
rect 10980 1426 11008 5630
rect 11072 5370 11100 6802
rect 11164 5642 11192 6938
rect 11348 6866 11376 6938
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11164 5166 11192 5306
rect 11152 5160 11204 5166
rect 11058 5128 11114 5137
rect 11152 5102 11204 5108
rect 11058 5063 11114 5072
rect 11072 3466 11100 5063
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11058 3360 11114 3369
rect 11058 3295 11114 3304
rect 11072 3074 11100 3295
rect 11072 3046 11192 3074
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11072 2582 11100 2790
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11164 2446 11192 3046
rect 11152 2440 11204 2446
rect 11072 2400 11152 2428
rect 11072 1970 11100 2400
rect 11152 2382 11204 2388
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11164 2106 11192 2246
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11060 1964 11112 1970
rect 11060 1906 11112 1912
rect 11256 1902 11284 6598
rect 11440 6322 11468 8774
rect 11532 8566 11560 10560
rect 11610 10296 11666 10305
rect 11716 10266 11744 11630
rect 11900 11558 11928 12786
rect 11992 12646 12020 14826
rect 13280 14278 13308 14894
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13280 13870 13308 14214
rect 13364 14172 13740 14181
rect 13420 14170 13444 14172
rect 13500 14170 13524 14172
rect 13580 14170 13604 14172
rect 13660 14170 13684 14172
rect 13420 14118 13430 14170
rect 13674 14118 13684 14170
rect 13420 14116 13444 14118
rect 13500 14116 13524 14118
rect 13580 14116 13604 14118
rect 13660 14116 13684 14118
rect 13364 14107 13740 14116
rect 13832 13977 13860 14758
rect 14752 14618 14780 15302
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14568 14074 14596 14418
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14188 14000 14240 14006
rect 13818 13968 13874 13977
rect 14188 13942 14240 13948
rect 13818 13903 13874 13912
rect 13832 13870 13860 13903
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 12084 11558 12112 13398
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12176 11830 12204 12106
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11610 10231 11666 10240
rect 11704 10260 11756 10266
rect 11624 9722 11652 10231
rect 11704 10202 11756 10208
rect 11808 9994 11836 10542
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11794 9072 11850 9081
rect 11794 9007 11796 9016
rect 11848 9007 11850 9016
rect 11796 8978 11848 8984
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11532 8022 11560 8366
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11624 7818 11652 8910
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8634 11836 8774
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11900 8514 11928 11086
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 11992 9042 12020 9658
rect 12176 9586 12204 10542
rect 12268 10441 12296 12038
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12254 10432 12310 10441
rect 12254 10367 12310 10376
rect 12452 9586 12480 10542
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11808 8486 11928 8514
rect 11992 8498 12020 8978
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11980 8492 12032 8498
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11716 7342 11744 8230
rect 11808 7342 11836 8486
rect 11980 8434 12032 8440
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11900 8090 11928 8366
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11900 7342 11928 7414
rect 11704 7336 11756 7342
rect 11796 7336 11848 7342
rect 11704 7278 11756 7284
rect 11794 7304 11796 7313
rect 11888 7336 11940 7342
rect 11848 7304 11850 7313
rect 11888 7278 11940 7284
rect 11794 7239 11850 7248
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11532 7041 11560 7142
rect 11518 7032 11574 7041
rect 11518 6967 11574 6976
rect 11518 6896 11574 6905
rect 11624 6866 11652 7142
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11518 6831 11574 6840
rect 11612 6860 11664 6866
rect 11532 6390 11560 6831
rect 11612 6802 11664 6808
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11348 5953 11376 6122
rect 11334 5944 11390 5953
rect 11334 5879 11390 5888
rect 11532 5846 11560 6190
rect 11624 5914 11652 6190
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11716 5370 11744 6938
rect 11808 5778 11836 7239
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11900 6866 11928 6967
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11900 6322 11928 6598
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11900 5828 11928 6258
rect 11992 6236 12020 7686
rect 12084 7002 12112 8910
rect 12176 7585 12204 9522
rect 12346 9344 12402 9353
rect 12346 9279 12402 9288
rect 12360 9110 12388 9279
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12452 9042 12480 9522
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12268 8894 12480 8922
rect 12268 8838 12296 8894
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12162 7576 12218 7585
rect 12162 7511 12218 7520
rect 12268 7290 12296 8570
rect 12360 7954 12388 8774
rect 12452 8265 12480 8894
rect 12544 8498 12572 11290
rect 12636 10810 12664 12174
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12532 8288 12584 8294
rect 12438 8256 12494 8265
rect 12532 8230 12584 8236
rect 12438 8191 12494 8200
rect 12544 8129 12572 8230
rect 12530 8120 12586 8129
rect 12440 8084 12492 8090
rect 12530 8055 12586 8064
rect 12440 8026 12492 8032
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12452 7410 12480 8026
rect 12544 8022 12572 8055
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12544 7410 12572 7958
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12268 7262 12480 7290
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 7041 12204 7142
rect 12162 7032 12218 7041
rect 12072 6996 12124 7002
rect 12162 6967 12218 6976
rect 12348 6996 12400 7002
rect 12072 6938 12124 6944
rect 12348 6938 12400 6944
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12084 6458 12112 6734
rect 12162 6624 12218 6633
rect 12162 6559 12218 6568
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 11992 6208 12112 6236
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 12084 6066 12112 6208
rect 12176 6186 12204 6559
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12256 6112 12308 6118
rect 11992 5953 12020 6054
rect 12084 6038 12204 6066
rect 12256 6054 12308 6060
rect 11978 5944 12034 5953
rect 11978 5879 12034 5888
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11980 5840 12032 5846
rect 11900 5800 11980 5828
rect 11980 5782 12032 5788
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11336 5296 11388 5302
rect 11808 5250 11836 5306
rect 11336 5238 11388 5244
rect 11348 5001 11376 5238
rect 11716 5234 11836 5250
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11704 5228 11836 5234
rect 11756 5222 11836 5228
rect 11704 5170 11756 5176
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11334 4992 11390 5001
rect 11334 4927 11390 4936
rect 11440 3942 11468 5102
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3670 11468 3878
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11532 2774 11560 4966
rect 11624 4282 11652 5034
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4690 11744 4966
rect 11900 4690 11928 5238
rect 11992 5166 12020 5782
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11808 3738 11836 4558
rect 11992 4554 12020 5102
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11808 3097 11836 3334
rect 11794 3088 11850 3097
rect 11794 3023 11850 3032
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11440 2746 11560 2774
rect 11334 2408 11390 2417
rect 11334 2343 11390 2352
rect 11348 1902 11376 2343
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 11336 1896 11388 1902
rect 11336 1838 11388 1844
rect 11060 1760 11112 1766
rect 11060 1702 11112 1708
rect 10968 1420 11020 1426
rect 10968 1362 11020 1368
rect 10508 1352 10560 1358
rect 10560 1312 10732 1340
rect 10508 1294 10560 1300
rect 10704 1306 10732 1312
rect 11072 1306 11100 1702
rect 11164 1562 11192 1838
rect 11152 1556 11204 1562
rect 11152 1498 11204 1504
rect 10704 1278 11100 1306
rect 11348 1290 11376 1838
rect 11440 1426 11468 2746
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11520 2304 11572 2310
rect 11716 2281 11744 2586
rect 11520 2246 11572 2252
rect 11702 2272 11758 2281
rect 11532 1902 11560 2246
rect 11702 2207 11758 2216
rect 11808 2145 11836 2790
rect 11794 2136 11850 2145
rect 11794 2071 11850 2080
rect 11520 1896 11572 1902
rect 11520 1838 11572 1844
rect 11612 1828 11664 1834
rect 11612 1770 11664 1776
rect 11518 1456 11574 1465
rect 11428 1420 11480 1426
rect 11624 1426 11652 1770
rect 11518 1391 11574 1400
rect 11612 1420 11664 1426
rect 11428 1362 11480 1368
rect 11336 1284 11388 1290
rect 11336 1226 11388 1232
rect 10784 1216 10836 1222
rect 10784 1158 10836 1164
rect 10796 1018 10824 1158
rect 10784 1012 10836 1018
rect 10784 954 10836 960
rect 11532 814 11560 1391
rect 11612 1362 11664 1368
rect 11612 1216 11664 1222
rect 11612 1158 11664 1164
rect 11624 882 11652 1158
rect 12084 1018 12112 5850
rect 12176 5166 12204 6038
rect 12268 5914 12296 6054
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12360 5794 12388 6938
rect 12268 5766 12388 5794
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12176 2774 12204 4966
rect 12268 2836 12296 5766
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12360 4826 12388 5646
rect 12452 5166 12480 7262
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12544 6905 12572 7210
rect 12636 6934 12664 10134
rect 12728 10062 12756 13126
rect 13004 12986 13032 13806
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12900 12912 12952 12918
rect 12898 12880 12900 12889
rect 12952 12880 12954 12889
rect 12898 12815 12954 12824
rect 13096 12782 13124 13466
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12808 12232 12860 12238
rect 12860 12180 12940 12186
rect 12808 12174 12940 12180
rect 12820 12158 12940 12174
rect 12912 11626 12940 12158
rect 13004 11801 13032 12242
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 12990 11792 13046 11801
rect 12990 11727 13046 11736
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12820 10674 12848 11154
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12912 9674 12940 11562
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13004 10130 13032 10542
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12728 9646 12940 9674
rect 12728 9353 12756 9646
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12714 9344 12770 9353
rect 12714 9279 12770 9288
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12728 8072 12756 8978
rect 12820 8294 12848 8978
rect 12912 8634 12940 9522
rect 13004 9110 13032 10066
rect 13096 9586 13124 12106
rect 13188 11218 13216 13806
rect 13364 13084 13740 13093
rect 13420 13082 13444 13084
rect 13500 13082 13524 13084
rect 13580 13082 13604 13084
rect 13660 13082 13684 13084
rect 13420 13030 13430 13082
rect 13674 13030 13684 13082
rect 13420 13028 13444 13030
rect 13500 13028 13524 13030
rect 13580 13028 13604 13030
rect 13660 13028 13684 13030
rect 13364 13019 13740 13028
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13726 12608 13782 12617
rect 13726 12543 13782 12552
rect 13740 12306 13768 12543
rect 13832 12442 13860 12786
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13280 11898 13308 12038
rect 13364 11996 13740 12005
rect 13420 11994 13444 11996
rect 13500 11994 13524 11996
rect 13580 11994 13604 11996
rect 13660 11994 13684 11996
rect 13420 11942 13430 11994
rect 13674 11942 13684 11994
rect 13420 11940 13444 11942
rect 13500 11940 13524 11942
rect 13580 11940 13604 11942
rect 13660 11940 13684 11942
rect 13364 11931 13740 11940
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13728 11688 13780 11694
rect 13832 11642 13860 12038
rect 13780 11636 13860 11642
rect 13728 11630 13860 11636
rect 13636 11620 13688 11626
rect 13740 11614 13860 11630
rect 13636 11562 13688 11568
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13648 11150 13676 11562
rect 13924 11393 13952 12718
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14108 11898 14136 12310
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13910 11384 13966 11393
rect 13910 11319 13966 11328
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13636 11144 13688 11150
rect 13832 11121 13860 11222
rect 13912 11212 13964 11218
rect 14016 11200 14044 11494
rect 14108 11354 14136 11630
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14096 11212 14148 11218
rect 14016 11172 14096 11200
rect 13912 11154 13964 11160
rect 14096 11154 14148 11160
rect 13636 11086 13688 11092
rect 13818 11112 13874 11121
rect 13268 11076 13320 11082
rect 13818 11047 13874 11056
rect 13268 11018 13320 11024
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13188 10606 13216 10746
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13188 10305 13216 10406
rect 13174 10296 13230 10305
rect 13174 10231 13230 10240
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13188 9586 13216 10066
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13096 9042 13124 9386
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13188 8498 13216 8774
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12728 8044 12848 8072
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12624 6928 12676 6934
rect 12530 6896 12586 6905
rect 12624 6870 12676 6876
rect 12530 6831 12586 6840
rect 12728 6798 12756 7890
rect 12820 7546 12848 8044
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12544 5914 12572 6054
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12728 5778 12756 6734
rect 12820 6458 12848 7278
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12820 5914 12848 6122
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12806 5672 12862 5681
rect 12806 5607 12862 5616
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12544 5166 12572 5510
rect 12820 5250 12848 5607
rect 12636 5222 12848 5250
rect 12636 5166 12664 5222
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12360 3602 12388 4422
rect 12452 4078 12480 5102
rect 12544 4146 12572 5102
rect 12820 4826 12848 5102
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12820 4078 12848 4558
rect 12912 4486 12940 8298
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13096 7460 13124 8230
rect 13188 7886 13216 8230
rect 13280 7954 13308 11018
rect 13364 10908 13740 10917
rect 13420 10906 13444 10908
rect 13500 10906 13524 10908
rect 13580 10906 13604 10908
rect 13660 10906 13684 10908
rect 13420 10854 13430 10906
rect 13674 10854 13684 10906
rect 13420 10852 13444 10854
rect 13500 10852 13524 10854
rect 13580 10852 13604 10854
rect 13660 10852 13684 10854
rect 13364 10843 13740 10852
rect 13832 10674 13860 11047
rect 13924 10742 13952 11154
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14200 10606 14228 13942
rect 14648 13864 14700 13870
rect 14646 13832 14648 13841
rect 14700 13832 14702 13841
rect 14646 13767 14702 13776
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14476 12782 14504 13126
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14292 12442 14320 12718
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14292 11354 14320 11562
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 13740 10266 13768 10542
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13364 9820 13740 9829
rect 13420 9818 13444 9820
rect 13500 9818 13524 9820
rect 13580 9818 13604 9820
rect 13660 9818 13684 9820
rect 13420 9766 13430 9818
rect 13674 9766 13684 9818
rect 13420 9764 13444 9766
rect 13500 9764 13524 9766
rect 13580 9764 13604 9766
rect 13660 9764 13684 9766
rect 13364 9755 13740 9764
rect 13832 9674 13860 10474
rect 13924 9926 13952 10542
rect 14108 10266 14136 10542
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13372 9646 13860 9674
rect 13372 9217 13400 9646
rect 13924 9602 13952 9862
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13832 9574 13952 9602
rect 14016 9586 14044 10066
rect 14200 9738 14228 10542
rect 14292 10130 14320 11290
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14200 9710 14320 9738
rect 14004 9580 14056 9586
rect 13358 9208 13414 9217
rect 13464 9178 13492 9522
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 9178 13768 9454
rect 13358 9143 13414 9152
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13634 9072 13690 9081
rect 13634 9007 13636 9016
rect 13688 9007 13690 9016
rect 13636 8978 13688 8984
rect 13648 8820 13676 8978
rect 13832 8888 13860 9574
rect 14004 9522 14056 9528
rect 14016 9058 14044 9522
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 13924 9042 14044 9058
rect 13912 9036 14044 9042
rect 13964 9030 14044 9036
rect 13912 8978 13964 8984
rect 13912 8900 13964 8906
rect 13832 8860 13912 8888
rect 13912 8842 13964 8848
rect 13648 8792 13860 8820
rect 13364 8732 13740 8741
rect 13420 8730 13444 8732
rect 13500 8730 13524 8732
rect 13580 8730 13604 8732
rect 13660 8730 13684 8732
rect 13420 8678 13430 8730
rect 13674 8678 13684 8730
rect 13420 8676 13444 8678
rect 13500 8676 13524 8678
rect 13580 8676 13604 8678
rect 13660 8676 13684 8678
rect 13364 8667 13740 8676
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13176 7880 13228 7886
rect 13372 7834 13400 8434
rect 13728 8356 13780 8362
rect 13648 8316 13728 8344
rect 13648 7868 13676 8316
rect 13728 8298 13780 8304
rect 13832 8090 13860 8792
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13740 7993 13768 8026
rect 13726 7984 13782 7993
rect 13726 7919 13782 7928
rect 13648 7840 13860 7868
rect 13176 7822 13228 7828
rect 13004 7432 13124 7460
rect 13280 7806 13400 7834
rect 13004 7342 13032 7432
rect 13280 7410 13308 7806
rect 13364 7644 13740 7653
rect 13420 7642 13444 7644
rect 13500 7642 13524 7644
rect 13580 7642 13604 7644
rect 13660 7642 13684 7644
rect 13420 7590 13430 7642
rect 13674 7590 13684 7642
rect 13420 7588 13444 7590
rect 13500 7588 13524 7590
rect 13580 7588 13604 7590
rect 13660 7588 13684 7590
rect 13364 7579 13740 7588
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13188 7002 13216 7346
rect 13556 7342 13584 7482
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13464 7002 13492 7210
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13004 4865 13032 6054
rect 12990 4856 13046 4865
rect 12990 4791 13046 4800
rect 13096 4690 13124 6666
rect 13188 5778 13216 6938
rect 13452 6724 13504 6730
rect 13556 6712 13584 7278
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13648 6848 13676 7210
rect 13740 7206 13768 7482
rect 13832 7410 13860 7840
rect 13924 7410 13952 8842
rect 14016 8362 14044 9030
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 14002 8120 14058 8129
rect 14002 8055 14058 8064
rect 14016 7954 14044 8055
rect 14108 7954 14136 8434
rect 14200 8294 14228 9386
rect 14292 9042 14320 9710
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14200 7954 14228 8230
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 7834 14228 7890
rect 14108 7806 14228 7834
rect 14108 7800 14136 7806
rect 14016 7772 14136 7800
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 6860 13780 6866
rect 13648 6820 13728 6848
rect 13648 6769 13676 6820
rect 13728 6802 13780 6808
rect 13504 6684 13584 6712
rect 13634 6760 13690 6769
rect 13634 6695 13690 6704
rect 13452 6666 13504 6672
rect 13364 6556 13740 6565
rect 13420 6554 13444 6556
rect 13500 6554 13524 6556
rect 13580 6554 13604 6556
rect 13660 6554 13684 6556
rect 13420 6502 13430 6554
rect 13674 6502 13684 6554
rect 13420 6500 13444 6502
rect 13500 6500 13524 6502
rect 13580 6500 13604 6502
rect 13660 6500 13684 6502
rect 13364 6491 13740 6500
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13740 6100 13768 6326
rect 13832 6254 13860 7142
rect 14016 6866 14044 7772
rect 14186 7576 14242 7585
rect 14108 7534 14186 7562
rect 14108 6866 14136 7534
rect 14186 7511 14242 7520
rect 14188 7336 14240 7342
rect 14186 7304 14188 7313
rect 14240 7304 14242 7313
rect 14186 7239 14242 7248
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13924 6497 13952 6666
rect 13910 6488 13966 6497
rect 13910 6423 13966 6432
rect 13924 6254 13952 6423
rect 14108 6361 14136 6802
rect 14188 6384 14240 6390
rect 14094 6352 14150 6361
rect 14188 6326 14240 6332
rect 14094 6287 14150 6296
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13740 6072 13860 6100
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13280 5681 13308 5714
rect 13266 5672 13322 5681
rect 13266 5607 13322 5616
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 5137 13216 5510
rect 13364 5468 13740 5477
rect 13420 5466 13444 5468
rect 13500 5466 13524 5468
rect 13580 5466 13604 5468
rect 13660 5466 13684 5468
rect 13420 5414 13430 5466
rect 13674 5414 13684 5466
rect 13420 5412 13444 5414
rect 13500 5412 13524 5414
rect 13580 5412 13604 5414
rect 13660 5412 13684 5414
rect 13364 5403 13740 5412
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13636 5160 13688 5166
rect 13174 5128 13230 5137
rect 13636 5102 13688 5108
rect 13174 5063 13230 5072
rect 13176 5024 13228 5030
rect 13648 5001 13676 5102
rect 13176 4966 13228 4972
rect 13634 4992 13690 5001
rect 13084 4684 13136 4690
rect 13004 4644 13084 4672
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12440 4072 12492 4078
rect 12808 4072 12860 4078
rect 12440 4014 12492 4020
rect 12806 4040 12808 4049
rect 12900 4072 12952 4078
rect 12860 4040 12862 4049
rect 12900 4014 12952 4020
rect 12806 3975 12862 3984
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 2961 12388 3538
rect 12820 3398 12848 3975
rect 12912 3738 12940 4014
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 13004 3194 13032 4644
rect 13084 4626 13136 4632
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 13096 3398 13124 4490
rect 13188 4078 13216 4966
rect 13634 4927 13690 4936
rect 13740 4672 13768 5306
rect 13832 5166 13860 6072
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13924 4758 13952 5646
rect 14016 4758 14044 5782
rect 14200 5166 14228 6326
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 14004 4752 14056 4758
rect 14004 4694 14056 4700
rect 13820 4684 13872 4690
rect 13740 4644 13820 4672
rect 14188 4684 14240 4690
rect 13820 4626 13872 4632
rect 14108 4644 14188 4672
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13280 4078 13308 4422
rect 13364 4380 13740 4389
rect 13420 4378 13444 4380
rect 13500 4378 13524 4380
rect 13580 4378 13604 4380
rect 13660 4378 13684 4380
rect 13420 4326 13430 4378
rect 13674 4326 13684 4378
rect 13420 4324 13444 4326
rect 13500 4324 13524 4326
rect 13580 4324 13604 4326
rect 13660 4324 13684 4326
rect 13364 4315 13740 4324
rect 13832 4264 13860 4626
rect 13556 4236 13860 4264
rect 13452 4208 13504 4214
rect 13450 4176 13452 4185
rect 13504 4176 13506 4185
rect 13360 4140 13412 4146
rect 13450 4111 13506 4120
rect 13360 4082 13412 4088
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13188 3602 13216 4014
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13084 3392 13136 3398
rect 13372 3380 13400 4082
rect 13452 3664 13504 3670
rect 13556 3652 13584 4236
rect 14108 4196 14136 4644
rect 14188 4626 14240 4632
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13504 3624 13584 3652
rect 13648 4168 14136 4196
rect 13452 3606 13504 3612
rect 13648 3602 13676 4168
rect 14200 4078 14228 4422
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14200 3670 14228 4014
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13084 3334 13136 3340
rect 13280 3352 13400 3380
rect 12992 3188 13044 3194
rect 13044 3148 13216 3176
rect 12992 3130 13044 3136
rect 12900 2984 12952 2990
rect 12346 2952 12402 2961
rect 12900 2926 12952 2932
rect 12346 2887 12402 2896
rect 12348 2848 12400 2854
rect 12268 2808 12348 2836
rect 12348 2790 12400 2796
rect 12176 2746 12296 2774
rect 12268 1426 12296 2746
rect 12912 2650 12940 2926
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 12990 2680 13046 2689
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12900 2644 12952 2650
rect 12990 2615 13046 2624
rect 12900 2586 12952 2592
rect 12820 2378 12848 2586
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 13004 1970 13032 2615
rect 13096 2428 13124 2790
rect 13188 2582 13216 3148
rect 13280 3040 13308 3352
rect 13364 3292 13740 3301
rect 13420 3290 13444 3292
rect 13500 3290 13524 3292
rect 13580 3290 13604 3292
rect 13660 3290 13684 3292
rect 13420 3238 13430 3290
rect 13674 3238 13684 3290
rect 13420 3236 13444 3238
rect 13500 3236 13524 3238
rect 13580 3236 13604 3238
rect 13660 3236 13684 3238
rect 13364 3227 13740 3236
rect 13636 3052 13688 3058
rect 13280 3012 13636 3040
rect 13636 2994 13688 3000
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13544 2848 13596 2854
rect 13740 2836 13768 2994
rect 13832 2990 13860 3470
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13924 2836 13952 3538
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14016 2990 14044 3130
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13596 2808 13952 2836
rect 14096 2848 14148 2854
rect 13544 2790 13596 2796
rect 14096 2790 14148 2796
rect 13542 2680 13598 2689
rect 13542 2615 13598 2624
rect 13820 2644 13872 2650
rect 13556 2582 13584 2615
rect 13820 2586 13872 2592
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 13096 2400 13308 2428
rect 13280 2310 13308 2400
rect 13832 2378 13860 2586
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 12992 1964 13044 1970
rect 12992 1906 13044 1912
rect 13096 1902 13124 2246
rect 13084 1896 13136 1902
rect 13084 1838 13136 1844
rect 13280 1834 13308 2246
rect 13364 2204 13740 2213
rect 13420 2202 13444 2204
rect 13500 2202 13524 2204
rect 13580 2202 13604 2204
rect 13660 2202 13684 2204
rect 13420 2150 13430 2202
rect 13674 2150 13684 2202
rect 13420 2148 13444 2150
rect 13500 2148 13524 2150
rect 13580 2148 13604 2150
rect 13660 2148 13684 2150
rect 13364 2139 13740 2148
rect 13820 1964 13872 1970
rect 13820 1906 13872 1912
rect 13268 1828 13320 1834
rect 13268 1770 13320 1776
rect 13452 1760 13504 1766
rect 13452 1702 13504 1708
rect 13358 1592 13414 1601
rect 13268 1556 13320 1562
rect 13320 1536 13358 1544
rect 13320 1527 13414 1536
rect 13320 1516 13400 1527
rect 13268 1498 13320 1504
rect 12256 1420 12308 1426
rect 12256 1362 12308 1368
rect 13464 1358 13492 1702
rect 13544 1556 13596 1562
rect 13544 1498 13596 1504
rect 12716 1352 12768 1358
rect 12716 1294 12768 1300
rect 13452 1352 13504 1358
rect 13452 1294 13504 1300
rect 12624 1216 12676 1222
rect 12624 1158 12676 1164
rect 12636 1018 12664 1158
rect 12072 1012 12124 1018
rect 12072 954 12124 960
rect 12624 1012 12676 1018
rect 12624 954 12676 960
rect 11612 876 11664 882
rect 11612 818 11664 824
rect 11520 808 11572 814
rect 11520 750 11572 756
rect 11152 672 11204 678
rect 11152 614 11204 620
rect 11612 672 11664 678
rect 11612 614 11664 620
rect 12624 672 12676 678
rect 12624 614 12676 620
rect 10364 572 10740 581
rect 10420 570 10444 572
rect 10500 570 10524 572
rect 10580 570 10604 572
rect 10660 570 10684 572
rect 10420 518 10430 570
rect 10674 518 10684 570
rect 10420 516 10444 518
rect 10500 516 10524 518
rect 10580 516 10604 518
rect 10660 516 10684 518
rect 10364 507 10740 516
rect 10796 462 10916 490
rect 10796 400 10824 462
rect 10232 264 10284 270
rect 10232 206 10284 212
rect 10782 0 10838 400
rect 10888 354 10916 462
rect 11164 354 11192 614
rect 11624 400 11652 614
rect 12636 490 12664 614
rect 12452 462 12664 490
rect 12452 400 12480 462
rect 10888 326 11192 354
rect 11610 0 11666 400
rect 12438 0 12494 400
rect 12728 270 12756 1294
rect 12992 1216 13044 1222
rect 12992 1158 13044 1164
rect 13452 1216 13504 1222
rect 13556 1204 13584 1498
rect 13832 1426 13860 1906
rect 14004 1828 14056 1834
rect 14004 1770 14056 1776
rect 14016 1494 14044 1770
rect 14004 1488 14056 1494
rect 14004 1430 14056 1436
rect 14108 1426 14136 2790
rect 14292 2650 14320 8978
rect 14384 2774 14412 12718
rect 14648 12640 14700 12646
rect 14646 12608 14648 12617
rect 14700 12608 14702 12617
rect 14646 12543 14702 12552
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14476 10470 14504 11290
rect 14568 10606 14596 11494
rect 14660 11393 14688 11562
rect 14646 11384 14702 11393
rect 14646 11319 14702 11328
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14554 10432 14610 10441
rect 14476 10130 14504 10406
rect 14554 10367 14610 10376
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 8498 14504 8774
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14476 7410 14504 8298
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14476 6662 14504 7210
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 4146 14504 5510
rect 14568 5216 14596 10367
rect 14660 9926 14688 10542
rect 14752 10305 14780 12310
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14936 11354 14964 11630
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14738 10296 14794 10305
rect 14738 10231 14794 10240
rect 14752 10198 14780 10231
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9722 14780 9862
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 15028 9654 15056 11494
rect 15120 11150 15148 12038
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 14646 9072 14702 9081
rect 14646 9007 14702 9016
rect 14660 8974 14688 9007
rect 15028 8974 15056 9590
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14660 8566 14688 8910
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14844 8566 14872 8774
rect 14936 8566 14964 8842
rect 15028 8809 15056 8910
rect 15014 8800 15070 8809
rect 15014 8735 15070 8744
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14844 8090 14872 8502
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14648 7948 14700 7954
rect 14700 7908 14872 7936
rect 14648 7890 14700 7896
rect 14844 7585 14872 7908
rect 14830 7576 14886 7585
rect 14830 7511 14886 7520
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14660 6746 14688 7142
rect 14752 6866 14780 7414
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14660 6718 14780 6746
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 5710 14688 6598
rect 14752 6089 14780 6718
rect 14738 6080 14794 6089
rect 14738 6015 14794 6024
rect 14738 5808 14794 5817
rect 14738 5743 14794 5752
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14568 5188 14688 5216
rect 14556 5092 14608 5098
rect 14556 5034 14608 5040
rect 14568 4486 14596 5034
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 4282 14596 4422
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3602 14504 3878
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 3058 14504 3334
rect 14660 3097 14688 5188
rect 14752 4826 14780 5743
rect 14844 5370 14872 7414
rect 14936 6662 14964 8026
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 15028 6390 15056 8570
rect 15120 7478 15148 11086
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 15120 6254 15148 6598
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15028 5914 15056 6190
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14936 5710 14964 5850
rect 15028 5778 15056 5850
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 14924 5704 14976 5710
rect 15212 5658 15240 14350
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15396 13938 15424 14214
rect 15764 13938 15792 14554
rect 15842 14376 15898 14385
rect 15842 14311 15844 14320
rect 15896 14311 15898 14320
rect 15844 14282 15896 14288
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15396 11694 15424 13874
rect 15764 12442 15792 13874
rect 15856 13705 15884 13874
rect 16132 13870 16160 14214
rect 16224 14074 16252 15370
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16364 14716 16740 14725
rect 16420 14714 16444 14716
rect 16500 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16420 14662 16430 14714
rect 16674 14662 16684 14714
rect 16420 14660 16444 14662
rect 16500 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16364 14651 16740 14660
rect 16776 14498 16804 14962
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16316 14476 16804 14498
rect 16316 14470 16488 14476
rect 16316 14414 16344 14470
rect 16540 14470 16804 14476
rect 16488 14418 16540 14424
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16868 14074 16896 14894
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16764 13728 16816 13734
rect 15842 13696 15898 13705
rect 16764 13670 16816 13676
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 15842 13631 15898 13640
rect 16364 13628 16740 13637
rect 16420 13626 16444 13628
rect 16500 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16420 13574 16430 13626
rect 16674 13574 16684 13626
rect 16420 13572 16444 13574
rect 16500 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16364 13563 16740 13572
rect 16776 13326 16804 13670
rect 16868 13394 16896 13670
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 15948 12986 15976 13262
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16408 12918 16436 13194
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16868 12714 16896 13330
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16364 12540 16740 12549
rect 16420 12538 16444 12540
rect 16500 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16420 12486 16430 12538
rect 16674 12486 16684 12538
rect 16420 12484 16444 12486
rect 16500 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 15842 12472 15898 12481
rect 16364 12475 16740 12484
rect 15752 12436 15804 12442
rect 15842 12407 15898 12416
rect 15752 12378 15804 12384
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11286 15424 11630
rect 15384 11280 15436 11286
rect 15304 11240 15384 11268
rect 15304 10606 15332 11240
rect 15384 11222 15436 11228
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15396 10674 15424 11086
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15304 9042 15332 10202
rect 15396 9081 15424 10406
rect 15488 10044 15516 10950
rect 15856 10810 15884 12407
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15948 12102 15976 12310
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16026 11792 16082 11801
rect 16132 11762 16160 12038
rect 16224 11898 16252 12242
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16762 11792 16818 11801
rect 16026 11727 16082 11736
rect 16120 11756 16172 11762
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 16040 10130 16068 11727
rect 16762 11727 16818 11736
rect 16120 11698 16172 11704
rect 16132 11354 16160 11698
rect 16364 11452 16740 11461
rect 16420 11450 16444 11452
rect 16500 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16420 11398 16430 11450
rect 16674 11398 16684 11450
rect 16420 11396 16444 11398
rect 16500 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16364 11387 16740 11396
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16132 11218 16160 11290
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16408 10810 16436 11222
rect 16776 11218 16804 11727
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16854 10568 16910 10577
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 15568 10056 15620 10062
rect 15488 10016 15568 10044
rect 15568 9998 15620 10004
rect 15580 9518 15608 9998
rect 16132 9926 16160 10542
rect 16224 10062 16252 10542
rect 16364 10364 16740 10373
rect 16420 10362 16444 10364
rect 16500 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16420 10310 16430 10362
rect 16674 10310 16684 10362
rect 16420 10308 16444 10310
rect 16500 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16364 10299 16740 10308
rect 16776 10266 16804 10542
rect 16854 10503 16910 10512
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16868 10130 16896 10503
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15580 9178 15608 9454
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15382 9072 15438 9081
rect 15292 9036 15344 9042
rect 15382 9007 15438 9016
rect 15292 8978 15344 8984
rect 15396 8498 15424 9007
rect 15488 8537 15516 9114
rect 15474 8528 15530 8537
rect 15384 8492 15436 8498
rect 15474 8463 15530 8472
rect 15384 8434 15436 8440
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15304 7954 15332 8230
rect 15292 7948 15344 7954
rect 15344 7908 15424 7936
rect 15292 7890 15344 7896
rect 15290 7304 15346 7313
rect 15290 7239 15346 7248
rect 15304 6322 15332 7239
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 14924 5646 14976 5652
rect 15028 5630 15240 5658
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14832 5092 14884 5098
rect 14832 5034 14884 5040
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14844 4554 14872 5034
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14646 3088 14702 3097
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14556 3052 14608 3058
rect 14608 3032 14646 3040
rect 14608 3023 14702 3032
rect 14608 3012 14688 3023
rect 14556 2994 14608 3000
rect 14384 2746 14688 2774
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14568 1834 14596 2382
rect 14556 1828 14608 1834
rect 14556 1770 14608 1776
rect 14660 1766 14688 2746
rect 14648 1760 14700 1766
rect 14648 1702 14700 1708
rect 14752 1426 14780 3130
rect 14844 3058 14872 3878
rect 14936 3738 14964 4966
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14830 2952 14886 2961
rect 14830 2887 14832 2896
rect 14884 2887 14886 2896
rect 14832 2858 14884 2864
rect 15028 2310 15056 5630
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5166 15240 5510
rect 15396 5234 15424 7908
rect 15488 7886 15516 8366
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15488 7410 15516 7686
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15580 5778 15608 9114
rect 15672 8265 15700 9386
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15658 8256 15714 8265
rect 15658 8191 15714 8200
rect 15672 7546 15700 8191
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15474 5264 15530 5273
rect 15384 5228 15436 5234
rect 15474 5199 15476 5208
rect 15384 5170 15436 5176
rect 15528 5199 15530 5208
rect 15476 5170 15528 5176
rect 15200 5160 15252 5166
rect 15252 5120 15332 5148
rect 15200 5102 15252 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15120 4282 15148 4626
rect 15212 4298 15240 4966
rect 15304 4622 15332 5120
rect 15396 4690 15424 5170
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15108 4276 15160 4282
rect 15212 4270 15332 4298
rect 15108 4218 15160 4224
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 14922 2136 14978 2145
rect 14922 2071 14978 2080
rect 14936 1426 14964 2071
rect 15028 1970 15056 2246
rect 15016 1964 15068 1970
rect 15016 1906 15068 1912
rect 15120 1850 15148 3946
rect 15304 3602 15332 4270
rect 15396 4214 15424 4626
rect 15488 4593 15516 5170
rect 15580 4690 15608 5306
rect 15672 5166 15700 6870
rect 15764 5846 15792 8774
rect 15856 8634 15884 9318
rect 15948 8838 15976 9522
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 16026 8800 16082 8809
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15856 7410 15884 8570
rect 15948 8276 15976 8774
rect 16026 8735 16082 8744
rect 16040 8430 16068 8735
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 15948 8248 16068 8276
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15934 6488 15990 6497
rect 15934 6423 15990 6432
rect 15948 6186 15976 6423
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15948 5914 15976 6122
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15764 5370 15792 5782
rect 15934 5536 15990 5545
rect 15934 5471 15990 5480
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15948 5234 15976 5471
rect 16040 5234 16068 8248
rect 16132 6934 16160 9862
rect 16592 9674 16620 9998
rect 16224 9646 16620 9674
rect 16224 9160 16252 9646
rect 16684 9518 16712 10066
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 9722 16804 9862
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16672 9512 16724 9518
rect 16670 9480 16672 9489
rect 16724 9480 16726 9489
rect 16670 9415 16726 9424
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16364 9276 16740 9285
rect 16420 9274 16444 9276
rect 16500 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16420 9222 16430 9274
rect 16674 9222 16684 9274
rect 16420 9220 16444 9222
rect 16500 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16364 9211 16740 9220
rect 16224 9132 16344 9160
rect 16316 8276 16344 9132
rect 16776 9110 16804 9318
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16684 8430 16712 8774
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16580 8424 16632 8430
rect 16578 8392 16580 8401
rect 16672 8424 16724 8430
rect 16632 8392 16634 8401
rect 16672 8366 16724 8372
rect 16776 8378 16804 8570
rect 16868 8498 16896 9386
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16776 8350 16896 8378
rect 16578 8327 16634 8336
rect 16316 8248 16804 8276
rect 16364 8188 16740 8197
rect 16420 8186 16444 8188
rect 16500 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16420 8134 16430 8186
rect 16674 8134 16684 8186
rect 16420 8132 16444 8134
rect 16500 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16364 8123 16740 8132
rect 16776 7886 16804 8248
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7410 16804 7686
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16364 7100 16740 7109
rect 16420 7098 16444 7100
rect 16500 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16420 7046 16430 7098
rect 16674 7046 16684 7098
rect 16420 7044 16444 7046
rect 16500 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16210 7032 16266 7041
rect 16364 7035 16740 7044
rect 16776 7002 16804 7346
rect 16868 7342 16896 8350
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16210 6967 16266 6976
rect 16764 6996 16816 7002
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15660 5024 15712 5030
rect 15712 4984 15884 5012
rect 15660 4966 15712 4972
rect 15568 4684 15620 4690
rect 15752 4684 15804 4690
rect 15620 4644 15700 4672
rect 15568 4626 15620 4632
rect 15474 4584 15530 4593
rect 15474 4519 15530 4528
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15568 4072 15620 4078
rect 15672 4060 15700 4644
rect 15752 4626 15804 4632
rect 15620 4032 15700 4060
rect 15568 4014 15620 4020
rect 15396 3738 15424 4014
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15764 3602 15792 4626
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15212 2650 15240 3470
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15488 2990 15516 3402
rect 15568 3392 15620 3398
rect 15566 3360 15568 3369
rect 15752 3392 15804 3398
rect 15620 3360 15622 3369
rect 15752 3334 15804 3340
rect 15566 3295 15622 3304
rect 15580 2990 15608 3295
rect 15764 3194 15792 3334
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15750 3088 15806 3097
rect 15750 3023 15806 3032
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15568 2984 15620 2990
rect 15620 2944 15700 2972
rect 15568 2926 15620 2932
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15488 1970 15516 2382
rect 15476 1964 15528 1970
rect 15476 1906 15528 1912
rect 15120 1834 15332 1850
rect 15120 1828 15344 1834
rect 15120 1822 15292 1828
rect 15292 1770 15344 1776
rect 15016 1760 15068 1766
rect 15016 1702 15068 1708
rect 15200 1760 15252 1766
rect 15200 1702 15252 1708
rect 15384 1760 15436 1766
rect 15384 1702 15436 1708
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 13820 1420 13872 1426
rect 13820 1362 13872 1368
rect 14096 1420 14148 1426
rect 14096 1362 14148 1368
rect 14740 1420 14792 1426
rect 14740 1362 14792 1368
rect 14924 1420 14976 1426
rect 14924 1362 14976 1368
rect 13504 1176 13584 1204
rect 13820 1216 13872 1222
rect 13452 1158 13504 1164
rect 13820 1158 13872 1164
rect 14372 1216 14424 1222
rect 14372 1158 14424 1164
rect 13004 1018 13032 1158
rect 13364 1116 13740 1125
rect 13420 1114 13444 1116
rect 13500 1114 13524 1116
rect 13580 1114 13604 1116
rect 13660 1114 13684 1116
rect 13420 1062 13430 1114
rect 13674 1062 13684 1114
rect 13420 1060 13444 1062
rect 13500 1060 13524 1062
rect 13580 1060 13604 1062
rect 13660 1060 13684 1062
rect 13364 1051 13740 1060
rect 12992 1012 13044 1018
rect 12992 954 13044 960
rect 13832 814 13860 1158
rect 14384 1018 14412 1158
rect 15028 1018 15056 1702
rect 15212 1426 15240 1702
rect 15200 1420 15252 1426
rect 15200 1362 15252 1368
rect 15108 1216 15160 1222
rect 15108 1158 15160 1164
rect 14372 1012 14424 1018
rect 14372 954 14424 960
rect 15016 1012 15068 1018
rect 15016 954 15068 960
rect 15120 814 15148 1158
rect 13820 808 13872 814
rect 13820 750 13872 756
rect 15108 808 15160 814
rect 15108 750 15160 756
rect 13268 672 13320 678
rect 13268 614 13320 620
rect 14280 672 14332 678
rect 14280 614 14332 620
rect 13280 400 13308 614
rect 14292 490 14320 614
rect 14108 462 14320 490
rect 14108 400 14136 462
rect 12716 264 12768 270
rect 12716 206 12768 212
rect 13266 0 13322 400
rect 14094 0 14150 400
rect 15396 338 15424 1702
rect 15488 1562 15516 1702
rect 15476 1556 15528 1562
rect 15476 1498 15528 1504
rect 15580 1426 15608 2790
rect 15672 2582 15700 2944
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15764 2394 15792 3023
rect 15672 2366 15792 2394
rect 15672 2145 15700 2366
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15658 2136 15714 2145
rect 15658 2071 15714 2080
rect 15658 1592 15714 1601
rect 15658 1527 15660 1536
rect 15712 1527 15714 1536
rect 15660 1498 15712 1504
rect 15764 1426 15792 2246
rect 15856 1902 15884 4984
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15948 4146 15976 4694
rect 16026 4584 16082 4593
rect 16026 4519 16082 4528
rect 16040 4146 16068 4519
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16040 3058 16068 3538
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15936 2848 15988 2854
rect 15988 2796 16068 2802
rect 15936 2790 16068 2796
rect 15948 2774 16068 2790
rect 15934 2272 15990 2281
rect 15934 2207 15990 2216
rect 15948 1902 15976 2207
rect 15844 1896 15896 1902
rect 15844 1838 15896 1844
rect 15936 1896 15988 1902
rect 15936 1838 15988 1844
rect 15948 1426 15976 1838
rect 15568 1420 15620 1426
rect 15568 1362 15620 1368
rect 15752 1420 15804 1426
rect 15752 1362 15804 1368
rect 15936 1420 15988 1426
rect 15936 1362 15988 1368
rect 15948 1306 15976 1362
rect 15752 1284 15804 1290
rect 15752 1226 15804 1232
rect 15856 1278 15976 1306
rect 15764 1018 15792 1226
rect 15752 1012 15804 1018
rect 15752 954 15804 960
rect 15856 814 15884 1278
rect 15936 1216 15988 1222
rect 15936 1158 15988 1164
rect 15948 1018 15976 1158
rect 16040 1018 16068 2774
rect 16132 2394 16160 6054
rect 16224 5370 16252 6967
rect 16764 6938 16816 6944
rect 16868 6254 16896 7278
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16364 6012 16740 6021
rect 16420 6010 16444 6012
rect 16500 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16420 5958 16430 6010
rect 16674 5958 16684 6010
rect 16420 5956 16444 5958
rect 16500 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16364 5947 16740 5956
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16868 5574 16896 5714
rect 16856 5568 16908 5574
rect 16960 5545 16988 14554
rect 17052 14414 17080 15030
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17130 14376 17186 14385
rect 17052 13938 17080 14350
rect 17130 14311 17132 14320
rect 17184 14311 17186 14320
rect 17132 14282 17184 14288
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17236 12782 17264 15370
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 17328 13734 17356 15030
rect 17696 14958 17724 15600
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 18064 14618 18092 15302
rect 18432 14958 18460 15600
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17958 14512 18014 14521
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17144 10713 17172 11698
rect 17236 11694 17264 12718
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17130 10704 17186 10713
rect 17040 10668 17092 10674
rect 17186 10662 17264 10690
rect 17130 10639 17186 10648
rect 17040 10610 17092 10616
rect 17052 9722 17080 10610
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17144 10266 17172 10542
rect 17236 10470 17264 10662
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17328 10146 17356 12582
rect 17420 12442 17448 14486
rect 17592 14476 17644 14482
rect 18248 14482 18276 14826
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 17958 14447 18014 14456
rect 18236 14476 18288 14482
rect 17592 14418 17644 14424
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17512 13530 17540 14282
rect 17604 14074 17632 14418
rect 17972 14414 18000 14447
rect 18236 14418 18288 14424
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 14074 17908 14214
rect 18432 14074 18460 14554
rect 17592 14068 17644 14074
rect 17868 14068 17920 14074
rect 17592 14010 17644 14016
rect 17788 14028 17868 14056
rect 17788 13530 17816 14028
rect 17868 14010 17920 14016
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17604 12986 17632 13126
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17406 12200 17462 12209
rect 17406 12135 17462 12144
rect 17592 12164 17644 12170
rect 17420 11898 17448 12135
rect 17592 12106 17644 12112
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17420 10248 17448 11834
rect 17604 11218 17632 12106
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17604 10606 17632 11154
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17420 10220 17724 10248
rect 17328 10118 17448 10146
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17052 8090 17080 9658
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 8974 17264 9318
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17222 8664 17278 8673
rect 17328 8634 17356 9998
rect 17222 8599 17224 8608
rect 17276 8599 17278 8608
rect 17316 8628 17368 8634
rect 17224 8570 17276 8576
rect 17316 8570 17368 8576
rect 17314 8528 17370 8537
rect 17314 8463 17370 8472
rect 17328 8430 17356 8463
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 7002 17080 7142
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17052 5778 17080 5850
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16856 5510 16908 5516
rect 16946 5536 17002 5545
rect 16946 5471 17002 5480
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16224 4758 16252 5170
rect 17040 5160 17092 5166
rect 16946 5128 17002 5137
rect 17040 5102 17092 5108
rect 16946 5063 17002 5072
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16364 4924 16740 4933
rect 16420 4922 16444 4924
rect 16500 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16420 4870 16430 4922
rect 16674 4870 16684 4922
rect 16420 4868 16444 4870
rect 16500 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16364 4859 16740 4868
rect 16868 4826 16896 4966
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 4078 16252 4422
rect 16408 4146 16436 4490
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16304 3936 16356 3942
rect 16224 3896 16304 3924
rect 16224 3482 16252 3896
rect 16304 3878 16356 3884
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16364 3836 16740 3845
rect 16420 3834 16444 3836
rect 16500 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16420 3782 16430 3834
rect 16674 3782 16684 3834
rect 16420 3780 16444 3782
rect 16500 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16364 3771 16740 3780
rect 16776 3670 16804 3878
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16224 3454 16344 3482
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16224 3194 16252 3334
rect 16316 3194 16344 3454
rect 16408 3369 16436 3538
rect 16578 3496 16634 3505
rect 16578 3431 16634 3440
rect 16856 3460 16908 3466
rect 16394 3360 16450 3369
rect 16394 3295 16450 3304
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16210 3088 16266 3097
rect 16304 3052 16356 3058
rect 16266 3032 16304 3040
rect 16210 3023 16304 3032
rect 16224 3012 16304 3023
rect 16304 2994 16356 3000
rect 16592 2990 16620 3431
rect 16856 3402 16908 3408
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16224 2514 16252 2790
rect 16364 2748 16740 2757
rect 16420 2746 16444 2748
rect 16500 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16420 2694 16430 2746
rect 16674 2694 16684 2746
rect 16420 2692 16444 2694
rect 16500 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16364 2683 16740 2692
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16672 2508 16724 2514
rect 16776 2496 16804 2858
rect 16868 2582 16896 3402
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 16724 2468 16804 2496
rect 16672 2450 16724 2456
rect 16132 2366 16252 2394
rect 16118 2136 16174 2145
rect 16118 2071 16174 2080
rect 16132 1970 16160 2071
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 16224 1426 16252 2366
rect 16776 1902 16804 2468
rect 16764 1896 16816 1902
rect 16764 1838 16816 1844
rect 16364 1660 16740 1669
rect 16420 1658 16444 1660
rect 16500 1658 16524 1660
rect 16580 1658 16604 1660
rect 16660 1658 16684 1660
rect 16420 1606 16430 1658
rect 16674 1606 16684 1658
rect 16420 1604 16444 1606
rect 16500 1604 16524 1606
rect 16580 1604 16604 1606
rect 16660 1604 16684 1606
rect 16364 1595 16740 1604
rect 16394 1456 16450 1465
rect 16212 1420 16264 1426
rect 16394 1391 16396 1400
rect 16212 1362 16264 1368
rect 16448 1391 16450 1400
rect 16764 1420 16816 1426
rect 16396 1362 16448 1368
rect 16960 1408 16988 5063
rect 17052 4729 17080 5102
rect 17038 4720 17094 4729
rect 17038 4655 17094 4664
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17052 2514 17080 2926
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17052 1970 17080 2246
rect 17144 2009 17172 7686
rect 17420 7562 17448 10118
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 8022 17540 10066
rect 17696 9722 17724 10220
rect 17788 10130 17816 10950
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17696 9382 17724 9658
rect 17788 9602 17816 10066
rect 17880 9674 17908 13806
rect 18524 13530 18552 14758
rect 18616 14482 18644 15098
rect 19168 14958 19196 15600
rect 19364 15260 19740 15269
rect 19420 15258 19444 15260
rect 19500 15258 19524 15260
rect 19580 15258 19604 15260
rect 19660 15258 19684 15260
rect 19420 15206 19430 15258
rect 19674 15206 19684 15258
rect 19420 15204 19444 15206
rect 19500 15204 19524 15206
rect 19580 15204 19604 15206
rect 19660 15204 19684 15206
rect 19364 15195 19740 15204
rect 20180 14958 20208 15694
rect 20626 15600 20682 16000
rect 21362 15600 21418 16000
rect 22098 15600 22154 16000
rect 22834 15600 22890 16000
rect 20640 14958 20668 15600
rect 21376 14958 21404 15600
rect 22112 14958 22140 15600
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22296 15094 22324 15302
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22848 14958 22876 15600
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 18892 14521 18920 14758
rect 19260 14618 19288 14758
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 18878 14512 18934 14521
rect 18604 14476 18656 14482
rect 19996 14482 20024 14758
rect 18878 14447 18934 14456
rect 19984 14476 20036 14482
rect 18604 14418 18656 14424
rect 18616 14362 18644 14418
rect 18788 14408 18840 14414
rect 18616 14334 18736 14362
rect 18788 14350 18840 14356
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18616 14074 18644 14214
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18616 13977 18644 14010
rect 18602 13968 18658 13977
rect 18602 13903 18658 13912
rect 18708 13870 18736 14334
rect 18696 13864 18748 13870
rect 18602 13832 18658 13841
rect 18658 13812 18696 13818
rect 18658 13806 18748 13812
rect 18658 13790 18736 13806
rect 18602 13767 18658 13776
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18708 13530 18736 13670
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17972 12434 18000 13398
rect 18064 12850 18092 13466
rect 18432 13326 18460 13466
rect 18524 13394 18552 13466
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18340 12850 18368 13262
rect 18800 12850 18828 14350
rect 18892 14346 18920 14447
rect 19984 14418 20036 14424
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 19364 14172 19740 14181
rect 19420 14170 19444 14172
rect 19500 14170 19524 14172
rect 19580 14170 19604 14172
rect 19660 14170 19684 14172
rect 19420 14118 19430 14170
rect 19674 14118 19684 14170
rect 19420 14116 19444 14118
rect 19500 14116 19524 14118
rect 19580 14116 19604 14118
rect 19660 14116 19684 14118
rect 19364 14107 19740 14116
rect 20088 14074 20116 14894
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20074 13968 20130 13977
rect 19156 13932 19208 13938
rect 20074 13903 20130 13912
rect 19156 13874 19208 13880
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18878 13424 18934 13433
rect 18984 13410 19012 13806
rect 19168 13530 19196 13874
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 18934 13382 19012 13410
rect 19800 13388 19852 13394
rect 18878 13359 18934 13368
rect 19800 13330 19852 13336
rect 19364 13084 19740 13093
rect 19420 13082 19444 13084
rect 19500 13082 19524 13084
rect 19580 13082 19604 13084
rect 19660 13082 19684 13084
rect 19420 13030 19430 13082
rect 19674 13030 19684 13082
rect 19420 13028 19444 13030
rect 19500 13028 19524 13030
rect 19580 13028 19604 13030
rect 19660 13028 19684 13030
rect 19364 13019 19740 13028
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 19812 12782 19840 13330
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18800 12434 18828 12582
rect 17972 12406 18092 12434
rect 18800 12406 19012 12434
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17972 11150 18000 11630
rect 17960 11144 18012 11150
rect 17958 11112 17960 11121
rect 18012 11112 18014 11121
rect 17958 11047 18014 11056
rect 17880 9646 18000 9674
rect 17788 9574 17908 9602
rect 17880 9518 17908 9574
rect 17868 9512 17920 9518
rect 17774 9480 17830 9489
rect 17868 9454 17920 9460
rect 17774 9415 17830 9424
rect 17788 9382 17816 9415
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9178 17816 9318
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17604 8634 17632 9046
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17696 8430 17724 8774
rect 17788 8673 17816 8774
rect 17774 8664 17830 8673
rect 17774 8599 17830 8608
rect 17774 8528 17830 8537
rect 17774 8463 17830 8472
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17500 8016 17552 8022
rect 17498 7984 17500 7993
rect 17552 7984 17554 7993
rect 17498 7919 17554 7928
rect 17420 7534 17540 7562
rect 17408 7472 17460 7478
rect 17406 7440 17408 7449
rect 17460 7440 17462 7449
rect 17406 7375 17462 7384
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 6798 17264 7142
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17314 6896 17370 6905
rect 17314 6831 17370 6840
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17236 5642 17264 5782
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17236 5234 17264 5578
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17236 3602 17264 4626
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17328 3482 17356 6831
rect 17236 3454 17356 3482
rect 17130 2000 17186 2009
rect 17040 1964 17092 1970
rect 17130 1935 17186 1944
rect 17040 1906 17092 1912
rect 17144 1562 17172 1935
rect 17132 1556 17184 1562
rect 17132 1498 17184 1504
rect 17236 1426 17264 3454
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17328 3194 17356 3334
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17420 1426 17448 6938
rect 17512 2281 17540 7534
rect 17604 6458 17632 8230
rect 17788 7886 17816 8463
rect 17880 8430 17908 9046
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17684 7336 17736 7342
rect 17682 7304 17684 7313
rect 17736 7304 17738 7313
rect 17682 7239 17738 7248
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17604 5914 17632 6394
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17498 2272 17554 2281
rect 17498 2207 17554 2216
rect 16816 1380 16988 1408
rect 17224 1420 17276 1426
rect 16764 1362 16816 1368
rect 17224 1362 17276 1368
rect 17408 1420 17460 1426
rect 17408 1362 17460 1368
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 15936 1012 15988 1018
rect 15936 954 15988 960
rect 16028 1012 16080 1018
rect 16028 954 16080 960
rect 16132 814 16160 1294
rect 16580 1216 16632 1222
rect 16580 1158 16632 1164
rect 17408 1216 17460 1222
rect 17408 1158 17460 1164
rect 16592 814 16620 1158
rect 17420 814 17448 1158
rect 17604 1018 17632 5306
rect 17696 4282 17724 7239
rect 17880 6866 17908 8366
rect 17972 7750 18000 9646
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17972 6934 18000 7142
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6254 17908 6802
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17788 5012 17816 6122
rect 17880 5710 17908 6190
rect 17972 5914 18000 6190
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17868 5024 17920 5030
rect 17788 4984 17868 5012
rect 17868 4966 17920 4972
rect 17880 4690 17908 4966
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17972 3505 18000 3538
rect 17958 3496 18014 3505
rect 17958 3431 18014 3440
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 17880 1902 17908 2518
rect 17868 1896 17920 1902
rect 18064 1850 18092 12406
rect 18326 12336 18382 12345
rect 18326 12271 18328 12280
rect 18380 12271 18382 12280
rect 18420 12300 18472 12306
rect 18328 12242 18380 12248
rect 18420 12242 18472 12248
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18340 11898 18368 12242
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18248 10810 18276 11222
rect 18432 11218 18460 12242
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18524 11898 18552 12038
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18616 11694 18644 12038
rect 18708 11898 18736 12242
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 8906 18184 9318
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18248 8106 18276 10746
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18340 9654 18368 10066
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18340 9042 18368 9590
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18432 8634 18460 11154
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 9466 18552 10406
rect 18616 9586 18644 11630
rect 18800 11218 18828 12174
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18524 9438 18644 9466
rect 18708 9450 18736 10202
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18156 8078 18276 8106
rect 18156 7342 18184 8078
rect 18326 7848 18382 7857
rect 18326 7783 18382 7792
rect 18340 7342 18368 7783
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18156 6118 18184 7278
rect 18340 6254 18368 7278
rect 18524 6644 18552 8978
rect 18616 8786 18644 9438
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18800 9178 18828 9318
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18892 9110 18920 9318
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18800 8786 18828 8842
rect 18616 8758 18828 8786
rect 18800 8401 18828 8758
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18786 8392 18842 8401
rect 18786 8327 18842 8336
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 7954 18736 8230
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 7546 18736 7890
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 7546 18828 7686
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18892 7342 18920 8570
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18708 6798 18736 7278
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18524 6616 18736 6644
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5778 18184 6054
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18248 5166 18276 5646
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18236 4752 18288 4758
rect 18236 4694 18288 4700
rect 18248 4282 18276 4694
rect 18432 4486 18460 5102
rect 18708 4622 18736 6616
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18800 5778 18828 6258
rect 18788 5772 18840 5778
rect 18788 5714 18840 5720
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18892 5302 18920 5714
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 18340 3058 18368 3402
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18234 2680 18290 2689
rect 18234 2615 18290 2624
rect 18248 2514 18276 2615
rect 18340 2514 18368 2994
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18248 1884 18276 2450
rect 18432 2310 18460 4422
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18524 4185 18552 4218
rect 18510 4176 18566 4185
rect 18708 4146 18736 4558
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18510 4111 18566 4120
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18510 4040 18566 4049
rect 18510 3975 18566 3984
rect 18604 4004 18656 4010
rect 18524 3398 18552 3975
rect 18604 3946 18656 3952
rect 18616 3738 18644 3946
rect 18604 3732 18656 3738
rect 18656 3692 18828 3720
rect 18604 3674 18656 3680
rect 18602 3496 18658 3505
rect 18696 3460 18748 3466
rect 18658 3440 18696 3448
rect 18602 3431 18696 3440
rect 18616 3420 18696 3431
rect 18696 3402 18748 3408
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18524 3126 18552 3334
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 18800 2990 18828 3692
rect 18892 3641 18920 4422
rect 18878 3632 18934 3641
rect 18878 3567 18934 3576
rect 18892 3194 18920 3567
rect 18880 3188 18932 3194
rect 18880 3130 18932 3136
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 17868 1838 17920 1844
rect 17972 1822 18092 1850
rect 18156 1856 18276 1884
rect 18432 1873 18460 2246
rect 18708 2106 18736 2790
rect 18984 2632 19012 12406
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 19076 10266 19104 12310
rect 19364 11996 19740 12005
rect 19420 11994 19444 11996
rect 19500 11994 19524 11996
rect 19580 11994 19604 11996
rect 19660 11994 19684 11996
rect 19420 11942 19430 11994
rect 19674 11942 19684 11994
rect 19420 11940 19444 11942
rect 19500 11940 19524 11942
rect 19580 11940 19604 11942
rect 19660 11940 19684 11942
rect 19364 11931 19740 11940
rect 19904 11694 19932 12650
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19168 11354 19196 11630
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19708 11144 19760 11150
rect 19706 11112 19708 11121
rect 19760 11112 19762 11121
rect 19706 11047 19762 11056
rect 19364 10908 19740 10917
rect 19420 10906 19444 10908
rect 19500 10906 19524 10908
rect 19580 10906 19604 10908
rect 19660 10906 19684 10908
rect 19420 10854 19430 10906
rect 19674 10854 19684 10906
rect 19420 10852 19444 10854
rect 19500 10852 19524 10854
rect 19580 10852 19604 10854
rect 19660 10852 19684 10854
rect 19364 10843 19740 10852
rect 19812 10810 19840 11222
rect 19904 10810 19932 11290
rect 19996 10962 20024 12650
rect 20088 11082 20116 13903
rect 20180 13870 20208 14758
rect 21468 14618 21496 14894
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21468 14074 21496 14554
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20180 12646 20208 13806
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 12782 20300 13262
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20456 12782 20484 13126
rect 21376 12986 21404 13330
rect 21468 13002 21496 13398
rect 21560 13258 21588 14758
rect 22364 14716 22740 14725
rect 22420 14714 22444 14716
rect 22500 14714 22524 14716
rect 22580 14714 22604 14716
rect 22660 14714 22684 14716
rect 22420 14662 22430 14714
rect 22674 14662 22684 14714
rect 22420 14660 22444 14662
rect 22500 14660 22524 14662
rect 22580 14660 22604 14662
rect 22660 14660 22684 14662
rect 22364 14651 22740 14660
rect 22364 13628 22740 13637
rect 22420 13626 22444 13628
rect 22500 13626 22524 13628
rect 22580 13626 22604 13628
rect 22660 13626 22684 13628
rect 22420 13574 22430 13626
rect 22674 13574 22684 13626
rect 22420 13572 22444 13574
rect 22500 13572 22524 13574
rect 22580 13572 22604 13574
rect 22660 13572 22684 13574
rect 22364 13563 22740 13572
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 21364 12980 21416 12986
rect 21468 12974 21680 13002
rect 21364 12922 21416 12928
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20272 12374 20300 12718
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20272 11762 20300 12310
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 20260 11008 20312 11014
rect 19996 10934 20208 10962
rect 20260 10950 20312 10956
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19340 10600 19392 10606
rect 19260 10560 19340 10588
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19062 10160 19118 10169
rect 19260 10146 19288 10560
rect 19340 10542 19392 10548
rect 19904 10554 19932 10746
rect 19904 10526 20116 10554
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19118 10118 19288 10146
rect 19062 10095 19118 10104
rect 19168 9586 19196 10118
rect 19352 10062 19380 10202
rect 19812 10130 19840 10406
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19340 10056 19392 10062
rect 19338 10024 19340 10033
rect 19392 10024 19394 10033
rect 19338 9959 19394 9968
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19812 9874 19840 10066
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19904 9897 19932 9998
rect 19890 9888 19946 9897
rect 19260 9704 19288 9862
rect 19812 9846 19849 9874
rect 19364 9820 19740 9829
rect 19420 9818 19444 9820
rect 19500 9818 19524 9820
rect 19580 9818 19604 9820
rect 19660 9818 19684 9820
rect 19420 9766 19430 9818
rect 19674 9766 19684 9818
rect 19420 9764 19444 9766
rect 19500 9764 19524 9766
rect 19580 9764 19604 9766
rect 19660 9764 19684 9766
rect 19364 9755 19740 9764
rect 19821 9738 19849 9846
rect 19890 9823 19946 9832
rect 19996 9738 20024 10406
rect 20088 10062 20116 10526
rect 20180 10266 20208 10934
rect 20272 10674 20300 10950
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20076 10056 20128 10062
rect 20128 10016 20208 10044
rect 20076 9998 20128 10004
rect 19812 9710 19849 9738
rect 19904 9710 20024 9738
rect 19260 9676 19472 9704
rect 19338 9616 19394 9625
rect 19156 9580 19208 9586
rect 19338 9551 19394 9560
rect 19156 9522 19208 9528
rect 19352 9042 19380 9551
rect 19444 9217 19472 9676
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19430 9208 19486 9217
rect 19430 9143 19486 9152
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19168 8922 19196 8978
rect 19536 8922 19564 9386
rect 19706 9072 19762 9081
rect 19812 9042 19840 9710
rect 19904 9654 19932 9710
rect 19892 9648 19944 9654
rect 19892 9590 19944 9596
rect 19982 9616 20038 9625
rect 19904 9484 19932 9590
rect 20038 9586 20116 9602
rect 20038 9580 20128 9586
rect 20038 9574 20076 9580
rect 19982 9551 20038 9560
rect 20076 9522 20128 9528
rect 19892 9478 19944 9484
rect 19892 9420 19944 9426
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 9042 20024 9318
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 19706 9007 19762 9016
rect 19800 9036 19852 9042
rect 19720 8974 19748 9007
rect 19800 8978 19852 8984
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19064 8900 19116 8906
rect 19168 8894 19564 8922
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19064 8842 19116 8848
rect 19076 8634 19104 8842
rect 19340 8832 19392 8838
rect 19260 8792 19340 8820
rect 19260 8634 19288 8792
rect 19340 8774 19392 8780
rect 19364 8732 19740 8741
rect 19420 8730 19444 8732
rect 19500 8730 19524 8732
rect 19580 8730 19604 8732
rect 19660 8730 19684 8732
rect 19420 8678 19430 8730
rect 19674 8678 19684 8730
rect 19420 8676 19444 8678
rect 19500 8676 19524 8678
rect 19580 8676 19604 8678
rect 19660 8676 19684 8678
rect 19364 8667 19740 8676
rect 19812 8634 19840 8978
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19352 7732 19380 8366
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19812 7954 19840 8230
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19260 7704 19380 7732
rect 19260 7528 19288 7704
rect 19364 7644 19740 7653
rect 19420 7642 19444 7644
rect 19500 7642 19524 7644
rect 19580 7642 19604 7644
rect 19660 7642 19684 7644
rect 19420 7590 19430 7642
rect 19674 7590 19684 7642
rect 19420 7588 19444 7590
rect 19500 7588 19524 7590
rect 19580 7588 19604 7590
rect 19660 7588 19684 7590
rect 19364 7579 19740 7588
rect 19340 7540 19392 7546
rect 19260 7500 19340 7528
rect 19340 7482 19392 7488
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19364 6556 19740 6565
rect 19420 6554 19444 6556
rect 19500 6554 19524 6556
rect 19580 6554 19604 6556
rect 19660 6554 19684 6556
rect 19420 6502 19430 6554
rect 19674 6502 19684 6554
rect 19420 6500 19444 6502
rect 19500 6500 19524 6502
rect 19580 6500 19604 6502
rect 19660 6500 19684 6502
rect 19364 6491 19740 6500
rect 19812 6254 19840 7278
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19076 5574 19104 6054
rect 19812 5778 19840 6190
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19168 5370 19196 5714
rect 19364 5468 19740 5477
rect 19420 5466 19444 5468
rect 19500 5466 19524 5468
rect 19580 5466 19604 5468
rect 19660 5466 19684 5468
rect 19420 5414 19430 5466
rect 19674 5414 19684 5466
rect 19420 5412 19444 5414
rect 19500 5412 19524 5414
rect 19580 5412 19604 5414
rect 19660 5412 19684 5414
rect 19364 5403 19740 5412
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 19614 4584 19670 4593
rect 19614 4519 19616 4528
rect 19668 4519 19670 4528
rect 19616 4490 19668 4496
rect 19364 4380 19740 4389
rect 19420 4378 19444 4380
rect 19500 4378 19524 4380
rect 19580 4378 19604 4380
rect 19660 4378 19684 4380
rect 19420 4326 19430 4378
rect 19674 4326 19684 4378
rect 19420 4324 19444 4326
rect 19500 4324 19524 4326
rect 19580 4324 19604 4326
rect 19660 4324 19684 4326
rect 19364 4315 19740 4324
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19628 3602 19656 3946
rect 19812 3602 19840 4694
rect 19904 3738 19932 8774
rect 19996 8566 20024 8978
rect 20088 8634 20116 9046
rect 20180 8974 20208 10016
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20272 9625 20300 9862
rect 20258 9616 20314 9625
rect 20258 9551 20314 9560
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20260 8832 20312 8838
rect 20180 8792 20260 8820
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20180 8378 20208 8792
rect 20260 8774 20312 8780
rect 19996 8362 20208 8378
rect 19984 8356 20208 8362
rect 20036 8350 20208 8356
rect 20260 8356 20312 8362
rect 19984 8298 20036 8304
rect 20260 8298 20312 8304
rect 20272 8265 20300 8298
rect 19982 8256 20038 8265
rect 19982 8191 20038 8200
rect 20258 8256 20314 8265
rect 20258 8191 20314 8200
rect 19996 7886 20024 8191
rect 20364 7970 20392 11630
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20456 9178 20484 11562
rect 20640 11354 20668 11698
rect 20732 11665 20760 12582
rect 21088 11688 21140 11694
rect 20718 11656 20774 11665
rect 20774 11614 20852 11642
rect 21088 11630 21140 11636
rect 20718 11591 20774 11600
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20548 9654 20576 11290
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20640 11121 20668 11154
rect 20626 11112 20682 11121
rect 20626 11047 20682 11056
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10606 20760 10950
rect 20824 10606 20852 11614
rect 20904 11620 20956 11626
rect 20904 11562 20956 11568
rect 20916 10810 20944 11562
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 21008 11354 21036 11494
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21100 11218 21128 11630
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 21560 10266 21588 12786
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21652 10130 21680 12974
rect 23294 12880 23350 12889
rect 23294 12815 23296 12824
rect 23348 12815 23350 12824
rect 23296 12786 23348 12792
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22112 10674 22140 11494
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20994 9888 21050 9897
rect 20640 9722 20668 9862
rect 20994 9823 21050 9832
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20088 7942 20392 7970
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19996 6225 20024 7686
rect 19982 6216 20038 6225
rect 19982 6151 20038 6160
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19996 4690 20024 5034
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19996 4078 20024 4422
rect 20088 4214 20116 7942
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 20180 4282 20208 4490
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20076 4208 20128 4214
rect 20076 4150 20128 4156
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19982 3632 20038 3641
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19800 3596 19852 3602
rect 19982 3567 20038 3576
rect 19800 3538 19852 3544
rect 19996 3534 20024 3567
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 19076 2990 19104 3334
rect 19364 3292 19740 3301
rect 19420 3290 19444 3292
rect 19500 3290 19524 3292
rect 19580 3290 19604 3292
rect 19660 3290 19684 3292
rect 19420 3238 19430 3290
rect 19674 3238 19684 3290
rect 19420 3236 19444 3238
rect 19500 3236 19524 3238
rect 19580 3236 19604 3238
rect 19660 3236 19684 3238
rect 19364 3227 19740 3236
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19352 2774 19380 2926
rect 18892 2604 19012 2632
rect 19260 2746 19380 2774
rect 18892 2417 18920 2604
rect 19260 2446 19288 2746
rect 19444 2632 19472 3062
rect 19706 2952 19762 2961
rect 19904 2938 19932 3334
rect 19762 2910 19932 2938
rect 20088 2922 20116 3334
rect 20272 2922 20300 7822
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20364 6866 20392 7482
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20364 5166 20392 5238
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20364 4146 20392 5102
rect 20456 4758 20484 9114
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20548 7954 20576 8366
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20548 7478 20576 7890
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20444 4752 20496 4758
rect 20444 4694 20496 4700
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20456 4078 20484 4694
rect 20640 4214 20668 9658
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20732 8634 20760 9318
rect 20824 8945 20852 9454
rect 21008 9042 21036 9823
rect 21192 9722 21220 9930
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21270 9616 21326 9625
rect 21270 9551 21326 9560
rect 21088 9512 21140 9518
rect 21086 9480 21088 9489
rect 21140 9480 21142 9489
rect 21086 9415 21142 9424
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 20904 8968 20956 8974
rect 20810 8936 20866 8945
rect 20904 8910 20956 8916
rect 20810 8871 20866 8880
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20718 8392 20774 8401
rect 20718 8327 20774 8336
rect 20732 7886 20760 8327
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20824 7546 20852 7890
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20732 6458 20760 6598
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20732 4486 20760 6394
rect 20916 6304 20944 8910
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21008 6322 21036 8774
rect 21284 8498 21312 9551
rect 21376 9081 21404 9658
rect 21456 9104 21508 9110
rect 21362 9072 21418 9081
rect 21456 9046 21508 9052
rect 21362 9007 21418 9016
rect 21376 8634 21404 9007
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21468 8566 21496 9046
rect 21456 8560 21508 8566
rect 21456 8502 21508 8508
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 7546 21128 7686
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20824 6276 20944 6304
rect 20996 6316 21048 6322
rect 20824 4826 20852 6276
rect 20996 6258 21048 6264
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20996 6180 21048 6186
rect 20996 6122 21048 6128
rect 20916 5370 20944 6122
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 21008 4690 21036 6122
rect 21088 5092 21140 5098
rect 21088 5034 21140 5040
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 21008 4554 21036 4626
rect 21100 4622 21128 5034
rect 21192 4826 21220 8298
rect 21284 8265 21312 8298
rect 21270 8256 21326 8265
rect 21270 8191 21326 8200
rect 21284 7002 21312 8191
rect 21376 7750 21404 8366
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21376 7342 21404 7686
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21284 4690 21312 6258
rect 21362 5672 21418 5681
rect 21362 5607 21364 5616
rect 21416 5607 21418 5616
rect 21364 5578 21416 5584
rect 21468 5166 21496 8502
rect 21560 6118 21588 9998
rect 21638 9616 21694 9625
rect 21638 9551 21694 9560
rect 21652 9518 21680 9551
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21652 8537 21680 9318
rect 21744 9178 21772 9998
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21638 8528 21694 8537
rect 21638 8463 21640 8472
rect 21692 8463 21694 8472
rect 21640 8434 21692 8440
rect 21836 6866 21864 10406
rect 22112 9722 22140 10610
rect 22204 10266 22232 12650
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22364 12540 22740 12549
rect 22420 12538 22444 12540
rect 22500 12538 22524 12540
rect 22580 12538 22604 12540
rect 22660 12538 22684 12540
rect 22420 12486 22430 12538
rect 22674 12486 22684 12538
rect 22420 12484 22444 12486
rect 22500 12484 22524 12486
rect 22580 12484 22604 12486
rect 22660 12484 22684 12486
rect 22364 12475 22740 12484
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22296 11014 22324 12038
rect 22364 11452 22740 11461
rect 22420 11450 22444 11452
rect 22500 11450 22524 11452
rect 22580 11450 22604 11452
rect 22660 11450 22684 11452
rect 22420 11398 22430 11450
rect 22674 11398 22684 11450
rect 22420 11396 22444 11398
rect 22500 11396 22524 11398
rect 22580 11396 22604 11398
rect 22660 11396 22684 11398
rect 22364 11387 22740 11396
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22296 10606 22324 10950
rect 22848 10674 22876 12582
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 22204 9722 22232 9998
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22192 9716 22244 9722
rect 22192 9658 22244 9664
rect 22008 9648 22060 9654
rect 22296 9602 22324 10542
rect 22364 10364 22740 10373
rect 22420 10362 22444 10364
rect 22500 10362 22524 10364
rect 22580 10362 22604 10364
rect 22660 10362 22684 10364
rect 22420 10310 22430 10362
rect 22674 10310 22684 10362
rect 22420 10308 22444 10310
rect 22500 10308 22524 10310
rect 22580 10308 22604 10310
rect 22660 10308 22684 10310
rect 22364 10299 22740 10308
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22480 9722 22508 10066
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22060 9596 22324 9602
rect 22008 9590 22324 9596
rect 22020 9574 22324 9590
rect 22192 9512 22244 9518
rect 22098 9480 22154 9489
rect 22192 9454 22244 9460
rect 22098 9415 22100 9424
rect 22152 9415 22154 9424
rect 22100 9386 22152 9392
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22020 8634 22048 9318
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21652 5370 21680 6598
rect 21744 5642 21772 6598
rect 21824 6452 21876 6458
rect 21928 6440 21956 6802
rect 21876 6412 21956 6440
rect 21824 6394 21876 6400
rect 21836 5778 21864 6394
rect 22112 5914 22140 9386
rect 22204 9178 22232 9454
rect 22756 9450 22784 9862
rect 22848 9518 22876 10610
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22836 9512 22888 9518
rect 22836 9454 22888 9460
rect 22744 9444 22796 9450
rect 22744 9386 22796 9392
rect 22364 9276 22740 9285
rect 22420 9274 22444 9276
rect 22500 9274 22524 9276
rect 22580 9274 22604 9276
rect 22660 9274 22684 9276
rect 22420 9222 22430 9274
rect 22674 9222 22684 9274
rect 22420 9220 22444 9222
rect 22500 9220 22524 9222
rect 22580 9220 22604 9222
rect 22660 9220 22684 9222
rect 22364 9211 22740 9220
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22940 8498 22968 10406
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22364 8188 22740 8197
rect 22420 8186 22444 8188
rect 22500 8186 22524 8188
rect 22580 8186 22604 8188
rect 22660 8186 22684 8188
rect 22420 8134 22430 8186
rect 22674 8134 22684 8186
rect 22420 8132 22444 8134
rect 22500 8132 22524 8134
rect 22580 8132 22604 8134
rect 22660 8132 22684 8134
rect 22364 8123 22740 8132
rect 22364 7100 22740 7109
rect 22420 7098 22444 7100
rect 22500 7098 22524 7100
rect 22580 7098 22604 7100
rect 22660 7098 22684 7100
rect 22420 7046 22430 7098
rect 22674 7046 22684 7098
rect 22420 7044 22444 7046
rect 22500 7044 22524 7046
rect 22580 7044 22604 7046
rect 22660 7044 22684 7046
rect 22364 7035 22740 7044
rect 22364 6012 22740 6021
rect 22420 6010 22444 6012
rect 22500 6010 22524 6012
rect 22580 6010 22604 6012
rect 22660 6010 22684 6012
rect 22420 5958 22430 6010
rect 22674 5958 22684 6010
rect 22420 5956 22444 5958
rect 22500 5956 22524 5958
rect 22580 5956 22604 5958
rect 22660 5956 22684 5958
rect 22364 5947 22740 5956
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21640 5364 21692 5370
rect 21640 5306 21692 5312
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20628 4208 20680 4214
rect 20824 4196 20852 4422
rect 20628 4150 20680 4156
rect 20732 4168 20852 4196
rect 20732 4078 20760 4168
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20076 2916 20128 2922
rect 19706 2887 19762 2896
rect 19352 2604 19472 2632
rect 19352 2514 19380 2604
rect 19720 2514 19748 2887
rect 20076 2858 20128 2864
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20272 2650 20300 2858
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 20640 2446 20668 4014
rect 20824 3738 20852 4014
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20904 3664 20956 3670
rect 20904 3606 20956 3612
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20824 2650 20852 3538
rect 20916 3194 20944 3606
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 19248 2440 19300 2446
rect 18878 2408 18934 2417
rect 18934 2366 19012 2394
rect 19248 2382 19300 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 18878 2343 18934 2352
rect 18696 2100 18748 2106
rect 18696 2042 18748 2048
rect 18880 2100 18932 2106
rect 18880 2042 18932 2048
rect 18418 1864 18474 1873
rect 17684 1420 17736 1426
rect 17972 1408 18000 1822
rect 18052 1760 18104 1766
rect 18052 1702 18104 1708
rect 18064 1494 18092 1702
rect 18052 1488 18104 1494
rect 18052 1430 18104 1436
rect 17736 1380 18000 1408
rect 17684 1362 17736 1368
rect 17960 1216 18012 1222
rect 17960 1158 18012 1164
rect 17592 1012 17644 1018
rect 17592 954 17644 960
rect 17972 882 18000 1158
rect 17960 876 18012 882
rect 17960 818 18012 824
rect 15844 808 15896 814
rect 15844 750 15896 756
rect 16120 808 16172 814
rect 16120 750 16172 756
rect 16580 808 16632 814
rect 16580 750 16632 756
rect 17408 808 17460 814
rect 17408 750 17460 756
rect 16764 672 16816 678
rect 16764 614 16816 620
rect 16856 672 16908 678
rect 16856 614 16908 620
rect 17408 672 17460 678
rect 17408 614 17460 620
rect 16364 572 16740 581
rect 16420 570 16444 572
rect 16500 570 16524 572
rect 16580 570 16604 572
rect 16660 570 16684 572
rect 16420 518 16430 570
rect 16674 518 16684 570
rect 16420 516 16444 518
rect 16500 516 16524 518
rect 16580 516 16604 518
rect 16660 516 16684 518
rect 16364 507 16740 516
rect 16592 428 16712 456
rect 16592 400 16620 428
rect 15384 332 15436 338
rect 15384 274 15436 280
rect 16578 0 16634 400
rect 16684 218 16712 428
rect 16776 406 16804 614
rect 16764 400 16816 406
rect 16764 342 16816 348
rect 16868 218 16896 614
rect 17420 400 17448 614
rect 16684 190 16896 218
rect 17406 0 17462 400
rect 18156 338 18184 1856
rect 18418 1799 18474 1808
rect 18892 1358 18920 2042
rect 18696 1352 18748 1358
rect 18696 1294 18748 1300
rect 18880 1352 18932 1358
rect 18880 1294 18932 1300
rect 18708 882 18736 1294
rect 18696 876 18748 882
rect 18696 818 18748 824
rect 18984 814 19012 2366
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 19364 2204 19740 2213
rect 19420 2202 19444 2204
rect 19500 2202 19524 2204
rect 19580 2202 19604 2204
rect 19660 2202 19684 2204
rect 19420 2150 19430 2202
rect 19674 2150 19684 2202
rect 19420 2148 19444 2150
rect 19500 2148 19524 2150
rect 19580 2148 19604 2150
rect 19660 2148 19684 2150
rect 19364 2139 19740 2148
rect 19340 1760 19392 1766
rect 19340 1702 19392 1708
rect 19352 1426 19380 1702
rect 19904 1562 19932 2246
rect 21100 1766 21128 4558
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21192 3738 21220 3878
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 21284 3602 21312 4626
rect 21376 4282 21404 5102
rect 21560 5030 21588 5306
rect 21836 5166 21864 5714
rect 21928 5166 21956 5714
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22112 5234 22140 5510
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21454 4584 21510 4593
rect 21454 4519 21510 4528
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21468 4078 21496 4519
rect 21560 4214 21588 4966
rect 21928 4826 21956 5102
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 21548 4208 21600 4214
rect 21548 4150 21600 4156
rect 21652 4078 21680 4694
rect 22112 4282 22140 5170
rect 22364 4924 22740 4933
rect 22420 4922 22444 4924
rect 22500 4922 22524 4924
rect 22580 4922 22604 4924
rect 22660 4922 22684 4924
rect 22420 4870 22430 4922
rect 22674 4870 22684 4922
rect 22420 4868 22444 4870
rect 22500 4868 22524 4870
rect 22580 4868 22604 4870
rect 22660 4868 22684 4870
rect 22364 4859 22740 4868
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 21546 3632 21602 3641
rect 21272 3596 21324 3602
rect 21324 3556 21404 3584
rect 21652 3618 21680 4014
rect 22020 4010 22048 4218
rect 22296 4078 22324 4762
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 21602 3590 21680 3618
rect 21546 3567 21602 3576
rect 21272 3538 21324 3544
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21284 2582 21312 2790
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 21376 2514 21404 3556
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 21454 2544 21510 2553
rect 21364 2508 21416 2514
rect 21454 2479 21510 2488
rect 21364 2450 21416 2456
rect 21088 1760 21140 1766
rect 21088 1702 21140 1708
rect 19892 1556 19944 1562
rect 19892 1498 19944 1504
rect 21376 1426 21404 2450
rect 21468 1426 21496 2479
rect 21744 2106 21772 3130
rect 21732 2100 21784 2106
rect 21732 2042 21784 2048
rect 22204 2038 22232 3946
rect 22364 3836 22740 3845
rect 22420 3834 22444 3836
rect 22500 3834 22524 3836
rect 22580 3834 22604 3836
rect 22660 3834 22684 3836
rect 22420 3782 22430 3834
rect 22674 3782 22684 3834
rect 22420 3780 22444 3782
rect 22500 3780 22524 3782
rect 22580 3780 22604 3782
rect 22660 3780 22684 3782
rect 22364 3771 22740 3780
rect 22848 3738 22876 4014
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22364 2748 22740 2757
rect 22420 2746 22444 2748
rect 22500 2746 22524 2748
rect 22580 2746 22604 2748
rect 22660 2746 22684 2748
rect 22420 2694 22430 2746
rect 22674 2694 22684 2746
rect 22420 2692 22444 2694
rect 22500 2692 22524 2694
rect 22580 2692 22604 2694
rect 22660 2692 22684 2694
rect 22364 2683 22740 2692
rect 22192 2032 22244 2038
rect 22192 1974 22244 1980
rect 22100 1964 22152 1970
rect 22100 1906 22152 1912
rect 21916 1896 21968 1902
rect 21916 1838 21968 1844
rect 19340 1420 19392 1426
rect 19340 1362 19392 1368
rect 19800 1420 19852 1426
rect 19800 1362 19852 1368
rect 21364 1420 21416 1426
rect 21364 1362 21416 1368
rect 21456 1420 21508 1426
rect 21456 1362 21508 1368
rect 19064 1284 19116 1290
rect 19064 1226 19116 1232
rect 19076 882 19104 1226
rect 19364 1116 19740 1125
rect 19420 1114 19444 1116
rect 19500 1114 19524 1116
rect 19580 1114 19604 1116
rect 19660 1114 19684 1116
rect 19420 1062 19430 1114
rect 19674 1062 19684 1114
rect 19420 1060 19444 1062
rect 19500 1060 19524 1062
rect 19580 1060 19604 1062
rect 19660 1060 19684 1062
rect 19364 1051 19740 1060
rect 19812 1018 19840 1362
rect 21928 1358 21956 1838
rect 22112 1494 22140 1906
rect 22100 1488 22152 1494
rect 22100 1430 22152 1436
rect 21916 1352 21968 1358
rect 21916 1294 21968 1300
rect 21640 1284 21692 1290
rect 21640 1226 21692 1232
rect 19800 1012 19852 1018
rect 19800 954 19852 960
rect 19064 876 19116 882
rect 19064 818 19116 824
rect 18972 808 19024 814
rect 18972 750 19024 756
rect 18420 672 18472 678
rect 18420 614 18472 620
rect 19064 672 19116 678
rect 19064 614 19116 620
rect 19892 672 19944 678
rect 19892 614 19944 620
rect 20720 672 20772 678
rect 20720 614 20772 620
rect 21548 672 21600 678
rect 21548 614 21600 620
rect 18432 490 18460 614
rect 18248 462 18460 490
rect 18248 400 18276 462
rect 19076 400 19104 614
rect 19904 400 19932 614
rect 20732 400 20760 614
rect 21560 400 21588 614
rect 21652 474 21680 1226
rect 22112 882 22140 1430
rect 22100 876 22152 882
rect 22100 818 22152 824
rect 22204 814 22232 1974
rect 22364 1660 22740 1669
rect 22420 1658 22444 1660
rect 22500 1658 22524 1660
rect 22580 1658 22604 1660
rect 22660 1658 22684 1660
rect 22420 1606 22430 1658
rect 22674 1606 22684 1658
rect 22420 1604 22444 1606
rect 22500 1604 22524 1606
rect 22580 1604 22604 1606
rect 22660 1604 22684 1606
rect 22364 1595 22740 1604
rect 22376 1556 22428 1562
rect 22376 1498 22428 1504
rect 22192 808 22244 814
rect 22388 762 22416 1498
rect 22192 750 22244 756
rect 22296 734 22416 762
rect 21640 468 21692 474
rect 22296 456 22324 734
rect 22364 572 22740 581
rect 22420 570 22444 572
rect 22500 570 22524 572
rect 22580 570 22604 572
rect 22660 570 22684 572
rect 22420 518 22430 570
rect 22674 518 22684 570
rect 22420 516 22444 518
rect 22500 516 22524 518
rect 22580 516 22604 518
rect 22660 516 22684 518
rect 22364 507 22740 516
rect 22296 428 22416 456
rect 21640 410 21692 416
rect 22388 400 22416 428
rect 18144 332 18196 338
rect 18144 274 18196 280
rect 18234 0 18290 400
rect 19062 0 19118 400
rect 19890 0 19946 400
rect 20718 0 20774 400
rect 21546 0 21602 400
rect 22374 0 22430 400
<< via2 >>
rect 1364 15258 1420 15260
rect 1444 15258 1500 15260
rect 1524 15258 1580 15260
rect 1604 15258 1660 15260
rect 1684 15258 1740 15260
rect 1364 15206 1366 15258
rect 1366 15206 1418 15258
rect 1418 15206 1420 15258
rect 1444 15206 1482 15258
rect 1482 15206 1494 15258
rect 1494 15206 1500 15258
rect 1524 15206 1546 15258
rect 1546 15206 1558 15258
rect 1558 15206 1580 15258
rect 1604 15206 1610 15258
rect 1610 15206 1622 15258
rect 1622 15206 1660 15258
rect 1684 15206 1686 15258
rect 1686 15206 1738 15258
rect 1738 15206 1740 15258
rect 1364 15204 1420 15206
rect 1444 15204 1500 15206
rect 1524 15204 1580 15206
rect 1604 15204 1660 15206
rect 1684 15204 1740 15206
rect 1364 14170 1420 14172
rect 1444 14170 1500 14172
rect 1524 14170 1580 14172
rect 1604 14170 1660 14172
rect 1684 14170 1740 14172
rect 1364 14118 1366 14170
rect 1366 14118 1418 14170
rect 1418 14118 1420 14170
rect 1444 14118 1482 14170
rect 1482 14118 1494 14170
rect 1494 14118 1500 14170
rect 1524 14118 1546 14170
rect 1546 14118 1558 14170
rect 1558 14118 1580 14170
rect 1604 14118 1610 14170
rect 1610 14118 1622 14170
rect 1622 14118 1660 14170
rect 1684 14118 1686 14170
rect 1686 14118 1738 14170
rect 1738 14118 1740 14170
rect 1364 14116 1420 14118
rect 1444 14116 1500 14118
rect 1524 14116 1580 14118
rect 1604 14116 1660 14118
rect 1684 14116 1740 14118
rect 4364 14714 4420 14716
rect 4444 14714 4500 14716
rect 4524 14714 4580 14716
rect 4604 14714 4660 14716
rect 4684 14714 4740 14716
rect 4364 14662 4366 14714
rect 4366 14662 4418 14714
rect 4418 14662 4420 14714
rect 4444 14662 4482 14714
rect 4482 14662 4494 14714
rect 4494 14662 4500 14714
rect 4524 14662 4546 14714
rect 4546 14662 4558 14714
rect 4558 14662 4580 14714
rect 4604 14662 4610 14714
rect 4610 14662 4622 14714
rect 4622 14662 4660 14714
rect 4684 14662 4686 14714
rect 4686 14662 4738 14714
rect 4738 14662 4740 14714
rect 4364 14660 4420 14662
rect 4444 14660 4500 14662
rect 4524 14660 4580 14662
rect 4604 14660 4660 14662
rect 4684 14660 4740 14662
rect 1364 13082 1420 13084
rect 1444 13082 1500 13084
rect 1524 13082 1580 13084
rect 1604 13082 1660 13084
rect 1684 13082 1740 13084
rect 1364 13030 1366 13082
rect 1366 13030 1418 13082
rect 1418 13030 1420 13082
rect 1444 13030 1482 13082
rect 1482 13030 1494 13082
rect 1494 13030 1500 13082
rect 1524 13030 1546 13082
rect 1546 13030 1558 13082
rect 1558 13030 1580 13082
rect 1604 13030 1610 13082
rect 1610 13030 1622 13082
rect 1622 13030 1660 13082
rect 1684 13030 1686 13082
rect 1686 13030 1738 13082
rect 1738 13030 1740 13082
rect 1364 13028 1420 13030
rect 1444 13028 1500 13030
rect 1524 13028 1580 13030
rect 1604 13028 1660 13030
rect 1684 13028 1740 13030
rect 1766 12688 1822 12744
rect 1858 12316 1860 12336
rect 1860 12316 1912 12336
rect 1912 12316 1914 12336
rect 1858 12280 1914 12316
rect 1364 11994 1420 11996
rect 1444 11994 1500 11996
rect 1524 11994 1580 11996
rect 1604 11994 1660 11996
rect 1684 11994 1740 11996
rect 1364 11942 1366 11994
rect 1366 11942 1418 11994
rect 1418 11942 1420 11994
rect 1444 11942 1482 11994
rect 1482 11942 1494 11994
rect 1494 11942 1500 11994
rect 1524 11942 1546 11994
rect 1546 11942 1558 11994
rect 1558 11942 1580 11994
rect 1604 11942 1610 11994
rect 1610 11942 1622 11994
rect 1622 11942 1660 11994
rect 1684 11942 1686 11994
rect 1686 11942 1738 11994
rect 1738 11942 1740 11994
rect 1364 11940 1420 11942
rect 1444 11940 1500 11942
rect 1524 11940 1580 11942
rect 1604 11940 1660 11942
rect 1684 11940 1740 11942
rect 1364 10906 1420 10908
rect 1444 10906 1500 10908
rect 1524 10906 1580 10908
rect 1604 10906 1660 10908
rect 1684 10906 1740 10908
rect 1364 10854 1366 10906
rect 1366 10854 1418 10906
rect 1418 10854 1420 10906
rect 1444 10854 1482 10906
rect 1482 10854 1494 10906
rect 1494 10854 1500 10906
rect 1524 10854 1546 10906
rect 1546 10854 1558 10906
rect 1558 10854 1580 10906
rect 1604 10854 1610 10906
rect 1610 10854 1622 10906
rect 1622 10854 1660 10906
rect 1684 10854 1686 10906
rect 1686 10854 1738 10906
rect 1738 10854 1740 10906
rect 1364 10852 1420 10854
rect 1444 10852 1500 10854
rect 1524 10852 1580 10854
rect 1604 10852 1660 10854
rect 1684 10852 1740 10854
rect 1674 10124 1730 10160
rect 1674 10104 1676 10124
rect 1676 10104 1728 10124
rect 1728 10104 1730 10124
rect 1364 9818 1420 9820
rect 1444 9818 1500 9820
rect 1524 9818 1580 9820
rect 1604 9818 1660 9820
rect 1684 9818 1740 9820
rect 1364 9766 1366 9818
rect 1366 9766 1418 9818
rect 1418 9766 1420 9818
rect 1444 9766 1482 9818
rect 1482 9766 1494 9818
rect 1494 9766 1500 9818
rect 1524 9766 1546 9818
rect 1546 9766 1558 9818
rect 1558 9766 1580 9818
rect 1604 9766 1610 9818
rect 1610 9766 1622 9818
rect 1622 9766 1660 9818
rect 1684 9766 1686 9818
rect 1686 9766 1738 9818
rect 1738 9766 1740 9818
rect 1364 9764 1420 9766
rect 1444 9764 1500 9766
rect 1524 9764 1580 9766
rect 1604 9764 1660 9766
rect 1684 9764 1740 9766
rect 1364 8730 1420 8732
rect 1444 8730 1500 8732
rect 1524 8730 1580 8732
rect 1604 8730 1660 8732
rect 1684 8730 1740 8732
rect 1364 8678 1366 8730
rect 1366 8678 1418 8730
rect 1418 8678 1420 8730
rect 1444 8678 1482 8730
rect 1482 8678 1494 8730
rect 1494 8678 1500 8730
rect 1524 8678 1546 8730
rect 1546 8678 1558 8730
rect 1558 8678 1580 8730
rect 1604 8678 1610 8730
rect 1610 8678 1622 8730
rect 1622 8678 1660 8730
rect 1684 8678 1686 8730
rect 1686 8678 1738 8730
rect 1738 8678 1740 8730
rect 1364 8676 1420 8678
rect 1444 8676 1500 8678
rect 1524 8676 1580 8678
rect 1604 8676 1660 8678
rect 1684 8676 1740 8678
rect 1364 7642 1420 7644
rect 1444 7642 1500 7644
rect 1524 7642 1580 7644
rect 1604 7642 1660 7644
rect 1684 7642 1740 7644
rect 1364 7590 1366 7642
rect 1366 7590 1418 7642
rect 1418 7590 1420 7642
rect 1444 7590 1482 7642
rect 1482 7590 1494 7642
rect 1494 7590 1500 7642
rect 1524 7590 1546 7642
rect 1546 7590 1558 7642
rect 1558 7590 1580 7642
rect 1604 7590 1610 7642
rect 1610 7590 1622 7642
rect 1622 7590 1660 7642
rect 1684 7590 1686 7642
rect 1686 7590 1738 7642
rect 1738 7590 1740 7642
rect 1364 7588 1420 7590
rect 1444 7588 1500 7590
rect 1524 7588 1580 7590
rect 1604 7588 1660 7590
rect 1684 7588 1740 7590
rect 2502 12300 2558 12336
rect 2502 12280 2504 12300
rect 2504 12280 2556 12300
rect 2556 12280 2558 12300
rect 2962 12724 2964 12744
rect 2964 12724 3016 12744
rect 3016 12724 3018 12744
rect 2962 12688 3018 12724
rect 1364 6554 1420 6556
rect 1444 6554 1500 6556
rect 1524 6554 1580 6556
rect 1604 6554 1660 6556
rect 1684 6554 1740 6556
rect 1364 6502 1366 6554
rect 1366 6502 1418 6554
rect 1418 6502 1420 6554
rect 1444 6502 1482 6554
rect 1482 6502 1494 6554
rect 1494 6502 1500 6554
rect 1524 6502 1546 6554
rect 1546 6502 1558 6554
rect 1558 6502 1580 6554
rect 1604 6502 1610 6554
rect 1610 6502 1622 6554
rect 1622 6502 1660 6554
rect 1684 6502 1686 6554
rect 1686 6502 1738 6554
rect 1738 6502 1740 6554
rect 1364 6500 1420 6502
rect 1444 6500 1500 6502
rect 1524 6500 1580 6502
rect 1604 6500 1660 6502
rect 1684 6500 1740 6502
rect 1364 5466 1420 5468
rect 1444 5466 1500 5468
rect 1524 5466 1580 5468
rect 1604 5466 1660 5468
rect 1684 5466 1740 5468
rect 1364 5414 1366 5466
rect 1366 5414 1418 5466
rect 1418 5414 1420 5466
rect 1444 5414 1482 5466
rect 1482 5414 1494 5466
rect 1494 5414 1500 5466
rect 1524 5414 1546 5466
rect 1546 5414 1558 5466
rect 1558 5414 1580 5466
rect 1604 5414 1610 5466
rect 1610 5414 1622 5466
rect 1622 5414 1660 5466
rect 1684 5414 1686 5466
rect 1686 5414 1738 5466
rect 1738 5414 1740 5466
rect 1364 5412 1420 5414
rect 1444 5412 1500 5414
rect 1524 5412 1580 5414
rect 1604 5412 1660 5414
rect 1684 5412 1740 5414
rect 2134 8608 2190 8664
rect 2594 11736 2650 11792
rect 3422 11736 3478 11792
rect 2962 11464 3018 11520
rect 2686 10512 2742 10568
rect 1364 4378 1420 4380
rect 1444 4378 1500 4380
rect 1524 4378 1580 4380
rect 1604 4378 1660 4380
rect 1684 4378 1740 4380
rect 1364 4326 1366 4378
rect 1366 4326 1418 4378
rect 1418 4326 1420 4378
rect 1444 4326 1482 4378
rect 1482 4326 1494 4378
rect 1494 4326 1500 4378
rect 1524 4326 1546 4378
rect 1546 4326 1558 4378
rect 1558 4326 1580 4378
rect 1604 4326 1610 4378
rect 1610 4326 1622 4378
rect 1622 4326 1660 4378
rect 1684 4326 1686 4378
rect 1686 4326 1738 4378
rect 1738 4326 1740 4378
rect 1364 4324 1420 4326
rect 1444 4324 1500 4326
rect 1524 4324 1580 4326
rect 1604 4324 1660 4326
rect 1684 4324 1740 4326
rect 1364 3290 1420 3292
rect 1444 3290 1500 3292
rect 1524 3290 1580 3292
rect 1604 3290 1660 3292
rect 1684 3290 1740 3292
rect 1364 3238 1366 3290
rect 1366 3238 1418 3290
rect 1418 3238 1420 3290
rect 1444 3238 1482 3290
rect 1482 3238 1494 3290
rect 1494 3238 1500 3290
rect 1524 3238 1546 3290
rect 1546 3238 1558 3290
rect 1558 3238 1580 3290
rect 1604 3238 1610 3290
rect 1610 3238 1622 3290
rect 1622 3238 1660 3290
rect 1684 3238 1686 3290
rect 1686 3238 1738 3290
rect 1738 3238 1740 3290
rect 1364 3236 1420 3238
rect 1444 3236 1500 3238
rect 1524 3236 1580 3238
rect 1604 3236 1660 3238
rect 1684 3236 1740 3238
rect 1582 2932 1584 2952
rect 1584 2932 1636 2952
rect 1636 2932 1638 2952
rect 1582 2896 1638 2932
rect 1364 2202 1420 2204
rect 1444 2202 1500 2204
rect 1524 2202 1580 2204
rect 1604 2202 1660 2204
rect 1684 2202 1740 2204
rect 1364 2150 1366 2202
rect 1366 2150 1418 2202
rect 1418 2150 1420 2202
rect 1444 2150 1482 2202
rect 1482 2150 1494 2202
rect 1494 2150 1500 2202
rect 1524 2150 1546 2202
rect 1546 2150 1558 2202
rect 1558 2150 1580 2202
rect 1604 2150 1610 2202
rect 1610 2150 1622 2202
rect 1622 2150 1660 2202
rect 1684 2150 1686 2202
rect 1686 2150 1738 2202
rect 1738 2150 1740 2202
rect 1364 2148 1420 2150
rect 1444 2148 1500 2150
rect 1524 2148 1580 2150
rect 1604 2148 1660 2150
rect 1684 2148 1740 2150
rect 1364 1114 1420 1116
rect 1444 1114 1500 1116
rect 1524 1114 1580 1116
rect 1604 1114 1660 1116
rect 1684 1114 1740 1116
rect 1364 1062 1366 1114
rect 1366 1062 1418 1114
rect 1418 1062 1420 1114
rect 1444 1062 1482 1114
rect 1482 1062 1494 1114
rect 1494 1062 1500 1114
rect 1524 1062 1546 1114
rect 1546 1062 1558 1114
rect 1558 1062 1580 1114
rect 1604 1062 1610 1114
rect 1610 1062 1622 1114
rect 1622 1062 1660 1114
rect 1684 1062 1686 1114
rect 1686 1062 1738 1114
rect 1738 1062 1740 1114
rect 1364 1060 1420 1062
rect 1444 1060 1500 1062
rect 1524 1060 1580 1062
rect 1604 1060 1660 1062
rect 1684 1060 1740 1062
rect 4364 13626 4420 13628
rect 4444 13626 4500 13628
rect 4524 13626 4580 13628
rect 4604 13626 4660 13628
rect 4684 13626 4740 13628
rect 4364 13574 4366 13626
rect 4366 13574 4418 13626
rect 4418 13574 4420 13626
rect 4444 13574 4482 13626
rect 4482 13574 4494 13626
rect 4494 13574 4500 13626
rect 4524 13574 4546 13626
rect 4546 13574 4558 13626
rect 4558 13574 4580 13626
rect 4604 13574 4610 13626
rect 4610 13574 4622 13626
rect 4622 13574 4660 13626
rect 4684 13574 4686 13626
rect 4686 13574 4738 13626
rect 4738 13574 4740 13626
rect 4364 13572 4420 13574
rect 4444 13572 4500 13574
rect 4524 13572 4580 13574
rect 4604 13572 4660 13574
rect 4684 13572 4740 13574
rect 4364 12538 4420 12540
rect 4444 12538 4500 12540
rect 4524 12538 4580 12540
rect 4604 12538 4660 12540
rect 4684 12538 4740 12540
rect 4364 12486 4366 12538
rect 4366 12486 4418 12538
rect 4418 12486 4420 12538
rect 4444 12486 4482 12538
rect 4482 12486 4494 12538
rect 4494 12486 4500 12538
rect 4524 12486 4546 12538
rect 4546 12486 4558 12538
rect 4558 12486 4580 12538
rect 4604 12486 4610 12538
rect 4610 12486 4622 12538
rect 4622 12486 4660 12538
rect 4684 12486 4686 12538
rect 4686 12486 4738 12538
rect 4738 12486 4740 12538
rect 4364 12484 4420 12486
rect 4444 12484 4500 12486
rect 4524 12484 4580 12486
rect 4604 12484 4660 12486
rect 4684 12484 4740 12486
rect 3054 8628 3110 8664
rect 3054 8608 3056 8628
rect 3056 8608 3108 8628
rect 3108 8608 3110 8628
rect 2870 7384 2926 7440
rect 3790 9560 3846 9616
rect 4364 11450 4420 11452
rect 4444 11450 4500 11452
rect 4524 11450 4580 11452
rect 4604 11450 4660 11452
rect 4684 11450 4740 11452
rect 4364 11398 4366 11450
rect 4366 11398 4418 11450
rect 4418 11398 4420 11450
rect 4444 11398 4482 11450
rect 4482 11398 4494 11450
rect 4494 11398 4500 11450
rect 4524 11398 4546 11450
rect 4546 11398 4558 11450
rect 4558 11398 4580 11450
rect 4604 11398 4610 11450
rect 4610 11398 4622 11450
rect 4622 11398 4660 11450
rect 4684 11398 4686 11450
rect 4686 11398 4738 11450
rect 4738 11398 4740 11450
rect 4364 11396 4420 11398
rect 4444 11396 4500 11398
rect 4524 11396 4580 11398
rect 4604 11396 4660 11398
rect 4684 11396 4740 11398
rect 4342 11076 4398 11112
rect 4342 11056 4344 11076
rect 4344 11056 4396 11076
rect 4396 11056 4398 11076
rect 4066 9968 4122 10024
rect 7364 15258 7420 15260
rect 7444 15258 7500 15260
rect 7524 15258 7580 15260
rect 7604 15258 7660 15260
rect 7684 15258 7740 15260
rect 7364 15206 7366 15258
rect 7366 15206 7418 15258
rect 7418 15206 7420 15258
rect 7444 15206 7482 15258
rect 7482 15206 7494 15258
rect 7494 15206 7500 15258
rect 7524 15206 7546 15258
rect 7546 15206 7558 15258
rect 7558 15206 7580 15258
rect 7604 15206 7610 15258
rect 7610 15206 7622 15258
rect 7622 15206 7660 15258
rect 7684 15206 7686 15258
rect 7686 15206 7738 15258
rect 7738 15206 7740 15258
rect 7364 15204 7420 15206
rect 7444 15204 7500 15206
rect 7524 15204 7580 15206
rect 7604 15204 7660 15206
rect 7684 15204 7740 15206
rect 13364 15258 13420 15260
rect 13444 15258 13500 15260
rect 13524 15258 13580 15260
rect 13604 15258 13660 15260
rect 13684 15258 13740 15260
rect 13364 15206 13366 15258
rect 13366 15206 13418 15258
rect 13418 15206 13420 15258
rect 13444 15206 13482 15258
rect 13482 15206 13494 15258
rect 13494 15206 13500 15258
rect 13524 15206 13546 15258
rect 13546 15206 13558 15258
rect 13558 15206 13580 15258
rect 13604 15206 13610 15258
rect 13610 15206 13622 15258
rect 13622 15206 13660 15258
rect 13684 15206 13686 15258
rect 13686 15206 13738 15258
rect 13738 15206 13740 15258
rect 13364 15204 13420 15206
rect 13444 15204 13500 15206
rect 13524 15204 13580 15206
rect 13604 15204 13660 15206
rect 13684 15204 13740 15206
rect 4894 11192 4950 11248
rect 4364 10362 4420 10364
rect 4444 10362 4500 10364
rect 4524 10362 4580 10364
rect 4604 10362 4660 10364
rect 4684 10362 4740 10364
rect 4364 10310 4366 10362
rect 4366 10310 4418 10362
rect 4418 10310 4420 10362
rect 4444 10310 4482 10362
rect 4482 10310 4494 10362
rect 4494 10310 4500 10362
rect 4524 10310 4546 10362
rect 4546 10310 4558 10362
rect 4558 10310 4580 10362
rect 4604 10310 4610 10362
rect 4610 10310 4622 10362
rect 4622 10310 4660 10362
rect 4684 10310 4686 10362
rect 4686 10310 4738 10362
rect 4738 10310 4740 10362
rect 4364 10308 4420 10310
rect 4444 10308 4500 10310
rect 4524 10308 4580 10310
rect 4604 10308 4660 10310
rect 4684 10308 4740 10310
rect 3514 7948 3570 7984
rect 3514 7928 3516 7948
rect 3516 7928 3568 7948
rect 3568 7928 3570 7948
rect 4364 9274 4420 9276
rect 4444 9274 4500 9276
rect 4524 9274 4580 9276
rect 4604 9274 4660 9276
rect 4684 9274 4740 9276
rect 4364 9222 4366 9274
rect 4366 9222 4418 9274
rect 4418 9222 4420 9274
rect 4444 9222 4482 9274
rect 4482 9222 4494 9274
rect 4494 9222 4500 9274
rect 4524 9222 4546 9274
rect 4546 9222 4558 9274
rect 4558 9222 4580 9274
rect 4604 9222 4610 9274
rect 4610 9222 4622 9274
rect 4622 9222 4660 9274
rect 4684 9222 4686 9274
rect 4686 9222 4738 9274
rect 4738 9222 4740 9274
rect 4364 9220 4420 9222
rect 4444 9220 4500 9222
rect 4524 9220 4580 9222
rect 4604 9220 4660 9222
rect 4684 9220 4740 9222
rect 4066 7420 4068 7440
rect 4068 7420 4120 7440
rect 4120 7420 4122 7440
rect 4066 7384 4122 7420
rect 4364 8186 4420 8188
rect 4444 8186 4500 8188
rect 4524 8186 4580 8188
rect 4604 8186 4660 8188
rect 4684 8186 4740 8188
rect 4364 8134 4366 8186
rect 4366 8134 4418 8186
rect 4418 8134 4420 8186
rect 4444 8134 4482 8186
rect 4482 8134 4494 8186
rect 4494 8134 4500 8186
rect 4524 8134 4546 8186
rect 4546 8134 4558 8186
rect 4558 8134 4580 8186
rect 4604 8134 4610 8186
rect 4610 8134 4622 8186
rect 4622 8134 4660 8186
rect 4684 8134 4686 8186
rect 4686 8134 4738 8186
rect 4738 8134 4740 8186
rect 4364 8132 4420 8134
rect 4444 8132 4500 8134
rect 4524 8132 4580 8134
rect 4604 8132 4660 8134
rect 4684 8132 4740 8134
rect 4364 7098 4420 7100
rect 4444 7098 4500 7100
rect 4524 7098 4580 7100
rect 4604 7098 4660 7100
rect 4684 7098 4740 7100
rect 4364 7046 4366 7098
rect 4366 7046 4418 7098
rect 4418 7046 4420 7098
rect 4444 7046 4482 7098
rect 4482 7046 4494 7098
rect 4494 7046 4500 7098
rect 4524 7046 4546 7098
rect 4546 7046 4558 7098
rect 4558 7046 4580 7098
rect 4604 7046 4610 7098
rect 4610 7046 4622 7098
rect 4622 7046 4660 7098
rect 4684 7046 4686 7098
rect 4686 7046 4738 7098
rect 4738 7046 4740 7098
rect 4364 7044 4420 7046
rect 4444 7044 4500 7046
rect 4524 7044 4580 7046
rect 4604 7044 4660 7046
rect 4684 7044 4740 7046
rect 5170 11600 5226 11656
rect 5354 11328 5410 11384
rect 5538 7384 5594 7440
rect 4364 6010 4420 6012
rect 4444 6010 4500 6012
rect 4524 6010 4580 6012
rect 4604 6010 4660 6012
rect 4684 6010 4740 6012
rect 4364 5958 4366 6010
rect 4366 5958 4418 6010
rect 4418 5958 4420 6010
rect 4444 5958 4482 6010
rect 4482 5958 4494 6010
rect 4494 5958 4500 6010
rect 4524 5958 4546 6010
rect 4546 5958 4558 6010
rect 4558 5958 4580 6010
rect 4604 5958 4610 6010
rect 4610 5958 4622 6010
rect 4622 5958 4660 6010
rect 4684 5958 4686 6010
rect 4686 5958 4738 6010
rect 4738 5958 4740 6010
rect 4364 5956 4420 5958
rect 4444 5956 4500 5958
rect 4524 5956 4580 5958
rect 4604 5956 4660 5958
rect 4684 5956 4740 5958
rect 4364 4922 4420 4924
rect 4444 4922 4500 4924
rect 4524 4922 4580 4924
rect 4604 4922 4660 4924
rect 4684 4922 4740 4924
rect 4364 4870 4366 4922
rect 4366 4870 4418 4922
rect 4418 4870 4420 4922
rect 4444 4870 4482 4922
rect 4482 4870 4494 4922
rect 4494 4870 4500 4922
rect 4524 4870 4546 4922
rect 4546 4870 4558 4922
rect 4558 4870 4580 4922
rect 4604 4870 4610 4922
rect 4610 4870 4622 4922
rect 4622 4870 4660 4922
rect 4684 4870 4686 4922
rect 4686 4870 4738 4922
rect 4738 4870 4740 4922
rect 4364 4868 4420 4870
rect 4444 4868 4500 4870
rect 4524 4868 4580 4870
rect 4604 4868 4660 4870
rect 4684 4868 4740 4870
rect 4364 3834 4420 3836
rect 4444 3834 4500 3836
rect 4524 3834 4580 3836
rect 4604 3834 4660 3836
rect 4684 3834 4740 3836
rect 4364 3782 4366 3834
rect 4366 3782 4418 3834
rect 4418 3782 4420 3834
rect 4444 3782 4482 3834
rect 4482 3782 4494 3834
rect 4494 3782 4500 3834
rect 4524 3782 4546 3834
rect 4546 3782 4558 3834
rect 4558 3782 4580 3834
rect 4604 3782 4610 3834
rect 4610 3782 4622 3834
rect 4622 3782 4660 3834
rect 4684 3782 4686 3834
rect 4686 3782 4738 3834
rect 4738 3782 4740 3834
rect 4364 3780 4420 3782
rect 4444 3780 4500 3782
rect 4524 3780 4580 3782
rect 4604 3780 4660 3782
rect 4684 3780 4740 3782
rect 7364 14170 7420 14172
rect 7444 14170 7500 14172
rect 7524 14170 7580 14172
rect 7604 14170 7660 14172
rect 7684 14170 7740 14172
rect 7364 14118 7366 14170
rect 7366 14118 7418 14170
rect 7418 14118 7420 14170
rect 7444 14118 7482 14170
rect 7482 14118 7494 14170
rect 7494 14118 7500 14170
rect 7524 14118 7546 14170
rect 7546 14118 7558 14170
rect 7558 14118 7580 14170
rect 7604 14118 7610 14170
rect 7610 14118 7622 14170
rect 7622 14118 7660 14170
rect 7684 14118 7686 14170
rect 7686 14118 7738 14170
rect 7738 14118 7740 14170
rect 7364 14116 7420 14118
rect 7444 14116 7500 14118
rect 7524 14116 7580 14118
rect 7604 14116 7660 14118
rect 7684 14116 7740 14118
rect 8114 13232 8170 13288
rect 7364 13082 7420 13084
rect 7444 13082 7500 13084
rect 7524 13082 7580 13084
rect 7604 13082 7660 13084
rect 7684 13082 7740 13084
rect 7364 13030 7366 13082
rect 7366 13030 7418 13082
rect 7418 13030 7420 13082
rect 7444 13030 7482 13082
rect 7482 13030 7494 13082
rect 7494 13030 7500 13082
rect 7524 13030 7546 13082
rect 7546 13030 7558 13082
rect 7558 13030 7580 13082
rect 7604 13030 7610 13082
rect 7610 13030 7622 13082
rect 7622 13030 7660 13082
rect 7684 13030 7686 13082
rect 7686 13030 7738 13082
rect 7738 13030 7740 13082
rect 7364 13028 7420 13030
rect 7444 13028 7500 13030
rect 7524 13028 7580 13030
rect 7604 13028 7660 13030
rect 7684 13028 7740 13030
rect 6826 11620 6882 11656
rect 6826 11600 6828 11620
rect 6828 11600 6880 11620
rect 6880 11600 6882 11620
rect 7194 11056 7250 11112
rect 6918 10376 6974 10432
rect 7364 11994 7420 11996
rect 7444 11994 7500 11996
rect 7524 11994 7580 11996
rect 7604 11994 7660 11996
rect 7684 11994 7740 11996
rect 7364 11942 7366 11994
rect 7366 11942 7418 11994
rect 7418 11942 7420 11994
rect 7444 11942 7482 11994
rect 7482 11942 7494 11994
rect 7494 11942 7500 11994
rect 7524 11942 7546 11994
rect 7546 11942 7558 11994
rect 7558 11942 7580 11994
rect 7604 11942 7610 11994
rect 7610 11942 7622 11994
rect 7622 11942 7660 11994
rect 7684 11942 7686 11994
rect 7686 11942 7738 11994
rect 7738 11942 7740 11994
rect 7364 11940 7420 11942
rect 7444 11940 7500 11942
rect 7524 11940 7580 11942
rect 7604 11940 7660 11942
rect 7684 11940 7740 11942
rect 7364 10906 7420 10908
rect 7444 10906 7500 10908
rect 7524 10906 7580 10908
rect 7604 10906 7660 10908
rect 7684 10906 7740 10908
rect 7364 10854 7366 10906
rect 7366 10854 7418 10906
rect 7418 10854 7420 10906
rect 7444 10854 7482 10906
rect 7482 10854 7494 10906
rect 7494 10854 7500 10906
rect 7524 10854 7546 10906
rect 7546 10854 7558 10906
rect 7558 10854 7580 10906
rect 7604 10854 7610 10906
rect 7610 10854 7622 10906
rect 7622 10854 7660 10906
rect 7684 10854 7686 10906
rect 7686 10854 7738 10906
rect 7738 10854 7740 10906
rect 7364 10852 7420 10854
rect 7444 10852 7500 10854
rect 7524 10852 7580 10854
rect 7604 10852 7660 10854
rect 7684 10852 7740 10854
rect 8206 10648 8262 10704
rect 7364 9818 7420 9820
rect 7444 9818 7500 9820
rect 7524 9818 7580 9820
rect 7604 9818 7660 9820
rect 7684 9818 7740 9820
rect 7364 9766 7366 9818
rect 7366 9766 7418 9818
rect 7418 9766 7420 9818
rect 7444 9766 7482 9818
rect 7482 9766 7494 9818
rect 7494 9766 7500 9818
rect 7524 9766 7546 9818
rect 7546 9766 7558 9818
rect 7558 9766 7580 9818
rect 7604 9766 7610 9818
rect 7610 9766 7622 9818
rect 7622 9766 7660 9818
rect 7684 9766 7686 9818
rect 7686 9766 7738 9818
rect 7738 9766 7740 9818
rect 7364 9764 7420 9766
rect 7444 9764 7500 9766
rect 7524 9764 7580 9766
rect 7604 9764 7660 9766
rect 7684 9764 7740 9766
rect 7364 8730 7420 8732
rect 7444 8730 7500 8732
rect 7524 8730 7580 8732
rect 7604 8730 7660 8732
rect 7684 8730 7740 8732
rect 7364 8678 7366 8730
rect 7366 8678 7418 8730
rect 7418 8678 7420 8730
rect 7444 8678 7482 8730
rect 7482 8678 7494 8730
rect 7494 8678 7500 8730
rect 7524 8678 7546 8730
rect 7546 8678 7558 8730
rect 7558 8678 7580 8730
rect 7604 8678 7610 8730
rect 7610 8678 7622 8730
rect 7622 8678 7660 8730
rect 7684 8678 7686 8730
rect 7686 8678 7738 8730
rect 7738 8678 7740 8730
rect 7364 8676 7420 8678
rect 7444 8676 7500 8678
rect 7524 8676 7580 8678
rect 7604 8676 7660 8678
rect 7684 8676 7740 8678
rect 7364 7642 7420 7644
rect 7444 7642 7500 7644
rect 7524 7642 7580 7644
rect 7604 7642 7660 7644
rect 7684 7642 7740 7644
rect 7364 7590 7366 7642
rect 7366 7590 7418 7642
rect 7418 7590 7420 7642
rect 7444 7590 7482 7642
rect 7482 7590 7494 7642
rect 7494 7590 7500 7642
rect 7524 7590 7546 7642
rect 7546 7590 7558 7642
rect 7558 7590 7580 7642
rect 7604 7590 7610 7642
rect 7610 7590 7622 7642
rect 7622 7590 7660 7642
rect 7684 7590 7686 7642
rect 7686 7590 7738 7642
rect 7738 7590 7740 7642
rect 7364 7588 7420 7590
rect 7444 7588 7500 7590
rect 7524 7588 7580 7590
rect 7604 7588 7660 7590
rect 7684 7588 7740 7590
rect 7364 6554 7420 6556
rect 7444 6554 7500 6556
rect 7524 6554 7580 6556
rect 7604 6554 7660 6556
rect 7684 6554 7740 6556
rect 7364 6502 7366 6554
rect 7366 6502 7418 6554
rect 7418 6502 7420 6554
rect 7444 6502 7482 6554
rect 7482 6502 7494 6554
rect 7494 6502 7500 6554
rect 7524 6502 7546 6554
rect 7546 6502 7558 6554
rect 7558 6502 7580 6554
rect 7604 6502 7610 6554
rect 7610 6502 7622 6554
rect 7622 6502 7660 6554
rect 7684 6502 7686 6554
rect 7686 6502 7738 6554
rect 7738 6502 7740 6554
rect 7364 6500 7420 6502
rect 7444 6500 7500 6502
rect 7524 6500 7580 6502
rect 7604 6500 7660 6502
rect 7684 6500 7740 6502
rect 6090 4548 6146 4584
rect 6090 4528 6092 4548
rect 6092 4528 6144 4548
rect 6144 4528 6146 4548
rect 6642 3576 6698 3632
rect 7364 5466 7420 5468
rect 7444 5466 7500 5468
rect 7524 5466 7580 5468
rect 7604 5466 7660 5468
rect 7684 5466 7740 5468
rect 7364 5414 7366 5466
rect 7366 5414 7418 5466
rect 7418 5414 7420 5466
rect 7444 5414 7482 5466
rect 7482 5414 7494 5466
rect 7494 5414 7500 5466
rect 7524 5414 7546 5466
rect 7546 5414 7558 5466
rect 7558 5414 7580 5466
rect 7604 5414 7610 5466
rect 7610 5414 7622 5466
rect 7622 5414 7660 5466
rect 7684 5414 7686 5466
rect 7686 5414 7738 5466
rect 7738 5414 7740 5466
rect 7364 5412 7420 5414
rect 7444 5412 7500 5414
rect 7524 5412 7580 5414
rect 7604 5412 7660 5414
rect 7684 5412 7740 5414
rect 7286 5208 7342 5264
rect 7746 4564 7748 4584
rect 7748 4564 7800 4584
rect 7800 4564 7802 4584
rect 7746 4528 7802 4564
rect 7364 4378 7420 4380
rect 7444 4378 7500 4380
rect 7524 4378 7580 4380
rect 7604 4378 7660 4380
rect 7684 4378 7740 4380
rect 7364 4326 7366 4378
rect 7366 4326 7418 4378
rect 7418 4326 7420 4378
rect 7444 4326 7482 4378
rect 7482 4326 7494 4378
rect 7494 4326 7500 4378
rect 7524 4326 7546 4378
rect 7546 4326 7558 4378
rect 7558 4326 7580 4378
rect 7604 4326 7610 4378
rect 7610 4326 7622 4378
rect 7622 4326 7660 4378
rect 7684 4326 7686 4378
rect 7686 4326 7738 4378
rect 7738 4326 7740 4378
rect 7364 4324 7420 4326
rect 7444 4324 7500 4326
rect 7524 4324 7580 4326
rect 7604 4324 7660 4326
rect 7684 4324 7740 4326
rect 7010 3440 7066 3496
rect 4364 2746 4420 2748
rect 4444 2746 4500 2748
rect 4524 2746 4580 2748
rect 4604 2746 4660 2748
rect 4684 2746 4740 2748
rect 4066 2488 4122 2544
rect 4364 2694 4366 2746
rect 4366 2694 4418 2746
rect 4418 2694 4420 2746
rect 4444 2694 4482 2746
rect 4482 2694 4494 2746
rect 4494 2694 4500 2746
rect 4524 2694 4546 2746
rect 4546 2694 4558 2746
rect 4558 2694 4580 2746
rect 4604 2694 4610 2746
rect 4610 2694 4622 2746
rect 4622 2694 4660 2746
rect 4684 2694 4686 2746
rect 4686 2694 4738 2746
rect 4738 2694 4740 2746
rect 4364 2692 4420 2694
rect 4444 2692 4500 2694
rect 4524 2692 4580 2694
rect 4604 2692 4660 2694
rect 4684 2692 4740 2694
rect 7364 3290 7420 3292
rect 7444 3290 7500 3292
rect 7524 3290 7580 3292
rect 7604 3290 7660 3292
rect 7684 3290 7740 3292
rect 7364 3238 7366 3290
rect 7366 3238 7418 3290
rect 7418 3238 7420 3290
rect 7444 3238 7482 3290
rect 7482 3238 7494 3290
rect 7494 3238 7500 3290
rect 7524 3238 7546 3290
rect 7546 3238 7558 3290
rect 7558 3238 7580 3290
rect 7604 3238 7610 3290
rect 7610 3238 7622 3290
rect 7622 3238 7660 3290
rect 7684 3238 7686 3290
rect 7686 3238 7738 3290
rect 7738 3238 7740 3290
rect 7364 3236 7420 3238
rect 7444 3236 7500 3238
rect 7524 3236 7580 3238
rect 7604 3236 7660 3238
rect 7684 3236 7740 3238
rect 8022 3712 8078 3768
rect 8206 5616 8262 5672
rect 8206 4664 8262 4720
rect 7838 2916 7894 2952
rect 7838 2896 7840 2916
rect 7840 2896 7892 2916
rect 7892 2896 7894 2916
rect 4342 1828 4398 1864
rect 4342 1808 4344 1828
rect 4344 1808 4396 1828
rect 4396 1808 4398 1828
rect 4364 1658 4420 1660
rect 4444 1658 4500 1660
rect 4524 1658 4580 1660
rect 4604 1658 4660 1660
rect 4684 1658 4740 1660
rect 4364 1606 4366 1658
rect 4366 1606 4418 1658
rect 4418 1606 4420 1658
rect 4444 1606 4482 1658
rect 4482 1606 4494 1658
rect 4494 1606 4500 1658
rect 4524 1606 4546 1658
rect 4546 1606 4558 1658
rect 4558 1606 4580 1658
rect 4604 1606 4610 1658
rect 4610 1606 4622 1658
rect 4622 1606 4660 1658
rect 4684 1606 4686 1658
rect 4686 1606 4738 1658
rect 4738 1606 4740 1658
rect 4364 1604 4420 1606
rect 4444 1604 4500 1606
rect 4524 1604 4580 1606
rect 4604 1604 4660 1606
rect 4684 1604 4740 1606
rect 7364 2202 7420 2204
rect 7444 2202 7500 2204
rect 7524 2202 7580 2204
rect 7604 2202 7660 2204
rect 7684 2202 7740 2204
rect 7364 2150 7366 2202
rect 7366 2150 7418 2202
rect 7418 2150 7420 2202
rect 7444 2150 7482 2202
rect 7482 2150 7494 2202
rect 7494 2150 7500 2202
rect 7524 2150 7546 2202
rect 7546 2150 7558 2202
rect 7558 2150 7580 2202
rect 7604 2150 7610 2202
rect 7610 2150 7622 2202
rect 7622 2150 7660 2202
rect 7684 2150 7686 2202
rect 7686 2150 7738 2202
rect 7738 2150 7740 2202
rect 7364 2148 7420 2150
rect 7444 2148 7500 2150
rect 7524 2148 7580 2150
rect 7604 2148 7660 2150
rect 7684 2148 7740 2150
rect 7562 1944 7618 2000
rect 4364 570 4420 572
rect 4444 570 4500 572
rect 4524 570 4580 572
rect 4604 570 4660 572
rect 4684 570 4740 572
rect 4364 518 4366 570
rect 4366 518 4418 570
rect 4418 518 4420 570
rect 4444 518 4482 570
rect 4482 518 4494 570
rect 4494 518 4500 570
rect 4524 518 4546 570
rect 4546 518 4558 570
rect 4558 518 4580 570
rect 4604 518 4610 570
rect 4610 518 4622 570
rect 4622 518 4660 570
rect 4684 518 4686 570
rect 4686 518 4738 570
rect 4738 518 4740 570
rect 4364 516 4420 518
rect 4444 516 4500 518
rect 4524 516 4580 518
rect 4604 516 4660 518
rect 4684 516 4740 518
rect 8574 2080 8630 2136
rect 9034 9696 9090 9752
rect 9494 12824 9550 12880
rect 9402 10376 9458 10432
rect 9494 8336 9550 8392
rect 9126 7928 9182 7984
rect 10364 14714 10420 14716
rect 10444 14714 10500 14716
rect 10524 14714 10580 14716
rect 10604 14714 10660 14716
rect 10684 14714 10740 14716
rect 10364 14662 10366 14714
rect 10366 14662 10418 14714
rect 10418 14662 10420 14714
rect 10444 14662 10482 14714
rect 10482 14662 10494 14714
rect 10494 14662 10500 14714
rect 10524 14662 10546 14714
rect 10546 14662 10558 14714
rect 10558 14662 10580 14714
rect 10604 14662 10610 14714
rect 10610 14662 10622 14714
rect 10622 14662 10660 14714
rect 10684 14662 10686 14714
rect 10686 14662 10738 14714
rect 10738 14662 10740 14714
rect 10364 14660 10420 14662
rect 10444 14660 10500 14662
rect 10524 14660 10580 14662
rect 10604 14660 10660 14662
rect 10684 14660 10740 14662
rect 9678 12688 9734 12744
rect 9770 12008 9826 12064
rect 10506 13776 10562 13832
rect 10364 13626 10420 13628
rect 10444 13626 10500 13628
rect 10524 13626 10580 13628
rect 10604 13626 10660 13628
rect 10684 13626 10740 13628
rect 10364 13574 10366 13626
rect 10366 13574 10418 13626
rect 10418 13574 10420 13626
rect 10444 13574 10482 13626
rect 10482 13574 10494 13626
rect 10494 13574 10500 13626
rect 10524 13574 10546 13626
rect 10546 13574 10558 13626
rect 10558 13574 10580 13626
rect 10604 13574 10610 13626
rect 10610 13574 10622 13626
rect 10622 13574 10660 13626
rect 10684 13574 10686 13626
rect 10686 13574 10738 13626
rect 10738 13574 10740 13626
rect 10364 13572 10420 13574
rect 10444 13572 10500 13574
rect 10524 13572 10580 13574
rect 10604 13572 10660 13574
rect 10684 13572 10740 13574
rect 9862 8744 9918 8800
rect 9126 3712 9182 3768
rect 9586 7384 9642 7440
rect 9678 6704 9734 6760
rect 9586 6160 9642 6216
rect 9586 3848 9642 3904
rect 9862 8472 9918 8528
rect 10138 12280 10194 12336
rect 10364 12538 10420 12540
rect 10444 12538 10500 12540
rect 10524 12538 10580 12540
rect 10604 12538 10660 12540
rect 10684 12538 10740 12540
rect 10364 12486 10366 12538
rect 10366 12486 10418 12538
rect 10418 12486 10420 12538
rect 10444 12486 10482 12538
rect 10482 12486 10494 12538
rect 10494 12486 10500 12538
rect 10524 12486 10546 12538
rect 10546 12486 10558 12538
rect 10558 12486 10580 12538
rect 10604 12486 10610 12538
rect 10610 12486 10622 12538
rect 10622 12486 10660 12538
rect 10684 12486 10686 12538
rect 10686 12486 10738 12538
rect 10738 12486 10740 12538
rect 10364 12484 10420 12486
rect 10444 12484 10500 12486
rect 10524 12484 10580 12486
rect 10604 12484 10660 12486
rect 10684 12484 10740 12486
rect 11794 13268 11796 13288
rect 11796 13268 11848 13288
rect 11848 13268 11850 13288
rect 11794 13232 11850 13268
rect 11150 12688 11206 12744
rect 11150 12552 11206 12608
rect 10598 12144 10654 12200
rect 10364 11450 10420 11452
rect 10444 11450 10500 11452
rect 10524 11450 10580 11452
rect 10604 11450 10660 11452
rect 10684 11450 10740 11452
rect 10364 11398 10366 11450
rect 10366 11398 10418 11450
rect 10418 11398 10420 11450
rect 10444 11398 10482 11450
rect 10482 11398 10494 11450
rect 10494 11398 10500 11450
rect 10524 11398 10546 11450
rect 10546 11398 10558 11450
rect 10558 11398 10580 11450
rect 10604 11398 10610 11450
rect 10610 11398 10622 11450
rect 10622 11398 10660 11450
rect 10684 11398 10686 11450
rect 10686 11398 10738 11450
rect 10738 11398 10740 11450
rect 10364 11396 10420 11398
rect 10444 11396 10500 11398
rect 10524 11396 10580 11398
rect 10604 11396 10660 11398
rect 10684 11396 10740 11398
rect 10364 10362 10420 10364
rect 10444 10362 10500 10364
rect 10524 10362 10580 10364
rect 10604 10362 10660 10364
rect 10684 10362 10740 10364
rect 10364 10310 10366 10362
rect 10366 10310 10418 10362
rect 10418 10310 10420 10362
rect 10444 10310 10482 10362
rect 10482 10310 10494 10362
rect 10494 10310 10500 10362
rect 10524 10310 10546 10362
rect 10546 10310 10558 10362
rect 10558 10310 10580 10362
rect 10604 10310 10610 10362
rect 10610 10310 10622 10362
rect 10622 10310 10660 10362
rect 10684 10310 10686 10362
rect 10686 10310 10738 10362
rect 10738 10310 10740 10362
rect 10364 10308 10420 10310
rect 10444 10308 10500 10310
rect 10524 10308 10580 10310
rect 10604 10308 10660 10310
rect 10684 10308 10740 10310
rect 11150 11328 11206 11384
rect 11518 12280 11574 12336
rect 11610 12008 11666 12064
rect 10690 9424 10746 9480
rect 10364 9274 10420 9276
rect 10444 9274 10500 9276
rect 10524 9274 10580 9276
rect 10604 9274 10660 9276
rect 10684 9274 10740 9276
rect 10364 9222 10366 9274
rect 10366 9222 10418 9274
rect 10418 9222 10420 9274
rect 10444 9222 10482 9274
rect 10482 9222 10494 9274
rect 10494 9222 10500 9274
rect 10524 9222 10546 9274
rect 10546 9222 10558 9274
rect 10558 9222 10580 9274
rect 10604 9222 10610 9274
rect 10610 9222 10622 9274
rect 10622 9222 10660 9274
rect 10684 9222 10686 9274
rect 10686 9222 10738 9274
rect 10738 9222 10740 9274
rect 10364 9220 10420 9222
rect 10444 9220 10500 9222
rect 10524 9220 10580 9222
rect 10604 9220 10660 9222
rect 10684 9220 10740 9222
rect 10230 8900 10286 8936
rect 10230 8880 10232 8900
rect 10232 8880 10284 8900
rect 10284 8880 10286 8900
rect 10364 8186 10420 8188
rect 10444 8186 10500 8188
rect 10524 8186 10580 8188
rect 10604 8186 10660 8188
rect 10684 8186 10740 8188
rect 10364 8134 10366 8186
rect 10366 8134 10418 8186
rect 10418 8134 10420 8186
rect 10444 8134 10482 8186
rect 10482 8134 10494 8186
rect 10494 8134 10500 8186
rect 10524 8134 10546 8186
rect 10546 8134 10558 8186
rect 10558 8134 10580 8186
rect 10604 8134 10610 8186
rect 10610 8134 10622 8186
rect 10622 8134 10660 8186
rect 10684 8134 10686 8186
rect 10686 8134 10738 8186
rect 10738 8134 10740 8186
rect 10364 8132 10420 8134
rect 10444 8132 10500 8134
rect 10524 8132 10580 8134
rect 10604 8132 10660 8134
rect 10684 8132 10740 8134
rect 10230 7520 10286 7576
rect 10364 7098 10420 7100
rect 10444 7098 10500 7100
rect 10524 7098 10580 7100
rect 10604 7098 10660 7100
rect 10684 7098 10740 7100
rect 10364 7046 10366 7098
rect 10366 7046 10418 7098
rect 10418 7046 10420 7098
rect 10444 7046 10482 7098
rect 10482 7046 10494 7098
rect 10494 7046 10500 7098
rect 10524 7046 10546 7098
rect 10546 7046 10558 7098
rect 10558 7046 10580 7098
rect 10604 7046 10610 7098
rect 10610 7046 10622 7098
rect 10622 7046 10660 7098
rect 10684 7046 10686 7098
rect 10686 7046 10738 7098
rect 10738 7046 10740 7098
rect 10364 7044 10420 7046
rect 10444 7044 10500 7046
rect 10524 7044 10580 7046
rect 10604 7044 10660 7046
rect 10684 7044 10740 7046
rect 10506 6568 10562 6624
rect 10046 5344 10102 5400
rect 10364 6010 10420 6012
rect 10444 6010 10500 6012
rect 10524 6010 10580 6012
rect 10604 6010 10660 6012
rect 10684 6010 10740 6012
rect 10364 5958 10366 6010
rect 10366 5958 10418 6010
rect 10418 5958 10420 6010
rect 10444 5958 10482 6010
rect 10482 5958 10494 6010
rect 10494 5958 10500 6010
rect 10524 5958 10546 6010
rect 10546 5958 10558 6010
rect 10558 5958 10580 6010
rect 10604 5958 10610 6010
rect 10610 5958 10622 6010
rect 10622 5958 10660 6010
rect 10684 5958 10686 6010
rect 10686 5958 10738 6010
rect 10738 5958 10740 6010
rect 10364 5956 10420 5958
rect 10444 5956 10500 5958
rect 10524 5956 10580 5958
rect 10604 5956 10660 5958
rect 10684 5956 10740 5958
rect 10874 6316 10930 6352
rect 10874 6296 10876 6316
rect 10876 6296 10928 6316
rect 10928 6296 10930 6316
rect 10874 6024 10930 6080
rect 10364 4922 10420 4924
rect 10444 4922 10500 4924
rect 10524 4922 10580 4924
rect 10604 4922 10660 4924
rect 10684 4922 10740 4924
rect 10364 4870 10366 4922
rect 10366 4870 10418 4922
rect 10418 4870 10420 4922
rect 10444 4870 10482 4922
rect 10482 4870 10494 4922
rect 10494 4870 10500 4922
rect 10524 4870 10546 4922
rect 10546 4870 10558 4922
rect 10558 4870 10580 4922
rect 10604 4870 10610 4922
rect 10610 4870 10622 4922
rect 10622 4870 10660 4922
rect 10684 4870 10686 4922
rect 10686 4870 10738 4922
rect 10738 4870 10740 4922
rect 10364 4868 10420 4870
rect 10444 4868 10500 4870
rect 10524 4868 10580 4870
rect 10604 4868 10660 4870
rect 10684 4868 10740 4870
rect 10506 4564 10508 4584
rect 10508 4564 10560 4584
rect 10560 4564 10562 4584
rect 10506 4528 10562 4564
rect 10046 3732 10102 3768
rect 10046 3712 10048 3732
rect 10048 3712 10100 3732
rect 10100 3712 10102 3732
rect 8758 2252 8760 2272
rect 8760 2252 8812 2272
rect 8812 2252 8814 2272
rect 8758 2216 8814 2252
rect 7364 1114 7420 1116
rect 7444 1114 7500 1116
rect 7524 1114 7580 1116
rect 7604 1114 7660 1116
rect 7684 1114 7740 1116
rect 7364 1062 7366 1114
rect 7366 1062 7418 1114
rect 7418 1062 7420 1114
rect 7444 1062 7482 1114
rect 7482 1062 7494 1114
rect 7494 1062 7500 1114
rect 7524 1062 7546 1114
rect 7546 1062 7558 1114
rect 7558 1062 7580 1114
rect 7604 1062 7610 1114
rect 7610 1062 7622 1114
rect 7622 1062 7660 1114
rect 7684 1062 7686 1114
rect 7686 1062 7738 1114
rect 7738 1062 7740 1114
rect 7364 1060 7420 1062
rect 7444 1060 7500 1062
rect 7524 1060 7580 1062
rect 7604 1060 7660 1062
rect 7684 1060 7740 1062
rect 8574 1420 8630 1456
rect 8574 1400 8576 1420
rect 8576 1400 8628 1420
rect 8628 1400 8630 1420
rect 10364 3834 10420 3836
rect 10444 3834 10500 3836
rect 10524 3834 10580 3836
rect 10604 3834 10660 3836
rect 10684 3834 10740 3836
rect 10364 3782 10366 3834
rect 10366 3782 10418 3834
rect 10418 3782 10420 3834
rect 10444 3782 10482 3834
rect 10482 3782 10494 3834
rect 10494 3782 10500 3834
rect 10524 3782 10546 3834
rect 10546 3782 10558 3834
rect 10558 3782 10580 3834
rect 10604 3782 10610 3834
rect 10610 3782 10622 3834
rect 10622 3782 10660 3834
rect 10684 3782 10686 3834
rect 10686 3782 10738 3834
rect 10738 3782 10740 3834
rect 10364 3780 10420 3782
rect 10444 3780 10500 3782
rect 10524 3780 10580 3782
rect 10604 3780 10660 3782
rect 10684 3780 10740 3782
rect 9586 3304 9642 3360
rect 9494 3168 9550 3224
rect 9954 3168 10010 3224
rect 9678 3032 9734 3088
rect 9310 2760 9366 2816
rect 9770 2796 9772 2816
rect 9772 2796 9824 2816
rect 9824 2796 9826 2816
rect 9770 2760 9826 2796
rect 9494 2624 9550 2680
rect 9770 2624 9826 2680
rect 10046 2624 10102 2680
rect 9402 2352 9458 2408
rect 9126 1944 9182 2000
rect 9494 1672 9550 1728
rect 10414 3168 10470 3224
rect 10364 2746 10420 2748
rect 10444 2746 10500 2748
rect 10524 2746 10580 2748
rect 10604 2746 10660 2748
rect 10684 2746 10740 2748
rect 10364 2694 10366 2746
rect 10366 2694 10418 2746
rect 10418 2694 10420 2746
rect 10444 2694 10482 2746
rect 10482 2694 10494 2746
rect 10494 2694 10500 2746
rect 10524 2694 10546 2746
rect 10546 2694 10558 2746
rect 10558 2694 10580 2746
rect 10604 2694 10610 2746
rect 10610 2694 10622 2746
rect 10622 2694 10660 2746
rect 10684 2694 10686 2746
rect 10686 2694 10738 2746
rect 10738 2694 10740 2746
rect 10364 2692 10420 2694
rect 10444 2692 10500 2694
rect 10524 2692 10580 2694
rect 10604 2692 10660 2694
rect 10684 2692 10740 2694
rect 10874 1944 10930 2000
rect 9770 856 9826 912
rect 10364 1658 10420 1660
rect 10444 1658 10500 1660
rect 10524 1658 10580 1660
rect 10604 1658 10660 1660
rect 10684 1658 10740 1660
rect 10364 1606 10366 1658
rect 10366 1606 10418 1658
rect 10418 1606 10420 1658
rect 10444 1606 10482 1658
rect 10482 1606 10494 1658
rect 10494 1606 10500 1658
rect 10524 1606 10546 1658
rect 10546 1606 10558 1658
rect 10558 1606 10580 1658
rect 10604 1606 10610 1658
rect 10610 1606 10622 1658
rect 10622 1606 10660 1658
rect 10684 1606 10686 1658
rect 10686 1606 10738 1658
rect 10738 1606 10740 1658
rect 10364 1604 10420 1606
rect 10444 1604 10500 1606
rect 10524 1604 10580 1606
rect 10604 1604 10660 1606
rect 10684 1604 10740 1606
rect 11058 5072 11114 5128
rect 11058 3304 11114 3360
rect 11610 10240 11666 10296
rect 13364 14170 13420 14172
rect 13444 14170 13500 14172
rect 13524 14170 13580 14172
rect 13604 14170 13660 14172
rect 13684 14170 13740 14172
rect 13364 14118 13366 14170
rect 13366 14118 13418 14170
rect 13418 14118 13420 14170
rect 13444 14118 13482 14170
rect 13482 14118 13494 14170
rect 13494 14118 13500 14170
rect 13524 14118 13546 14170
rect 13546 14118 13558 14170
rect 13558 14118 13580 14170
rect 13604 14118 13610 14170
rect 13610 14118 13622 14170
rect 13622 14118 13660 14170
rect 13684 14118 13686 14170
rect 13686 14118 13738 14170
rect 13738 14118 13740 14170
rect 13364 14116 13420 14118
rect 13444 14116 13500 14118
rect 13524 14116 13580 14118
rect 13604 14116 13660 14118
rect 13684 14116 13740 14118
rect 13818 13912 13874 13968
rect 11794 9036 11850 9072
rect 11794 9016 11796 9036
rect 11796 9016 11848 9036
rect 11848 9016 11850 9036
rect 12254 10376 12310 10432
rect 11794 7284 11796 7304
rect 11796 7284 11848 7304
rect 11848 7284 11850 7304
rect 11794 7248 11850 7284
rect 11518 6976 11574 7032
rect 11518 6840 11574 6896
rect 11334 5888 11390 5944
rect 11886 6976 11942 7032
rect 12346 9288 12402 9344
rect 12162 7520 12218 7576
rect 12438 8200 12494 8256
rect 12530 8064 12586 8120
rect 12162 6976 12218 7032
rect 12162 6568 12218 6624
rect 11978 5888 12034 5944
rect 11334 4936 11390 4992
rect 11794 3032 11850 3088
rect 11334 2352 11390 2408
rect 11702 2216 11758 2272
rect 11794 2080 11850 2136
rect 11518 1400 11574 1456
rect 12898 12860 12900 12880
rect 12900 12860 12952 12880
rect 12952 12860 12954 12880
rect 12898 12824 12954 12860
rect 12990 11736 13046 11792
rect 12714 9288 12770 9344
rect 13364 13082 13420 13084
rect 13444 13082 13500 13084
rect 13524 13082 13580 13084
rect 13604 13082 13660 13084
rect 13684 13082 13740 13084
rect 13364 13030 13366 13082
rect 13366 13030 13418 13082
rect 13418 13030 13420 13082
rect 13444 13030 13482 13082
rect 13482 13030 13494 13082
rect 13494 13030 13500 13082
rect 13524 13030 13546 13082
rect 13546 13030 13558 13082
rect 13558 13030 13580 13082
rect 13604 13030 13610 13082
rect 13610 13030 13622 13082
rect 13622 13030 13660 13082
rect 13684 13030 13686 13082
rect 13686 13030 13738 13082
rect 13738 13030 13740 13082
rect 13364 13028 13420 13030
rect 13444 13028 13500 13030
rect 13524 13028 13580 13030
rect 13604 13028 13660 13030
rect 13684 13028 13740 13030
rect 13726 12552 13782 12608
rect 13364 11994 13420 11996
rect 13444 11994 13500 11996
rect 13524 11994 13580 11996
rect 13604 11994 13660 11996
rect 13684 11994 13740 11996
rect 13364 11942 13366 11994
rect 13366 11942 13418 11994
rect 13418 11942 13420 11994
rect 13444 11942 13482 11994
rect 13482 11942 13494 11994
rect 13494 11942 13500 11994
rect 13524 11942 13546 11994
rect 13546 11942 13558 11994
rect 13558 11942 13580 11994
rect 13604 11942 13610 11994
rect 13610 11942 13622 11994
rect 13622 11942 13660 11994
rect 13684 11942 13686 11994
rect 13686 11942 13738 11994
rect 13738 11942 13740 11994
rect 13364 11940 13420 11942
rect 13444 11940 13500 11942
rect 13524 11940 13580 11942
rect 13604 11940 13660 11942
rect 13684 11940 13740 11942
rect 13910 11328 13966 11384
rect 13818 11056 13874 11112
rect 13174 10240 13230 10296
rect 12530 6840 12586 6896
rect 12806 5616 12862 5672
rect 13364 10906 13420 10908
rect 13444 10906 13500 10908
rect 13524 10906 13580 10908
rect 13604 10906 13660 10908
rect 13684 10906 13740 10908
rect 13364 10854 13366 10906
rect 13366 10854 13418 10906
rect 13418 10854 13420 10906
rect 13444 10854 13482 10906
rect 13482 10854 13494 10906
rect 13494 10854 13500 10906
rect 13524 10854 13546 10906
rect 13546 10854 13558 10906
rect 13558 10854 13580 10906
rect 13604 10854 13610 10906
rect 13610 10854 13622 10906
rect 13622 10854 13660 10906
rect 13684 10854 13686 10906
rect 13686 10854 13738 10906
rect 13738 10854 13740 10906
rect 13364 10852 13420 10854
rect 13444 10852 13500 10854
rect 13524 10852 13580 10854
rect 13604 10852 13660 10854
rect 13684 10852 13740 10854
rect 14646 13812 14648 13832
rect 14648 13812 14700 13832
rect 14700 13812 14702 13832
rect 14646 13776 14702 13812
rect 13364 9818 13420 9820
rect 13444 9818 13500 9820
rect 13524 9818 13580 9820
rect 13604 9818 13660 9820
rect 13684 9818 13740 9820
rect 13364 9766 13366 9818
rect 13366 9766 13418 9818
rect 13418 9766 13420 9818
rect 13444 9766 13482 9818
rect 13482 9766 13494 9818
rect 13494 9766 13500 9818
rect 13524 9766 13546 9818
rect 13546 9766 13558 9818
rect 13558 9766 13580 9818
rect 13604 9766 13610 9818
rect 13610 9766 13622 9818
rect 13622 9766 13660 9818
rect 13684 9766 13686 9818
rect 13686 9766 13738 9818
rect 13738 9766 13740 9818
rect 13364 9764 13420 9766
rect 13444 9764 13500 9766
rect 13524 9764 13580 9766
rect 13604 9764 13660 9766
rect 13684 9764 13740 9766
rect 13358 9152 13414 9208
rect 13634 9036 13690 9072
rect 13634 9016 13636 9036
rect 13636 9016 13688 9036
rect 13688 9016 13690 9036
rect 13364 8730 13420 8732
rect 13444 8730 13500 8732
rect 13524 8730 13580 8732
rect 13604 8730 13660 8732
rect 13684 8730 13740 8732
rect 13364 8678 13366 8730
rect 13366 8678 13418 8730
rect 13418 8678 13420 8730
rect 13444 8678 13482 8730
rect 13482 8678 13494 8730
rect 13494 8678 13500 8730
rect 13524 8678 13546 8730
rect 13546 8678 13558 8730
rect 13558 8678 13580 8730
rect 13604 8678 13610 8730
rect 13610 8678 13622 8730
rect 13622 8678 13660 8730
rect 13684 8678 13686 8730
rect 13686 8678 13738 8730
rect 13738 8678 13740 8730
rect 13364 8676 13420 8678
rect 13444 8676 13500 8678
rect 13524 8676 13580 8678
rect 13604 8676 13660 8678
rect 13684 8676 13740 8678
rect 13726 7928 13782 7984
rect 13364 7642 13420 7644
rect 13444 7642 13500 7644
rect 13524 7642 13580 7644
rect 13604 7642 13660 7644
rect 13684 7642 13740 7644
rect 13364 7590 13366 7642
rect 13366 7590 13418 7642
rect 13418 7590 13420 7642
rect 13444 7590 13482 7642
rect 13482 7590 13494 7642
rect 13494 7590 13500 7642
rect 13524 7590 13546 7642
rect 13546 7590 13558 7642
rect 13558 7590 13580 7642
rect 13604 7590 13610 7642
rect 13610 7590 13622 7642
rect 13622 7590 13660 7642
rect 13684 7590 13686 7642
rect 13686 7590 13738 7642
rect 13738 7590 13740 7642
rect 13364 7588 13420 7590
rect 13444 7588 13500 7590
rect 13524 7588 13580 7590
rect 13604 7588 13660 7590
rect 13684 7588 13740 7590
rect 12990 4800 13046 4856
rect 14002 8064 14058 8120
rect 13634 6704 13690 6760
rect 13364 6554 13420 6556
rect 13444 6554 13500 6556
rect 13524 6554 13580 6556
rect 13604 6554 13660 6556
rect 13684 6554 13740 6556
rect 13364 6502 13366 6554
rect 13366 6502 13418 6554
rect 13418 6502 13420 6554
rect 13444 6502 13482 6554
rect 13482 6502 13494 6554
rect 13494 6502 13500 6554
rect 13524 6502 13546 6554
rect 13546 6502 13558 6554
rect 13558 6502 13580 6554
rect 13604 6502 13610 6554
rect 13610 6502 13622 6554
rect 13622 6502 13660 6554
rect 13684 6502 13686 6554
rect 13686 6502 13738 6554
rect 13738 6502 13740 6554
rect 13364 6500 13420 6502
rect 13444 6500 13500 6502
rect 13524 6500 13580 6502
rect 13604 6500 13660 6502
rect 13684 6500 13740 6502
rect 14186 7520 14242 7576
rect 14186 7284 14188 7304
rect 14188 7284 14240 7304
rect 14240 7284 14242 7304
rect 14186 7248 14242 7284
rect 13910 6432 13966 6488
rect 14094 6296 14150 6352
rect 13266 5616 13322 5672
rect 13364 5466 13420 5468
rect 13444 5466 13500 5468
rect 13524 5466 13580 5468
rect 13604 5466 13660 5468
rect 13684 5466 13740 5468
rect 13364 5414 13366 5466
rect 13366 5414 13418 5466
rect 13418 5414 13420 5466
rect 13444 5414 13482 5466
rect 13482 5414 13494 5466
rect 13494 5414 13500 5466
rect 13524 5414 13546 5466
rect 13546 5414 13558 5466
rect 13558 5414 13580 5466
rect 13604 5414 13610 5466
rect 13610 5414 13622 5466
rect 13622 5414 13660 5466
rect 13684 5414 13686 5466
rect 13686 5414 13738 5466
rect 13738 5414 13740 5466
rect 13364 5412 13420 5414
rect 13444 5412 13500 5414
rect 13524 5412 13580 5414
rect 13604 5412 13660 5414
rect 13684 5412 13740 5414
rect 13174 5072 13230 5128
rect 12806 4020 12808 4040
rect 12808 4020 12860 4040
rect 12860 4020 12862 4040
rect 12806 3984 12862 4020
rect 13634 4936 13690 4992
rect 13364 4378 13420 4380
rect 13444 4378 13500 4380
rect 13524 4378 13580 4380
rect 13604 4378 13660 4380
rect 13684 4378 13740 4380
rect 13364 4326 13366 4378
rect 13366 4326 13418 4378
rect 13418 4326 13420 4378
rect 13444 4326 13482 4378
rect 13482 4326 13494 4378
rect 13494 4326 13500 4378
rect 13524 4326 13546 4378
rect 13546 4326 13558 4378
rect 13558 4326 13580 4378
rect 13604 4326 13610 4378
rect 13610 4326 13622 4378
rect 13622 4326 13660 4378
rect 13684 4326 13686 4378
rect 13686 4326 13738 4378
rect 13738 4326 13740 4378
rect 13364 4324 13420 4326
rect 13444 4324 13500 4326
rect 13524 4324 13580 4326
rect 13604 4324 13660 4326
rect 13684 4324 13740 4326
rect 13450 4156 13452 4176
rect 13452 4156 13504 4176
rect 13504 4156 13506 4176
rect 13450 4120 13506 4156
rect 12346 2896 12402 2952
rect 12990 2624 13046 2680
rect 13364 3290 13420 3292
rect 13444 3290 13500 3292
rect 13524 3290 13580 3292
rect 13604 3290 13660 3292
rect 13684 3290 13740 3292
rect 13364 3238 13366 3290
rect 13366 3238 13418 3290
rect 13418 3238 13420 3290
rect 13444 3238 13482 3290
rect 13482 3238 13494 3290
rect 13494 3238 13500 3290
rect 13524 3238 13546 3290
rect 13546 3238 13558 3290
rect 13558 3238 13580 3290
rect 13604 3238 13610 3290
rect 13610 3238 13622 3290
rect 13622 3238 13660 3290
rect 13684 3238 13686 3290
rect 13686 3238 13738 3290
rect 13738 3238 13740 3290
rect 13364 3236 13420 3238
rect 13444 3236 13500 3238
rect 13524 3236 13580 3238
rect 13604 3236 13660 3238
rect 13684 3236 13740 3238
rect 13542 2624 13598 2680
rect 13364 2202 13420 2204
rect 13444 2202 13500 2204
rect 13524 2202 13580 2204
rect 13604 2202 13660 2204
rect 13684 2202 13740 2204
rect 13364 2150 13366 2202
rect 13366 2150 13418 2202
rect 13418 2150 13420 2202
rect 13444 2150 13482 2202
rect 13482 2150 13494 2202
rect 13494 2150 13500 2202
rect 13524 2150 13546 2202
rect 13546 2150 13558 2202
rect 13558 2150 13580 2202
rect 13604 2150 13610 2202
rect 13610 2150 13622 2202
rect 13622 2150 13660 2202
rect 13684 2150 13686 2202
rect 13686 2150 13738 2202
rect 13738 2150 13740 2202
rect 13364 2148 13420 2150
rect 13444 2148 13500 2150
rect 13524 2148 13580 2150
rect 13604 2148 13660 2150
rect 13684 2148 13740 2150
rect 13358 1536 13414 1592
rect 10364 570 10420 572
rect 10444 570 10500 572
rect 10524 570 10580 572
rect 10604 570 10660 572
rect 10684 570 10740 572
rect 10364 518 10366 570
rect 10366 518 10418 570
rect 10418 518 10420 570
rect 10444 518 10482 570
rect 10482 518 10494 570
rect 10494 518 10500 570
rect 10524 518 10546 570
rect 10546 518 10558 570
rect 10558 518 10580 570
rect 10604 518 10610 570
rect 10610 518 10622 570
rect 10622 518 10660 570
rect 10684 518 10686 570
rect 10686 518 10738 570
rect 10738 518 10740 570
rect 10364 516 10420 518
rect 10444 516 10500 518
rect 10524 516 10580 518
rect 10604 516 10660 518
rect 10684 516 10740 518
rect 14646 12588 14648 12608
rect 14648 12588 14700 12608
rect 14700 12588 14702 12608
rect 14646 12552 14702 12588
rect 14646 11328 14702 11384
rect 14554 10376 14610 10432
rect 14738 10240 14794 10296
rect 14646 9016 14702 9072
rect 15014 8744 15070 8800
rect 14830 7520 14886 7576
rect 14738 6024 14794 6080
rect 14738 5752 14794 5808
rect 15842 14340 15898 14376
rect 15842 14320 15844 14340
rect 15844 14320 15896 14340
rect 15896 14320 15898 14340
rect 16364 14714 16420 14716
rect 16444 14714 16500 14716
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16364 14662 16366 14714
rect 16366 14662 16418 14714
rect 16418 14662 16420 14714
rect 16444 14662 16482 14714
rect 16482 14662 16494 14714
rect 16494 14662 16500 14714
rect 16524 14662 16546 14714
rect 16546 14662 16558 14714
rect 16558 14662 16580 14714
rect 16604 14662 16610 14714
rect 16610 14662 16622 14714
rect 16622 14662 16660 14714
rect 16684 14662 16686 14714
rect 16686 14662 16738 14714
rect 16738 14662 16740 14714
rect 16364 14660 16420 14662
rect 16444 14660 16500 14662
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 15842 13640 15898 13696
rect 16364 13626 16420 13628
rect 16444 13626 16500 13628
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16364 13574 16366 13626
rect 16366 13574 16418 13626
rect 16418 13574 16420 13626
rect 16444 13574 16482 13626
rect 16482 13574 16494 13626
rect 16494 13574 16500 13626
rect 16524 13574 16546 13626
rect 16546 13574 16558 13626
rect 16558 13574 16580 13626
rect 16604 13574 16610 13626
rect 16610 13574 16622 13626
rect 16622 13574 16660 13626
rect 16684 13574 16686 13626
rect 16686 13574 16738 13626
rect 16738 13574 16740 13626
rect 16364 13572 16420 13574
rect 16444 13572 16500 13574
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16364 12538 16420 12540
rect 16444 12538 16500 12540
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16364 12486 16366 12538
rect 16366 12486 16418 12538
rect 16418 12486 16420 12538
rect 16444 12486 16482 12538
rect 16482 12486 16494 12538
rect 16494 12486 16500 12538
rect 16524 12486 16546 12538
rect 16546 12486 16558 12538
rect 16558 12486 16580 12538
rect 16604 12486 16610 12538
rect 16610 12486 16622 12538
rect 16622 12486 16660 12538
rect 16684 12486 16686 12538
rect 16686 12486 16738 12538
rect 16738 12486 16740 12538
rect 16364 12484 16420 12486
rect 16444 12484 16500 12486
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 15842 12416 15898 12472
rect 16026 11736 16082 11792
rect 16762 11736 16818 11792
rect 16364 11450 16420 11452
rect 16444 11450 16500 11452
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16364 11398 16366 11450
rect 16366 11398 16418 11450
rect 16418 11398 16420 11450
rect 16444 11398 16482 11450
rect 16482 11398 16494 11450
rect 16494 11398 16500 11450
rect 16524 11398 16546 11450
rect 16546 11398 16558 11450
rect 16558 11398 16580 11450
rect 16604 11398 16610 11450
rect 16610 11398 16622 11450
rect 16622 11398 16660 11450
rect 16684 11398 16686 11450
rect 16686 11398 16738 11450
rect 16738 11398 16740 11450
rect 16364 11396 16420 11398
rect 16444 11396 16500 11398
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16364 10362 16420 10364
rect 16444 10362 16500 10364
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16364 10310 16366 10362
rect 16366 10310 16418 10362
rect 16418 10310 16420 10362
rect 16444 10310 16482 10362
rect 16482 10310 16494 10362
rect 16494 10310 16500 10362
rect 16524 10310 16546 10362
rect 16546 10310 16558 10362
rect 16558 10310 16580 10362
rect 16604 10310 16610 10362
rect 16610 10310 16622 10362
rect 16622 10310 16660 10362
rect 16684 10310 16686 10362
rect 16686 10310 16738 10362
rect 16738 10310 16740 10362
rect 16364 10308 16420 10310
rect 16444 10308 16500 10310
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16854 10512 16910 10568
rect 15382 9016 15438 9072
rect 15474 8472 15530 8528
rect 15290 7248 15346 7304
rect 14646 3032 14702 3088
rect 14830 2916 14886 2952
rect 14830 2896 14832 2916
rect 14832 2896 14884 2916
rect 14884 2896 14886 2916
rect 15658 8200 15714 8256
rect 15474 5228 15530 5264
rect 15474 5208 15476 5228
rect 15476 5208 15528 5228
rect 15528 5208 15530 5228
rect 14922 2080 14978 2136
rect 16026 8744 16082 8800
rect 15934 6432 15990 6488
rect 15934 5480 15990 5536
rect 16670 9460 16672 9480
rect 16672 9460 16724 9480
rect 16724 9460 16726 9480
rect 16670 9424 16726 9460
rect 16364 9274 16420 9276
rect 16444 9274 16500 9276
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16364 9222 16366 9274
rect 16366 9222 16418 9274
rect 16418 9222 16420 9274
rect 16444 9222 16482 9274
rect 16482 9222 16494 9274
rect 16494 9222 16500 9274
rect 16524 9222 16546 9274
rect 16546 9222 16558 9274
rect 16558 9222 16580 9274
rect 16604 9222 16610 9274
rect 16610 9222 16622 9274
rect 16622 9222 16660 9274
rect 16684 9222 16686 9274
rect 16686 9222 16738 9274
rect 16738 9222 16740 9274
rect 16364 9220 16420 9222
rect 16444 9220 16500 9222
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16578 8372 16580 8392
rect 16580 8372 16632 8392
rect 16632 8372 16634 8392
rect 16578 8336 16634 8372
rect 16364 8186 16420 8188
rect 16444 8186 16500 8188
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16364 8134 16366 8186
rect 16366 8134 16418 8186
rect 16418 8134 16420 8186
rect 16444 8134 16482 8186
rect 16482 8134 16494 8186
rect 16494 8134 16500 8186
rect 16524 8134 16546 8186
rect 16546 8134 16558 8186
rect 16558 8134 16580 8186
rect 16604 8134 16610 8186
rect 16610 8134 16622 8186
rect 16622 8134 16660 8186
rect 16684 8134 16686 8186
rect 16686 8134 16738 8186
rect 16738 8134 16740 8186
rect 16364 8132 16420 8134
rect 16444 8132 16500 8134
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16364 7098 16420 7100
rect 16444 7098 16500 7100
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16364 7046 16366 7098
rect 16366 7046 16418 7098
rect 16418 7046 16420 7098
rect 16444 7046 16482 7098
rect 16482 7046 16494 7098
rect 16494 7046 16500 7098
rect 16524 7046 16546 7098
rect 16546 7046 16558 7098
rect 16558 7046 16580 7098
rect 16604 7046 16610 7098
rect 16610 7046 16622 7098
rect 16622 7046 16660 7098
rect 16684 7046 16686 7098
rect 16686 7046 16738 7098
rect 16738 7046 16740 7098
rect 16364 7044 16420 7046
rect 16444 7044 16500 7046
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16210 6976 16266 7032
rect 15474 4528 15530 4584
rect 15566 3340 15568 3360
rect 15568 3340 15620 3360
rect 15620 3340 15622 3360
rect 15566 3304 15622 3340
rect 15750 3032 15806 3088
rect 13364 1114 13420 1116
rect 13444 1114 13500 1116
rect 13524 1114 13580 1116
rect 13604 1114 13660 1116
rect 13684 1114 13740 1116
rect 13364 1062 13366 1114
rect 13366 1062 13418 1114
rect 13418 1062 13420 1114
rect 13444 1062 13482 1114
rect 13482 1062 13494 1114
rect 13494 1062 13500 1114
rect 13524 1062 13546 1114
rect 13546 1062 13558 1114
rect 13558 1062 13580 1114
rect 13604 1062 13610 1114
rect 13610 1062 13622 1114
rect 13622 1062 13660 1114
rect 13684 1062 13686 1114
rect 13686 1062 13738 1114
rect 13738 1062 13740 1114
rect 13364 1060 13420 1062
rect 13444 1060 13500 1062
rect 13524 1060 13580 1062
rect 13604 1060 13660 1062
rect 13684 1060 13740 1062
rect 15658 2080 15714 2136
rect 15658 1556 15714 1592
rect 15658 1536 15660 1556
rect 15660 1536 15712 1556
rect 15712 1536 15714 1556
rect 16026 4528 16082 4584
rect 15934 2216 15990 2272
rect 16364 6010 16420 6012
rect 16444 6010 16500 6012
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16364 5958 16366 6010
rect 16366 5958 16418 6010
rect 16418 5958 16420 6010
rect 16444 5958 16482 6010
rect 16482 5958 16494 6010
rect 16494 5958 16500 6010
rect 16524 5958 16546 6010
rect 16546 5958 16558 6010
rect 16558 5958 16580 6010
rect 16604 5958 16610 6010
rect 16610 5958 16622 6010
rect 16622 5958 16660 6010
rect 16684 5958 16686 6010
rect 16686 5958 16738 6010
rect 16738 5958 16740 6010
rect 16364 5956 16420 5958
rect 16444 5956 16500 5958
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 17130 14340 17186 14376
rect 17130 14320 17132 14340
rect 17132 14320 17184 14340
rect 17184 14320 17186 14340
rect 17130 10648 17186 10704
rect 17958 14456 18014 14512
rect 17406 12144 17462 12200
rect 17222 8628 17278 8664
rect 17222 8608 17224 8628
rect 17224 8608 17276 8628
rect 17276 8608 17278 8628
rect 17314 8472 17370 8528
rect 16946 5480 17002 5536
rect 16946 5072 17002 5128
rect 16364 4922 16420 4924
rect 16444 4922 16500 4924
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16364 4870 16366 4922
rect 16366 4870 16418 4922
rect 16418 4870 16420 4922
rect 16444 4870 16482 4922
rect 16482 4870 16494 4922
rect 16494 4870 16500 4922
rect 16524 4870 16546 4922
rect 16546 4870 16558 4922
rect 16558 4870 16580 4922
rect 16604 4870 16610 4922
rect 16610 4870 16622 4922
rect 16622 4870 16660 4922
rect 16684 4870 16686 4922
rect 16686 4870 16738 4922
rect 16738 4870 16740 4922
rect 16364 4868 16420 4870
rect 16444 4868 16500 4870
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16364 3834 16420 3836
rect 16444 3834 16500 3836
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16364 3782 16366 3834
rect 16366 3782 16418 3834
rect 16418 3782 16420 3834
rect 16444 3782 16482 3834
rect 16482 3782 16494 3834
rect 16494 3782 16500 3834
rect 16524 3782 16546 3834
rect 16546 3782 16558 3834
rect 16558 3782 16580 3834
rect 16604 3782 16610 3834
rect 16610 3782 16622 3834
rect 16622 3782 16660 3834
rect 16684 3782 16686 3834
rect 16686 3782 16738 3834
rect 16738 3782 16740 3834
rect 16364 3780 16420 3782
rect 16444 3780 16500 3782
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16578 3440 16634 3496
rect 16394 3304 16450 3360
rect 16210 3032 16266 3088
rect 16364 2746 16420 2748
rect 16444 2746 16500 2748
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16364 2694 16366 2746
rect 16366 2694 16418 2746
rect 16418 2694 16420 2746
rect 16444 2694 16482 2746
rect 16482 2694 16494 2746
rect 16494 2694 16500 2746
rect 16524 2694 16546 2746
rect 16546 2694 16558 2746
rect 16558 2694 16580 2746
rect 16604 2694 16610 2746
rect 16610 2694 16622 2746
rect 16622 2694 16660 2746
rect 16684 2694 16686 2746
rect 16686 2694 16738 2746
rect 16738 2694 16740 2746
rect 16364 2692 16420 2694
rect 16444 2692 16500 2694
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16118 2080 16174 2136
rect 16364 1658 16420 1660
rect 16444 1658 16500 1660
rect 16524 1658 16580 1660
rect 16604 1658 16660 1660
rect 16684 1658 16740 1660
rect 16364 1606 16366 1658
rect 16366 1606 16418 1658
rect 16418 1606 16420 1658
rect 16444 1606 16482 1658
rect 16482 1606 16494 1658
rect 16494 1606 16500 1658
rect 16524 1606 16546 1658
rect 16546 1606 16558 1658
rect 16558 1606 16580 1658
rect 16604 1606 16610 1658
rect 16610 1606 16622 1658
rect 16622 1606 16660 1658
rect 16684 1606 16686 1658
rect 16686 1606 16738 1658
rect 16738 1606 16740 1658
rect 16364 1604 16420 1606
rect 16444 1604 16500 1606
rect 16524 1604 16580 1606
rect 16604 1604 16660 1606
rect 16684 1604 16740 1606
rect 16394 1420 16450 1456
rect 16394 1400 16396 1420
rect 16396 1400 16448 1420
rect 16448 1400 16450 1420
rect 17038 4664 17094 4720
rect 19364 15258 19420 15260
rect 19444 15258 19500 15260
rect 19524 15258 19580 15260
rect 19604 15258 19660 15260
rect 19684 15258 19740 15260
rect 19364 15206 19366 15258
rect 19366 15206 19418 15258
rect 19418 15206 19420 15258
rect 19444 15206 19482 15258
rect 19482 15206 19494 15258
rect 19494 15206 19500 15258
rect 19524 15206 19546 15258
rect 19546 15206 19558 15258
rect 19558 15206 19580 15258
rect 19604 15206 19610 15258
rect 19610 15206 19622 15258
rect 19622 15206 19660 15258
rect 19684 15206 19686 15258
rect 19686 15206 19738 15258
rect 19738 15206 19740 15258
rect 19364 15204 19420 15206
rect 19444 15204 19500 15206
rect 19524 15204 19580 15206
rect 19604 15204 19660 15206
rect 19684 15204 19740 15206
rect 18878 14456 18934 14512
rect 18602 13912 18658 13968
rect 18602 13776 18658 13832
rect 19364 14170 19420 14172
rect 19444 14170 19500 14172
rect 19524 14170 19580 14172
rect 19604 14170 19660 14172
rect 19684 14170 19740 14172
rect 19364 14118 19366 14170
rect 19366 14118 19418 14170
rect 19418 14118 19420 14170
rect 19444 14118 19482 14170
rect 19482 14118 19494 14170
rect 19494 14118 19500 14170
rect 19524 14118 19546 14170
rect 19546 14118 19558 14170
rect 19558 14118 19580 14170
rect 19604 14118 19610 14170
rect 19610 14118 19622 14170
rect 19622 14118 19660 14170
rect 19684 14118 19686 14170
rect 19686 14118 19738 14170
rect 19738 14118 19740 14170
rect 19364 14116 19420 14118
rect 19444 14116 19500 14118
rect 19524 14116 19580 14118
rect 19604 14116 19660 14118
rect 19684 14116 19740 14118
rect 20074 13912 20130 13968
rect 18878 13368 18934 13424
rect 19364 13082 19420 13084
rect 19444 13082 19500 13084
rect 19524 13082 19580 13084
rect 19604 13082 19660 13084
rect 19684 13082 19740 13084
rect 19364 13030 19366 13082
rect 19366 13030 19418 13082
rect 19418 13030 19420 13082
rect 19444 13030 19482 13082
rect 19482 13030 19494 13082
rect 19494 13030 19500 13082
rect 19524 13030 19546 13082
rect 19546 13030 19558 13082
rect 19558 13030 19580 13082
rect 19604 13030 19610 13082
rect 19610 13030 19622 13082
rect 19622 13030 19660 13082
rect 19684 13030 19686 13082
rect 19686 13030 19738 13082
rect 19738 13030 19740 13082
rect 19364 13028 19420 13030
rect 19444 13028 19500 13030
rect 19524 13028 19580 13030
rect 19604 13028 19660 13030
rect 19684 13028 19740 13030
rect 17958 11092 17960 11112
rect 17960 11092 18012 11112
rect 18012 11092 18014 11112
rect 17958 11056 18014 11092
rect 17774 9424 17830 9480
rect 17774 8608 17830 8664
rect 17774 8472 17830 8528
rect 17498 7964 17500 7984
rect 17500 7964 17552 7984
rect 17552 7964 17554 7984
rect 17498 7928 17554 7964
rect 17406 7420 17408 7440
rect 17408 7420 17460 7440
rect 17460 7420 17462 7440
rect 17406 7384 17462 7420
rect 17314 6840 17370 6896
rect 17130 1944 17186 2000
rect 17682 7284 17684 7304
rect 17684 7284 17736 7304
rect 17736 7284 17738 7304
rect 17682 7248 17738 7284
rect 17498 2216 17554 2272
rect 17958 3440 18014 3496
rect 18326 12300 18382 12336
rect 18326 12280 18328 12300
rect 18328 12280 18380 12300
rect 18380 12280 18382 12300
rect 18326 7792 18382 7848
rect 18786 8336 18842 8392
rect 18234 2624 18290 2680
rect 18510 4120 18566 4176
rect 18510 3984 18566 4040
rect 18602 3440 18658 3496
rect 18878 3576 18934 3632
rect 19364 11994 19420 11996
rect 19444 11994 19500 11996
rect 19524 11994 19580 11996
rect 19604 11994 19660 11996
rect 19684 11994 19740 11996
rect 19364 11942 19366 11994
rect 19366 11942 19418 11994
rect 19418 11942 19420 11994
rect 19444 11942 19482 11994
rect 19482 11942 19494 11994
rect 19494 11942 19500 11994
rect 19524 11942 19546 11994
rect 19546 11942 19558 11994
rect 19558 11942 19580 11994
rect 19604 11942 19610 11994
rect 19610 11942 19622 11994
rect 19622 11942 19660 11994
rect 19684 11942 19686 11994
rect 19686 11942 19738 11994
rect 19738 11942 19740 11994
rect 19364 11940 19420 11942
rect 19444 11940 19500 11942
rect 19524 11940 19580 11942
rect 19604 11940 19660 11942
rect 19684 11940 19740 11942
rect 19706 11092 19708 11112
rect 19708 11092 19760 11112
rect 19760 11092 19762 11112
rect 19706 11056 19762 11092
rect 19364 10906 19420 10908
rect 19444 10906 19500 10908
rect 19524 10906 19580 10908
rect 19604 10906 19660 10908
rect 19684 10906 19740 10908
rect 19364 10854 19366 10906
rect 19366 10854 19418 10906
rect 19418 10854 19420 10906
rect 19444 10854 19482 10906
rect 19482 10854 19494 10906
rect 19494 10854 19500 10906
rect 19524 10854 19546 10906
rect 19546 10854 19558 10906
rect 19558 10854 19580 10906
rect 19604 10854 19610 10906
rect 19610 10854 19622 10906
rect 19622 10854 19660 10906
rect 19684 10854 19686 10906
rect 19686 10854 19738 10906
rect 19738 10854 19740 10906
rect 19364 10852 19420 10854
rect 19444 10852 19500 10854
rect 19524 10852 19580 10854
rect 19604 10852 19660 10854
rect 19684 10852 19740 10854
rect 22364 14714 22420 14716
rect 22444 14714 22500 14716
rect 22524 14714 22580 14716
rect 22604 14714 22660 14716
rect 22684 14714 22740 14716
rect 22364 14662 22366 14714
rect 22366 14662 22418 14714
rect 22418 14662 22420 14714
rect 22444 14662 22482 14714
rect 22482 14662 22494 14714
rect 22494 14662 22500 14714
rect 22524 14662 22546 14714
rect 22546 14662 22558 14714
rect 22558 14662 22580 14714
rect 22604 14662 22610 14714
rect 22610 14662 22622 14714
rect 22622 14662 22660 14714
rect 22684 14662 22686 14714
rect 22686 14662 22738 14714
rect 22738 14662 22740 14714
rect 22364 14660 22420 14662
rect 22444 14660 22500 14662
rect 22524 14660 22580 14662
rect 22604 14660 22660 14662
rect 22684 14660 22740 14662
rect 22364 13626 22420 13628
rect 22444 13626 22500 13628
rect 22524 13626 22580 13628
rect 22604 13626 22660 13628
rect 22684 13626 22740 13628
rect 22364 13574 22366 13626
rect 22366 13574 22418 13626
rect 22418 13574 22420 13626
rect 22444 13574 22482 13626
rect 22482 13574 22494 13626
rect 22494 13574 22500 13626
rect 22524 13574 22546 13626
rect 22546 13574 22558 13626
rect 22558 13574 22580 13626
rect 22604 13574 22610 13626
rect 22610 13574 22622 13626
rect 22622 13574 22660 13626
rect 22684 13574 22686 13626
rect 22686 13574 22738 13626
rect 22738 13574 22740 13626
rect 22364 13572 22420 13574
rect 22444 13572 22500 13574
rect 22524 13572 22580 13574
rect 22604 13572 22660 13574
rect 22684 13572 22740 13574
rect 19062 10104 19118 10160
rect 19338 10004 19340 10024
rect 19340 10004 19392 10024
rect 19392 10004 19394 10024
rect 19338 9968 19394 10004
rect 19364 9818 19420 9820
rect 19444 9818 19500 9820
rect 19524 9818 19580 9820
rect 19604 9818 19660 9820
rect 19684 9818 19740 9820
rect 19364 9766 19366 9818
rect 19366 9766 19418 9818
rect 19418 9766 19420 9818
rect 19444 9766 19482 9818
rect 19482 9766 19494 9818
rect 19494 9766 19500 9818
rect 19524 9766 19546 9818
rect 19546 9766 19558 9818
rect 19558 9766 19580 9818
rect 19604 9766 19610 9818
rect 19610 9766 19622 9818
rect 19622 9766 19660 9818
rect 19684 9766 19686 9818
rect 19686 9766 19738 9818
rect 19738 9766 19740 9818
rect 19364 9764 19420 9766
rect 19444 9764 19500 9766
rect 19524 9764 19580 9766
rect 19604 9764 19660 9766
rect 19684 9764 19740 9766
rect 19890 9832 19946 9888
rect 19338 9560 19394 9616
rect 19430 9152 19486 9208
rect 19706 9016 19762 9072
rect 19982 9560 20038 9616
rect 19364 8730 19420 8732
rect 19444 8730 19500 8732
rect 19524 8730 19580 8732
rect 19604 8730 19660 8732
rect 19684 8730 19740 8732
rect 19364 8678 19366 8730
rect 19366 8678 19418 8730
rect 19418 8678 19420 8730
rect 19444 8678 19482 8730
rect 19482 8678 19494 8730
rect 19494 8678 19500 8730
rect 19524 8678 19546 8730
rect 19546 8678 19558 8730
rect 19558 8678 19580 8730
rect 19604 8678 19610 8730
rect 19610 8678 19622 8730
rect 19622 8678 19660 8730
rect 19684 8678 19686 8730
rect 19686 8678 19738 8730
rect 19738 8678 19740 8730
rect 19364 8676 19420 8678
rect 19444 8676 19500 8678
rect 19524 8676 19580 8678
rect 19604 8676 19660 8678
rect 19684 8676 19740 8678
rect 19364 7642 19420 7644
rect 19444 7642 19500 7644
rect 19524 7642 19580 7644
rect 19604 7642 19660 7644
rect 19684 7642 19740 7644
rect 19364 7590 19366 7642
rect 19366 7590 19418 7642
rect 19418 7590 19420 7642
rect 19444 7590 19482 7642
rect 19482 7590 19494 7642
rect 19494 7590 19500 7642
rect 19524 7590 19546 7642
rect 19546 7590 19558 7642
rect 19558 7590 19580 7642
rect 19604 7590 19610 7642
rect 19610 7590 19622 7642
rect 19622 7590 19660 7642
rect 19684 7590 19686 7642
rect 19686 7590 19738 7642
rect 19738 7590 19740 7642
rect 19364 7588 19420 7590
rect 19444 7588 19500 7590
rect 19524 7588 19580 7590
rect 19604 7588 19660 7590
rect 19684 7588 19740 7590
rect 19364 6554 19420 6556
rect 19444 6554 19500 6556
rect 19524 6554 19580 6556
rect 19604 6554 19660 6556
rect 19684 6554 19740 6556
rect 19364 6502 19366 6554
rect 19366 6502 19418 6554
rect 19418 6502 19420 6554
rect 19444 6502 19482 6554
rect 19482 6502 19494 6554
rect 19494 6502 19500 6554
rect 19524 6502 19546 6554
rect 19546 6502 19558 6554
rect 19558 6502 19580 6554
rect 19604 6502 19610 6554
rect 19610 6502 19622 6554
rect 19622 6502 19660 6554
rect 19684 6502 19686 6554
rect 19686 6502 19738 6554
rect 19738 6502 19740 6554
rect 19364 6500 19420 6502
rect 19444 6500 19500 6502
rect 19524 6500 19580 6502
rect 19604 6500 19660 6502
rect 19684 6500 19740 6502
rect 19364 5466 19420 5468
rect 19444 5466 19500 5468
rect 19524 5466 19580 5468
rect 19604 5466 19660 5468
rect 19684 5466 19740 5468
rect 19364 5414 19366 5466
rect 19366 5414 19418 5466
rect 19418 5414 19420 5466
rect 19444 5414 19482 5466
rect 19482 5414 19494 5466
rect 19494 5414 19500 5466
rect 19524 5414 19546 5466
rect 19546 5414 19558 5466
rect 19558 5414 19580 5466
rect 19604 5414 19610 5466
rect 19610 5414 19622 5466
rect 19622 5414 19660 5466
rect 19684 5414 19686 5466
rect 19686 5414 19738 5466
rect 19738 5414 19740 5466
rect 19364 5412 19420 5414
rect 19444 5412 19500 5414
rect 19524 5412 19580 5414
rect 19604 5412 19660 5414
rect 19684 5412 19740 5414
rect 19614 4548 19670 4584
rect 19614 4528 19616 4548
rect 19616 4528 19668 4548
rect 19668 4528 19670 4548
rect 19364 4378 19420 4380
rect 19444 4378 19500 4380
rect 19524 4378 19580 4380
rect 19604 4378 19660 4380
rect 19684 4378 19740 4380
rect 19364 4326 19366 4378
rect 19366 4326 19418 4378
rect 19418 4326 19420 4378
rect 19444 4326 19482 4378
rect 19482 4326 19494 4378
rect 19494 4326 19500 4378
rect 19524 4326 19546 4378
rect 19546 4326 19558 4378
rect 19558 4326 19580 4378
rect 19604 4326 19610 4378
rect 19610 4326 19622 4378
rect 19622 4326 19660 4378
rect 19684 4326 19686 4378
rect 19686 4326 19738 4378
rect 19738 4326 19740 4378
rect 19364 4324 19420 4326
rect 19444 4324 19500 4326
rect 19524 4324 19580 4326
rect 19604 4324 19660 4326
rect 19684 4324 19740 4326
rect 20258 9560 20314 9616
rect 19982 8200 20038 8256
rect 20258 8200 20314 8256
rect 20718 11600 20774 11656
rect 20626 11056 20682 11112
rect 23294 12844 23350 12880
rect 23294 12824 23296 12844
rect 23296 12824 23348 12844
rect 23348 12824 23350 12844
rect 20994 9832 21050 9888
rect 19982 6160 20038 6216
rect 19982 3576 20038 3632
rect 19364 3290 19420 3292
rect 19444 3290 19500 3292
rect 19524 3290 19580 3292
rect 19604 3290 19660 3292
rect 19684 3290 19740 3292
rect 19364 3238 19366 3290
rect 19366 3238 19418 3290
rect 19418 3238 19420 3290
rect 19444 3238 19482 3290
rect 19482 3238 19494 3290
rect 19494 3238 19500 3290
rect 19524 3238 19546 3290
rect 19546 3238 19558 3290
rect 19558 3238 19580 3290
rect 19604 3238 19610 3290
rect 19610 3238 19622 3290
rect 19622 3238 19660 3290
rect 19684 3238 19686 3290
rect 19686 3238 19738 3290
rect 19738 3238 19740 3290
rect 19364 3236 19420 3238
rect 19444 3236 19500 3238
rect 19524 3236 19580 3238
rect 19604 3236 19660 3238
rect 19684 3236 19740 3238
rect 19706 2896 19762 2952
rect 21270 9560 21326 9616
rect 21086 9460 21088 9480
rect 21088 9460 21140 9480
rect 21140 9460 21142 9480
rect 21086 9424 21142 9460
rect 20810 8880 20866 8936
rect 20718 8336 20774 8392
rect 21362 9016 21418 9072
rect 21270 8200 21326 8256
rect 21362 5636 21418 5672
rect 21362 5616 21364 5636
rect 21364 5616 21416 5636
rect 21416 5616 21418 5636
rect 21638 9560 21694 9616
rect 21638 8492 21694 8528
rect 21638 8472 21640 8492
rect 21640 8472 21692 8492
rect 21692 8472 21694 8492
rect 22364 12538 22420 12540
rect 22444 12538 22500 12540
rect 22524 12538 22580 12540
rect 22604 12538 22660 12540
rect 22684 12538 22740 12540
rect 22364 12486 22366 12538
rect 22366 12486 22418 12538
rect 22418 12486 22420 12538
rect 22444 12486 22482 12538
rect 22482 12486 22494 12538
rect 22494 12486 22500 12538
rect 22524 12486 22546 12538
rect 22546 12486 22558 12538
rect 22558 12486 22580 12538
rect 22604 12486 22610 12538
rect 22610 12486 22622 12538
rect 22622 12486 22660 12538
rect 22684 12486 22686 12538
rect 22686 12486 22738 12538
rect 22738 12486 22740 12538
rect 22364 12484 22420 12486
rect 22444 12484 22500 12486
rect 22524 12484 22580 12486
rect 22604 12484 22660 12486
rect 22684 12484 22740 12486
rect 22364 11450 22420 11452
rect 22444 11450 22500 11452
rect 22524 11450 22580 11452
rect 22604 11450 22660 11452
rect 22684 11450 22740 11452
rect 22364 11398 22366 11450
rect 22366 11398 22418 11450
rect 22418 11398 22420 11450
rect 22444 11398 22482 11450
rect 22482 11398 22494 11450
rect 22494 11398 22500 11450
rect 22524 11398 22546 11450
rect 22546 11398 22558 11450
rect 22558 11398 22580 11450
rect 22604 11398 22610 11450
rect 22610 11398 22622 11450
rect 22622 11398 22660 11450
rect 22684 11398 22686 11450
rect 22686 11398 22738 11450
rect 22738 11398 22740 11450
rect 22364 11396 22420 11398
rect 22444 11396 22500 11398
rect 22524 11396 22580 11398
rect 22604 11396 22660 11398
rect 22684 11396 22740 11398
rect 22364 10362 22420 10364
rect 22444 10362 22500 10364
rect 22524 10362 22580 10364
rect 22604 10362 22660 10364
rect 22684 10362 22740 10364
rect 22364 10310 22366 10362
rect 22366 10310 22418 10362
rect 22418 10310 22420 10362
rect 22444 10310 22482 10362
rect 22482 10310 22494 10362
rect 22494 10310 22500 10362
rect 22524 10310 22546 10362
rect 22546 10310 22558 10362
rect 22558 10310 22580 10362
rect 22604 10310 22610 10362
rect 22610 10310 22622 10362
rect 22622 10310 22660 10362
rect 22684 10310 22686 10362
rect 22686 10310 22738 10362
rect 22738 10310 22740 10362
rect 22364 10308 22420 10310
rect 22444 10308 22500 10310
rect 22524 10308 22580 10310
rect 22604 10308 22660 10310
rect 22684 10308 22740 10310
rect 22098 9444 22154 9480
rect 22098 9424 22100 9444
rect 22100 9424 22152 9444
rect 22152 9424 22154 9444
rect 22364 9274 22420 9276
rect 22444 9274 22500 9276
rect 22524 9274 22580 9276
rect 22604 9274 22660 9276
rect 22684 9274 22740 9276
rect 22364 9222 22366 9274
rect 22366 9222 22418 9274
rect 22418 9222 22420 9274
rect 22444 9222 22482 9274
rect 22482 9222 22494 9274
rect 22494 9222 22500 9274
rect 22524 9222 22546 9274
rect 22546 9222 22558 9274
rect 22558 9222 22580 9274
rect 22604 9222 22610 9274
rect 22610 9222 22622 9274
rect 22622 9222 22660 9274
rect 22684 9222 22686 9274
rect 22686 9222 22738 9274
rect 22738 9222 22740 9274
rect 22364 9220 22420 9222
rect 22444 9220 22500 9222
rect 22524 9220 22580 9222
rect 22604 9220 22660 9222
rect 22684 9220 22740 9222
rect 22364 8186 22420 8188
rect 22444 8186 22500 8188
rect 22524 8186 22580 8188
rect 22604 8186 22660 8188
rect 22684 8186 22740 8188
rect 22364 8134 22366 8186
rect 22366 8134 22418 8186
rect 22418 8134 22420 8186
rect 22444 8134 22482 8186
rect 22482 8134 22494 8186
rect 22494 8134 22500 8186
rect 22524 8134 22546 8186
rect 22546 8134 22558 8186
rect 22558 8134 22580 8186
rect 22604 8134 22610 8186
rect 22610 8134 22622 8186
rect 22622 8134 22660 8186
rect 22684 8134 22686 8186
rect 22686 8134 22738 8186
rect 22738 8134 22740 8186
rect 22364 8132 22420 8134
rect 22444 8132 22500 8134
rect 22524 8132 22580 8134
rect 22604 8132 22660 8134
rect 22684 8132 22740 8134
rect 22364 7098 22420 7100
rect 22444 7098 22500 7100
rect 22524 7098 22580 7100
rect 22604 7098 22660 7100
rect 22684 7098 22740 7100
rect 22364 7046 22366 7098
rect 22366 7046 22418 7098
rect 22418 7046 22420 7098
rect 22444 7046 22482 7098
rect 22482 7046 22494 7098
rect 22494 7046 22500 7098
rect 22524 7046 22546 7098
rect 22546 7046 22558 7098
rect 22558 7046 22580 7098
rect 22604 7046 22610 7098
rect 22610 7046 22622 7098
rect 22622 7046 22660 7098
rect 22684 7046 22686 7098
rect 22686 7046 22738 7098
rect 22738 7046 22740 7098
rect 22364 7044 22420 7046
rect 22444 7044 22500 7046
rect 22524 7044 22580 7046
rect 22604 7044 22660 7046
rect 22684 7044 22740 7046
rect 22364 6010 22420 6012
rect 22444 6010 22500 6012
rect 22524 6010 22580 6012
rect 22604 6010 22660 6012
rect 22684 6010 22740 6012
rect 22364 5958 22366 6010
rect 22366 5958 22418 6010
rect 22418 5958 22420 6010
rect 22444 5958 22482 6010
rect 22482 5958 22494 6010
rect 22494 5958 22500 6010
rect 22524 5958 22546 6010
rect 22546 5958 22558 6010
rect 22558 5958 22580 6010
rect 22604 5958 22610 6010
rect 22610 5958 22622 6010
rect 22622 5958 22660 6010
rect 22684 5958 22686 6010
rect 22686 5958 22738 6010
rect 22738 5958 22740 6010
rect 22364 5956 22420 5958
rect 22444 5956 22500 5958
rect 22524 5956 22580 5958
rect 22604 5956 22660 5958
rect 22684 5956 22740 5958
rect 18878 2352 18934 2408
rect 16364 570 16420 572
rect 16444 570 16500 572
rect 16524 570 16580 572
rect 16604 570 16660 572
rect 16684 570 16740 572
rect 16364 518 16366 570
rect 16366 518 16418 570
rect 16418 518 16420 570
rect 16444 518 16482 570
rect 16482 518 16494 570
rect 16494 518 16500 570
rect 16524 518 16546 570
rect 16546 518 16558 570
rect 16558 518 16580 570
rect 16604 518 16610 570
rect 16610 518 16622 570
rect 16622 518 16660 570
rect 16684 518 16686 570
rect 16686 518 16738 570
rect 16738 518 16740 570
rect 16364 516 16420 518
rect 16444 516 16500 518
rect 16524 516 16580 518
rect 16604 516 16660 518
rect 16684 516 16740 518
rect 18418 1808 18474 1864
rect 19364 2202 19420 2204
rect 19444 2202 19500 2204
rect 19524 2202 19580 2204
rect 19604 2202 19660 2204
rect 19684 2202 19740 2204
rect 19364 2150 19366 2202
rect 19366 2150 19418 2202
rect 19418 2150 19420 2202
rect 19444 2150 19482 2202
rect 19482 2150 19494 2202
rect 19494 2150 19500 2202
rect 19524 2150 19546 2202
rect 19546 2150 19558 2202
rect 19558 2150 19580 2202
rect 19604 2150 19610 2202
rect 19610 2150 19622 2202
rect 19622 2150 19660 2202
rect 19684 2150 19686 2202
rect 19686 2150 19738 2202
rect 19738 2150 19740 2202
rect 19364 2148 19420 2150
rect 19444 2148 19500 2150
rect 19524 2148 19580 2150
rect 19604 2148 19660 2150
rect 19684 2148 19740 2150
rect 21454 4528 21510 4584
rect 22364 4922 22420 4924
rect 22444 4922 22500 4924
rect 22524 4922 22580 4924
rect 22604 4922 22660 4924
rect 22684 4922 22740 4924
rect 22364 4870 22366 4922
rect 22366 4870 22418 4922
rect 22418 4870 22420 4922
rect 22444 4870 22482 4922
rect 22482 4870 22494 4922
rect 22494 4870 22500 4922
rect 22524 4870 22546 4922
rect 22546 4870 22558 4922
rect 22558 4870 22580 4922
rect 22604 4870 22610 4922
rect 22610 4870 22622 4922
rect 22622 4870 22660 4922
rect 22684 4870 22686 4922
rect 22686 4870 22738 4922
rect 22738 4870 22740 4922
rect 22364 4868 22420 4870
rect 22444 4868 22500 4870
rect 22524 4868 22580 4870
rect 22604 4868 22660 4870
rect 22684 4868 22740 4870
rect 21546 3576 21602 3632
rect 21454 2488 21510 2544
rect 22364 3834 22420 3836
rect 22444 3834 22500 3836
rect 22524 3834 22580 3836
rect 22604 3834 22660 3836
rect 22684 3834 22740 3836
rect 22364 3782 22366 3834
rect 22366 3782 22418 3834
rect 22418 3782 22420 3834
rect 22444 3782 22482 3834
rect 22482 3782 22494 3834
rect 22494 3782 22500 3834
rect 22524 3782 22546 3834
rect 22546 3782 22558 3834
rect 22558 3782 22580 3834
rect 22604 3782 22610 3834
rect 22610 3782 22622 3834
rect 22622 3782 22660 3834
rect 22684 3782 22686 3834
rect 22686 3782 22738 3834
rect 22738 3782 22740 3834
rect 22364 3780 22420 3782
rect 22444 3780 22500 3782
rect 22524 3780 22580 3782
rect 22604 3780 22660 3782
rect 22684 3780 22740 3782
rect 22364 2746 22420 2748
rect 22444 2746 22500 2748
rect 22524 2746 22580 2748
rect 22604 2746 22660 2748
rect 22684 2746 22740 2748
rect 22364 2694 22366 2746
rect 22366 2694 22418 2746
rect 22418 2694 22420 2746
rect 22444 2694 22482 2746
rect 22482 2694 22494 2746
rect 22494 2694 22500 2746
rect 22524 2694 22546 2746
rect 22546 2694 22558 2746
rect 22558 2694 22580 2746
rect 22604 2694 22610 2746
rect 22610 2694 22622 2746
rect 22622 2694 22660 2746
rect 22684 2694 22686 2746
rect 22686 2694 22738 2746
rect 22738 2694 22740 2746
rect 22364 2692 22420 2694
rect 22444 2692 22500 2694
rect 22524 2692 22580 2694
rect 22604 2692 22660 2694
rect 22684 2692 22740 2694
rect 19364 1114 19420 1116
rect 19444 1114 19500 1116
rect 19524 1114 19580 1116
rect 19604 1114 19660 1116
rect 19684 1114 19740 1116
rect 19364 1062 19366 1114
rect 19366 1062 19418 1114
rect 19418 1062 19420 1114
rect 19444 1062 19482 1114
rect 19482 1062 19494 1114
rect 19494 1062 19500 1114
rect 19524 1062 19546 1114
rect 19546 1062 19558 1114
rect 19558 1062 19580 1114
rect 19604 1062 19610 1114
rect 19610 1062 19622 1114
rect 19622 1062 19660 1114
rect 19684 1062 19686 1114
rect 19686 1062 19738 1114
rect 19738 1062 19740 1114
rect 19364 1060 19420 1062
rect 19444 1060 19500 1062
rect 19524 1060 19580 1062
rect 19604 1060 19660 1062
rect 19684 1060 19740 1062
rect 22364 1658 22420 1660
rect 22444 1658 22500 1660
rect 22524 1658 22580 1660
rect 22604 1658 22660 1660
rect 22684 1658 22740 1660
rect 22364 1606 22366 1658
rect 22366 1606 22418 1658
rect 22418 1606 22420 1658
rect 22444 1606 22482 1658
rect 22482 1606 22494 1658
rect 22494 1606 22500 1658
rect 22524 1606 22546 1658
rect 22546 1606 22558 1658
rect 22558 1606 22580 1658
rect 22604 1606 22610 1658
rect 22610 1606 22622 1658
rect 22622 1606 22660 1658
rect 22684 1606 22686 1658
rect 22686 1606 22738 1658
rect 22738 1606 22740 1658
rect 22364 1604 22420 1606
rect 22444 1604 22500 1606
rect 22524 1604 22580 1606
rect 22604 1604 22660 1606
rect 22684 1604 22740 1606
rect 22364 570 22420 572
rect 22444 570 22500 572
rect 22524 570 22580 572
rect 22604 570 22660 572
rect 22684 570 22740 572
rect 22364 518 22366 570
rect 22366 518 22418 570
rect 22418 518 22420 570
rect 22444 518 22482 570
rect 22482 518 22494 570
rect 22494 518 22500 570
rect 22524 518 22546 570
rect 22546 518 22558 570
rect 22558 518 22580 570
rect 22604 518 22610 570
rect 22610 518 22622 570
rect 22622 518 22660 570
rect 22684 518 22686 570
rect 22686 518 22738 570
rect 22738 518 22740 570
rect 22364 516 22420 518
rect 22444 516 22500 518
rect 22524 516 22580 518
rect 22604 516 22660 518
rect 22684 516 22740 518
<< metal3 >>
rect 1354 15264 1750 15265
rect 1354 15200 1360 15264
rect 1424 15200 1440 15264
rect 1504 15200 1520 15264
rect 1584 15200 1600 15264
rect 1664 15200 1680 15264
rect 1744 15200 1750 15264
rect 1354 15199 1750 15200
rect 7354 15264 7750 15265
rect 7354 15200 7360 15264
rect 7424 15200 7440 15264
rect 7504 15200 7520 15264
rect 7584 15200 7600 15264
rect 7664 15200 7680 15264
rect 7744 15200 7750 15264
rect 7354 15199 7750 15200
rect 13354 15264 13750 15265
rect 13354 15200 13360 15264
rect 13424 15200 13440 15264
rect 13504 15200 13520 15264
rect 13584 15200 13600 15264
rect 13664 15200 13680 15264
rect 13744 15200 13750 15264
rect 13354 15199 13750 15200
rect 19354 15264 19750 15265
rect 19354 15200 19360 15264
rect 19424 15200 19440 15264
rect 19504 15200 19520 15264
rect 19584 15200 19600 15264
rect 19664 15200 19680 15264
rect 19744 15200 19750 15264
rect 19354 15199 19750 15200
rect 4354 14720 4750 14721
rect 4354 14656 4360 14720
rect 4424 14656 4440 14720
rect 4504 14656 4520 14720
rect 4584 14656 4600 14720
rect 4664 14656 4680 14720
rect 4744 14656 4750 14720
rect 4354 14655 4750 14656
rect 10354 14720 10750 14721
rect 10354 14656 10360 14720
rect 10424 14656 10440 14720
rect 10504 14656 10520 14720
rect 10584 14656 10600 14720
rect 10664 14656 10680 14720
rect 10744 14656 10750 14720
rect 10354 14655 10750 14656
rect 16354 14720 16750 14721
rect 16354 14656 16360 14720
rect 16424 14656 16440 14720
rect 16504 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16750 14720
rect 16354 14655 16750 14656
rect 22354 14720 22750 14721
rect 22354 14656 22360 14720
rect 22424 14656 22440 14720
rect 22504 14656 22520 14720
rect 22584 14656 22600 14720
rect 22664 14656 22680 14720
rect 22744 14656 22750 14720
rect 22354 14655 22750 14656
rect 17953 14514 18019 14517
rect 18873 14514 18939 14517
rect 17953 14512 18939 14514
rect 17953 14456 17958 14512
rect 18014 14456 18878 14512
rect 18934 14456 18939 14512
rect 17953 14454 18939 14456
rect 17953 14451 18019 14454
rect 18873 14451 18939 14454
rect 15837 14378 15903 14381
rect 17125 14378 17191 14381
rect 15837 14376 17191 14378
rect 15837 14320 15842 14376
rect 15898 14320 17130 14376
rect 17186 14320 17191 14376
rect 15837 14318 17191 14320
rect 15837 14315 15903 14318
rect 17125 14315 17191 14318
rect 1354 14176 1750 14177
rect 1354 14112 1360 14176
rect 1424 14112 1440 14176
rect 1504 14112 1520 14176
rect 1584 14112 1600 14176
rect 1664 14112 1680 14176
rect 1744 14112 1750 14176
rect 1354 14111 1750 14112
rect 7354 14176 7750 14177
rect 7354 14112 7360 14176
rect 7424 14112 7440 14176
rect 7504 14112 7520 14176
rect 7584 14112 7600 14176
rect 7664 14112 7680 14176
rect 7744 14112 7750 14176
rect 7354 14111 7750 14112
rect 13354 14176 13750 14177
rect 13354 14112 13360 14176
rect 13424 14112 13440 14176
rect 13504 14112 13520 14176
rect 13584 14112 13600 14176
rect 13664 14112 13680 14176
rect 13744 14112 13750 14176
rect 13354 14111 13750 14112
rect 19354 14176 19750 14177
rect 19354 14112 19360 14176
rect 19424 14112 19440 14176
rect 19504 14112 19520 14176
rect 19584 14112 19600 14176
rect 19664 14112 19680 14176
rect 19744 14112 19750 14176
rect 19354 14111 19750 14112
rect 13813 13970 13879 13973
rect 18597 13970 18663 13973
rect 13813 13968 18663 13970
rect 13813 13912 13818 13968
rect 13874 13912 18602 13968
rect 18658 13912 18663 13968
rect 13813 13910 18663 13912
rect 13813 13907 13879 13910
rect 18597 13907 18663 13910
rect 20069 13970 20135 13973
rect 23600 13970 24000 14000
rect 20069 13968 24000 13970
rect 20069 13912 20074 13968
rect 20130 13912 24000 13968
rect 20069 13910 24000 13912
rect 20069 13907 20135 13910
rect 23600 13880 24000 13910
rect 10501 13834 10567 13837
rect 14641 13834 14707 13837
rect 18597 13834 18663 13837
rect 10501 13832 14474 13834
rect 10501 13776 10506 13832
rect 10562 13776 14474 13832
rect 10501 13774 14474 13776
rect 10501 13771 10567 13774
rect 14414 13698 14474 13774
rect 14641 13832 18663 13834
rect 14641 13776 14646 13832
rect 14702 13776 18602 13832
rect 18658 13776 18663 13832
rect 14641 13774 18663 13776
rect 14641 13771 14707 13774
rect 18597 13771 18663 13774
rect 15837 13698 15903 13701
rect 14414 13696 15903 13698
rect 14414 13640 15842 13696
rect 15898 13640 15903 13696
rect 14414 13638 15903 13640
rect 15837 13635 15903 13638
rect 4354 13632 4750 13633
rect 4354 13568 4360 13632
rect 4424 13568 4440 13632
rect 4504 13568 4520 13632
rect 4584 13568 4600 13632
rect 4664 13568 4680 13632
rect 4744 13568 4750 13632
rect 4354 13567 4750 13568
rect 10354 13632 10750 13633
rect 10354 13568 10360 13632
rect 10424 13568 10440 13632
rect 10504 13568 10520 13632
rect 10584 13568 10600 13632
rect 10664 13568 10680 13632
rect 10744 13568 10750 13632
rect 10354 13567 10750 13568
rect 16354 13632 16750 13633
rect 16354 13568 16360 13632
rect 16424 13568 16440 13632
rect 16504 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16750 13632
rect 16354 13567 16750 13568
rect 22354 13632 22750 13633
rect 22354 13568 22360 13632
rect 22424 13568 22440 13632
rect 22504 13568 22520 13632
rect 22584 13568 22600 13632
rect 22664 13568 22680 13632
rect 22744 13568 22750 13632
rect 22354 13567 22750 13568
rect 13118 13364 13124 13428
rect 13188 13426 13194 13428
rect 18873 13426 18939 13429
rect 13188 13424 18939 13426
rect 13188 13368 18878 13424
rect 18934 13368 18939 13424
rect 13188 13366 18939 13368
rect 13188 13364 13194 13366
rect 18873 13363 18939 13366
rect 8109 13290 8175 13293
rect 11789 13290 11855 13293
rect 8109 13288 11855 13290
rect 8109 13232 8114 13288
rect 8170 13232 11794 13288
rect 11850 13232 11855 13288
rect 8109 13230 11855 13232
rect 8109 13227 8175 13230
rect 11789 13227 11855 13230
rect 1354 13088 1750 13089
rect 1354 13024 1360 13088
rect 1424 13024 1440 13088
rect 1504 13024 1520 13088
rect 1584 13024 1600 13088
rect 1664 13024 1680 13088
rect 1744 13024 1750 13088
rect 1354 13023 1750 13024
rect 7354 13088 7750 13089
rect 7354 13024 7360 13088
rect 7424 13024 7440 13088
rect 7504 13024 7520 13088
rect 7584 13024 7600 13088
rect 7664 13024 7680 13088
rect 7744 13024 7750 13088
rect 7354 13023 7750 13024
rect 13354 13088 13750 13089
rect 13354 13024 13360 13088
rect 13424 13024 13440 13088
rect 13504 13024 13520 13088
rect 13584 13024 13600 13088
rect 13664 13024 13680 13088
rect 13744 13024 13750 13088
rect 13354 13023 13750 13024
rect 19354 13088 19750 13089
rect 19354 13024 19360 13088
rect 19424 13024 19440 13088
rect 19504 13024 19520 13088
rect 19584 13024 19600 13088
rect 19664 13024 19680 13088
rect 19744 13024 19750 13088
rect 19354 13023 19750 13024
rect 9489 12882 9555 12885
rect 12893 12882 12959 12885
rect 15694 12882 15700 12884
rect 9489 12880 15700 12882
rect 9489 12824 9494 12880
rect 9550 12824 12898 12880
rect 12954 12824 15700 12880
rect 9489 12822 15700 12824
rect 9489 12819 9555 12822
rect 12893 12819 12959 12822
rect 15694 12820 15700 12822
rect 15764 12820 15770 12884
rect 23289 12882 23355 12885
rect 23600 12882 24000 12912
rect 23289 12880 24000 12882
rect 23289 12824 23294 12880
rect 23350 12824 24000 12880
rect 23289 12822 24000 12824
rect 23289 12819 23355 12822
rect 23600 12792 24000 12822
rect 1761 12746 1827 12749
rect 2957 12746 3023 12749
rect 1761 12744 3023 12746
rect 1761 12688 1766 12744
rect 1822 12688 2962 12744
rect 3018 12688 3023 12744
rect 1761 12686 3023 12688
rect 1761 12683 1827 12686
rect 2957 12683 3023 12686
rect 9673 12746 9739 12749
rect 11145 12746 11211 12749
rect 9673 12744 11211 12746
rect 9673 12688 9678 12744
rect 9734 12688 11150 12744
rect 11206 12688 11211 12744
rect 9673 12686 11211 12688
rect 9673 12683 9739 12686
rect 11145 12683 11211 12686
rect 11145 12610 11211 12613
rect 13721 12610 13787 12613
rect 11145 12608 13787 12610
rect 11145 12552 11150 12608
rect 11206 12552 13726 12608
rect 13782 12552 13787 12608
rect 11145 12550 13787 12552
rect 11145 12547 11211 12550
rect 13721 12547 13787 12550
rect 14641 12610 14707 12613
rect 14958 12610 14964 12612
rect 14641 12608 14964 12610
rect 14641 12552 14646 12608
rect 14702 12552 14964 12608
rect 14641 12550 14964 12552
rect 14641 12547 14707 12550
rect 14958 12548 14964 12550
rect 15028 12548 15034 12612
rect 4354 12544 4750 12545
rect 4354 12480 4360 12544
rect 4424 12480 4440 12544
rect 4504 12480 4520 12544
rect 4584 12480 4600 12544
rect 4664 12480 4680 12544
rect 4744 12480 4750 12544
rect 4354 12479 4750 12480
rect 10354 12544 10750 12545
rect 10354 12480 10360 12544
rect 10424 12480 10440 12544
rect 10504 12480 10520 12544
rect 10584 12480 10600 12544
rect 10664 12480 10680 12544
rect 10744 12480 10750 12544
rect 10354 12479 10750 12480
rect 16354 12544 16750 12545
rect 16354 12480 16360 12544
rect 16424 12480 16440 12544
rect 16504 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16750 12544
rect 16354 12479 16750 12480
rect 22354 12544 22750 12545
rect 22354 12480 22360 12544
rect 22424 12480 22440 12544
rect 22504 12480 22520 12544
rect 22584 12480 22600 12544
rect 22664 12480 22680 12544
rect 22744 12480 22750 12544
rect 22354 12479 22750 12480
rect 15837 12474 15903 12477
rect 11286 12472 15903 12474
rect 11286 12416 15842 12472
rect 15898 12416 15903 12472
rect 11286 12414 15903 12416
rect 1853 12338 1919 12341
rect 2497 12338 2563 12341
rect 1853 12336 2563 12338
rect 1853 12280 1858 12336
rect 1914 12280 2502 12336
rect 2558 12280 2563 12336
rect 1853 12278 2563 12280
rect 1853 12275 1919 12278
rect 2497 12275 2563 12278
rect 10133 12338 10199 12341
rect 11286 12338 11346 12414
rect 15837 12411 15903 12414
rect 10133 12336 11346 12338
rect 10133 12280 10138 12336
rect 10194 12280 11346 12336
rect 10133 12278 11346 12280
rect 11513 12338 11579 12341
rect 18321 12338 18387 12341
rect 11513 12336 18387 12338
rect 11513 12280 11518 12336
rect 11574 12280 18326 12336
rect 18382 12280 18387 12336
rect 11513 12278 18387 12280
rect 10133 12275 10199 12278
rect 11513 12275 11579 12278
rect 18321 12275 18387 12278
rect 10593 12202 10659 12205
rect 17401 12202 17467 12205
rect 10593 12200 17467 12202
rect 10593 12144 10598 12200
rect 10654 12144 17406 12200
rect 17462 12144 17467 12200
rect 10593 12142 17467 12144
rect 10593 12139 10659 12142
rect 17401 12139 17467 12142
rect 9765 12066 9831 12069
rect 11605 12066 11671 12069
rect 9765 12064 11671 12066
rect 9765 12008 9770 12064
rect 9826 12008 11610 12064
rect 11666 12008 11671 12064
rect 9765 12006 11671 12008
rect 9765 12003 9831 12006
rect 11605 12003 11671 12006
rect 1354 12000 1750 12001
rect 1354 11936 1360 12000
rect 1424 11936 1440 12000
rect 1504 11936 1520 12000
rect 1584 11936 1600 12000
rect 1664 11936 1680 12000
rect 1744 11936 1750 12000
rect 1354 11935 1750 11936
rect 7354 12000 7750 12001
rect 7354 11936 7360 12000
rect 7424 11936 7440 12000
rect 7504 11936 7520 12000
rect 7584 11936 7600 12000
rect 7664 11936 7680 12000
rect 7744 11936 7750 12000
rect 7354 11935 7750 11936
rect 13354 12000 13750 12001
rect 13354 11936 13360 12000
rect 13424 11936 13440 12000
rect 13504 11936 13520 12000
rect 13584 11936 13600 12000
rect 13664 11936 13680 12000
rect 13744 11936 13750 12000
rect 13354 11935 13750 11936
rect 19354 12000 19750 12001
rect 19354 11936 19360 12000
rect 19424 11936 19440 12000
rect 19504 11936 19520 12000
rect 19584 11936 19600 12000
rect 19664 11936 19680 12000
rect 19744 11936 19750 12000
rect 19354 11935 19750 11936
rect 2589 11794 2655 11797
rect 3417 11794 3483 11797
rect 2589 11792 3483 11794
rect 2589 11736 2594 11792
rect 2650 11736 3422 11792
rect 3478 11736 3483 11792
rect 2589 11734 3483 11736
rect 2589 11731 2655 11734
rect 3417 11731 3483 11734
rect 12985 11794 13051 11797
rect 16021 11794 16087 11797
rect 16757 11794 16823 11797
rect 12985 11792 16823 11794
rect 12985 11736 12990 11792
rect 13046 11736 16026 11792
rect 16082 11736 16762 11792
rect 16818 11736 16823 11792
rect 12985 11734 16823 11736
rect 12985 11731 13051 11734
rect 16021 11731 16087 11734
rect 16757 11731 16823 11734
rect 5165 11658 5231 11661
rect 6821 11658 6887 11661
rect 20713 11658 20779 11661
rect 5165 11656 20779 11658
rect 5165 11600 5170 11656
rect 5226 11600 6826 11656
rect 6882 11600 20718 11656
rect 20774 11600 20779 11656
rect 5165 11598 20779 11600
rect 5165 11595 5231 11598
rect 6821 11595 6887 11598
rect 20713 11595 20779 11598
rect 2957 11522 3023 11525
rect 4102 11522 4108 11524
rect 2957 11520 4108 11522
rect 2957 11464 2962 11520
rect 3018 11464 4108 11520
rect 2957 11462 4108 11464
rect 2957 11459 3023 11462
rect 4102 11460 4108 11462
rect 4172 11460 4178 11524
rect 4354 11456 4750 11457
rect 4354 11392 4360 11456
rect 4424 11392 4440 11456
rect 4504 11392 4520 11456
rect 4584 11392 4600 11456
rect 4664 11392 4680 11456
rect 4744 11392 4750 11456
rect 4354 11391 4750 11392
rect 10354 11456 10750 11457
rect 10354 11392 10360 11456
rect 10424 11392 10440 11456
rect 10504 11392 10520 11456
rect 10584 11392 10600 11456
rect 10664 11392 10680 11456
rect 10744 11392 10750 11456
rect 10354 11391 10750 11392
rect 16354 11456 16750 11457
rect 16354 11392 16360 11456
rect 16424 11392 16440 11456
rect 16504 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16750 11456
rect 16354 11391 16750 11392
rect 22354 11456 22750 11457
rect 22354 11392 22360 11456
rect 22424 11392 22440 11456
rect 22504 11392 22520 11456
rect 22584 11392 22600 11456
rect 22664 11392 22680 11456
rect 22744 11392 22750 11456
rect 22354 11391 22750 11392
rect 5349 11386 5415 11389
rect 4892 11384 5415 11386
rect 4892 11328 5354 11384
rect 5410 11328 5415 11384
rect 4892 11326 5415 11328
rect 4892 11253 4952 11326
rect 5349 11323 5415 11326
rect 11145 11386 11211 11389
rect 13905 11386 13971 11389
rect 14641 11386 14707 11389
rect 11145 11384 14707 11386
rect 11145 11328 11150 11384
rect 11206 11328 13910 11384
rect 13966 11328 14646 11384
rect 14702 11328 14707 11384
rect 11145 11326 14707 11328
rect 11145 11323 11211 11326
rect 13905 11323 13971 11326
rect 14641 11323 14707 11326
rect 4889 11248 4955 11253
rect 4889 11192 4894 11248
rect 4950 11192 4955 11248
rect 4889 11187 4955 11192
rect 4337 11114 4403 11117
rect 7189 11114 7255 11117
rect 4337 11112 7255 11114
rect 4337 11056 4342 11112
rect 4398 11056 7194 11112
rect 7250 11056 7255 11112
rect 4337 11054 7255 11056
rect 4337 11051 4403 11054
rect 7189 11051 7255 11054
rect 13813 11114 13879 11117
rect 17953 11114 18019 11117
rect 13813 11112 18019 11114
rect 13813 11056 13818 11112
rect 13874 11056 17958 11112
rect 18014 11056 18019 11112
rect 13813 11054 18019 11056
rect 13813 11051 13879 11054
rect 17953 11051 18019 11054
rect 19701 11114 19767 11117
rect 20621 11114 20687 11117
rect 19701 11112 20687 11114
rect 19701 11056 19706 11112
rect 19762 11056 20626 11112
rect 20682 11056 20687 11112
rect 19701 11054 20687 11056
rect 19701 11051 19767 11054
rect 20621 11051 20687 11054
rect 1354 10912 1750 10913
rect 1354 10848 1360 10912
rect 1424 10848 1440 10912
rect 1504 10848 1520 10912
rect 1584 10848 1600 10912
rect 1664 10848 1680 10912
rect 1744 10848 1750 10912
rect 1354 10847 1750 10848
rect 7354 10912 7750 10913
rect 7354 10848 7360 10912
rect 7424 10848 7440 10912
rect 7504 10848 7520 10912
rect 7584 10848 7600 10912
rect 7664 10848 7680 10912
rect 7744 10848 7750 10912
rect 7354 10847 7750 10848
rect 13354 10912 13750 10913
rect 13354 10848 13360 10912
rect 13424 10848 13440 10912
rect 13504 10848 13520 10912
rect 13584 10848 13600 10912
rect 13664 10848 13680 10912
rect 13744 10848 13750 10912
rect 13354 10847 13750 10848
rect 19354 10912 19750 10913
rect 19354 10848 19360 10912
rect 19424 10848 19440 10912
rect 19504 10848 19520 10912
rect 19584 10848 19600 10912
rect 19664 10848 19680 10912
rect 19744 10848 19750 10912
rect 19354 10847 19750 10848
rect 8201 10706 8267 10709
rect 17125 10706 17191 10709
rect 8201 10704 17191 10706
rect 8201 10648 8206 10704
rect 8262 10648 17130 10704
rect 17186 10648 17191 10704
rect 8201 10646 17191 10648
rect 8201 10643 8267 10646
rect 17125 10643 17191 10646
rect 2681 10570 2747 10573
rect 16849 10570 16915 10573
rect 2681 10568 16915 10570
rect 2681 10512 2686 10568
rect 2742 10512 16854 10568
rect 16910 10512 16915 10568
rect 2681 10510 16915 10512
rect 2681 10507 2747 10510
rect 16849 10507 16915 10510
rect 6913 10434 6979 10437
rect 9397 10434 9463 10437
rect 6913 10432 9463 10434
rect 6913 10376 6918 10432
rect 6974 10376 9402 10432
rect 9458 10376 9463 10432
rect 6913 10374 9463 10376
rect 6913 10371 6979 10374
rect 9397 10371 9463 10374
rect 12249 10434 12315 10437
rect 14549 10434 14615 10437
rect 12249 10432 14615 10434
rect 12249 10376 12254 10432
rect 12310 10376 14554 10432
rect 14610 10376 14615 10432
rect 12249 10374 14615 10376
rect 12249 10371 12315 10374
rect 14549 10371 14615 10374
rect 4354 10368 4750 10369
rect 4354 10304 4360 10368
rect 4424 10304 4440 10368
rect 4504 10304 4520 10368
rect 4584 10304 4600 10368
rect 4664 10304 4680 10368
rect 4744 10304 4750 10368
rect 4354 10303 4750 10304
rect 10354 10368 10750 10369
rect 10354 10304 10360 10368
rect 10424 10304 10440 10368
rect 10504 10304 10520 10368
rect 10584 10304 10600 10368
rect 10664 10304 10680 10368
rect 10744 10304 10750 10368
rect 10354 10303 10750 10304
rect 16354 10368 16750 10369
rect 16354 10304 16360 10368
rect 16424 10304 16440 10368
rect 16504 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16750 10368
rect 16354 10303 16750 10304
rect 22354 10368 22750 10369
rect 22354 10304 22360 10368
rect 22424 10304 22440 10368
rect 22504 10304 22520 10368
rect 22584 10304 22600 10368
rect 22664 10304 22680 10368
rect 22744 10304 22750 10368
rect 22354 10303 22750 10304
rect 11605 10298 11671 10301
rect 13169 10298 13235 10301
rect 11605 10296 13235 10298
rect 11605 10240 11610 10296
rect 11666 10240 13174 10296
rect 13230 10240 13235 10296
rect 11605 10238 13235 10240
rect 11605 10235 11671 10238
rect 13169 10235 13235 10238
rect 14733 10298 14799 10301
rect 15142 10298 15148 10300
rect 14733 10296 15148 10298
rect 14733 10240 14738 10296
rect 14794 10240 15148 10296
rect 14733 10238 15148 10240
rect 14733 10235 14799 10238
rect 15142 10236 15148 10238
rect 15212 10236 15218 10300
rect 1669 10162 1735 10165
rect 19057 10162 19123 10165
rect 1669 10160 19123 10162
rect 1669 10104 1674 10160
rect 1730 10104 19062 10160
rect 19118 10104 19123 10160
rect 1669 10102 19123 10104
rect 1669 10099 1735 10102
rect 19057 10099 19123 10102
rect 4061 10026 4127 10029
rect 19333 10026 19399 10029
rect 4061 10024 19399 10026
rect 4061 9968 4066 10024
rect 4122 9968 19338 10024
rect 19394 9968 19399 10024
rect 4061 9966 19399 9968
rect 4061 9963 4127 9966
rect 19333 9963 19399 9966
rect 19885 9890 19951 9893
rect 20989 9890 21055 9893
rect 19885 9888 21055 9890
rect 19885 9832 19890 9888
rect 19946 9832 20994 9888
rect 21050 9832 21055 9888
rect 19885 9830 21055 9832
rect 19885 9827 19951 9830
rect 20989 9827 21055 9830
rect 1354 9824 1750 9825
rect 1354 9760 1360 9824
rect 1424 9760 1440 9824
rect 1504 9760 1520 9824
rect 1584 9760 1600 9824
rect 1664 9760 1680 9824
rect 1744 9760 1750 9824
rect 1354 9759 1750 9760
rect 7354 9824 7750 9825
rect 7354 9760 7360 9824
rect 7424 9760 7440 9824
rect 7504 9760 7520 9824
rect 7584 9760 7600 9824
rect 7664 9760 7680 9824
rect 7744 9760 7750 9824
rect 7354 9759 7750 9760
rect 13354 9824 13750 9825
rect 13354 9760 13360 9824
rect 13424 9760 13440 9824
rect 13504 9760 13520 9824
rect 13584 9760 13600 9824
rect 13664 9760 13680 9824
rect 13744 9760 13750 9824
rect 13354 9759 13750 9760
rect 19354 9824 19750 9825
rect 19354 9760 19360 9824
rect 19424 9760 19440 9824
rect 19504 9760 19520 9824
rect 19584 9760 19600 9824
rect 19664 9760 19680 9824
rect 19744 9760 19750 9824
rect 19354 9759 19750 9760
rect 9029 9754 9095 9757
rect 9806 9754 9812 9756
rect 9029 9752 9812 9754
rect 9029 9696 9034 9752
rect 9090 9696 9812 9752
rect 9029 9694 9812 9696
rect 9029 9691 9095 9694
rect 9806 9692 9812 9694
rect 9876 9692 9882 9756
rect 3785 9618 3851 9621
rect 19333 9618 19399 9621
rect 19977 9618 20043 9621
rect 3785 9616 20043 9618
rect 3785 9560 3790 9616
rect 3846 9560 19338 9616
rect 19394 9560 19982 9616
rect 20038 9560 20043 9616
rect 3785 9558 20043 9560
rect 3785 9555 3851 9558
rect 19333 9555 19399 9558
rect 19977 9555 20043 9558
rect 20253 9618 20319 9621
rect 21265 9618 21331 9621
rect 21633 9618 21699 9621
rect 20253 9616 21699 9618
rect 20253 9560 20258 9616
rect 20314 9560 21270 9616
rect 21326 9560 21638 9616
rect 21694 9560 21699 9616
rect 20253 9558 21699 9560
rect 20253 9555 20319 9558
rect 21265 9555 21331 9558
rect 21633 9555 21699 9558
rect 10685 9482 10751 9485
rect 11094 9482 11100 9484
rect 10685 9480 11100 9482
rect 10685 9424 10690 9480
rect 10746 9424 11100 9480
rect 10685 9422 11100 9424
rect 10685 9419 10751 9422
rect 11094 9420 11100 9422
rect 11164 9420 11170 9484
rect 16665 9482 16731 9485
rect 17769 9482 17835 9485
rect 16665 9480 17835 9482
rect 16665 9424 16670 9480
rect 16726 9424 17774 9480
rect 17830 9424 17835 9480
rect 16665 9422 17835 9424
rect 16665 9419 16731 9422
rect 17769 9419 17835 9422
rect 21081 9482 21147 9485
rect 22093 9482 22159 9485
rect 21081 9480 22159 9482
rect 21081 9424 21086 9480
rect 21142 9424 22098 9480
rect 22154 9424 22159 9480
rect 21081 9422 22159 9424
rect 21081 9419 21147 9422
rect 22093 9419 22159 9422
rect 12341 9346 12407 9349
rect 12709 9346 12775 9349
rect 12341 9344 12775 9346
rect 12341 9288 12346 9344
rect 12402 9288 12714 9344
rect 12770 9288 12775 9344
rect 12341 9286 12775 9288
rect 12341 9283 12407 9286
rect 12709 9283 12775 9286
rect 4354 9280 4750 9281
rect 4354 9216 4360 9280
rect 4424 9216 4440 9280
rect 4504 9216 4520 9280
rect 4584 9216 4600 9280
rect 4664 9216 4680 9280
rect 4744 9216 4750 9280
rect 4354 9215 4750 9216
rect 10354 9280 10750 9281
rect 10354 9216 10360 9280
rect 10424 9216 10440 9280
rect 10504 9216 10520 9280
rect 10584 9216 10600 9280
rect 10664 9216 10680 9280
rect 10744 9216 10750 9280
rect 10354 9215 10750 9216
rect 16354 9280 16750 9281
rect 16354 9216 16360 9280
rect 16424 9216 16440 9280
rect 16504 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16750 9280
rect 16354 9215 16750 9216
rect 22354 9280 22750 9281
rect 22354 9216 22360 9280
rect 22424 9216 22440 9280
rect 22504 9216 22520 9280
rect 22584 9216 22600 9280
rect 22664 9216 22680 9280
rect 22744 9216 22750 9280
rect 22354 9215 22750 9216
rect 13353 9210 13419 9213
rect 14774 9210 14780 9212
rect 13353 9208 14780 9210
rect 13353 9152 13358 9208
rect 13414 9152 14780 9208
rect 13353 9150 14780 9152
rect 13353 9147 13419 9150
rect 14774 9148 14780 9150
rect 14844 9148 14850 9212
rect 19425 9210 19491 9213
rect 19926 9210 19932 9212
rect 19425 9208 19932 9210
rect 19425 9152 19430 9208
rect 19486 9152 19932 9208
rect 19425 9150 19932 9152
rect 19425 9147 19491 9150
rect 19926 9148 19932 9150
rect 19996 9148 20002 9212
rect 11789 9074 11855 9077
rect 13629 9074 13695 9077
rect 11789 9072 13695 9074
rect 11789 9016 11794 9072
rect 11850 9016 13634 9072
rect 13690 9016 13695 9072
rect 11789 9014 13695 9016
rect 11789 9011 11855 9014
rect 13629 9011 13695 9014
rect 14641 9074 14707 9077
rect 15377 9074 15443 9077
rect 14641 9072 15443 9074
rect 14641 9016 14646 9072
rect 14702 9016 15382 9072
rect 15438 9016 15443 9072
rect 14641 9014 15443 9016
rect 14641 9011 14707 9014
rect 15377 9011 15443 9014
rect 19701 9074 19767 9077
rect 21357 9074 21423 9077
rect 19701 9072 21423 9074
rect 19701 9016 19706 9072
rect 19762 9016 21362 9072
rect 21418 9016 21423 9072
rect 19701 9014 21423 9016
rect 19701 9011 19767 9014
rect 21357 9011 21423 9014
rect 10225 8938 10291 8941
rect 20805 8938 20871 8941
rect 10225 8936 20871 8938
rect 10225 8880 10230 8936
rect 10286 8880 20810 8936
rect 20866 8880 20871 8936
rect 10225 8878 20871 8880
rect 10225 8875 10291 8878
rect 20805 8875 20871 8878
rect 9857 8802 9923 8805
rect 9814 8800 9923 8802
rect 9814 8744 9862 8800
rect 9918 8744 9923 8800
rect 9814 8739 9923 8744
rect 15009 8802 15075 8805
rect 16021 8802 16087 8805
rect 15009 8800 16087 8802
rect 15009 8744 15014 8800
rect 15070 8744 16026 8800
rect 16082 8744 16087 8800
rect 15009 8742 16087 8744
rect 15009 8739 15075 8742
rect 16021 8739 16087 8742
rect 1354 8736 1750 8737
rect 1354 8672 1360 8736
rect 1424 8672 1440 8736
rect 1504 8672 1520 8736
rect 1584 8672 1600 8736
rect 1664 8672 1680 8736
rect 1744 8672 1750 8736
rect 1354 8671 1750 8672
rect 7354 8736 7750 8737
rect 7354 8672 7360 8736
rect 7424 8672 7440 8736
rect 7504 8672 7520 8736
rect 7584 8672 7600 8736
rect 7664 8672 7680 8736
rect 7744 8672 7750 8736
rect 7354 8671 7750 8672
rect 2129 8666 2195 8669
rect 3049 8666 3115 8669
rect 2129 8664 3115 8666
rect 2129 8608 2134 8664
rect 2190 8608 3054 8664
rect 3110 8608 3115 8664
rect 2129 8606 3115 8608
rect 2129 8603 2195 8606
rect 3049 8603 3115 8606
rect 9814 8533 9874 8739
rect 13354 8736 13750 8737
rect 13354 8672 13360 8736
rect 13424 8672 13440 8736
rect 13504 8672 13520 8736
rect 13584 8672 13600 8736
rect 13664 8672 13680 8736
rect 13744 8672 13750 8736
rect 13354 8671 13750 8672
rect 19354 8736 19750 8737
rect 19354 8672 19360 8736
rect 19424 8672 19440 8736
rect 19504 8672 19520 8736
rect 19584 8672 19600 8736
rect 19664 8672 19680 8736
rect 19744 8672 19750 8736
rect 19354 8671 19750 8672
rect 17217 8666 17283 8669
rect 17769 8666 17835 8669
rect 17217 8664 17835 8666
rect 17217 8608 17222 8664
rect 17278 8608 17774 8664
rect 17830 8608 17835 8664
rect 17217 8606 17835 8608
rect 17217 8603 17283 8606
rect 17769 8603 17835 8606
rect 9814 8528 9923 8533
rect 9814 8472 9862 8528
rect 9918 8472 9923 8528
rect 9814 8470 9923 8472
rect 9857 8467 9923 8470
rect 15469 8530 15535 8533
rect 17309 8530 17375 8533
rect 15469 8528 17375 8530
rect 15469 8472 15474 8528
rect 15530 8472 17314 8528
rect 17370 8472 17375 8528
rect 15469 8470 17375 8472
rect 15469 8467 15535 8470
rect 17309 8467 17375 8470
rect 17769 8530 17835 8533
rect 21633 8530 21699 8533
rect 17769 8528 21699 8530
rect 17769 8472 17774 8528
rect 17830 8472 21638 8528
rect 21694 8472 21699 8528
rect 17769 8470 21699 8472
rect 17769 8467 17835 8470
rect 21633 8467 21699 8470
rect 9489 8394 9555 8397
rect 16573 8394 16639 8397
rect 9489 8392 16639 8394
rect 9489 8336 9494 8392
rect 9550 8336 16578 8392
rect 16634 8336 16639 8392
rect 9489 8334 16639 8336
rect 9489 8331 9555 8334
rect 16573 8331 16639 8334
rect 18781 8394 18847 8397
rect 20713 8394 20779 8397
rect 18781 8392 20779 8394
rect 18781 8336 18786 8392
rect 18842 8336 20718 8392
rect 20774 8336 20779 8392
rect 18781 8334 20779 8336
rect 18781 8331 18847 8334
rect 20713 8331 20779 8334
rect 12433 8258 12499 8261
rect 15653 8258 15719 8261
rect 19977 8260 20043 8261
rect 19926 8258 19932 8260
rect 12433 8256 15719 8258
rect 12433 8200 12438 8256
rect 12494 8200 15658 8256
rect 15714 8200 15719 8256
rect 12433 8198 15719 8200
rect 19886 8198 19932 8258
rect 19996 8256 20043 8260
rect 20038 8200 20043 8256
rect 12433 8195 12499 8198
rect 15653 8195 15719 8198
rect 19926 8196 19932 8198
rect 19996 8196 20043 8200
rect 19977 8195 20043 8196
rect 20253 8258 20319 8261
rect 21265 8258 21331 8261
rect 20253 8256 21331 8258
rect 20253 8200 20258 8256
rect 20314 8200 21270 8256
rect 21326 8200 21331 8256
rect 20253 8198 21331 8200
rect 20253 8195 20319 8198
rect 21265 8195 21331 8198
rect 4354 8192 4750 8193
rect 4354 8128 4360 8192
rect 4424 8128 4440 8192
rect 4504 8128 4520 8192
rect 4584 8128 4600 8192
rect 4664 8128 4680 8192
rect 4744 8128 4750 8192
rect 4354 8127 4750 8128
rect 10354 8192 10750 8193
rect 10354 8128 10360 8192
rect 10424 8128 10440 8192
rect 10504 8128 10520 8192
rect 10584 8128 10600 8192
rect 10664 8128 10680 8192
rect 10744 8128 10750 8192
rect 10354 8127 10750 8128
rect 16354 8192 16750 8193
rect 16354 8128 16360 8192
rect 16424 8128 16440 8192
rect 16504 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16750 8192
rect 16354 8127 16750 8128
rect 22354 8192 22750 8193
rect 22354 8128 22360 8192
rect 22424 8128 22440 8192
rect 22504 8128 22520 8192
rect 22584 8128 22600 8192
rect 22664 8128 22680 8192
rect 22744 8128 22750 8192
rect 22354 8127 22750 8128
rect 12525 8122 12591 8125
rect 13997 8122 14063 8125
rect 12525 8120 14063 8122
rect 12525 8064 12530 8120
rect 12586 8064 14002 8120
rect 14058 8064 14063 8120
rect 12525 8062 14063 8064
rect 12525 8059 12591 8062
rect 13997 8059 14063 8062
rect 3509 7986 3575 7989
rect 9121 7986 9187 7989
rect 3509 7984 9187 7986
rect 3509 7928 3514 7984
rect 3570 7928 9126 7984
rect 9182 7928 9187 7984
rect 3509 7926 9187 7928
rect 3509 7923 3575 7926
rect 9121 7923 9187 7926
rect 13721 7986 13787 7989
rect 17493 7986 17559 7989
rect 13721 7984 17559 7986
rect 13721 7928 13726 7984
rect 13782 7928 17498 7984
rect 17554 7928 17559 7984
rect 13721 7926 17559 7928
rect 13721 7923 13787 7926
rect 17493 7923 17559 7926
rect 4102 7788 4108 7852
rect 4172 7850 4178 7852
rect 18321 7850 18387 7853
rect 4172 7848 18387 7850
rect 4172 7792 18326 7848
rect 18382 7792 18387 7848
rect 4172 7790 18387 7792
rect 4172 7788 4178 7790
rect 18321 7787 18387 7790
rect 1354 7648 1750 7649
rect 1354 7584 1360 7648
rect 1424 7584 1440 7648
rect 1504 7584 1520 7648
rect 1584 7584 1600 7648
rect 1664 7584 1680 7648
rect 1744 7584 1750 7648
rect 1354 7583 1750 7584
rect 7354 7648 7750 7649
rect 7354 7584 7360 7648
rect 7424 7584 7440 7648
rect 7504 7584 7520 7648
rect 7584 7584 7600 7648
rect 7664 7584 7680 7648
rect 7744 7584 7750 7648
rect 7354 7583 7750 7584
rect 13354 7648 13750 7649
rect 13354 7584 13360 7648
rect 13424 7584 13440 7648
rect 13504 7584 13520 7648
rect 13584 7584 13600 7648
rect 13664 7584 13680 7648
rect 13744 7584 13750 7648
rect 13354 7583 13750 7584
rect 19354 7648 19750 7649
rect 19354 7584 19360 7648
rect 19424 7584 19440 7648
rect 19504 7584 19520 7648
rect 19584 7584 19600 7648
rect 19664 7584 19680 7648
rect 19744 7584 19750 7648
rect 19354 7583 19750 7584
rect 10225 7578 10291 7581
rect 12157 7578 12223 7581
rect 10225 7576 12223 7578
rect 10225 7520 10230 7576
rect 10286 7520 12162 7576
rect 12218 7520 12223 7576
rect 10225 7518 12223 7520
rect 10225 7515 10291 7518
rect 12157 7515 12223 7518
rect 14181 7578 14247 7581
rect 14825 7578 14891 7581
rect 14181 7576 14891 7578
rect 14181 7520 14186 7576
rect 14242 7520 14830 7576
rect 14886 7520 14891 7576
rect 14181 7518 14891 7520
rect 14181 7515 14247 7518
rect 14825 7515 14891 7518
rect 2865 7442 2931 7445
rect 4061 7442 4127 7445
rect 5533 7442 5599 7445
rect 2865 7440 5599 7442
rect 2865 7384 2870 7440
rect 2926 7384 4066 7440
rect 4122 7384 5538 7440
rect 5594 7384 5599 7440
rect 2865 7382 5599 7384
rect 2865 7379 2931 7382
rect 4061 7379 4127 7382
rect 5533 7379 5599 7382
rect 9581 7442 9647 7445
rect 17401 7442 17467 7445
rect 9581 7440 17467 7442
rect 9581 7384 9586 7440
rect 9642 7384 17406 7440
rect 17462 7384 17467 7440
rect 9581 7382 17467 7384
rect 9581 7379 9647 7382
rect 17401 7379 17467 7382
rect 9806 7244 9812 7308
rect 9876 7306 9882 7308
rect 11789 7306 11855 7309
rect 14181 7306 14247 7309
rect 15285 7306 15351 7309
rect 17677 7306 17743 7309
rect 9876 7246 11714 7306
rect 9876 7244 9882 7246
rect 11654 7170 11714 7246
rect 11789 7304 15351 7306
rect 11789 7248 11794 7304
rect 11850 7248 14186 7304
rect 14242 7248 15290 7304
rect 15346 7248 15351 7304
rect 11789 7246 15351 7248
rect 11789 7243 11855 7246
rect 14181 7243 14247 7246
rect 15285 7243 15351 7246
rect 16208 7304 17743 7306
rect 16208 7248 17682 7304
rect 17738 7248 17743 7304
rect 16208 7246 17743 7248
rect 16208 7170 16268 7246
rect 17677 7243 17743 7246
rect 11654 7110 16268 7170
rect 4354 7104 4750 7105
rect 4354 7040 4360 7104
rect 4424 7040 4440 7104
rect 4504 7040 4520 7104
rect 4584 7040 4600 7104
rect 4664 7040 4680 7104
rect 4744 7040 4750 7104
rect 4354 7039 4750 7040
rect 10354 7104 10750 7105
rect 10354 7040 10360 7104
rect 10424 7040 10440 7104
rect 10504 7040 10520 7104
rect 10584 7040 10600 7104
rect 10664 7040 10680 7104
rect 10744 7040 10750 7104
rect 10354 7039 10750 7040
rect 16354 7104 16750 7105
rect 16354 7040 16360 7104
rect 16424 7040 16440 7104
rect 16504 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16750 7104
rect 16354 7039 16750 7040
rect 22354 7104 22750 7105
rect 22354 7040 22360 7104
rect 22424 7040 22440 7104
rect 22504 7040 22520 7104
rect 22584 7040 22600 7104
rect 22664 7040 22680 7104
rect 22744 7040 22750 7104
rect 22354 7039 22750 7040
rect 11513 7034 11579 7037
rect 11881 7034 11947 7037
rect 11513 7032 11947 7034
rect 11513 6976 11518 7032
rect 11574 6976 11886 7032
rect 11942 6976 11947 7032
rect 11513 6974 11947 6976
rect 11513 6971 11579 6974
rect 11881 6971 11947 6974
rect 12157 7034 12223 7037
rect 16205 7034 16271 7037
rect 12157 7032 16271 7034
rect 12157 6976 12162 7032
rect 12218 6976 16210 7032
rect 16266 6976 16271 7032
rect 12157 6974 16271 6976
rect 12157 6971 12223 6974
rect 16205 6971 16271 6974
rect 11513 6898 11579 6901
rect 12525 6898 12591 6901
rect 11513 6896 12591 6898
rect 11513 6840 11518 6896
rect 11574 6840 12530 6896
rect 12586 6840 12591 6896
rect 11513 6838 12591 6840
rect 11513 6835 11579 6838
rect 12525 6835 12591 6838
rect 15694 6836 15700 6900
rect 15764 6898 15770 6900
rect 17309 6898 17375 6901
rect 15764 6896 17375 6898
rect 15764 6840 17314 6896
rect 17370 6840 17375 6896
rect 15764 6838 17375 6840
rect 15764 6836 15770 6838
rect 17309 6835 17375 6838
rect 9673 6762 9739 6765
rect 13629 6762 13695 6765
rect 9673 6760 13695 6762
rect 9673 6704 9678 6760
rect 9734 6704 13634 6760
rect 13690 6704 13695 6760
rect 9673 6702 13695 6704
rect 9673 6699 9739 6702
rect 13629 6699 13695 6702
rect 10501 6626 10567 6629
rect 12157 6626 12223 6629
rect 10501 6624 12223 6626
rect 10501 6568 10506 6624
rect 10562 6568 12162 6624
rect 12218 6568 12223 6624
rect 10501 6566 12223 6568
rect 10501 6563 10567 6566
rect 12157 6563 12223 6566
rect 1354 6560 1750 6561
rect 1354 6496 1360 6560
rect 1424 6496 1440 6560
rect 1504 6496 1520 6560
rect 1584 6496 1600 6560
rect 1664 6496 1680 6560
rect 1744 6496 1750 6560
rect 1354 6495 1750 6496
rect 7354 6560 7750 6561
rect 7354 6496 7360 6560
rect 7424 6496 7440 6560
rect 7504 6496 7520 6560
rect 7584 6496 7600 6560
rect 7664 6496 7680 6560
rect 7744 6496 7750 6560
rect 7354 6495 7750 6496
rect 13354 6560 13750 6561
rect 13354 6496 13360 6560
rect 13424 6496 13440 6560
rect 13504 6496 13520 6560
rect 13584 6496 13600 6560
rect 13664 6496 13680 6560
rect 13744 6496 13750 6560
rect 13354 6495 13750 6496
rect 19354 6560 19750 6561
rect 19354 6496 19360 6560
rect 19424 6496 19440 6560
rect 19504 6496 19520 6560
rect 19584 6496 19600 6560
rect 19664 6496 19680 6560
rect 19744 6496 19750 6560
rect 19354 6495 19750 6496
rect 13905 6490 13971 6493
rect 15929 6490 15995 6493
rect 13905 6488 15995 6490
rect 13905 6432 13910 6488
rect 13966 6432 15934 6488
rect 15990 6432 15995 6488
rect 13905 6430 15995 6432
rect 13905 6427 13971 6430
rect 15929 6427 15995 6430
rect 10869 6354 10935 6357
rect 14089 6354 14155 6357
rect 10869 6352 14155 6354
rect 10869 6296 10874 6352
rect 10930 6296 14094 6352
rect 14150 6296 14155 6352
rect 10869 6294 14155 6296
rect 10869 6291 10935 6294
rect 14089 6291 14155 6294
rect 9581 6218 9647 6221
rect 19977 6218 20043 6221
rect 9581 6216 20043 6218
rect 9581 6160 9586 6216
rect 9642 6160 19982 6216
rect 20038 6160 20043 6216
rect 9581 6158 20043 6160
rect 9581 6155 9647 6158
rect 19977 6155 20043 6158
rect 10869 6082 10935 6085
rect 14733 6082 14799 6085
rect 10869 6080 14799 6082
rect 10869 6024 10874 6080
rect 10930 6024 14738 6080
rect 14794 6024 14799 6080
rect 10869 6022 14799 6024
rect 10869 6019 10935 6022
rect 14733 6019 14799 6022
rect 4354 6016 4750 6017
rect 4354 5952 4360 6016
rect 4424 5952 4440 6016
rect 4504 5952 4520 6016
rect 4584 5952 4600 6016
rect 4664 5952 4680 6016
rect 4744 5952 4750 6016
rect 4354 5951 4750 5952
rect 10354 6016 10750 6017
rect 10354 5952 10360 6016
rect 10424 5952 10440 6016
rect 10504 5952 10520 6016
rect 10584 5952 10600 6016
rect 10664 5952 10680 6016
rect 10744 5952 10750 6016
rect 10354 5951 10750 5952
rect 16354 6016 16750 6017
rect 16354 5952 16360 6016
rect 16424 5952 16440 6016
rect 16504 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16750 6016
rect 16354 5951 16750 5952
rect 22354 6016 22750 6017
rect 22354 5952 22360 6016
rect 22424 5952 22440 6016
rect 22504 5952 22520 6016
rect 22584 5952 22600 6016
rect 22664 5952 22680 6016
rect 22744 5952 22750 6016
rect 22354 5951 22750 5952
rect 11329 5946 11395 5949
rect 11973 5946 12039 5949
rect 11329 5944 12039 5946
rect 11329 5888 11334 5944
rect 11390 5888 11978 5944
rect 12034 5888 12039 5944
rect 11329 5886 12039 5888
rect 11329 5883 11395 5886
rect 11973 5883 12039 5886
rect 14733 5812 14799 5813
rect 14733 5810 14780 5812
rect 14688 5808 14780 5810
rect 14688 5752 14738 5808
rect 14688 5750 14780 5752
rect 14733 5748 14780 5750
rect 14844 5748 14850 5812
rect 14733 5747 14799 5748
rect 8201 5674 8267 5677
rect 12801 5674 12867 5677
rect 13261 5674 13327 5677
rect 8201 5672 13327 5674
rect 8201 5616 8206 5672
rect 8262 5616 12806 5672
rect 12862 5616 13266 5672
rect 13322 5616 13327 5672
rect 8201 5614 13327 5616
rect 8201 5611 8267 5614
rect 12801 5611 12867 5614
rect 13261 5611 13327 5614
rect 20662 5612 20668 5676
rect 20732 5674 20738 5676
rect 21357 5674 21423 5677
rect 20732 5672 21423 5674
rect 20732 5616 21362 5672
rect 21418 5616 21423 5672
rect 20732 5614 21423 5616
rect 20732 5612 20738 5614
rect 21357 5611 21423 5614
rect 15142 5476 15148 5540
rect 15212 5538 15218 5540
rect 15929 5538 15995 5541
rect 15212 5536 15995 5538
rect 15212 5480 15934 5536
rect 15990 5480 15995 5536
rect 15212 5478 15995 5480
rect 15212 5476 15218 5478
rect 15929 5475 15995 5478
rect 16062 5476 16068 5540
rect 16132 5538 16138 5540
rect 16941 5538 17007 5541
rect 16132 5536 17007 5538
rect 16132 5480 16946 5536
rect 17002 5480 17007 5536
rect 16132 5478 17007 5480
rect 16132 5476 16138 5478
rect 16941 5475 17007 5478
rect 1354 5472 1750 5473
rect 1354 5408 1360 5472
rect 1424 5408 1440 5472
rect 1504 5408 1520 5472
rect 1584 5408 1600 5472
rect 1664 5408 1680 5472
rect 1744 5408 1750 5472
rect 1354 5407 1750 5408
rect 7354 5472 7750 5473
rect 7354 5408 7360 5472
rect 7424 5408 7440 5472
rect 7504 5408 7520 5472
rect 7584 5408 7600 5472
rect 7664 5408 7680 5472
rect 7744 5408 7750 5472
rect 7354 5407 7750 5408
rect 13354 5472 13750 5473
rect 13354 5408 13360 5472
rect 13424 5408 13440 5472
rect 13504 5408 13520 5472
rect 13584 5408 13600 5472
rect 13664 5408 13680 5472
rect 13744 5408 13750 5472
rect 13354 5407 13750 5408
rect 19354 5472 19750 5473
rect 19354 5408 19360 5472
rect 19424 5408 19440 5472
rect 19504 5408 19520 5472
rect 19584 5408 19600 5472
rect 19664 5408 19680 5472
rect 19744 5408 19750 5472
rect 19354 5407 19750 5408
rect 10041 5404 10107 5405
rect 9990 5340 9996 5404
rect 10060 5402 10107 5404
rect 10060 5400 10152 5402
rect 10102 5344 10152 5400
rect 10060 5342 10152 5344
rect 10060 5340 10107 5342
rect 10041 5339 10107 5340
rect 7281 5266 7347 5269
rect 15469 5266 15535 5269
rect 7281 5264 15535 5266
rect 7281 5208 7286 5264
rect 7342 5208 15474 5264
rect 15530 5208 15535 5264
rect 7281 5206 15535 5208
rect 7281 5203 7347 5206
rect 15469 5203 15535 5206
rect 9806 5068 9812 5132
rect 9876 5130 9882 5132
rect 11053 5130 11119 5133
rect 9876 5128 11119 5130
rect 9876 5072 11058 5128
rect 11114 5072 11119 5128
rect 9876 5070 11119 5072
rect 9876 5068 9882 5070
rect 11053 5067 11119 5070
rect 13169 5130 13235 5133
rect 16941 5130 17007 5133
rect 13169 5128 17007 5130
rect 13169 5072 13174 5128
rect 13230 5072 16946 5128
rect 17002 5072 17007 5128
rect 13169 5070 17007 5072
rect 13169 5067 13235 5070
rect 16941 5067 17007 5070
rect 11329 4994 11395 4997
rect 13629 4994 13695 4997
rect 11329 4992 13695 4994
rect 11329 4936 11334 4992
rect 11390 4936 13634 4992
rect 13690 4936 13695 4992
rect 11329 4934 13695 4936
rect 11329 4931 11395 4934
rect 13629 4931 13695 4934
rect 4354 4928 4750 4929
rect 4354 4864 4360 4928
rect 4424 4864 4440 4928
rect 4504 4864 4520 4928
rect 4584 4864 4600 4928
rect 4664 4864 4680 4928
rect 4744 4864 4750 4928
rect 4354 4863 4750 4864
rect 10354 4928 10750 4929
rect 10354 4864 10360 4928
rect 10424 4864 10440 4928
rect 10504 4864 10520 4928
rect 10584 4864 10600 4928
rect 10664 4864 10680 4928
rect 10744 4864 10750 4928
rect 10354 4863 10750 4864
rect 16354 4928 16750 4929
rect 16354 4864 16360 4928
rect 16424 4864 16440 4928
rect 16504 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16750 4928
rect 16354 4863 16750 4864
rect 22354 4928 22750 4929
rect 22354 4864 22360 4928
rect 22424 4864 22440 4928
rect 22504 4864 22520 4928
rect 22584 4864 22600 4928
rect 22664 4864 22680 4928
rect 22744 4864 22750 4928
rect 22354 4863 22750 4864
rect 12985 4858 13051 4861
rect 12390 4856 13051 4858
rect 12390 4800 12990 4856
rect 13046 4800 13051 4856
rect 12390 4798 13051 4800
rect 8201 4722 8267 4725
rect 12390 4722 12450 4798
rect 12985 4795 13051 4798
rect 17033 4722 17099 4725
rect 8201 4720 12450 4722
rect 8201 4664 8206 4720
rect 8262 4664 12450 4720
rect 8201 4662 12450 4664
rect 15334 4720 17099 4722
rect 15334 4664 17038 4720
rect 17094 4664 17099 4720
rect 15334 4662 17099 4664
rect 8201 4659 8267 4662
rect 6085 4586 6151 4589
rect 7741 4586 7807 4589
rect 6085 4584 7807 4586
rect 6085 4528 6090 4584
rect 6146 4528 7746 4584
rect 7802 4528 7807 4584
rect 6085 4526 7807 4528
rect 6085 4523 6151 4526
rect 7741 4523 7807 4526
rect 10501 4586 10567 4589
rect 15334 4586 15394 4662
rect 17033 4659 17099 4662
rect 10501 4584 15394 4586
rect 10501 4528 10506 4584
rect 10562 4528 15394 4584
rect 10501 4526 15394 4528
rect 15469 4586 15535 4589
rect 16021 4586 16087 4589
rect 15469 4584 16087 4586
rect 15469 4528 15474 4584
rect 15530 4528 16026 4584
rect 16082 4528 16087 4584
rect 15469 4526 16087 4528
rect 10501 4523 10567 4526
rect 15469 4523 15535 4526
rect 16021 4523 16087 4526
rect 19609 4586 19675 4589
rect 21449 4586 21515 4589
rect 19609 4584 21515 4586
rect 19609 4528 19614 4584
rect 19670 4528 21454 4584
rect 21510 4528 21515 4584
rect 19609 4526 21515 4528
rect 19609 4523 19675 4526
rect 21449 4523 21515 4526
rect 1354 4384 1750 4385
rect 1354 4320 1360 4384
rect 1424 4320 1440 4384
rect 1504 4320 1520 4384
rect 1584 4320 1600 4384
rect 1664 4320 1680 4384
rect 1744 4320 1750 4384
rect 1354 4319 1750 4320
rect 7354 4384 7750 4385
rect 7354 4320 7360 4384
rect 7424 4320 7440 4384
rect 7504 4320 7520 4384
rect 7584 4320 7600 4384
rect 7664 4320 7680 4384
rect 7744 4320 7750 4384
rect 7354 4319 7750 4320
rect 13354 4384 13750 4385
rect 13354 4320 13360 4384
rect 13424 4320 13440 4384
rect 13504 4320 13520 4384
rect 13584 4320 13600 4384
rect 13664 4320 13680 4384
rect 13744 4320 13750 4384
rect 13354 4319 13750 4320
rect 19354 4384 19750 4385
rect 19354 4320 19360 4384
rect 19424 4320 19440 4384
rect 19504 4320 19520 4384
rect 19584 4320 19600 4384
rect 19664 4320 19680 4384
rect 19744 4320 19750 4384
rect 19354 4319 19750 4320
rect 13445 4178 13511 4181
rect 18505 4178 18571 4181
rect 13445 4176 18571 4178
rect 13445 4120 13450 4176
rect 13506 4120 18510 4176
rect 18566 4120 18571 4176
rect 13445 4118 18571 4120
rect 13445 4115 13511 4118
rect 18505 4115 18571 4118
rect 12801 4042 12867 4045
rect 18505 4042 18571 4045
rect 12801 4040 18571 4042
rect 12801 3984 12806 4040
rect 12862 3984 18510 4040
rect 18566 3984 18571 4040
rect 12801 3982 18571 3984
rect 12801 3979 12867 3982
rect 18505 3979 18571 3982
rect 9438 3844 9444 3908
rect 9508 3906 9514 3908
rect 9581 3906 9647 3909
rect 9508 3904 9647 3906
rect 9508 3848 9586 3904
rect 9642 3848 9647 3904
rect 9508 3846 9647 3848
rect 9508 3844 9514 3846
rect 9581 3843 9647 3846
rect 4354 3840 4750 3841
rect 4354 3776 4360 3840
rect 4424 3776 4440 3840
rect 4504 3776 4520 3840
rect 4584 3776 4600 3840
rect 4664 3776 4680 3840
rect 4744 3776 4750 3840
rect 4354 3775 4750 3776
rect 10354 3840 10750 3841
rect 10354 3776 10360 3840
rect 10424 3776 10440 3840
rect 10504 3776 10520 3840
rect 10584 3776 10600 3840
rect 10664 3776 10680 3840
rect 10744 3776 10750 3840
rect 10354 3775 10750 3776
rect 16354 3840 16750 3841
rect 16354 3776 16360 3840
rect 16424 3776 16440 3840
rect 16504 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16750 3840
rect 16354 3775 16750 3776
rect 22354 3840 22750 3841
rect 22354 3776 22360 3840
rect 22424 3776 22440 3840
rect 22504 3776 22520 3840
rect 22584 3776 22600 3840
rect 22664 3776 22680 3840
rect 22744 3776 22750 3840
rect 22354 3775 22750 3776
rect 8017 3770 8083 3773
rect 9121 3770 9187 3773
rect 8017 3768 9187 3770
rect 8017 3712 8022 3768
rect 8078 3712 9126 3768
rect 9182 3712 9187 3768
rect 8017 3710 9187 3712
rect 8017 3707 8083 3710
rect 9121 3707 9187 3710
rect 9806 3708 9812 3772
rect 9876 3770 9882 3772
rect 10041 3770 10107 3773
rect 9876 3768 10107 3770
rect 9876 3712 10046 3768
rect 10102 3712 10107 3768
rect 9876 3710 10107 3712
rect 9876 3708 9882 3710
rect 10041 3707 10107 3710
rect 6637 3634 6703 3637
rect 18873 3634 18939 3637
rect 6637 3632 18939 3634
rect 6637 3576 6642 3632
rect 6698 3576 18878 3632
rect 18934 3576 18939 3632
rect 6637 3574 18939 3576
rect 6637 3571 6703 3574
rect 18873 3571 18939 3574
rect 19977 3634 20043 3637
rect 21541 3634 21607 3637
rect 19977 3632 21607 3634
rect 19977 3576 19982 3632
rect 20038 3576 21546 3632
rect 21602 3576 21607 3632
rect 19977 3574 21607 3576
rect 19977 3571 20043 3574
rect 21541 3571 21607 3574
rect 7005 3498 7071 3501
rect 16573 3498 16639 3501
rect 7005 3496 16639 3498
rect 7005 3440 7010 3496
rect 7066 3440 16578 3496
rect 16634 3440 16639 3496
rect 7005 3438 16639 3440
rect 7005 3435 7071 3438
rect 16573 3435 16639 3438
rect 17953 3498 18019 3501
rect 18597 3498 18663 3501
rect 17953 3496 18663 3498
rect 17953 3440 17958 3496
rect 18014 3440 18602 3496
rect 18658 3440 18663 3496
rect 17953 3438 18663 3440
rect 17953 3435 18019 3438
rect 18597 3435 18663 3438
rect 9070 3300 9076 3364
rect 9140 3362 9146 3364
rect 9581 3362 9647 3365
rect 11053 3364 11119 3365
rect 11053 3362 11100 3364
rect 9140 3360 9647 3362
rect 9140 3304 9586 3360
rect 9642 3304 9647 3360
rect 9140 3302 9647 3304
rect 11008 3360 11100 3362
rect 11008 3304 11058 3360
rect 11008 3302 11100 3304
rect 9140 3300 9146 3302
rect 9581 3299 9647 3302
rect 11053 3300 11100 3302
rect 11164 3300 11170 3364
rect 15561 3362 15627 3365
rect 16389 3362 16455 3365
rect 15561 3360 16455 3362
rect 15561 3304 15566 3360
rect 15622 3304 16394 3360
rect 16450 3304 16455 3360
rect 15561 3302 16455 3304
rect 11053 3299 11119 3300
rect 15561 3299 15627 3302
rect 16389 3299 16455 3302
rect 1354 3296 1750 3297
rect 1354 3232 1360 3296
rect 1424 3232 1440 3296
rect 1504 3232 1520 3296
rect 1584 3232 1600 3296
rect 1664 3232 1680 3296
rect 1744 3232 1750 3296
rect 1354 3231 1750 3232
rect 7354 3296 7750 3297
rect 7354 3232 7360 3296
rect 7424 3232 7440 3296
rect 7504 3232 7520 3296
rect 7584 3232 7600 3296
rect 7664 3232 7680 3296
rect 7744 3232 7750 3296
rect 7354 3231 7750 3232
rect 13354 3296 13750 3297
rect 13354 3232 13360 3296
rect 13424 3232 13440 3296
rect 13504 3232 13520 3296
rect 13584 3232 13600 3296
rect 13664 3232 13680 3296
rect 13744 3232 13750 3296
rect 13354 3231 13750 3232
rect 19354 3296 19750 3297
rect 19354 3232 19360 3296
rect 19424 3232 19440 3296
rect 19504 3232 19520 3296
rect 19584 3232 19600 3296
rect 19664 3232 19680 3296
rect 19744 3232 19750 3296
rect 19354 3231 19750 3232
rect 9489 3224 9555 3229
rect 9489 3168 9494 3224
rect 9550 3168 9555 3224
rect 9489 3163 9555 3168
rect 9949 3226 10015 3229
rect 10409 3226 10475 3229
rect 9949 3224 10475 3226
rect 9949 3168 9954 3224
rect 10010 3168 10414 3224
rect 10470 3168 10475 3224
rect 9949 3166 10475 3168
rect 9949 3163 10015 3166
rect 10409 3163 10475 3166
rect 9254 3028 9260 3092
rect 9324 3090 9330 3092
rect 9492 3090 9552 3163
rect 9324 3030 9552 3090
rect 9673 3090 9739 3093
rect 11789 3090 11855 3093
rect 9673 3088 11855 3090
rect 9673 3032 9678 3088
rect 9734 3032 11794 3088
rect 11850 3032 11855 3088
rect 9673 3030 11855 3032
rect 9324 3028 9330 3030
rect 9673 3027 9739 3030
rect 11789 3027 11855 3030
rect 14641 3090 14707 3093
rect 15745 3090 15811 3093
rect 16205 3090 16271 3093
rect 14641 3088 16271 3090
rect 14641 3032 14646 3088
rect 14702 3032 15750 3088
rect 15806 3032 16210 3088
rect 16266 3032 16271 3088
rect 14641 3030 16271 3032
rect 14641 3027 14707 3030
rect 15745 3027 15811 3030
rect 16205 3027 16271 3030
rect 1577 2954 1643 2957
rect 7833 2954 7899 2957
rect 12341 2954 12407 2957
rect 14825 2954 14891 2957
rect 19701 2954 19767 2957
rect 1577 2952 7666 2954
rect 1577 2896 1582 2952
rect 1638 2896 7666 2952
rect 1577 2894 7666 2896
rect 1577 2891 1643 2894
rect 7606 2818 7666 2894
rect 7833 2952 9552 2954
rect 7833 2896 7838 2952
rect 7894 2920 9552 2952
rect 9630 2920 10978 2954
rect 7894 2896 10978 2920
rect 7833 2894 10978 2896
rect 7833 2891 7899 2894
rect 9492 2860 9690 2894
rect 9305 2818 9371 2821
rect 7606 2816 9371 2818
rect 7606 2760 9310 2816
rect 9366 2760 9371 2816
rect 7606 2758 9371 2760
rect 9305 2755 9371 2758
rect 9765 2820 9831 2821
rect 9765 2816 9812 2820
rect 9876 2818 9882 2820
rect 10918 2818 10978 2894
rect 12341 2952 14891 2954
rect 12341 2896 12346 2952
rect 12402 2896 14830 2952
rect 14886 2896 14891 2952
rect 12341 2894 14891 2896
rect 12341 2891 12407 2894
rect 14825 2891 14891 2894
rect 16070 2952 19767 2954
rect 16070 2896 19706 2952
rect 19762 2896 19767 2952
rect 16070 2894 19767 2896
rect 16070 2818 16130 2894
rect 19701 2891 19767 2894
rect 9765 2760 9770 2816
rect 9765 2756 9812 2760
rect 9876 2758 9922 2818
rect 10918 2758 16130 2818
rect 9876 2756 9882 2758
rect 9765 2755 9831 2756
rect 4354 2752 4750 2753
rect 4354 2688 4360 2752
rect 4424 2688 4440 2752
rect 4504 2688 4520 2752
rect 4584 2688 4600 2752
rect 4664 2688 4680 2752
rect 4744 2688 4750 2752
rect 4354 2687 4750 2688
rect 10354 2752 10750 2753
rect 10354 2688 10360 2752
rect 10424 2688 10440 2752
rect 10504 2688 10520 2752
rect 10584 2688 10600 2752
rect 10664 2688 10680 2752
rect 10744 2688 10750 2752
rect 10354 2687 10750 2688
rect 16354 2752 16750 2753
rect 16354 2688 16360 2752
rect 16424 2688 16440 2752
rect 16504 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16750 2752
rect 16354 2687 16750 2688
rect 22354 2752 22750 2753
rect 22354 2688 22360 2752
rect 22424 2688 22440 2752
rect 22504 2688 22520 2752
rect 22584 2688 22600 2752
rect 22664 2688 22680 2752
rect 22744 2688 22750 2752
rect 22354 2687 22750 2688
rect 9070 2620 9076 2684
rect 9140 2682 9146 2684
rect 9489 2682 9555 2685
rect 9140 2680 9555 2682
rect 9140 2624 9494 2680
rect 9550 2624 9555 2680
rect 9140 2622 9555 2624
rect 9140 2620 9146 2622
rect 9489 2619 9555 2622
rect 9765 2682 9831 2685
rect 10041 2682 10107 2685
rect 9765 2680 10107 2682
rect 9765 2624 9770 2680
rect 9826 2624 10046 2680
rect 10102 2624 10107 2680
rect 9765 2622 10107 2624
rect 9765 2619 9831 2622
rect 10041 2619 10107 2622
rect 12985 2682 13051 2685
rect 13118 2682 13124 2684
rect 12985 2680 13124 2682
rect 12985 2624 12990 2680
rect 13046 2624 13124 2680
rect 12985 2622 13124 2624
rect 12985 2619 13051 2622
rect 13118 2620 13124 2622
rect 13188 2682 13194 2684
rect 13537 2682 13603 2685
rect 13188 2680 13603 2682
rect 13188 2624 13542 2680
rect 13598 2624 13603 2680
rect 13188 2622 13603 2624
rect 13188 2620 13194 2622
rect 13537 2619 13603 2622
rect 18229 2682 18295 2685
rect 20662 2682 20668 2684
rect 18229 2680 20668 2682
rect 18229 2624 18234 2680
rect 18290 2624 20668 2680
rect 18229 2622 20668 2624
rect 18229 2619 18295 2622
rect 20662 2620 20668 2622
rect 20732 2620 20738 2684
rect 4061 2546 4127 2549
rect 21449 2546 21515 2549
rect 4061 2544 21515 2546
rect 4061 2488 4066 2544
rect 4122 2488 21454 2544
rect 21510 2488 21515 2544
rect 4061 2486 21515 2488
rect 4061 2483 4127 2486
rect 21449 2483 21515 2486
rect 9254 2348 9260 2412
rect 9324 2410 9330 2412
rect 9397 2410 9463 2413
rect 9324 2408 9463 2410
rect 9324 2352 9402 2408
rect 9458 2352 9463 2408
rect 9324 2350 9463 2352
rect 9324 2348 9330 2350
rect 9397 2347 9463 2350
rect 11329 2410 11395 2413
rect 18873 2410 18939 2413
rect 11329 2408 18939 2410
rect 11329 2352 11334 2408
rect 11390 2352 18878 2408
rect 18934 2352 18939 2408
rect 11329 2350 18939 2352
rect 11329 2347 11395 2350
rect 18873 2347 18939 2350
rect 8753 2274 8819 2277
rect 11697 2274 11763 2277
rect 8753 2272 11763 2274
rect 8753 2216 8758 2272
rect 8814 2216 11702 2272
rect 11758 2216 11763 2272
rect 8753 2214 11763 2216
rect 8753 2211 8819 2214
rect 11697 2211 11763 2214
rect 15929 2274 15995 2277
rect 17493 2274 17559 2277
rect 15929 2272 17559 2274
rect 15929 2216 15934 2272
rect 15990 2216 17498 2272
rect 17554 2216 17559 2272
rect 15929 2214 17559 2216
rect 15929 2211 15995 2214
rect 17493 2211 17559 2214
rect 1354 2208 1750 2209
rect 1354 2144 1360 2208
rect 1424 2144 1440 2208
rect 1504 2144 1520 2208
rect 1584 2144 1600 2208
rect 1664 2144 1680 2208
rect 1744 2144 1750 2208
rect 1354 2143 1750 2144
rect 7354 2208 7750 2209
rect 7354 2144 7360 2208
rect 7424 2144 7440 2208
rect 7504 2144 7520 2208
rect 7584 2144 7600 2208
rect 7664 2144 7680 2208
rect 7744 2144 7750 2208
rect 7354 2143 7750 2144
rect 13354 2208 13750 2209
rect 13354 2144 13360 2208
rect 13424 2144 13440 2208
rect 13504 2144 13520 2208
rect 13584 2144 13600 2208
rect 13664 2144 13680 2208
rect 13744 2144 13750 2208
rect 13354 2143 13750 2144
rect 19354 2208 19750 2209
rect 19354 2144 19360 2208
rect 19424 2144 19440 2208
rect 19504 2144 19520 2208
rect 19584 2144 19600 2208
rect 19664 2144 19680 2208
rect 19744 2144 19750 2208
rect 19354 2143 19750 2144
rect 8569 2138 8635 2141
rect 11789 2138 11855 2141
rect 8569 2136 11855 2138
rect 8569 2080 8574 2136
rect 8630 2080 11794 2136
rect 11850 2080 11855 2136
rect 8569 2078 11855 2080
rect 8569 2075 8635 2078
rect 11789 2075 11855 2078
rect 14917 2140 14983 2141
rect 14917 2136 14964 2140
rect 15028 2138 15034 2140
rect 15653 2138 15719 2141
rect 16113 2138 16179 2141
rect 14917 2080 14922 2136
rect 14917 2076 14964 2080
rect 15028 2078 15074 2138
rect 15653 2136 16179 2138
rect 15653 2080 15658 2136
rect 15714 2080 16118 2136
rect 16174 2080 16179 2136
rect 15653 2078 16179 2080
rect 15028 2076 15034 2078
rect 14917 2075 14983 2076
rect 15653 2075 15719 2078
rect 16113 2075 16179 2078
rect 7557 2002 7623 2005
rect 9121 2002 9187 2005
rect 7557 2000 9187 2002
rect 7557 1944 7562 2000
rect 7618 1944 9126 2000
rect 9182 1944 9187 2000
rect 7557 1942 9187 1944
rect 7557 1939 7623 1942
rect 9121 1939 9187 1942
rect 10869 2002 10935 2005
rect 17125 2002 17191 2005
rect 10869 2000 17191 2002
rect 10869 1944 10874 2000
rect 10930 1944 17130 2000
rect 17186 1944 17191 2000
rect 10869 1942 17191 1944
rect 10869 1939 10935 1942
rect 17125 1939 17191 1942
rect 4337 1866 4403 1869
rect 18413 1866 18479 1869
rect 4337 1864 18479 1866
rect 4337 1808 4342 1864
rect 4398 1808 18418 1864
rect 18474 1808 18479 1864
rect 4337 1806 18479 1808
rect 4337 1803 4403 1806
rect 18413 1803 18479 1806
rect 9489 1732 9555 1733
rect 9438 1668 9444 1732
rect 9508 1730 9555 1732
rect 9508 1728 9600 1730
rect 9550 1672 9600 1728
rect 9508 1670 9600 1672
rect 9508 1668 9555 1670
rect 9489 1667 9555 1668
rect 4354 1664 4750 1665
rect 4354 1600 4360 1664
rect 4424 1600 4440 1664
rect 4504 1600 4520 1664
rect 4584 1600 4600 1664
rect 4664 1600 4680 1664
rect 4744 1600 4750 1664
rect 4354 1599 4750 1600
rect 10354 1664 10750 1665
rect 10354 1600 10360 1664
rect 10424 1600 10440 1664
rect 10504 1600 10520 1664
rect 10584 1600 10600 1664
rect 10664 1600 10680 1664
rect 10744 1600 10750 1664
rect 10354 1599 10750 1600
rect 16354 1664 16750 1665
rect 16354 1600 16360 1664
rect 16424 1600 16440 1664
rect 16504 1600 16520 1664
rect 16584 1600 16600 1664
rect 16664 1600 16680 1664
rect 16744 1600 16750 1664
rect 16354 1599 16750 1600
rect 22354 1664 22750 1665
rect 22354 1600 22360 1664
rect 22424 1600 22440 1664
rect 22504 1600 22520 1664
rect 22584 1600 22600 1664
rect 22664 1600 22680 1664
rect 22744 1600 22750 1664
rect 22354 1599 22750 1600
rect 13353 1594 13419 1597
rect 15653 1594 15719 1597
rect 13353 1592 15719 1594
rect 13353 1536 13358 1592
rect 13414 1536 15658 1592
rect 15714 1536 15719 1592
rect 13353 1534 15719 1536
rect 13353 1531 13419 1534
rect 15653 1531 15719 1534
rect 8569 1458 8635 1461
rect 11513 1458 11579 1461
rect 16062 1458 16068 1460
rect 8569 1456 16068 1458
rect 8569 1400 8574 1456
rect 8630 1400 11518 1456
rect 11574 1400 16068 1456
rect 8569 1398 16068 1400
rect 8569 1395 8635 1398
rect 11513 1395 11579 1398
rect 16062 1396 16068 1398
rect 16132 1458 16138 1460
rect 16389 1458 16455 1461
rect 16132 1456 16455 1458
rect 16132 1400 16394 1456
rect 16450 1400 16455 1456
rect 16132 1398 16455 1400
rect 16132 1396 16138 1398
rect 16389 1395 16455 1398
rect 1354 1120 1750 1121
rect 1354 1056 1360 1120
rect 1424 1056 1440 1120
rect 1504 1056 1520 1120
rect 1584 1056 1600 1120
rect 1664 1056 1680 1120
rect 1744 1056 1750 1120
rect 1354 1055 1750 1056
rect 7354 1120 7750 1121
rect 7354 1056 7360 1120
rect 7424 1056 7440 1120
rect 7504 1056 7520 1120
rect 7584 1056 7600 1120
rect 7664 1056 7680 1120
rect 7744 1056 7750 1120
rect 7354 1055 7750 1056
rect 13354 1120 13750 1121
rect 13354 1056 13360 1120
rect 13424 1056 13440 1120
rect 13504 1056 13520 1120
rect 13584 1056 13600 1120
rect 13664 1056 13680 1120
rect 13744 1056 13750 1120
rect 13354 1055 13750 1056
rect 19354 1120 19750 1121
rect 19354 1056 19360 1120
rect 19424 1056 19440 1120
rect 19504 1056 19520 1120
rect 19584 1056 19600 1120
rect 19664 1056 19680 1120
rect 19744 1056 19750 1120
rect 19354 1055 19750 1056
rect 9765 914 9831 917
rect 9990 914 9996 916
rect 9765 912 9996 914
rect 9765 856 9770 912
rect 9826 856 9996 912
rect 9765 854 9996 856
rect 9765 851 9831 854
rect 9990 852 9996 854
rect 10060 852 10066 916
rect 4354 576 4750 577
rect 4354 512 4360 576
rect 4424 512 4440 576
rect 4504 512 4520 576
rect 4584 512 4600 576
rect 4664 512 4680 576
rect 4744 512 4750 576
rect 4354 511 4750 512
rect 10354 576 10750 577
rect 10354 512 10360 576
rect 10424 512 10440 576
rect 10504 512 10520 576
rect 10584 512 10600 576
rect 10664 512 10680 576
rect 10744 512 10750 576
rect 10354 511 10750 512
rect 16354 576 16750 577
rect 16354 512 16360 576
rect 16424 512 16440 576
rect 16504 512 16520 576
rect 16584 512 16600 576
rect 16664 512 16680 576
rect 16744 512 16750 576
rect 16354 511 16750 512
rect 22354 576 22750 577
rect 22354 512 22360 576
rect 22424 512 22440 576
rect 22504 512 22520 576
rect 22584 512 22600 576
rect 22664 512 22680 576
rect 22744 512 22750 576
rect 22354 511 22750 512
<< via3 >>
rect 1360 15260 1424 15264
rect 1360 15204 1364 15260
rect 1364 15204 1420 15260
rect 1420 15204 1424 15260
rect 1360 15200 1424 15204
rect 1440 15260 1504 15264
rect 1440 15204 1444 15260
rect 1444 15204 1500 15260
rect 1500 15204 1504 15260
rect 1440 15200 1504 15204
rect 1520 15260 1584 15264
rect 1520 15204 1524 15260
rect 1524 15204 1580 15260
rect 1580 15204 1584 15260
rect 1520 15200 1584 15204
rect 1600 15260 1664 15264
rect 1600 15204 1604 15260
rect 1604 15204 1660 15260
rect 1660 15204 1664 15260
rect 1600 15200 1664 15204
rect 1680 15260 1744 15264
rect 1680 15204 1684 15260
rect 1684 15204 1740 15260
rect 1740 15204 1744 15260
rect 1680 15200 1744 15204
rect 7360 15260 7424 15264
rect 7360 15204 7364 15260
rect 7364 15204 7420 15260
rect 7420 15204 7424 15260
rect 7360 15200 7424 15204
rect 7440 15260 7504 15264
rect 7440 15204 7444 15260
rect 7444 15204 7500 15260
rect 7500 15204 7504 15260
rect 7440 15200 7504 15204
rect 7520 15260 7584 15264
rect 7520 15204 7524 15260
rect 7524 15204 7580 15260
rect 7580 15204 7584 15260
rect 7520 15200 7584 15204
rect 7600 15260 7664 15264
rect 7600 15204 7604 15260
rect 7604 15204 7660 15260
rect 7660 15204 7664 15260
rect 7600 15200 7664 15204
rect 7680 15260 7744 15264
rect 7680 15204 7684 15260
rect 7684 15204 7740 15260
rect 7740 15204 7744 15260
rect 7680 15200 7744 15204
rect 13360 15260 13424 15264
rect 13360 15204 13364 15260
rect 13364 15204 13420 15260
rect 13420 15204 13424 15260
rect 13360 15200 13424 15204
rect 13440 15260 13504 15264
rect 13440 15204 13444 15260
rect 13444 15204 13500 15260
rect 13500 15204 13504 15260
rect 13440 15200 13504 15204
rect 13520 15260 13584 15264
rect 13520 15204 13524 15260
rect 13524 15204 13580 15260
rect 13580 15204 13584 15260
rect 13520 15200 13584 15204
rect 13600 15260 13664 15264
rect 13600 15204 13604 15260
rect 13604 15204 13660 15260
rect 13660 15204 13664 15260
rect 13600 15200 13664 15204
rect 13680 15260 13744 15264
rect 13680 15204 13684 15260
rect 13684 15204 13740 15260
rect 13740 15204 13744 15260
rect 13680 15200 13744 15204
rect 19360 15260 19424 15264
rect 19360 15204 19364 15260
rect 19364 15204 19420 15260
rect 19420 15204 19424 15260
rect 19360 15200 19424 15204
rect 19440 15260 19504 15264
rect 19440 15204 19444 15260
rect 19444 15204 19500 15260
rect 19500 15204 19504 15260
rect 19440 15200 19504 15204
rect 19520 15260 19584 15264
rect 19520 15204 19524 15260
rect 19524 15204 19580 15260
rect 19580 15204 19584 15260
rect 19520 15200 19584 15204
rect 19600 15260 19664 15264
rect 19600 15204 19604 15260
rect 19604 15204 19660 15260
rect 19660 15204 19664 15260
rect 19600 15200 19664 15204
rect 19680 15260 19744 15264
rect 19680 15204 19684 15260
rect 19684 15204 19740 15260
rect 19740 15204 19744 15260
rect 19680 15200 19744 15204
rect 4360 14716 4424 14720
rect 4360 14660 4364 14716
rect 4364 14660 4420 14716
rect 4420 14660 4424 14716
rect 4360 14656 4424 14660
rect 4440 14716 4504 14720
rect 4440 14660 4444 14716
rect 4444 14660 4500 14716
rect 4500 14660 4504 14716
rect 4440 14656 4504 14660
rect 4520 14716 4584 14720
rect 4520 14660 4524 14716
rect 4524 14660 4580 14716
rect 4580 14660 4584 14716
rect 4520 14656 4584 14660
rect 4600 14716 4664 14720
rect 4600 14660 4604 14716
rect 4604 14660 4660 14716
rect 4660 14660 4664 14716
rect 4600 14656 4664 14660
rect 4680 14716 4744 14720
rect 4680 14660 4684 14716
rect 4684 14660 4740 14716
rect 4740 14660 4744 14716
rect 4680 14656 4744 14660
rect 10360 14716 10424 14720
rect 10360 14660 10364 14716
rect 10364 14660 10420 14716
rect 10420 14660 10424 14716
rect 10360 14656 10424 14660
rect 10440 14716 10504 14720
rect 10440 14660 10444 14716
rect 10444 14660 10500 14716
rect 10500 14660 10504 14716
rect 10440 14656 10504 14660
rect 10520 14716 10584 14720
rect 10520 14660 10524 14716
rect 10524 14660 10580 14716
rect 10580 14660 10584 14716
rect 10520 14656 10584 14660
rect 10600 14716 10664 14720
rect 10600 14660 10604 14716
rect 10604 14660 10660 14716
rect 10660 14660 10664 14716
rect 10600 14656 10664 14660
rect 10680 14716 10744 14720
rect 10680 14660 10684 14716
rect 10684 14660 10740 14716
rect 10740 14660 10744 14716
rect 10680 14656 10744 14660
rect 16360 14716 16424 14720
rect 16360 14660 16364 14716
rect 16364 14660 16420 14716
rect 16420 14660 16424 14716
rect 16360 14656 16424 14660
rect 16440 14716 16504 14720
rect 16440 14660 16444 14716
rect 16444 14660 16500 14716
rect 16500 14660 16504 14716
rect 16440 14656 16504 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 22360 14716 22424 14720
rect 22360 14660 22364 14716
rect 22364 14660 22420 14716
rect 22420 14660 22424 14716
rect 22360 14656 22424 14660
rect 22440 14716 22504 14720
rect 22440 14660 22444 14716
rect 22444 14660 22500 14716
rect 22500 14660 22504 14716
rect 22440 14656 22504 14660
rect 22520 14716 22584 14720
rect 22520 14660 22524 14716
rect 22524 14660 22580 14716
rect 22580 14660 22584 14716
rect 22520 14656 22584 14660
rect 22600 14716 22664 14720
rect 22600 14660 22604 14716
rect 22604 14660 22660 14716
rect 22660 14660 22664 14716
rect 22600 14656 22664 14660
rect 22680 14716 22744 14720
rect 22680 14660 22684 14716
rect 22684 14660 22740 14716
rect 22740 14660 22744 14716
rect 22680 14656 22744 14660
rect 1360 14172 1424 14176
rect 1360 14116 1364 14172
rect 1364 14116 1420 14172
rect 1420 14116 1424 14172
rect 1360 14112 1424 14116
rect 1440 14172 1504 14176
rect 1440 14116 1444 14172
rect 1444 14116 1500 14172
rect 1500 14116 1504 14172
rect 1440 14112 1504 14116
rect 1520 14172 1584 14176
rect 1520 14116 1524 14172
rect 1524 14116 1580 14172
rect 1580 14116 1584 14172
rect 1520 14112 1584 14116
rect 1600 14172 1664 14176
rect 1600 14116 1604 14172
rect 1604 14116 1660 14172
rect 1660 14116 1664 14172
rect 1600 14112 1664 14116
rect 1680 14172 1744 14176
rect 1680 14116 1684 14172
rect 1684 14116 1740 14172
rect 1740 14116 1744 14172
rect 1680 14112 1744 14116
rect 7360 14172 7424 14176
rect 7360 14116 7364 14172
rect 7364 14116 7420 14172
rect 7420 14116 7424 14172
rect 7360 14112 7424 14116
rect 7440 14172 7504 14176
rect 7440 14116 7444 14172
rect 7444 14116 7500 14172
rect 7500 14116 7504 14172
rect 7440 14112 7504 14116
rect 7520 14172 7584 14176
rect 7520 14116 7524 14172
rect 7524 14116 7580 14172
rect 7580 14116 7584 14172
rect 7520 14112 7584 14116
rect 7600 14172 7664 14176
rect 7600 14116 7604 14172
rect 7604 14116 7660 14172
rect 7660 14116 7664 14172
rect 7600 14112 7664 14116
rect 7680 14172 7744 14176
rect 7680 14116 7684 14172
rect 7684 14116 7740 14172
rect 7740 14116 7744 14172
rect 7680 14112 7744 14116
rect 13360 14172 13424 14176
rect 13360 14116 13364 14172
rect 13364 14116 13420 14172
rect 13420 14116 13424 14172
rect 13360 14112 13424 14116
rect 13440 14172 13504 14176
rect 13440 14116 13444 14172
rect 13444 14116 13500 14172
rect 13500 14116 13504 14172
rect 13440 14112 13504 14116
rect 13520 14172 13584 14176
rect 13520 14116 13524 14172
rect 13524 14116 13580 14172
rect 13580 14116 13584 14172
rect 13520 14112 13584 14116
rect 13600 14172 13664 14176
rect 13600 14116 13604 14172
rect 13604 14116 13660 14172
rect 13660 14116 13664 14172
rect 13600 14112 13664 14116
rect 13680 14172 13744 14176
rect 13680 14116 13684 14172
rect 13684 14116 13740 14172
rect 13740 14116 13744 14172
rect 13680 14112 13744 14116
rect 19360 14172 19424 14176
rect 19360 14116 19364 14172
rect 19364 14116 19420 14172
rect 19420 14116 19424 14172
rect 19360 14112 19424 14116
rect 19440 14172 19504 14176
rect 19440 14116 19444 14172
rect 19444 14116 19500 14172
rect 19500 14116 19504 14172
rect 19440 14112 19504 14116
rect 19520 14172 19584 14176
rect 19520 14116 19524 14172
rect 19524 14116 19580 14172
rect 19580 14116 19584 14172
rect 19520 14112 19584 14116
rect 19600 14172 19664 14176
rect 19600 14116 19604 14172
rect 19604 14116 19660 14172
rect 19660 14116 19664 14172
rect 19600 14112 19664 14116
rect 19680 14172 19744 14176
rect 19680 14116 19684 14172
rect 19684 14116 19740 14172
rect 19740 14116 19744 14172
rect 19680 14112 19744 14116
rect 4360 13628 4424 13632
rect 4360 13572 4364 13628
rect 4364 13572 4420 13628
rect 4420 13572 4424 13628
rect 4360 13568 4424 13572
rect 4440 13628 4504 13632
rect 4440 13572 4444 13628
rect 4444 13572 4500 13628
rect 4500 13572 4504 13628
rect 4440 13568 4504 13572
rect 4520 13628 4584 13632
rect 4520 13572 4524 13628
rect 4524 13572 4580 13628
rect 4580 13572 4584 13628
rect 4520 13568 4584 13572
rect 4600 13628 4664 13632
rect 4600 13572 4604 13628
rect 4604 13572 4660 13628
rect 4660 13572 4664 13628
rect 4600 13568 4664 13572
rect 4680 13628 4744 13632
rect 4680 13572 4684 13628
rect 4684 13572 4740 13628
rect 4740 13572 4744 13628
rect 4680 13568 4744 13572
rect 10360 13628 10424 13632
rect 10360 13572 10364 13628
rect 10364 13572 10420 13628
rect 10420 13572 10424 13628
rect 10360 13568 10424 13572
rect 10440 13628 10504 13632
rect 10440 13572 10444 13628
rect 10444 13572 10500 13628
rect 10500 13572 10504 13628
rect 10440 13568 10504 13572
rect 10520 13628 10584 13632
rect 10520 13572 10524 13628
rect 10524 13572 10580 13628
rect 10580 13572 10584 13628
rect 10520 13568 10584 13572
rect 10600 13628 10664 13632
rect 10600 13572 10604 13628
rect 10604 13572 10660 13628
rect 10660 13572 10664 13628
rect 10600 13568 10664 13572
rect 10680 13628 10744 13632
rect 10680 13572 10684 13628
rect 10684 13572 10740 13628
rect 10740 13572 10744 13628
rect 10680 13568 10744 13572
rect 16360 13628 16424 13632
rect 16360 13572 16364 13628
rect 16364 13572 16420 13628
rect 16420 13572 16424 13628
rect 16360 13568 16424 13572
rect 16440 13628 16504 13632
rect 16440 13572 16444 13628
rect 16444 13572 16500 13628
rect 16500 13572 16504 13628
rect 16440 13568 16504 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 22360 13628 22424 13632
rect 22360 13572 22364 13628
rect 22364 13572 22420 13628
rect 22420 13572 22424 13628
rect 22360 13568 22424 13572
rect 22440 13628 22504 13632
rect 22440 13572 22444 13628
rect 22444 13572 22500 13628
rect 22500 13572 22504 13628
rect 22440 13568 22504 13572
rect 22520 13628 22584 13632
rect 22520 13572 22524 13628
rect 22524 13572 22580 13628
rect 22580 13572 22584 13628
rect 22520 13568 22584 13572
rect 22600 13628 22664 13632
rect 22600 13572 22604 13628
rect 22604 13572 22660 13628
rect 22660 13572 22664 13628
rect 22600 13568 22664 13572
rect 22680 13628 22744 13632
rect 22680 13572 22684 13628
rect 22684 13572 22740 13628
rect 22740 13572 22744 13628
rect 22680 13568 22744 13572
rect 13124 13364 13188 13428
rect 1360 13084 1424 13088
rect 1360 13028 1364 13084
rect 1364 13028 1420 13084
rect 1420 13028 1424 13084
rect 1360 13024 1424 13028
rect 1440 13084 1504 13088
rect 1440 13028 1444 13084
rect 1444 13028 1500 13084
rect 1500 13028 1504 13084
rect 1440 13024 1504 13028
rect 1520 13084 1584 13088
rect 1520 13028 1524 13084
rect 1524 13028 1580 13084
rect 1580 13028 1584 13084
rect 1520 13024 1584 13028
rect 1600 13084 1664 13088
rect 1600 13028 1604 13084
rect 1604 13028 1660 13084
rect 1660 13028 1664 13084
rect 1600 13024 1664 13028
rect 1680 13084 1744 13088
rect 1680 13028 1684 13084
rect 1684 13028 1740 13084
rect 1740 13028 1744 13084
rect 1680 13024 1744 13028
rect 7360 13084 7424 13088
rect 7360 13028 7364 13084
rect 7364 13028 7420 13084
rect 7420 13028 7424 13084
rect 7360 13024 7424 13028
rect 7440 13084 7504 13088
rect 7440 13028 7444 13084
rect 7444 13028 7500 13084
rect 7500 13028 7504 13084
rect 7440 13024 7504 13028
rect 7520 13084 7584 13088
rect 7520 13028 7524 13084
rect 7524 13028 7580 13084
rect 7580 13028 7584 13084
rect 7520 13024 7584 13028
rect 7600 13084 7664 13088
rect 7600 13028 7604 13084
rect 7604 13028 7660 13084
rect 7660 13028 7664 13084
rect 7600 13024 7664 13028
rect 7680 13084 7744 13088
rect 7680 13028 7684 13084
rect 7684 13028 7740 13084
rect 7740 13028 7744 13084
rect 7680 13024 7744 13028
rect 13360 13084 13424 13088
rect 13360 13028 13364 13084
rect 13364 13028 13420 13084
rect 13420 13028 13424 13084
rect 13360 13024 13424 13028
rect 13440 13084 13504 13088
rect 13440 13028 13444 13084
rect 13444 13028 13500 13084
rect 13500 13028 13504 13084
rect 13440 13024 13504 13028
rect 13520 13084 13584 13088
rect 13520 13028 13524 13084
rect 13524 13028 13580 13084
rect 13580 13028 13584 13084
rect 13520 13024 13584 13028
rect 13600 13084 13664 13088
rect 13600 13028 13604 13084
rect 13604 13028 13660 13084
rect 13660 13028 13664 13084
rect 13600 13024 13664 13028
rect 13680 13084 13744 13088
rect 13680 13028 13684 13084
rect 13684 13028 13740 13084
rect 13740 13028 13744 13084
rect 13680 13024 13744 13028
rect 19360 13084 19424 13088
rect 19360 13028 19364 13084
rect 19364 13028 19420 13084
rect 19420 13028 19424 13084
rect 19360 13024 19424 13028
rect 19440 13084 19504 13088
rect 19440 13028 19444 13084
rect 19444 13028 19500 13084
rect 19500 13028 19504 13084
rect 19440 13024 19504 13028
rect 19520 13084 19584 13088
rect 19520 13028 19524 13084
rect 19524 13028 19580 13084
rect 19580 13028 19584 13084
rect 19520 13024 19584 13028
rect 19600 13084 19664 13088
rect 19600 13028 19604 13084
rect 19604 13028 19660 13084
rect 19660 13028 19664 13084
rect 19600 13024 19664 13028
rect 19680 13084 19744 13088
rect 19680 13028 19684 13084
rect 19684 13028 19740 13084
rect 19740 13028 19744 13084
rect 19680 13024 19744 13028
rect 15700 12820 15764 12884
rect 14964 12548 15028 12612
rect 4360 12540 4424 12544
rect 4360 12484 4364 12540
rect 4364 12484 4420 12540
rect 4420 12484 4424 12540
rect 4360 12480 4424 12484
rect 4440 12540 4504 12544
rect 4440 12484 4444 12540
rect 4444 12484 4500 12540
rect 4500 12484 4504 12540
rect 4440 12480 4504 12484
rect 4520 12540 4584 12544
rect 4520 12484 4524 12540
rect 4524 12484 4580 12540
rect 4580 12484 4584 12540
rect 4520 12480 4584 12484
rect 4600 12540 4664 12544
rect 4600 12484 4604 12540
rect 4604 12484 4660 12540
rect 4660 12484 4664 12540
rect 4600 12480 4664 12484
rect 4680 12540 4744 12544
rect 4680 12484 4684 12540
rect 4684 12484 4740 12540
rect 4740 12484 4744 12540
rect 4680 12480 4744 12484
rect 10360 12540 10424 12544
rect 10360 12484 10364 12540
rect 10364 12484 10420 12540
rect 10420 12484 10424 12540
rect 10360 12480 10424 12484
rect 10440 12540 10504 12544
rect 10440 12484 10444 12540
rect 10444 12484 10500 12540
rect 10500 12484 10504 12540
rect 10440 12480 10504 12484
rect 10520 12540 10584 12544
rect 10520 12484 10524 12540
rect 10524 12484 10580 12540
rect 10580 12484 10584 12540
rect 10520 12480 10584 12484
rect 10600 12540 10664 12544
rect 10600 12484 10604 12540
rect 10604 12484 10660 12540
rect 10660 12484 10664 12540
rect 10600 12480 10664 12484
rect 10680 12540 10744 12544
rect 10680 12484 10684 12540
rect 10684 12484 10740 12540
rect 10740 12484 10744 12540
rect 10680 12480 10744 12484
rect 16360 12540 16424 12544
rect 16360 12484 16364 12540
rect 16364 12484 16420 12540
rect 16420 12484 16424 12540
rect 16360 12480 16424 12484
rect 16440 12540 16504 12544
rect 16440 12484 16444 12540
rect 16444 12484 16500 12540
rect 16500 12484 16504 12540
rect 16440 12480 16504 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 22360 12540 22424 12544
rect 22360 12484 22364 12540
rect 22364 12484 22420 12540
rect 22420 12484 22424 12540
rect 22360 12480 22424 12484
rect 22440 12540 22504 12544
rect 22440 12484 22444 12540
rect 22444 12484 22500 12540
rect 22500 12484 22504 12540
rect 22440 12480 22504 12484
rect 22520 12540 22584 12544
rect 22520 12484 22524 12540
rect 22524 12484 22580 12540
rect 22580 12484 22584 12540
rect 22520 12480 22584 12484
rect 22600 12540 22664 12544
rect 22600 12484 22604 12540
rect 22604 12484 22660 12540
rect 22660 12484 22664 12540
rect 22600 12480 22664 12484
rect 22680 12540 22744 12544
rect 22680 12484 22684 12540
rect 22684 12484 22740 12540
rect 22740 12484 22744 12540
rect 22680 12480 22744 12484
rect 1360 11996 1424 12000
rect 1360 11940 1364 11996
rect 1364 11940 1420 11996
rect 1420 11940 1424 11996
rect 1360 11936 1424 11940
rect 1440 11996 1504 12000
rect 1440 11940 1444 11996
rect 1444 11940 1500 11996
rect 1500 11940 1504 11996
rect 1440 11936 1504 11940
rect 1520 11996 1584 12000
rect 1520 11940 1524 11996
rect 1524 11940 1580 11996
rect 1580 11940 1584 11996
rect 1520 11936 1584 11940
rect 1600 11996 1664 12000
rect 1600 11940 1604 11996
rect 1604 11940 1660 11996
rect 1660 11940 1664 11996
rect 1600 11936 1664 11940
rect 1680 11996 1744 12000
rect 1680 11940 1684 11996
rect 1684 11940 1740 11996
rect 1740 11940 1744 11996
rect 1680 11936 1744 11940
rect 7360 11996 7424 12000
rect 7360 11940 7364 11996
rect 7364 11940 7420 11996
rect 7420 11940 7424 11996
rect 7360 11936 7424 11940
rect 7440 11996 7504 12000
rect 7440 11940 7444 11996
rect 7444 11940 7500 11996
rect 7500 11940 7504 11996
rect 7440 11936 7504 11940
rect 7520 11996 7584 12000
rect 7520 11940 7524 11996
rect 7524 11940 7580 11996
rect 7580 11940 7584 11996
rect 7520 11936 7584 11940
rect 7600 11996 7664 12000
rect 7600 11940 7604 11996
rect 7604 11940 7660 11996
rect 7660 11940 7664 11996
rect 7600 11936 7664 11940
rect 7680 11996 7744 12000
rect 7680 11940 7684 11996
rect 7684 11940 7740 11996
rect 7740 11940 7744 11996
rect 7680 11936 7744 11940
rect 13360 11996 13424 12000
rect 13360 11940 13364 11996
rect 13364 11940 13420 11996
rect 13420 11940 13424 11996
rect 13360 11936 13424 11940
rect 13440 11996 13504 12000
rect 13440 11940 13444 11996
rect 13444 11940 13500 11996
rect 13500 11940 13504 11996
rect 13440 11936 13504 11940
rect 13520 11996 13584 12000
rect 13520 11940 13524 11996
rect 13524 11940 13580 11996
rect 13580 11940 13584 11996
rect 13520 11936 13584 11940
rect 13600 11996 13664 12000
rect 13600 11940 13604 11996
rect 13604 11940 13660 11996
rect 13660 11940 13664 11996
rect 13600 11936 13664 11940
rect 13680 11996 13744 12000
rect 13680 11940 13684 11996
rect 13684 11940 13740 11996
rect 13740 11940 13744 11996
rect 13680 11936 13744 11940
rect 19360 11996 19424 12000
rect 19360 11940 19364 11996
rect 19364 11940 19420 11996
rect 19420 11940 19424 11996
rect 19360 11936 19424 11940
rect 19440 11996 19504 12000
rect 19440 11940 19444 11996
rect 19444 11940 19500 11996
rect 19500 11940 19504 11996
rect 19440 11936 19504 11940
rect 19520 11996 19584 12000
rect 19520 11940 19524 11996
rect 19524 11940 19580 11996
rect 19580 11940 19584 11996
rect 19520 11936 19584 11940
rect 19600 11996 19664 12000
rect 19600 11940 19604 11996
rect 19604 11940 19660 11996
rect 19660 11940 19664 11996
rect 19600 11936 19664 11940
rect 19680 11996 19744 12000
rect 19680 11940 19684 11996
rect 19684 11940 19740 11996
rect 19740 11940 19744 11996
rect 19680 11936 19744 11940
rect 4108 11460 4172 11524
rect 4360 11452 4424 11456
rect 4360 11396 4364 11452
rect 4364 11396 4420 11452
rect 4420 11396 4424 11452
rect 4360 11392 4424 11396
rect 4440 11452 4504 11456
rect 4440 11396 4444 11452
rect 4444 11396 4500 11452
rect 4500 11396 4504 11452
rect 4440 11392 4504 11396
rect 4520 11452 4584 11456
rect 4520 11396 4524 11452
rect 4524 11396 4580 11452
rect 4580 11396 4584 11452
rect 4520 11392 4584 11396
rect 4600 11452 4664 11456
rect 4600 11396 4604 11452
rect 4604 11396 4660 11452
rect 4660 11396 4664 11452
rect 4600 11392 4664 11396
rect 4680 11452 4744 11456
rect 4680 11396 4684 11452
rect 4684 11396 4740 11452
rect 4740 11396 4744 11452
rect 4680 11392 4744 11396
rect 10360 11452 10424 11456
rect 10360 11396 10364 11452
rect 10364 11396 10420 11452
rect 10420 11396 10424 11452
rect 10360 11392 10424 11396
rect 10440 11452 10504 11456
rect 10440 11396 10444 11452
rect 10444 11396 10500 11452
rect 10500 11396 10504 11452
rect 10440 11392 10504 11396
rect 10520 11452 10584 11456
rect 10520 11396 10524 11452
rect 10524 11396 10580 11452
rect 10580 11396 10584 11452
rect 10520 11392 10584 11396
rect 10600 11452 10664 11456
rect 10600 11396 10604 11452
rect 10604 11396 10660 11452
rect 10660 11396 10664 11452
rect 10600 11392 10664 11396
rect 10680 11452 10744 11456
rect 10680 11396 10684 11452
rect 10684 11396 10740 11452
rect 10740 11396 10744 11452
rect 10680 11392 10744 11396
rect 16360 11452 16424 11456
rect 16360 11396 16364 11452
rect 16364 11396 16420 11452
rect 16420 11396 16424 11452
rect 16360 11392 16424 11396
rect 16440 11452 16504 11456
rect 16440 11396 16444 11452
rect 16444 11396 16500 11452
rect 16500 11396 16504 11452
rect 16440 11392 16504 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 22360 11452 22424 11456
rect 22360 11396 22364 11452
rect 22364 11396 22420 11452
rect 22420 11396 22424 11452
rect 22360 11392 22424 11396
rect 22440 11452 22504 11456
rect 22440 11396 22444 11452
rect 22444 11396 22500 11452
rect 22500 11396 22504 11452
rect 22440 11392 22504 11396
rect 22520 11452 22584 11456
rect 22520 11396 22524 11452
rect 22524 11396 22580 11452
rect 22580 11396 22584 11452
rect 22520 11392 22584 11396
rect 22600 11452 22664 11456
rect 22600 11396 22604 11452
rect 22604 11396 22660 11452
rect 22660 11396 22664 11452
rect 22600 11392 22664 11396
rect 22680 11452 22744 11456
rect 22680 11396 22684 11452
rect 22684 11396 22740 11452
rect 22740 11396 22744 11452
rect 22680 11392 22744 11396
rect 1360 10908 1424 10912
rect 1360 10852 1364 10908
rect 1364 10852 1420 10908
rect 1420 10852 1424 10908
rect 1360 10848 1424 10852
rect 1440 10908 1504 10912
rect 1440 10852 1444 10908
rect 1444 10852 1500 10908
rect 1500 10852 1504 10908
rect 1440 10848 1504 10852
rect 1520 10908 1584 10912
rect 1520 10852 1524 10908
rect 1524 10852 1580 10908
rect 1580 10852 1584 10908
rect 1520 10848 1584 10852
rect 1600 10908 1664 10912
rect 1600 10852 1604 10908
rect 1604 10852 1660 10908
rect 1660 10852 1664 10908
rect 1600 10848 1664 10852
rect 1680 10908 1744 10912
rect 1680 10852 1684 10908
rect 1684 10852 1740 10908
rect 1740 10852 1744 10908
rect 1680 10848 1744 10852
rect 7360 10908 7424 10912
rect 7360 10852 7364 10908
rect 7364 10852 7420 10908
rect 7420 10852 7424 10908
rect 7360 10848 7424 10852
rect 7440 10908 7504 10912
rect 7440 10852 7444 10908
rect 7444 10852 7500 10908
rect 7500 10852 7504 10908
rect 7440 10848 7504 10852
rect 7520 10908 7584 10912
rect 7520 10852 7524 10908
rect 7524 10852 7580 10908
rect 7580 10852 7584 10908
rect 7520 10848 7584 10852
rect 7600 10908 7664 10912
rect 7600 10852 7604 10908
rect 7604 10852 7660 10908
rect 7660 10852 7664 10908
rect 7600 10848 7664 10852
rect 7680 10908 7744 10912
rect 7680 10852 7684 10908
rect 7684 10852 7740 10908
rect 7740 10852 7744 10908
rect 7680 10848 7744 10852
rect 13360 10908 13424 10912
rect 13360 10852 13364 10908
rect 13364 10852 13420 10908
rect 13420 10852 13424 10908
rect 13360 10848 13424 10852
rect 13440 10908 13504 10912
rect 13440 10852 13444 10908
rect 13444 10852 13500 10908
rect 13500 10852 13504 10908
rect 13440 10848 13504 10852
rect 13520 10908 13584 10912
rect 13520 10852 13524 10908
rect 13524 10852 13580 10908
rect 13580 10852 13584 10908
rect 13520 10848 13584 10852
rect 13600 10908 13664 10912
rect 13600 10852 13604 10908
rect 13604 10852 13660 10908
rect 13660 10852 13664 10908
rect 13600 10848 13664 10852
rect 13680 10908 13744 10912
rect 13680 10852 13684 10908
rect 13684 10852 13740 10908
rect 13740 10852 13744 10908
rect 13680 10848 13744 10852
rect 19360 10908 19424 10912
rect 19360 10852 19364 10908
rect 19364 10852 19420 10908
rect 19420 10852 19424 10908
rect 19360 10848 19424 10852
rect 19440 10908 19504 10912
rect 19440 10852 19444 10908
rect 19444 10852 19500 10908
rect 19500 10852 19504 10908
rect 19440 10848 19504 10852
rect 19520 10908 19584 10912
rect 19520 10852 19524 10908
rect 19524 10852 19580 10908
rect 19580 10852 19584 10908
rect 19520 10848 19584 10852
rect 19600 10908 19664 10912
rect 19600 10852 19604 10908
rect 19604 10852 19660 10908
rect 19660 10852 19664 10908
rect 19600 10848 19664 10852
rect 19680 10908 19744 10912
rect 19680 10852 19684 10908
rect 19684 10852 19740 10908
rect 19740 10852 19744 10908
rect 19680 10848 19744 10852
rect 4360 10364 4424 10368
rect 4360 10308 4364 10364
rect 4364 10308 4420 10364
rect 4420 10308 4424 10364
rect 4360 10304 4424 10308
rect 4440 10364 4504 10368
rect 4440 10308 4444 10364
rect 4444 10308 4500 10364
rect 4500 10308 4504 10364
rect 4440 10304 4504 10308
rect 4520 10364 4584 10368
rect 4520 10308 4524 10364
rect 4524 10308 4580 10364
rect 4580 10308 4584 10364
rect 4520 10304 4584 10308
rect 4600 10364 4664 10368
rect 4600 10308 4604 10364
rect 4604 10308 4660 10364
rect 4660 10308 4664 10364
rect 4600 10304 4664 10308
rect 4680 10364 4744 10368
rect 4680 10308 4684 10364
rect 4684 10308 4740 10364
rect 4740 10308 4744 10364
rect 4680 10304 4744 10308
rect 10360 10364 10424 10368
rect 10360 10308 10364 10364
rect 10364 10308 10420 10364
rect 10420 10308 10424 10364
rect 10360 10304 10424 10308
rect 10440 10364 10504 10368
rect 10440 10308 10444 10364
rect 10444 10308 10500 10364
rect 10500 10308 10504 10364
rect 10440 10304 10504 10308
rect 10520 10364 10584 10368
rect 10520 10308 10524 10364
rect 10524 10308 10580 10364
rect 10580 10308 10584 10364
rect 10520 10304 10584 10308
rect 10600 10364 10664 10368
rect 10600 10308 10604 10364
rect 10604 10308 10660 10364
rect 10660 10308 10664 10364
rect 10600 10304 10664 10308
rect 10680 10364 10744 10368
rect 10680 10308 10684 10364
rect 10684 10308 10740 10364
rect 10740 10308 10744 10364
rect 10680 10304 10744 10308
rect 16360 10364 16424 10368
rect 16360 10308 16364 10364
rect 16364 10308 16420 10364
rect 16420 10308 16424 10364
rect 16360 10304 16424 10308
rect 16440 10364 16504 10368
rect 16440 10308 16444 10364
rect 16444 10308 16500 10364
rect 16500 10308 16504 10364
rect 16440 10304 16504 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 22360 10364 22424 10368
rect 22360 10308 22364 10364
rect 22364 10308 22420 10364
rect 22420 10308 22424 10364
rect 22360 10304 22424 10308
rect 22440 10364 22504 10368
rect 22440 10308 22444 10364
rect 22444 10308 22500 10364
rect 22500 10308 22504 10364
rect 22440 10304 22504 10308
rect 22520 10364 22584 10368
rect 22520 10308 22524 10364
rect 22524 10308 22580 10364
rect 22580 10308 22584 10364
rect 22520 10304 22584 10308
rect 22600 10364 22664 10368
rect 22600 10308 22604 10364
rect 22604 10308 22660 10364
rect 22660 10308 22664 10364
rect 22600 10304 22664 10308
rect 22680 10364 22744 10368
rect 22680 10308 22684 10364
rect 22684 10308 22740 10364
rect 22740 10308 22744 10364
rect 22680 10304 22744 10308
rect 15148 10236 15212 10300
rect 1360 9820 1424 9824
rect 1360 9764 1364 9820
rect 1364 9764 1420 9820
rect 1420 9764 1424 9820
rect 1360 9760 1424 9764
rect 1440 9820 1504 9824
rect 1440 9764 1444 9820
rect 1444 9764 1500 9820
rect 1500 9764 1504 9820
rect 1440 9760 1504 9764
rect 1520 9820 1584 9824
rect 1520 9764 1524 9820
rect 1524 9764 1580 9820
rect 1580 9764 1584 9820
rect 1520 9760 1584 9764
rect 1600 9820 1664 9824
rect 1600 9764 1604 9820
rect 1604 9764 1660 9820
rect 1660 9764 1664 9820
rect 1600 9760 1664 9764
rect 1680 9820 1744 9824
rect 1680 9764 1684 9820
rect 1684 9764 1740 9820
rect 1740 9764 1744 9820
rect 1680 9760 1744 9764
rect 7360 9820 7424 9824
rect 7360 9764 7364 9820
rect 7364 9764 7420 9820
rect 7420 9764 7424 9820
rect 7360 9760 7424 9764
rect 7440 9820 7504 9824
rect 7440 9764 7444 9820
rect 7444 9764 7500 9820
rect 7500 9764 7504 9820
rect 7440 9760 7504 9764
rect 7520 9820 7584 9824
rect 7520 9764 7524 9820
rect 7524 9764 7580 9820
rect 7580 9764 7584 9820
rect 7520 9760 7584 9764
rect 7600 9820 7664 9824
rect 7600 9764 7604 9820
rect 7604 9764 7660 9820
rect 7660 9764 7664 9820
rect 7600 9760 7664 9764
rect 7680 9820 7744 9824
rect 7680 9764 7684 9820
rect 7684 9764 7740 9820
rect 7740 9764 7744 9820
rect 7680 9760 7744 9764
rect 13360 9820 13424 9824
rect 13360 9764 13364 9820
rect 13364 9764 13420 9820
rect 13420 9764 13424 9820
rect 13360 9760 13424 9764
rect 13440 9820 13504 9824
rect 13440 9764 13444 9820
rect 13444 9764 13500 9820
rect 13500 9764 13504 9820
rect 13440 9760 13504 9764
rect 13520 9820 13584 9824
rect 13520 9764 13524 9820
rect 13524 9764 13580 9820
rect 13580 9764 13584 9820
rect 13520 9760 13584 9764
rect 13600 9820 13664 9824
rect 13600 9764 13604 9820
rect 13604 9764 13660 9820
rect 13660 9764 13664 9820
rect 13600 9760 13664 9764
rect 13680 9820 13744 9824
rect 13680 9764 13684 9820
rect 13684 9764 13740 9820
rect 13740 9764 13744 9820
rect 13680 9760 13744 9764
rect 19360 9820 19424 9824
rect 19360 9764 19364 9820
rect 19364 9764 19420 9820
rect 19420 9764 19424 9820
rect 19360 9760 19424 9764
rect 19440 9820 19504 9824
rect 19440 9764 19444 9820
rect 19444 9764 19500 9820
rect 19500 9764 19504 9820
rect 19440 9760 19504 9764
rect 19520 9820 19584 9824
rect 19520 9764 19524 9820
rect 19524 9764 19580 9820
rect 19580 9764 19584 9820
rect 19520 9760 19584 9764
rect 19600 9820 19664 9824
rect 19600 9764 19604 9820
rect 19604 9764 19660 9820
rect 19660 9764 19664 9820
rect 19600 9760 19664 9764
rect 19680 9820 19744 9824
rect 19680 9764 19684 9820
rect 19684 9764 19740 9820
rect 19740 9764 19744 9820
rect 19680 9760 19744 9764
rect 9812 9692 9876 9756
rect 11100 9420 11164 9484
rect 4360 9276 4424 9280
rect 4360 9220 4364 9276
rect 4364 9220 4420 9276
rect 4420 9220 4424 9276
rect 4360 9216 4424 9220
rect 4440 9276 4504 9280
rect 4440 9220 4444 9276
rect 4444 9220 4500 9276
rect 4500 9220 4504 9276
rect 4440 9216 4504 9220
rect 4520 9276 4584 9280
rect 4520 9220 4524 9276
rect 4524 9220 4580 9276
rect 4580 9220 4584 9276
rect 4520 9216 4584 9220
rect 4600 9276 4664 9280
rect 4600 9220 4604 9276
rect 4604 9220 4660 9276
rect 4660 9220 4664 9276
rect 4600 9216 4664 9220
rect 4680 9276 4744 9280
rect 4680 9220 4684 9276
rect 4684 9220 4740 9276
rect 4740 9220 4744 9276
rect 4680 9216 4744 9220
rect 10360 9276 10424 9280
rect 10360 9220 10364 9276
rect 10364 9220 10420 9276
rect 10420 9220 10424 9276
rect 10360 9216 10424 9220
rect 10440 9276 10504 9280
rect 10440 9220 10444 9276
rect 10444 9220 10500 9276
rect 10500 9220 10504 9276
rect 10440 9216 10504 9220
rect 10520 9276 10584 9280
rect 10520 9220 10524 9276
rect 10524 9220 10580 9276
rect 10580 9220 10584 9276
rect 10520 9216 10584 9220
rect 10600 9276 10664 9280
rect 10600 9220 10604 9276
rect 10604 9220 10660 9276
rect 10660 9220 10664 9276
rect 10600 9216 10664 9220
rect 10680 9276 10744 9280
rect 10680 9220 10684 9276
rect 10684 9220 10740 9276
rect 10740 9220 10744 9276
rect 10680 9216 10744 9220
rect 16360 9276 16424 9280
rect 16360 9220 16364 9276
rect 16364 9220 16420 9276
rect 16420 9220 16424 9276
rect 16360 9216 16424 9220
rect 16440 9276 16504 9280
rect 16440 9220 16444 9276
rect 16444 9220 16500 9276
rect 16500 9220 16504 9276
rect 16440 9216 16504 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 22360 9276 22424 9280
rect 22360 9220 22364 9276
rect 22364 9220 22420 9276
rect 22420 9220 22424 9276
rect 22360 9216 22424 9220
rect 22440 9276 22504 9280
rect 22440 9220 22444 9276
rect 22444 9220 22500 9276
rect 22500 9220 22504 9276
rect 22440 9216 22504 9220
rect 22520 9276 22584 9280
rect 22520 9220 22524 9276
rect 22524 9220 22580 9276
rect 22580 9220 22584 9276
rect 22520 9216 22584 9220
rect 22600 9276 22664 9280
rect 22600 9220 22604 9276
rect 22604 9220 22660 9276
rect 22660 9220 22664 9276
rect 22600 9216 22664 9220
rect 22680 9276 22744 9280
rect 22680 9220 22684 9276
rect 22684 9220 22740 9276
rect 22740 9220 22744 9276
rect 22680 9216 22744 9220
rect 14780 9148 14844 9212
rect 19932 9148 19996 9212
rect 1360 8732 1424 8736
rect 1360 8676 1364 8732
rect 1364 8676 1420 8732
rect 1420 8676 1424 8732
rect 1360 8672 1424 8676
rect 1440 8732 1504 8736
rect 1440 8676 1444 8732
rect 1444 8676 1500 8732
rect 1500 8676 1504 8732
rect 1440 8672 1504 8676
rect 1520 8732 1584 8736
rect 1520 8676 1524 8732
rect 1524 8676 1580 8732
rect 1580 8676 1584 8732
rect 1520 8672 1584 8676
rect 1600 8732 1664 8736
rect 1600 8676 1604 8732
rect 1604 8676 1660 8732
rect 1660 8676 1664 8732
rect 1600 8672 1664 8676
rect 1680 8732 1744 8736
rect 1680 8676 1684 8732
rect 1684 8676 1740 8732
rect 1740 8676 1744 8732
rect 1680 8672 1744 8676
rect 7360 8732 7424 8736
rect 7360 8676 7364 8732
rect 7364 8676 7420 8732
rect 7420 8676 7424 8732
rect 7360 8672 7424 8676
rect 7440 8732 7504 8736
rect 7440 8676 7444 8732
rect 7444 8676 7500 8732
rect 7500 8676 7504 8732
rect 7440 8672 7504 8676
rect 7520 8732 7584 8736
rect 7520 8676 7524 8732
rect 7524 8676 7580 8732
rect 7580 8676 7584 8732
rect 7520 8672 7584 8676
rect 7600 8732 7664 8736
rect 7600 8676 7604 8732
rect 7604 8676 7660 8732
rect 7660 8676 7664 8732
rect 7600 8672 7664 8676
rect 7680 8732 7744 8736
rect 7680 8676 7684 8732
rect 7684 8676 7740 8732
rect 7740 8676 7744 8732
rect 7680 8672 7744 8676
rect 13360 8732 13424 8736
rect 13360 8676 13364 8732
rect 13364 8676 13420 8732
rect 13420 8676 13424 8732
rect 13360 8672 13424 8676
rect 13440 8732 13504 8736
rect 13440 8676 13444 8732
rect 13444 8676 13500 8732
rect 13500 8676 13504 8732
rect 13440 8672 13504 8676
rect 13520 8732 13584 8736
rect 13520 8676 13524 8732
rect 13524 8676 13580 8732
rect 13580 8676 13584 8732
rect 13520 8672 13584 8676
rect 13600 8732 13664 8736
rect 13600 8676 13604 8732
rect 13604 8676 13660 8732
rect 13660 8676 13664 8732
rect 13600 8672 13664 8676
rect 13680 8732 13744 8736
rect 13680 8676 13684 8732
rect 13684 8676 13740 8732
rect 13740 8676 13744 8732
rect 13680 8672 13744 8676
rect 19360 8732 19424 8736
rect 19360 8676 19364 8732
rect 19364 8676 19420 8732
rect 19420 8676 19424 8732
rect 19360 8672 19424 8676
rect 19440 8732 19504 8736
rect 19440 8676 19444 8732
rect 19444 8676 19500 8732
rect 19500 8676 19504 8732
rect 19440 8672 19504 8676
rect 19520 8732 19584 8736
rect 19520 8676 19524 8732
rect 19524 8676 19580 8732
rect 19580 8676 19584 8732
rect 19520 8672 19584 8676
rect 19600 8732 19664 8736
rect 19600 8676 19604 8732
rect 19604 8676 19660 8732
rect 19660 8676 19664 8732
rect 19600 8672 19664 8676
rect 19680 8732 19744 8736
rect 19680 8676 19684 8732
rect 19684 8676 19740 8732
rect 19740 8676 19744 8732
rect 19680 8672 19744 8676
rect 19932 8256 19996 8260
rect 19932 8200 19982 8256
rect 19982 8200 19996 8256
rect 19932 8196 19996 8200
rect 4360 8188 4424 8192
rect 4360 8132 4364 8188
rect 4364 8132 4420 8188
rect 4420 8132 4424 8188
rect 4360 8128 4424 8132
rect 4440 8188 4504 8192
rect 4440 8132 4444 8188
rect 4444 8132 4500 8188
rect 4500 8132 4504 8188
rect 4440 8128 4504 8132
rect 4520 8188 4584 8192
rect 4520 8132 4524 8188
rect 4524 8132 4580 8188
rect 4580 8132 4584 8188
rect 4520 8128 4584 8132
rect 4600 8188 4664 8192
rect 4600 8132 4604 8188
rect 4604 8132 4660 8188
rect 4660 8132 4664 8188
rect 4600 8128 4664 8132
rect 4680 8188 4744 8192
rect 4680 8132 4684 8188
rect 4684 8132 4740 8188
rect 4740 8132 4744 8188
rect 4680 8128 4744 8132
rect 10360 8188 10424 8192
rect 10360 8132 10364 8188
rect 10364 8132 10420 8188
rect 10420 8132 10424 8188
rect 10360 8128 10424 8132
rect 10440 8188 10504 8192
rect 10440 8132 10444 8188
rect 10444 8132 10500 8188
rect 10500 8132 10504 8188
rect 10440 8128 10504 8132
rect 10520 8188 10584 8192
rect 10520 8132 10524 8188
rect 10524 8132 10580 8188
rect 10580 8132 10584 8188
rect 10520 8128 10584 8132
rect 10600 8188 10664 8192
rect 10600 8132 10604 8188
rect 10604 8132 10660 8188
rect 10660 8132 10664 8188
rect 10600 8128 10664 8132
rect 10680 8188 10744 8192
rect 10680 8132 10684 8188
rect 10684 8132 10740 8188
rect 10740 8132 10744 8188
rect 10680 8128 10744 8132
rect 16360 8188 16424 8192
rect 16360 8132 16364 8188
rect 16364 8132 16420 8188
rect 16420 8132 16424 8188
rect 16360 8128 16424 8132
rect 16440 8188 16504 8192
rect 16440 8132 16444 8188
rect 16444 8132 16500 8188
rect 16500 8132 16504 8188
rect 16440 8128 16504 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 22360 8188 22424 8192
rect 22360 8132 22364 8188
rect 22364 8132 22420 8188
rect 22420 8132 22424 8188
rect 22360 8128 22424 8132
rect 22440 8188 22504 8192
rect 22440 8132 22444 8188
rect 22444 8132 22500 8188
rect 22500 8132 22504 8188
rect 22440 8128 22504 8132
rect 22520 8188 22584 8192
rect 22520 8132 22524 8188
rect 22524 8132 22580 8188
rect 22580 8132 22584 8188
rect 22520 8128 22584 8132
rect 22600 8188 22664 8192
rect 22600 8132 22604 8188
rect 22604 8132 22660 8188
rect 22660 8132 22664 8188
rect 22600 8128 22664 8132
rect 22680 8188 22744 8192
rect 22680 8132 22684 8188
rect 22684 8132 22740 8188
rect 22740 8132 22744 8188
rect 22680 8128 22744 8132
rect 4108 7788 4172 7852
rect 1360 7644 1424 7648
rect 1360 7588 1364 7644
rect 1364 7588 1420 7644
rect 1420 7588 1424 7644
rect 1360 7584 1424 7588
rect 1440 7644 1504 7648
rect 1440 7588 1444 7644
rect 1444 7588 1500 7644
rect 1500 7588 1504 7644
rect 1440 7584 1504 7588
rect 1520 7644 1584 7648
rect 1520 7588 1524 7644
rect 1524 7588 1580 7644
rect 1580 7588 1584 7644
rect 1520 7584 1584 7588
rect 1600 7644 1664 7648
rect 1600 7588 1604 7644
rect 1604 7588 1660 7644
rect 1660 7588 1664 7644
rect 1600 7584 1664 7588
rect 1680 7644 1744 7648
rect 1680 7588 1684 7644
rect 1684 7588 1740 7644
rect 1740 7588 1744 7644
rect 1680 7584 1744 7588
rect 7360 7644 7424 7648
rect 7360 7588 7364 7644
rect 7364 7588 7420 7644
rect 7420 7588 7424 7644
rect 7360 7584 7424 7588
rect 7440 7644 7504 7648
rect 7440 7588 7444 7644
rect 7444 7588 7500 7644
rect 7500 7588 7504 7644
rect 7440 7584 7504 7588
rect 7520 7644 7584 7648
rect 7520 7588 7524 7644
rect 7524 7588 7580 7644
rect 7580 7588 7584 7644
rect 7520 7584 7584 7588
rect 7600 7644 7664 7648
rect 7600 7588 7604 7644
rect 7604 7588 7660 7644
rect 7660 7588 7664 7644
rect 7600 7584 7664 7588
rect 7680 7644 7744 7648
rect 7680 7588 7684 7644
rect 7684 7588 7740 7644
rect 7740 7588 7744 7644
rect 7680 7584 7744 7588
rect 13360 7644 13424 7648
rect 13360 7588 13364 7644
rect 13364 7588 13420 7644
rect 13420 7588 13424 7644
rect 13360 7584 13424 7588
rect 13440 7644 13504 7648
rect 13440 7588 13444 7644
rect 13444 7588 13500 7644
rect 13500 7588 13504 7644
rect 13440 7584 13504 7588
rect 13520 7644 13584 7648
rect 13520 7588 13524 7644
rect 13524 7588 13580 7644
rect 13580 7588 13584 7644
rect 13520 7584 13584 7588
rect 13600 7644 13664 7648
rect 13600 7588 13604 7644
rect 13604 7588 13660 7644
rect 13660 7588 13664 7644
rect 13600 7584 13664 7588
rect 13680 7644 13744 7648
rect 13680 7588 13684 7644
rect 13684 7588 13740 7644
rect 13740 7588 13744 7644
rect 13680 7584 13744 7588
rect 19360 7644 19424 7648
rect 19360 7588 19364 7644
rect 19364 7588 19420 7644
rect 19420 7588 19424 7644
rect 19360 7584 19424 7588
rect 19440 7644 19504 7648
rect 19440 7588 19444 7644
rect 19444 7588 19500 7644
rect 19500 7588 19504 7644
rect 19440 7584 19504 7588
rect 19520 7644 19584 7648
rect 19520 7588 19524 7644
rect 19524 7588 19580 7644
rect 19580 7588 19584 7644
rect 19520 7584 19584 7588
rect 19600 7644 19664 7648
rect 19600 7588 19604 7644
rect 19604 7588 19660 7644
rect 19660 7588 19664 7644
rect 19600 7584 19664 7588
rect 19680 7644 19744 7648
rect 19680 7588 19684 7644
rect 19684 7588 19740 7644
rect 19740 7588 19744 7644
rect 19680 7584 19744 7588
rect 9812 7244 9876 7308
rect 4360 7100 4424 7104
rect 4360 7044 4364 7100
rect 4364 7044 4420 7100
rect 4420 7044 4424 7100
rect 4360 7040 4424 7044
rect 4440 7100 4504 7104
rect 4440 7044 4444 7100
rect 4444 7044 4500 7100
rect 4500 7044 4504 7100
rect 4440 7040 4504 7044
rect 4520 7100 4584 7104
rect 4520 7044 4524 7100
rect 4524 7044 4580 7100
rect 4580 7044 4584 7100
rect 4520 7040 4584 7044
rect 4600 7100 4664 7104
rect 4600 7044 4604 7100
rect 4604 7044 4660 7100
rect 4660 7044 4664 7100
rect 4600 7040 4664 7044
rect 4680 7100 4744 7104
rect 4680 7044 4684 7100
rect 4684 7044 4740 7100
rect 4740 7044 4744 7100
rect 4680 7040 4744 7044
rect 10360 7100 10424 7104
rect 10360 7044 10364 7100
rect 10364 7044 10420 7100
rect 10420 7044 10424 7100
rect 10360 7040 10424 7044
rect 10440 7100 10504 7104
rect 10440 7044 10444 7100
rect 10444 7044 10500 7100
rect 10500 7044 10504 7100
rect 10440 7040 10504 7044
rect 10520 7100 10584 7104
rect 10520 7044 10524 7100
rect 10524 7044 10580 7100
rect 10580 7044 10584 7100
rect 10520 7040 10584 7044
rect 10600 7100 10664 7104
rect 10600 7044 10604 7100
rect 10604 7044 10660 7100
rect 10660 7044 10664 7100
rect 10600 7040 10664 7044
rect 10680 7100 10744 7104
rect 10680 7044 10684 7100
rect 10684 7044 10740 7100
rect 10740 7044 10744 7100
rect 10680 7040 10744 7044
rect 16360 7100 16424 7104
rect 16360 7044 16364 7100
rect 16364 7044 16420 7100
rect 16420 7044 16424 7100
rect 16360 7040 16424 7044
rect 16440 7100 16504 7104
rect 16440 7044 16444 7100
rect 16444 7044 16500 7100
rect 16500 7044 16504 7100
rect 16440 7040 16504 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 22360 7100 22424 7104
rect 22360 7044 22364 7100
rect 22364 7044 22420 7100
rect 22420 7044 22424 7100
rect 22360 7040 22424 7044
rect 22440 7100 22504 7104
rect 22440 7044 22444 7100
rect 22444 7044 22500 7100
rect 22500 7044 22504 7100
rect 22440 7040 22504 7044
rect 22520 7100 22584 7104
rect 22520 7044 22524 7100
rect 22524 7044 22580 7100
rect 22580 7044 22584 7100
rect 22520 7040 22584 7044
rect 22600 7100 22664 7104
rect 22600 7044 22604 7100
rect 22604 7044 22660 7100
rect 22660 7044 22664 7100
rect 22600 7040 22664 7044
rect 22680 7100 22744 7104
rect 22680 7044 22684 7100
rect 22684 7044 22740 7100
rect 22740 7044 22744 7100
rect 22680 7040 22744 7044
rect 15700 6836 15764 6900
rect 1360 6556 1424 6560
rect 1360 6500 1364 6556
rect 1364 6500 1420 6556
rect 1420 6500 1424 6556
rect 1360 6496 1424 6500
rect 1440 6556 1504 6560
rect 1440 6500 1444 6556
rect 1444 6500 1500 6556
rect 1500 6500 1504 6556
rect 1440 6496 1504 6500
rect 1520 6556 1584 6560
rect 1520 6500 1524 6556
rect 1524 6500 1580 6556
rect 1580 6500 1584 6556
rect 1520 6496 1584 6500
rect 1600 6556 1664 6560
rect 1600 6500 1604 6556
rect 1604 6500 1660 6556
rect 1660 6500 1664 6556
rect 1600 6496 1664 6500
rect 1680 6556 1744 6560
rect 1680 6500 1684 6556
rect 1684 6500 1740 6556
rect 1740 6500 1744 6556
rect 1680 6496 1744 6500
rect 7360 6556 7424 6560
rect 7360 6500 7364 6556
rect 7364 6500 7420 6556
rect 7420 6500 7424 6556
rect 7360 6496 7424 6500
rect 7440 6556 7504 6560
rect 7440 6500 7444 6556
rect 7444 6500 7500 6556
rect 7500 6500 7504 6556
rect 7440 6496 7504 6500
rect 7520 6556 7584 6560
rect 7520 6500 7524 6556
rect 7524 6500 7580 6556
rect 7580 6500 7584 6556
rect 7520 6496 7584 6500
rect 7600 6556 7664 6560
rect 7600 6500 7604 6556
rect 7604 6500 7660 6556
rect 7660 6500 7664 6556
rect 7600 6496 7664 6500
rect 7680 6556 7744 6560
rect 7680 6500 7684 6556
rect 7684 6500 7740 6556
rect 7740 6500 7744 6556
rect 7680 6496 7744 6500
rect 13360 6556 13424 6560
rect 13360 6500 13364 6556
rect 13364 6500 13420 6556
rect 13420 6500 13424 6556
rect 13360 6496 13424 6500
rect 13440 6556 13504 6560
rect 13440 6500 13444 6556
rect 13444 6500 13500 6556
rect 13500 6500 13504 6556
rect 13440 6496 13504 6500
rect 13520 6556 13584 6560
rect 13520 6500 13524 6556
rect 13524 6500 13580 6556
rect 13580 6500 13584 6556
rect 13520 6496 13584 6500
rect 13600 6556 13664 6560
rect 13600 6500 13604 6556
rect 13604 6500 13660 6556
rect 13660 6500 13664 6556
rect 13600 6496 13664 6500
rect 13680 6556 13744 6560
rect 13680 6500 13684 6556
rect 13684 6500 13740 6556
rect 13740 6500 13744 6556
rect 13680 6496 13744 6500
rect 19360 6556 19424 6560
rect 19360 6500 19364 6556
rect 19364 6500 19420 6556
rect 19420 6500 19424 6556
rect 19360 6496 19424 6500
rect 19440 6556 19504 6560
rect 19440 6500 19444 6556
rect 19444 6500 19500 6556
rect 19500 6500 19504 6556
rect 19440 6496 19504 6500
rect 19520 6556 19584 6560
rect 19520 6500 19524 6556
rect 19524 6500 19580 6556
rect 19580 6500 19584 6556
rect 19520 6496 19584 6500
rect 19600 6556 19664 6560
rect 19600 6500 19604 6556
rect 19604 6500 19660 6556
rect 19660 6500 19664 6556
rect 19600 6496 19664 6500
rect 19680 6556 19744 6560
rect 19680 6500 19684 6556
rect 19684 6500 19740 6556
rect 19740 6500 19744 6556
rect 19680 6496 19744 6500
rect 4360 6012 4424 6016
rect 4360 5956 4364 6012
rect 4364 5956 4420 6012
rect 4420 5956 4424 6012
rect 4360 5952 4424 5956
rect 4440 6012 4504 6016
rect 4440 5956 4444 6012
rect 4444 5956 4500 6012
rect 4500 5956 4504 6012
rect 4440 5952 4504 5956
rect 4520 6012 4584 6016
rect 4520 5956 4524 6012
rect 4524 5956 4580 6012
rect 4580 5956 4584 6012
rect 4520 5952 4584 5956
rect 4600 6012 4664 6016
rect 4600 5956 4604 6012
rect 4604 5956 4660 6012
rect 4660 5956 4664 6012
rect 4600 5952 4664 5956
rect 4680 6012 4744 6016
rect 4680 5956 4684 6012
rect 4684 5956 4740 6012
rect 4740 5956 4744 6012
rect 4680 5952 4744 5956
rect 10360 6012 10424 6016
rect 10360 5956 10364 6012
rect 10364 5956 10420 6012
rect 10420 5956 10424 6012
rect 10360 5952 10424 5956
rect 10440 6012 10504 6016
rect 10440 5956 10444 6012
rect 10444 5956 10500 6012
rect 10500 5956 10504 6012
rect 10440 5952 10504 5956
rect 10520 6012 10584 6016
rect 10520 5956 10524 6012
rect 10524 5956 10580 6012
rect 10580 5956 10584 6012
rect 10520 5952 10584 5956
rect 10600 6012 10664 6016
rect 10600 5956 10604 6012
rect 10604 5956 10660 6012
rect 10660 5956 10664 6012
rect 10600 5952 10664 5956
rect 10680 6012 10744 6016
rect 10680 5956 10684 6012
rect 10684 5956 10740 6012
rect 10740 5956 10744 6012
rect 10680 5952 10744 5956
rect 16360 6012 16424 6016
rect 16360 5956 16364 6012
rect 16364 5956 16420 6012
rect 16420 5956 16424 6012
rect 16360 5952 16424 5956
rect 16440 6012 16504 6016
rect 16440 5956 16444 6012
rect 16444 5956 16500 6012
rect 16500 5956 16504 6012
rect 16440 5952 16504 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 22360 6012 22424 6016
rect 22360 5956 22364 6012
rect 22364 5956 22420 6012
rect 22420 5956 22424 6012
rect 22360 5952 22424 5956
rect 22440 6012 22504 6016
rect 22440 5956 22444 6012
rect 22444 5956 22500 6012
rect 22500 5956 22504 6012
rect 22440 5952 22504 5956
rect 22520 6012 22584 6016
rect 22520 5956 22524 6012
rect 22524 5956 22580 6012
rect 22580 5956 22584 6012
rect 22520 5952 22584 5956
rect 22600 6012 22664 6016
rect 22600 5956 22604 6012
rect 22604 5956 22660 6012
rect 22660 5956 22664 6012
rect 22600 5952 22664 5956
rect 22680 6012 22744 6016
rect 22680 5956 22684 6012
rect 22684 5956 22740 6012
rect 22740 5956 22744 6012
rect 22680 5952 22744 5956
rect 14780 5808 14844 5812
rect 14780 5752 14794 5808
rect 14794 5752 14844 5808
rect 14780 5748 14844 5752
rect 20668 5612 20732 5676
rect 15148 5476 15212 5540
rect 16068 5476 16132 5540
rect 1360 5468 1424 5472
rect 1360 5412 1364 5468
rect 1364 5412 1420 5468
rect 1420 5412 1424 5468
rect 1360 5408 1424 5412
rect 1440 5468 1504 5472
rect 1440 5412 1444 5468
rect 1444 5412 1500 5468
rect 1500 5412 1504 5468
rect 1440 5408 1504 5412
rect 1520 5468 1584 5472
rect 1520 5412 1524 5468
rect 1524 5412 1580 5468
rect 1580 5412 1584 5468
rect 1520 5408 1584 5412
rect 1600 5468 1664 5472
rect 1600 5412 1604 5468
rect 1604 5412 1660 5468
rect 1660 5412 1664 5468
rect 1600 5408 1664 5412
rect 1680 5468 1744 5472
rect 1680 5412 1684 5468
rect 1684 5412 1740 5468
rect 1740 5412 1744 5468
rect 1680 5408 1744 5412
rect 7360 5468 7424 5472
rect 7360 5412 7364 5468
rect 7364 5412 7420 5468
rect 7420 5412 7424 5468
rect 7360 5408 7424 5412
rect 7440 5468 7504 5472
rect 7440 5412 7444 5468
rect 7444 5412 7500 5468
rect 7500 5412 7504 5468
rect 7440 5408 7504 5412
rect 7520 5468 7584 5472
rect 7520 5412 7524 5468
rect 7524 5412 7580 5468
rect 7580 5412 7584 5468
rect 7520 5408 7584 5412
rect 7600 5468 7664 5472
rect 7600 5412 7604 5468
rect 7604 5412 7660 5468
rect 7660 5412 7664 5468
rect 7600 5408 7664 5412
rect 7680 5468 7744 5472
rect 7680 5412 7684 5468
rect 7684 5412 7740 5468
rect 7740 5412 7744 5468
rect 7680 5408 7744 5412
rect 13360 5468 13424 5472
rect 13360 5412 13364 5468
rect 13364 5412 13420 5468
rect 13420 5412 13424 5468
rect 13360 5408 13424 5412
rect 13440 5468 13504 5472
rect 13440 5412 13444 5468
rect 13444 5412 13500 5468
rect 13500 5412 13504 5468
rect 13440 5408 13504 5412
rect 13520 5468 13584 5472
rect 13520 5412 13524 5468
rect 13524 5412 13580 5468
rect 13580 5412 13584 5468
rect 13520 5408 13584 5412
rect 13600 5468 13664 5472
rect 13600 5412 13604 5468
rect 13604 5412 13660 5468
rect 13660 5412 13664 5468
rect 13600 5408 13664 5412
rect 13680 5468 13744 5472
rect 13680 5412 13684 5468
rect 13684 5412 13740 5468
rect 13740 5412 13744 5468
rect 13680 5408 13744 5412
rect 19360 5468 19424 5472
rect 19360 5412 19364 5468
rect 19364 5412 19420 5468
rect 19420 5412 19424 5468
rect 19360 5408 19424 5412
rect 19440 5468 19504 5472
rect 19440 5412 19444 5468
rect 19444 5412 19500 5468
rect 19500 5412 19504 5468
rect 19440 5408 19504 5412
rect 19520 5468 19584 5472
rect 19520 5412 19524 5468
rect 19524 5412 19580 5468
rect 19580 5412 19584 5468
rect 19520 5408 19584 5412
rect 19600 5468 19664 5472
rect 19600 5412 19604 5468
rect 19604 5412 19660 5468
rect 19660 5412 19664 5468
rect 19600 5408 19664 5412
rect 19680 5468 19744 5472
rect 19680 5412 19684 5468
rect 19684 5412 19740 5468
rect 19740 5412 19744 5468
rect 19680 5408 19744 5412
rect 9996 5400 10060 5404
rect 9996 5344 10046 5400
rect 10046 5344 10060 5400
rect 9996 5340 10060 5344
rect 9812 5068 9876 5132
rect 4360 4924 4424 4928
rect 4360 4868 4364 4924
rect 4364 4868 4420 4924
rect 4420 4868 4424 4924
rect 4360 4864 4424 4868
rect 4440 4924 4504 4928
rect 4440 4868 4444 4924
rect 4444 4868 4500 4924
rect 4500 4868 4504 4924
rect 4440 4864 4504 4868
rect 4520 4924 4584 4928
rect 4520 4868 4524 4924
rect 4524 4868 4580 4924
rect 4580 4868 4584 4924
rect 4520 4864 4584 4868
rect 4600 4924 4664 4928
rect 4600 4868 4604 4924
rect 4604 4868 4660 4924
rect 4660 4868 4664 4924
rect 4600 4864 4664 4868
rect 4680 4924 4744 4928
rect 4680 4868 4684 4924
rect 4684 4868 4740 4924
rect 4740 4868 4744 4924
rect 4680 4864 4744 4868
rect 10360 4924 10424 4928
rect 10360 4868 10364 4924
rect 10364 4868 10420 4924
rect 10420 4868 10424 4924
rect 10360 4864 10424 4868
rect 10440 4924 10504 4928
rect 10440 4868 10444 4924
rect 10444 4868 10500 4924
rect 10500 4868 10504 4924
rect 10440 4864 10504 4868
rect 10520 4924 10584 4928
rect 10520 4868 10524 4924
rect 10524 4868 10580 4924
rect 10580 4868 10584 4924
rect 10520 4864 10584 4868
rect 10600 4924 10664 4928
rect 10600 4868 10604 4924
rect 10604 4868 10660 4924
rect 10660 4868 10664 4924
rect 10600 4864 10664 4868
rect 10680 4924 10744 4928
rect 10680 4868 10684 4924
rect 10684 4868 10740 4924
rect 10740 4868 10744 4924
rect 10680 4864 10744 4868
rect 16360 4924 16424 4928
rect 16360 4868 16364 4924
rect 16364 4868 16420 4924
rect 16420 4868 16424 4924
rect 16360 4864 16424 4868
rect 16440 4924 16504 4928
rect 16440 4868 16444 4924
rect 16444 4868 16500 4924
rect 16500 4868 16504 4924
rect 16440 4864 16504 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 22360 4924 22424 4928
rect 22360 4868 22364 4924
rect 22364 4868 22420 4924
rect 22420 4868 22424 4924
rect 22360 4864 22424 4868
rect 22440 4924 22504 4928
rect 22440 4868 22444 4924
rect 22444 4868 22500 4924
rect 22500 4868 22504 4924
rect 22440 4864 22504 4868
rect 22520 4924 22584 4928
rect 22520 4868 22524 4924
rect 22524 4868 22580 4924
rect 22580 4868 22584 4924
rect 22520 4864 22584 4868
rect 22600 4924 22664 4928
rect 22600 4868 22604 4924
rect 22604 4868 22660 4924
rect 22660 4868 22664 4924
rect 22600 4864 22664 4868
rect 22680 4924 22744 4928
rect 22680 4868 22684 4924
rect 22684 4868 22740 4924
rect 22740 4868 22744 4924
rect 22680 4864 22744 4868
rect 1360 4380 1424 4384
rect 1360 4324 1364 4380
rect 1364 4324 1420 4380
rect 1420 4324 1424 4380
rect 1360 4320 1424 4324
rect 1440 4380 1504 4384
rect 1440 4324 1444 4380
rect 1444 4324 1500 4380
rect 1500 4324 1504 4380
rect 1440 4320 1504 4324
rect 1520 4380 1584 4384
rect 1520 4324 1524 4380
rect 1524 4324 1580 4380
rect 1580 4324 1584 4380
rect 1520 4320 1584 4324
rect 1600 4380 1664 4384
rect 1600 4324 1604 4380
rect 1604 4324 1660 4380
rect 1660 4324 1664 4380
rect 1600 4320 1664 4324
rect 1680 4380 1744 4384
rect 1680 4324 1684 4380
rect 1684 4324 1740 4380
rect 1740 4324 1744 4380
rect 1680 4320 1744 4324
rect 7360 4380 7424 4384
rect 7360 4324 7364 4380
rect 7364 4324 7420 4380
rect 7420 4324 7424 4380
rect 7360 4320 7424 4324
rect 7440 4380 7504 4384
rect 7440 4324 7444 4380
rect 7444 4324 7500 4380
rect 7500 4324 7504 4380
rect 7440 4320 7504 4324
rect 7520 4380 7584 4384
rect 7520 4324 7524 4380
rect 7524 4324 7580 4380
rect 7580 4324 7584 4380
rect 7520 4320 7584 4324
rect 7600 4380 7664 4384
rect 7600 4324 7604 4380
rect 7604 4324 7660 4380
rect 7660 4324 7664 4380
rect 7600 4320 7664 4324
rect 7680 4380 7744 4384
rect 7680 4324 7684 4380
rect 7684 4324 7740 4380
rect 7740 4324 7744 4380
rect 7680 4320 7744 4324
rect 13360 4380 13424 4384
rect 13360 4324 13364 4380
rect 13364 4324 13420 4380
rect 13420 4324 13424 4380
rect 13360 4320 13424 4324
rect 13440 4380 13504 4384
rect 13440 4324 13444 4380
rect 13444 4324 13500 4380
rect 13500 4324 13504 4380
rect 13440 4320 13504 4324
rect 13520 4380 13584 4384
rect 13520 4324 13524 4380
rect 13524 4324 13580 4380
rect 13580 4324 13584 4380
rect 13520 4320 13584 4324
rect 13600 4380 13664 4384
rect 13600 4324 13604 4380
rect 13604 4324 13660 4380
rect 13660 4324 13664 4380
rect 13600 4320 13664 4324
rect 13680 4380 13744 4384
rect 13680 4324 13684 4380
rect 13684 4324 13740 4380
rect 13740 4324 13744 4380
rect 13680 4320 13744 4324
rect 19360 4380 19424 4384
rect 19360 4324 19364 4380
rect 19364 4324 19420 4380
rect 19420 4324 19424 4380
rect 19360 4320 19424 4324
rect 19440 4380 19504 4384
rect 19440 4324 19444 4380
rect 19444 4324 19500 4380
rect 19500 4324 19504 4380
rect 19440 4320 19504 4324
rect 19520 4380 19584 4384
rect 19520 4324 19524 4380
rect 19524 4324 19580 4380
rect 19580 4324 19584 4380
rect 19520 4320 19584 4324
rect 19600 4380 19664 4384
rect 19600 4324 19604 4380
rect 19604 4324 19660 4380
rect 19660 4324 19664 4380
rect 19600 4320 19664 4324
rect 19680 4380 19744 4384
rect 19680 4324 19684 4380
rect 19684 4324 19740 4380
rect 19740 4324 19744 4380
rect 19680 4320 19744 4324
rect 9444 3844 9508 3908
rect 4360 3836 4424 3840
rect 4360 3780 4364 3836
rect 4364 3780 4420 3836
rect 4420 3780 4424 3836
rect 4360 3776 4424 3780
rect 4440 3836 4504 3840
rect 4440 3780 4444 3836
rect 4444 3780 4500 3836
rect 4500 3780 4504 3836
rect 4440 3776 4504 3780
rect 4520 3836 4584 3840
rect 4520 3780 4524 3836
rect 4524 3780 4580 3836
rect 4580 3780 4584 3836
rect 4520 3776 4584 3780
rect 4600 3836 4664 3840
rect 4600 3780 4604 3836
rect 4604 3780 4660 3836
rect 4660 3780 4664 3836
rect 4600 3776 4664 3780
rect 4680 3836 4744 3840
rect 4680 3780 4684 3836
rect 4684 3780 4740 3836
rect 4740 3780 4744 3836
rect 4680 3776 4744 3780
rect 10360 3836 10424 3840
rect 10360 3780 10364 3836
rect 10364 3780 10420 3836
rect 10420 3780 10424 3836
rect 10360 3776 10424 3780
rect 10440 3836 10504 3840
rect 10440 3780 10444 3836
rect 10444 3780 10500 3836
rect 10500 3780 10504 3836
rect 10440 3776 10504 3780
rect 10520 3836 10584 3840
rect 10520 3780 10524 3836
rect 10524 3780 10580 3836
rect 10580 3780 10584 3836
rect 10520 3776 10584 3780
rect 10600 3836 10664 3840
rect 10600 3780 10604 3836
rect 10604 3780 10660 3836
rect 10660 3780 10664 3836
rect 10600 3776 10664 3780
rect 10680 3836 10744 3840
rect 10680 3780 10684 3836
rect 10684 3780 10740 3836
rect 10740 3780 10744 3836
rect 10680 3776 10744 3780
rect 16360 3836 16424 3840
rect 16360 3780 16364 3836
rect 16364 3780 16420 3836
rect 16420 3780 16424 3836
rect 16360 3776 16424 3780
rect 16440 3836 16504 3840
rect 16440 3780 16444 3836
rect 16444 3780 16500 3836
rect 16500 3780 16504 3836
rect 16440 3776 16504 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 22360 3836 22424 3840
rect 22360 3780 22364 3836
rect 22364 3780 22420 3836
rect 22420 3780 22424 3836
rect 22360 3776 22424 3780
rect 22440 3836 22504 3840
rect 22440 3780 22444 3836
rect 22444 3780 22500 3836
rect 22500 3780 22504 3836
rect 22440 3776 22504 3780
rect 22520 3836 22584 3840
rect 22520 3780 22524 3836
rect 22524 3780 22580 3836
rect 22580 3780 22584 3836
rect 22520 3776 22584 3780
rect 22600 3836 22664 3840
rect 22600 3780 22604 3836
rect 22604 3780 22660 3836
rect 22660 3780 22664 3836
rect 22600 3776 22664 3780
rect 22680 3836 22744 3840
rect 22680 3780 22684 3836
rect 22684 3780 22740 3836
rect 22740 3780 22744 3836
rect 22680 3776 22744 3780
rect 9812 3708 9876 3772
rect 9076 3300 9140 3364
rect 11100 3360 11164 3364
rect 11100 3304 11114 3360
rect 11114 3304 11164 3360
rect 11100 3300 11164 3304
rect 1360 3292 1424 3296
rect 1360 3236 1364 3292
rect 1364 3236 1420 3292
rect 1420 3236 1424 3292
rect 1360 3232 1424 3236
rect 1440 3292 1504 3296
rect 1440 3236 1444 3292
rect 1444 3236 1500 3292
rect 1500 3236 1504 3292
rect 1440 3232 1504 3236
rect 1520 3292 1584 3296
rect 1520 3236 1524 3292
rect 1524 3236 1580 3292
rect 1580 3236 1584 3292
rect 1520 3232 1584 3236
rect 1600 3292 1664 3296
rect 1600 3236 1604 3292
rect 1604 3236 1660 3292
rect 1660 3236 1664 3292
rect 1600 3232 1664 3236
rect 1680 3292 1744 3296
rect 1680 3236 1684 3292
rect 1684 3236 1740 3292
rect 1740 3236 1744 3292
rect 1680 3232 1744 3236
rect 7360 3292 7424 3296
rect 7360 3236 7364 3292
rect 7364 3236 7420 3292
rect 7420 3236 7424 3292
rect 7360 3232 7424 3236
rect 7440 3292 7504 3296
rect 7440 3236 7444 3292
rect 7444 3236 7500 3292
rect 7500 3236 7504 3292
rect 7440 3232 7504 3236
rect 7520 3292 7584 3296
rect 7520 3236 7524 3292
rect 7524 3236 7580 3292
rect 7580 3236 7584 3292
rect 7520 3232 7584 3236
rect 7600 3292 7664 3296
rect 7600 3236 7604 3292
rect 7604 3236 7660 3292
rect 7660 3236 7664 3292
rect 7600 3232 7664 3236
rect 7680 3292 7744 3296
rect 7680 3236 7684 3292
rect 7684 3236 7740 3292
rect 7740 3236 7744 3292
rect 7680 3232 7744 3236
rect 13360 3292 13424 3296
rect 13360 3236 13364 3292
rect 13364 3236 13420 3292
rect 13420 3236 13424 3292
rect 13360 3232 13424 3236
rect 13440 3292 13504 3296
rect 13440 3236 13444 3292
rect 13444 3236 13500 3292
rect 13500 3236 13504 3292
rect 13440 3232 13504 3236
rect 13520 3292 13584 3296
rect 13520 3236 13524 3292
rect 13524 3236 13580 3292
rect 13580 3236 13584 3292
rect 13520 3232 13584 3236
rect 13600 3292 13664 3296
rect 13600 3236 13604 3292
rect 13604 3236 13660 3292
rect 13660 3236 13664 3292
rect 13600 3232 13664 3236
rect 13680 3292 13744 3296
rect 13680 3236 13684 3292
rect 13684 3236 13740 3292
rect 13740 3236 13744 3292
rect 13680 3232 13744 3236
rect 19360 3292 19424 3296
rect 19360 3236 19364 3292
rect 19364 3236 19420 3292
rect 19420 3236 19424 3292
rect 19360 3232 19424 3236
rect 19440 3292 19504 3296
rect 19440 3236 19444 3292
rect 19444 3236 19500 3292
rect 19500 3236 19504 3292
rect 19440 3232 19504 3236
rect 19520 3292 19584 3296
rect 19520 3236 19524 3292
rect 19524 3236 19580 3292
rect 19580 3236 19584 3292
rect 19520 3232 19584 3236
rect 19600 3292 19664 3296
rect 19600 3236 19604 3292
rect 19604 3236 19660 3292
rect 19660 3236 19664 3292
rect 19600 3232 19664 3236
rect 19680 3292 19744 3296
rect 19680 3236 19684 3292
rect 19684 3236 19740 3292
rect 19740 3236 19744 3292
rect 19680 3232 19744 3236
rect 9260 3028 9324 3092
rect 9812 2816 9876 2820
rect 9812 2760 9826 2816
rect 9826 2760 9876 2816
rect 9812 2756 9876 2760
rect 4360 2748 4424 2752
rect 4360 2692 4364 2748
rect 4364 2692 4420 2748
rect 4420 2692 4424 2748
rect 4360 2688 4424 2692
rect 4440 2748 4504 2752
rect 4440 2692 4444 2748
rect 4444 2692 4500 2748
rect 4500 2692 4504 2748
rect 4440 2688 4504 2692
rect 4520 2748 4584 2752
rect 4520 2692 4524 2748
rect 4524 2692 4580 2748
rect 4580 2692 4584 2748
rect 4520 2688 4584 2692
rect 4600 2748 4664 2752
rect 4600 2692 4604 2748
rect 4604 2692 4660 2748
rect 4660 2692 4664 2748
rect 4600 2688 4664 2692
rect 4680 2748 4744 2752
rect 4680 2692 4684 2748
rect 4684 2692 4740 2748
rect 4740 2692 4744 2748
rect 4680 2688 4744 2692
rect 10360 2748 10424 2752
rect 10360 2692 10364 2748
rect 10364 2692 10420 2748
rect 10420 2692 10424 2748
rect 10360 2688 10424 2692
rect 10440 2748 10504 2752
rect 10440 2692 10444 2748
rect 10444 2692 10500 2748
rect 10500 2692 10504 2748
rect 10440 2688 10504 2692
rect 10520 2748 10584 2752
rect 10520 2692 10524 2748
rect 10524 2692 10580 2748
rect 10580 2692 10584 2748
rect 10520 2688 10584 2692
rect 10600 2748 10664 2752
rect 10600 2692 10604 2748
rect 10604 2692 10660 2748
rect 10660 2692 10664 2748
rect 10600 2688 10664 2692
rect 10680 2748 10744 2752
rect 10680 2692 10684 2748
rect 10684 2692 10740 2748
rect 10740 2692 10744 2748
rect 10680 2688 10744 2692
rect 16360 2748 16424 2752
rect 16360 2692 16364 2748
rect 16364 2692 16420 2748
rect 16420 2692 16424 2748
rect 16360 2688 16424 2692
rect 16440 2748 16504 2752
rect 16440 2692 16444 2748
rect 16444 2692 16500 2748
rect 16500 2692 16504 2748
rect 16440 2688 16504 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 22360 2748 22424 2752
rect 22360 2692 22364 2748
rect 22364 2692 22420 2748
rect 22420 2692 22424 2748
rect 22360 2688 22424 2692
rect 22440 2748 22504 2752
rect 22440 2692 22444 2748
rect 22444 2692 22500 2748
rect 22500 2692 22504 2748
rect 22440 2688 22504 2692
rect 22520 2748 22584 2752
rect 22520 2692 22524 2748
rect 22524 2692 22580 2748
rect 22580 2692 22584 2748
rect 22520 2688 22584 2692
rect 22600 2748 22664 2752
rect 22600 2692 22604 2748
rect 22604 2692 22660 2748
rect 22660 2692 22664 2748
rect 22600 2688 22664 2692
rect 22680 2748 22744 2752
rect 22680 2692 22684 2748
rect 22684 2692 22740 2748
rect 22740 2692 22744 2748
rect 22680 2688 22744 2692
rect 9076 2620 9140 2684
rect 13124 2620 13188 2684
rect 20668 2620 20732 2684
rect 9260 2348 9324 2412
rect 1360 2204 1424 2208
rect 1360 2148 1364 2204
rect 1364 2148 1420 2204
rect 1420 2148 1424 2204
rect 1360 2144 1424 2148
rect 1440 2204 1504 2208
rect 1440 2148 1444 2204
rect 1444 2148 1500 2204
rect 1500 2148 1504 2204
rect 1440 2144 1504 2148
rect 1520 2204 1584 2208
rect 1520 2148 1524 2204
rect 1524 2148 1580 2204
rect 1580 2148 1584 2204
rect 1520 2144 1584 2148
rect 1600 2204 1664 2208
rect 1600 2148 1604 2204
rect 1604 2148 1660 2204
rect 1660 2148 1664 2204
rect 1600 2144 1664 2148
rect 1680 2204 1744 2208
rect 1680 2148 1684 2204
rect 1684 2148 1740 2204
rect 1740 2148 1744 2204
rect 1680 2144 1744 2148
rect 7360 2204 7424 2208
rect 7360 2148 7364 2204
rect 7364 2148 7420 2204
rect 7420 2148 7424 2204
rect 7360 2144 7424 2148
rect 7440 2204 7504 2208
rect 7440 2148 7444 2204
rect 7444 2148 7500 2204
rect 7500 2148 7504 2204
rect 7440 2144 7504 2148
rect 7520 2204 7584 2208
rect 7520 2148 7524 2204
rect 7524 2148 7580 2204
rect 7580 2148 7584 2204
rect 7520 2144 7584 2148
rect 7600 2204 7664 2208
rect 7600 2148 7604 2204
rect 7604 2148 7660 2204
rect 7660 2148 7664 2204
rect 7600 2144 7664 2148
rect 7680 2204 7744 2208
rect 7680 2148 7684 2204
rect 7684 2148 7740 2204
rect 7740 2148 7744 2204
rect 7680 2144 7744 2148
rect 13360 2204 13424 2208
rect 13360 2148 13364 2204
rect 13364 2148 13420 2204
rect 13420 2148 13424 2204
rect 13360 2144 13424 2148
rect 13440 2204 13504 2208
rect 13440 2148 13444 2204
rect 13444 2148 13500 2204
rect 13500 2148 13504 2204
rect 13440 2144 13504 2148
rect 13520 2204 13584 2208
rect 13520 2148 13524 2204
rect 13524 2148 13580 2204
rect 13580 2148 13584 2204
rect 13520 2144 13584 2148
rect 13600 2204 13664 2208
rect 13600 2148 13604 2204
rect 13604 2148 13660 2204
rect 13660 2148 13664 2204
rect 13600 2144 13664 2148
rect 13680 2204 13744 2208
rect 13680 2148 13684 2204
rect 13684 2148 13740 2204
rect 13740 2148 13744 2204
rect 13680 2144 13744 2148
rect 19360 2204 19424 2208
rect 19360 2148 19364 2204
rect 19364 2148 19420 2204
rect 19420 2148 19424 2204
rect 19360 2144 19424 2148
rect 19440 2204 19504 2208
rect 19440 2148 19444 2204
rect 19444 2148 19500 2204
rect 19500 2148 19504 2204
rect 19440 2144 19504 2148
rect 19520 2204 19584 2208
rect 19520 2148 19524 2204
rect 19524 2148 19580 2204
rect 19580 2148 19584 2204
rect 19520 2144 19584 2148
rect 19600 2204 19664 2208
rect 19600 2148 19604 2204
rect 19604 2148 19660 2204
rect 19660 2148 19664 2204
rect 19600 2144 19664 2148
rect 19680 2204 19744 2208
rect 19680 2148 19684 2204
rect 19684 2148 19740 2204
rect 19740 2148 19744 2204
rect 19680 2144 19744 2148
rect 14964 2136 15028 2140
rect 14964 2080 14978 2136
rect 14978 2080 15028 2136
rect 14964 2076 15028 2080
rect 9444 1728 9508 1732
rect 9444 1672 9494 1728
rect 9494 1672 9508 1728
rect 9444 1668 9508 1672
rect 4360 1660 4424 1664
rect 4360 1604 4364 1660
rect 4364 1604 4420 1660
rect 4420 1604 4424 1660
rect 4360 1600 4424 1604
rect 4440 1660 4504 1664
rect 4440 1604 4444 1660
rect 4444 1604 4500 1660
rect 4500 1604 4504 1660
rect 4440 1600 4504 1604
rect 4520 1660 4584 1664
rect 4520 1604 4524 1660
rect 4524 1604 4580 1660
rect 4580 1604 4584 1660
rect 4520 1600 4584 1604
rect 4600 1660 4664 1664
rect 4600 1604 4604 1660
rect 4604 1604 4660 1660
rect 4660 1604 4664 1660
rect 4600 1600 4664 1604
rect 4680 1660 4744 1664
rect 4680 1604 4684 1660
rect 4684 1604 4740 1660
rect 4740 1604 4744 1660
rect 4680 1600 4744 1604
rect 10360 1660 10424 1664
rect 10360 1604 10364 1660
rect 10364 1604 10420 1660
rect 10420 1604 10424 1660
rect 10360 1600 10424 1604
rect 10440 1660 10504 1664
rect 10440 1604 10444 1660
rect 10444 1604 10500 1660
rect 10500 1604 10504 1660
rect 10440 1600 10504 1604
rect 10520 1660 10584 1664
rect 10520 1604 10524 1660
rect 10524 1604 10580 1660
rect 10580 1604 10584 1660
rect 10520 1600 10584 1604
rect 10600 1660 10664 1664
rect 10600 1604 10604 1660
rect 10604 1604 10660 1660
rect 10660 1604 10664 1660
rect 10600 1600 10664 1604
rect 10680 1660 10744 1664
rect 10680 1604 10684 1660
rect 10684 1604 10740 1660
rect 10740 1604 10744 1660
rect 10680 1600 10744 1604
rect 16360 1660 16424 1664
rect 16360 1604 16364 1660
rect 16364 1604 16420 1660
rect 16420 1604 16424 1660
rect 16360 1600 16424 1604
rect 16440 1660 16504 1664
rect 16440 1604 16444 1660
rect 16444 1604 16500 1660
rect 16500 1604 16504 1660
rect 16440 1600 16504 1604
rect 16520 1660 16584 1664
rect 16520 1604 16524 1660
rect 16524 1604 16580 1660
rect 16580 1604 16584 1660
rect 16520 1600 16584 1604
rect 16600 1660 16664 1664
rect 16600 1604 16604 1660
rect 16604 1604 16660 1660
rect 16660 1604 16664 1660
rect 16600 1600 16664 1604
rect 16680 1660 16744 1664
rect 16680 1604 16684 1660
rect 16684 1604 16740 1660
rect 16740 1604 16744 1660
rect 16680 1600 16744 1604
rect 22360 1660 22424 1664
rect 22360 1604 22364 1660
rect 22364 1604 22420 1660
rect 22420 1604 22424 1660
rect 22360 1600 22424 1604
rect 22440 1660 22504 1664
rect 22440 1604 22444 1660
rect 22444 1604 22500 1660
rect 22500 1604 22504 1660
rect 22440 1600 22504 1604
rect 22520 1660 22584 1664
rect 22520 1604 22524 1660
rect 22524 1604 22580 1660
rect 22580 1604 22584 1660
rect 22520 1600 22584 1604
rect 22600 1660 22664 1664
rect 22600 1604 22604 1660
rect 22604 1604 22660 1660
rect 22660 1604 22664 1660
rect 22600 1600 22664 1604
rect 22680 1660 22744 1664
rect 22680 1604 22684 1660
rect 22684 1604 22740 1660
rect 22740 1604 22744 1660
rect 22680 1600 22744 1604
rect 16068 1396 16132 1460
rect 1360 1116 1424 1120
rect 1360 1060 1364 1116
rect 1364 1060 1420 1116
rect 1420 1060 1424 1116
rect 1360 1056 1424 1060
rect 1440 1116 1504 1120
rect 1440 1060 1444 1116
rect 1444 1060 1500 1116
rect 1500 1060 1504 1116
rect 1440 1056 1504 1060
rect 1520 1116 1584 1120
rect 1520 1060 1524 1116
rect 1524 1060 1580 1116
rect 1580 1060 1584 1116
rect 1520 1056 1584 1060
rect 1600 1116 1664 1120
rect 1600 1060 1604 1116
rect 1604 1060 1660 1116
rect 1660 1060 1664 1116
rect 1600 1056 1664 1060
rect 1680 1116 1744 1120
rect 1680 1060 1684 1116
rect 1684 1060 1740 1116
rect 1740 1060 1744 1116
rect 1680 1056 1744 1060
rect 7360 1116 7424 1120
rect 7360 1060 7364 1116
rect 7364 1060 7420 1116
rect 7420 1060 7424 1116
rect 7360 1056 7424 1060
rect 7440 1116 7504 1120
rect 7440 1060 7444 1116
rect 7444 1060 7500 1116
rect 7500 1060 7504 1116
rect 7440 1056 7504 1060
rect 7520 1116 7584 1120
rect 7520 1060 7524 1116
rect 7524 1060 7580 1116
rect 7580 1060 7584 1116
rect 7520 1056 7584 1060
rect 7600 1116 7664 1120
rect 7600 1060 7604 1116
rect 7604 1060 7660 1116
rect 7660 1060 7664 1116
rect 7600 1056 7664 1060
rect 7680 1116 7744 1120
rect 7680 1060 7684 1116
rect 7684 1060 7740 1116
rect 7740 1060 7744 1116
rect 7680 1056 7744 1060
rect 13360 1116 13424 1120
rect 13360 1060 13364 1116
rect 13364 1060 13420 1116
rect 13420 1060 13424 1116
rect 13360 1056 13424 1060
rect 13440 1116 13504 1120
rect 13440 1060 13444 1116
rect 13444 1060 13500 1116
rect 13500 1060 13504 1116
rect 13440 1056 13504 1060
rect 13520 1116 13584 1120
rect 13520 1060 13524 1116
rect 13524 1060 13580 1116
rect 13580 1060 13584 1116
rect 13520 1056 13584 1060
rect 13600 1116 13664 1120
rect 13600 1060 13604 1116
rect 13604 1060 13660 1116
rect 13660 1060 13664 1116
rect 13600 1056 13664 1060
rect 13680 1116 13744 1120
rect 13680 1060 13684 1116
rect 13684 1060 13740 1116
rect 13740 1060 13744 1116
rect 13680 1056 13744 1060
rect 19360 1116 19424 1120
rect 19360 1060 19364 1116
rect 19364 1060 19420 1116
rect 19420 1060 19424 1116
rect 19360 1056 19424 1060
rect 19440 1116 19504 1120
rect 19440 1060 19444 1116
rect 19444 1060 19500 1116
rect 19500 1060 19504 1116
rect 19440 1056 19504 1060
rect 19520 1116 19584 1120
rect 19520 1060 19524 1116
rect 19524 1060 19580 1116
rect 19580 1060 19584 1116
rect 19520 1056 19584 1060
rect 19600 1116 19664 1120
rect 19600 1060 19604 1116
rect 19604 1060 19660 1116
rect 19660 1060 19664 1116
rect 19600 1056 19664 1060
rect 19680 1116 19744 1120
rect 19680 1060 19684 1116
rect 19684 1060 19740 1116
rect 19740 1060 19744 1116
rect 19680 1056 19744 1060
rect 9996 852 10060 916
rect 4360 572 4424 576
rect 4360 516 4364 572
rect 4364 516 4420 572
rect 4420 516 4424 572
rect 4360 512 4424 516
rect 4440 572 4504 576
rect 4440 516 4444 572
rect 4444 516 4500 572
rect 4500 516 4504 572
rect 4440 512 4504 516
rect 4520 572 4584 576
rect 4520 516 4524 572
rect 4524 516 4580 572
rect 4580 516 4584 572
rect 4520 512 4584 516
rect 4600 572 4664 576
rect 4600 516 4604 572
rect 4604 516 4660 572
rect 4660 516 4664 572
rect 4600 512 4664 516
rect 4680 572 4744 576
rect 4680 516 4684 572
rect 4684 516 4740 572
rect 4740 516 4744 572
rect 4680 512 4744 516
rect 10360 572 10424 576
rect 10360 516 10364 572
rect 10364 516 10420 572
rect 10420 516 10424 572
rect 10360 512 10424 516
rect 10440 572 10504 576
rect 10440 516 10444 572
rect 10444 516 10500 572
rect 10500 516 10504 572
rect 10440 512 10504 516
rect 10520 572 10584 576
rect 10520 516 10524 572
rect 10524 516 10580 572
rect 10580 516 10584 572
rect 10520 512 10584 516
rect 10600 572 10664 576
rect 10600 516 10604 572
rect 10604 516 10660 572
rect 10660 516 10664 572
rect 10600 512 10664 516
rect 10680 572 10744 576
rect 10680 516 10684 572
rect 10684 516 10740 572
rect 10740 516 10744 572
rect 10680 512 10744 516
rect 16360 572 16424 576
rect 16360 516 16364 572
rect 16364 516 16420 572
rect 16420 516 16424 572
rect 16360 512 16424 516
rect 16440 572 16504 576
rect 16440 516 16444 572
rect 16444 516 16500 572
rect 16500 516 16504 572
rect 16440 512 16504 516
rect 16520 572 16584 576
rect 16520 516 16524 572
rect 16524 516 16580 572
rect 16580 516 16584 572
rect 16520 512 16584 516
rect 16600 572 16664 576
rect 16600 516 16604 572
rect 16604 516 16660 572
rect 16660 516 16664 572
rect 16600 512 16664 516
rect 16680 572 16744 576
rect 16680 516 16684 572
rect 16684 516 16740 572
rect 16740 516 16744 572
rect 16680 512 16744 516
rect 22360 572 22424 576
rect 22360 516 22364 572
rect 22364 516 22420 572
rect 22420 516 22424 572
rect 22360 512 22424 516
rect 22440 572 22504 576
rect 22440 516 22444 572
rect 22444 516 22500 572
rect 22500 516 22504 572
rect 22440 512 22504 516
rect 22520 572 22584 576
rect 22520 516 22524 572
rect 22524 516 22580 572
rect 22580 516 22584 572
rect 22520 512 22584 516
rect 22600 572 22664 576
rect 22600 516 22604 572
rect 22604 516 22660 572
rect 22660 516 22664 572
rect 22600 512 22664 516
rect 22680 572 22744 576
rect 22680 516 22684 572
rect 22684 516 22740 572
rect 22740 516 22744 572
rect 22680 512 22744 516
<< metal4 >>
rect 1352 15264 1752 15280
rect 1352 15200 1360 15264
rect 1424 15200 1440 15264
rect 1504 15200 1520 15264
rect 1584 15200 1600 15264
rect 1664 15200 1680 15264
rect 1744 15200 1752 15264
rect 1352 14176 1752 15200
rect 1352 14112 1360 14176
rect 1424 14112 1440 14176
rect 1504 14112 1520 14176
rect 1584 14112 1600 14176
rect 1664 14112 1680 14176
rect 1744 14112 1752 14176
rect 1352 13088 1752 14112
rect 1352 13024 1360 13088
rect 1424 13024 1440 13088
rect 1504 13024 1520 13088
rect 1584 13024 1600 13088
rect 1664 13024 1680 13088
rect 1744 13024 1752 13088
rect 1352 12000 1752 13024
rect 1352 11936 1360 12000
rect 1424 11936 1440 12000
rect 1504 11936 1520 12000
rect 1584 11936 1600 12000
rect 1664 11936 1680 12000
rect 1744 11936 1752 12000
rect 1352 10912 1752 11936
rect 4352 14720 4752 15280
rect 4352 14656 4360 14720
rect 4424 14656 4440 14720
rect 4504 14656 4520 14720
rect 4584 14656 4600 14720
rect 4664 14656 4680 14720
rect 4744 14656 4752 14720
rect 4352 13632 4752 14656
rect 4352 13568 4360 13632
rect 4424 13568 4440 13632
rect 4504 13568 4520 13632
rect 4584 13568 4600 13632
rect 4664 13568 4680 13632
rect 4744 13568 4752 13632
rect 4352 12544 4752 13568
rect 4352 12480 4360 12544
rect 4424 12480 4440 12544
rect 4504 12480 4520 12544
rect 4584 12480 4600 12544
rect 4664 12480 4680 12544
rect 4744 12480 4752 12544
rect 4107 11524 4173 11525
rect 4107 11460 4108 11524
rect 4172 11460 4173 11524
rect 4107 11459 4173 11460
rect 1352 10848 1360 10912
rect 1424 10848 1440 10912
rect 1504 10848 1520 10912
rect 1584 10848 1600 10912
rect 1664 10848 1680 10912
rect 1744 10848 1752 10912
rect 1352 9824 1752 10848
rect 1352 9760 1360 9824
rect 1424 9760 1440 9824
rect 1504 9760 1520 9824
rect 1584 9760 1600 9824
rect 1664 9760 1680 9824
rect 1744 9760 1752 9824
rect 1352 8736 1752 9760
rect 1352 8672 1360 8736
rect 1424 8672 1440 8736
rect 1504 8672 1520 8736
rect 1584 8672 1600 8736
rect 1664 8672 1680 8736
rect 1744 8672 1752 8736
rect 1352 7648 1752 8672
rect 4110 7853 4170 11459
rect 4352 11456 4752 12480
rect 4352 11392 4360 11456
rect 4424 11392 4440 11456
rect 4504 11392 4520 11456
rect 4584 11392 4600 11456
rect 4664 11392 4680 11456
rect 4744 11392 4752 11456
rect 4352 10368 4752 11392
rect 4352 10304 4360 10368
rect 4424 10304 4440 10368
rect 4504 10304 4520 10368
rect 4584 10304 4600 10368
rect 4664 10304 4680 10368
rect 4744 10304 4752 10368
rect 4352 9280 4752 10304
rect 4352 9216 4360 9280
rect 4424 9216 4440 9280
rect 4504 9216 4520 9280
rect 4584 9216 4600 9280
rect 4664 9216 4680 9280
rect 4744 9216 4752 9280
rect 4352 8192 4752 9216
rect 4352 8128 4360 8192
rect 4424 8128 4440 8192
rect 4504 8128 4520 8192
rect 4584 8128 4600 8192
rect 4664 8128 4680 8192
rect 4744 8128 4752 8192
rect 4107 7852 4173 7853
rect 4107 7788 4108 7852
rect 4172 7788 4173 7852
rect 4107 7787 4173 7788
rect 1352 7584 1360 7648
rect 1424 7584 1440 7648
rect 1504 7584 1520 7648
rect 1584 7584 1600 7648
rect 1664 7584 1680 7648
rect 1744 7584 1752 7648
rect 1352 6560 1752 7584
rect 1352 6496 1360 6560
rect 1424 6496 1440 6560
rect 1504 6496 1520 6560
rect 1584 6496 1600 6560
rect 1664 6496 1680 6560
rect 1744 6496 1752 6560
rect 1352 5472 1752 6496
rect 1352 5408 1360 5472
rect 1424 5408 1440 5472
rect 1504 5408 1520 5472
rect 1584 5408 1600 5472
rect 1664 5408 1680 5472
rect 1744 5408 1752 5472
rect 1352 4384 1752 5408
rect 1352 4320 1360 4384
rect 1424 4320 1440 4384
rect 1504 4320 1520 4384
rect 1584 4320 1600 4384
rect 1664 4320 1680 4384
rect 1744 4320 1752 4384
rect 1352 3296 1752 4320
rect 1352 3232 1360 3296
rect 1424 3232 1440 3296
rect 1504 3232 1520 3296
rect 1584 3232 1600 3296
rect 1664 3232 1680 3296
rect 1744 3232 1752 3296
rect 1352 2208 1752 3232
rect 1352 2144 1360 2208
rect 1424 2144 1440 2208
rect 1504 2144 1520 2208
rect 1584 2144 1600 2208
rect 1664 2144 1680 2208
rect 1744 2144 1752 2208
rect 1352 1120 1752 2144
rect 1352 1056 1360 1120
rect 1424 1056 1440 1120
rect 1504 1056 1520 1120
rect 1584 1056 1600 1120
rect 1664 1056 1680 1120
rect 1744 1056 1752 1120
rect 1352 496 1752 1056
rect 4352 7104 4752 8128
rect 4352 7040 4360 7104
rect 4424 7040 4440 7104
rect 4504 7040 4520 7104
rect 4584 7040 4600 7104
rect 4664 7040 4680 7104
rect 4744 7040 4752 7104
rect 4352 6016 4752 7040
rect 4352 5952 4360 6016
rect 4424 5952 4440 6016
rect 4504 5952 4520 6016
rect 4584 5952 4600 6016
rect 4664 5952 4680 6016
rect 4744 5952 4752 6016
rect 4352 4928 4752 5952
rect 4352 4864 4360 4928
rect 4424 4864 4440 4928
rect 4504 4864 4520 4928
rect 4584 4864 4600 4928
rect 4664 4864 4680 4928
rect 4744 4864 4752 4928
rect 4352 3840 4752 4864
rect 4352 3776 4360 3840
rect 4424 3776 4440 3840
rect 4504 3776 4520 3840
rect 4584 3776 4600 3840
rect 4664 3776 4680 3840
rect 4744 3776 4752 3840
rect 4352 2752 4752 3776
rect 4352 2688 4360 2752
rect 4424 2688 4440 2752
rect 4504 2688 4520 2752
rect 4584 2688 4600 2752
rect 4664 2688 4680 2752
rect 4744 2688 4752 2752
rect 4352 1664 4752 2688
rect 4352 1600 4360 1664
rect 4424 1600 4440 1664
rect 4504 1600 4520 1664
rect 4584 1600 4600 1664
rect 4664 1600 4680 1664
rect 4744 1600 4752 1664
rect 4352 576 4752 1600
rect 4352 512 4360 576
rect 4424 512 4440 576
rect 4504 512 4520 576
rect 4584 512 4600 576
rect 4664 512 4680 576
rect 4744 512 4752 576
rect 4352 496 4752 512
rect 7352 15264 7752 15280
rect 7352 15200 7360 15264
rect 7424 15200 7440 15264
rect 7504 15200 7520 15264
rect 7584 15200 7600 15264
rect 7664 15200 7680 15264
rect 7744 15200 7752 15264
rect 7352 14176 7752 15200
rect 7352 14112 7360 14176
rect 7424 14112 7440 14176
rect 7504 14112 7520 14176
rect 7584 14112 7600 14176
rect 7664 14112 7680 14176
rect 7744 14112 7752 14176
rect 7352 13088 7752 14112
rect 7352 13024 7360 13088
rect 7424 13024 7440 13088
rect 7504 13024 7520 13088
rect 7584 13024 7600 13088
rect 7664 13024 7680 13088
rect 7744 13024 7752 13088
rect 7352 12000 7752 13024
rect 7352 11936 7360 12000
rect 7424 11936 7440 12000
rect 7504 11936 7520 12000
rect 7584 11936 7600 12000
rect 7664 11936 7680 12000
rect 7744 11936 7752 12000
rect 7352 10912 7752 11936
rect 7352 10848 7360 10912
rect 7424 10848 7440 10912
rect 7504 10848 7520 10912
rect 7584 10848 7600 10912
rect 7664 10848 7680 10912
rect 7744 10848 7752 10912
rect 7352 9824 7752 10848
rect 7352 9760 7360 9824
rect 7424 9760 7440 9824
rect 7504 9760 7520 9824
rect 7584 9760 7600 9824
rect 7664 9760 7680 9824
rect 7744 9760 7752 9824
rect 7352 8736 7752 9760
rect 10352 14720 10752 15280
rect 10352 14656 10360 14720
rect 10424 14656 10440 14720
rect 10504 14656 10520 14720
rect 10584 14656 10600 14720
rect 10664 14656 10680 14720
rect 10744 14656 10752 14720
rect 10352 13632 10752 14656
rect 10352 13568 10360 13632
rect 10424 13568 10440 13632
rect 10504 13568 10520 13632
rect 10584 13568 10600 13632
rect 10664 13568 10680 13632
rect 10744 13568 10752 13632
rect 10352 12544 10752 13568
rect 13352 15264 13752 15280
rect 13352 15200 13360 15264
rect 13424 15200 13440 15264
rect 13504 15200 13520 15264
rect 13584 15200 13600 15264
rect 13664 15200 13680 15264
rect 13744 15200 13752 15264
rect 13352 14176 13752 15200
rect 13352 14112 13360 14176
rect 13424 14112 13440 14176
rect 13504 14112 13520 14176
rect 13584 14112 13600 14176
rect 13664 14112 13680 14176
rect 13744 14112 13752 14176
rect 13123 13428 13189 13429
rect 13123 13364 13124 13428
rect 13188 13364 13189 13428
rect 13123 13363 13189 13364
rect 10352 12480 10360 12544
rect 10424 12480 10440 12544
rect 10504 12480 10520 12544
rect 10584 12480 10600 12544
rect 10664 12480 10680 12544
rect 10744 12480 10752 12544
rect 10352 11456 10752 12480
rect 10352 11392 10360 11456
rect 10424 11392 10440 11456
rect 10504 11392 10520 11456
rect 10584 11392 10600 11456
rect 10664 11392 10680 11456
rect 10744 11392 10752 11456
rect 10352 10368 10752 11392
rect 10352 10304 10360 10368
rect 10424 10304 10440 10368
rect 10504 10304 10520 10368
rect 10584 10304 10600 10368
rect 10664 10304 10680 10368
rect 10744 10304 10752 10368
rect 9811 9756 9877 9757
rect 9811 9692 9812 9756
rect 9876 9692 9877 9756
rect 9811 9691 9877 9692
rect 7352 8672 7360 8736
rect 7424 8672 7440 8736
rect 7504 8672 7520 8736
rect 7584 8672 7600 8736
rect 7664 8672 7680 8736
rect 7744 8672 7752 8736
rect 7352 7648 7752 8672
rect 7352 7584 7360 7648
rect 7424 7584 7440 7648
rect 7504 7584 7520 7648
rect 7584 7584 7600 7648
rect 7664 7584 7680 7648
rect 7744 7584 7752 7648
rect 7352 6560 7752 7584
rect 9814 7309 9874 9691
rect 10352 9280 10752 10304
rect 11099 9484 11165 9485
rect 11099 9420 11100 9484
rect 11164 9420 11165 9484
rect 11099 9419 11165 9420
rect 10352 9216 10360 9280
rect 10424 9216 10440 9280
rect 10504 9216 10520 9280
rect 10584 9216 10600 9280
rect 10664 9216 10680 9280
rect 10744 9216 10752 9280
rect 10352 8192 10752 9216
rect 10352 8128 10360 8192
rect 10424 8128 10440 8192
rect 10504 8128 10520 8192
rect 10584 8128 10600 8192
rect 10664 8128 10680 8192
rect 10744 8128 10752 8192
rect 9811 7308 9877 7309
rect 9811 7244 9812 7308
rect 9876 7244 9877 7308
rect 9811 7243 9877 7244
rect 7352 6496 7360 6560
rect 7424 6496 7440 6560
rect 7504 6496 7520 6560
rect 7584 6496 7600 6560
rect 7664 6496 7680 6560
rect 7744 6496 7752 6560
rect 7352 5472 7752 6496
rect 7352 5408 7360 5472
rect 7424 5408 7440 5472
rect 7504 5408 7520 5472
rect 7584 5408 7600 5472
rect 7664 5408 7680 5472
rect 7744 5408 7752 5472
rect 7352 4384 7752 5408
rect 9814 5133 9874 7243
rect 10352 7104 10752 8128
rect 10352 7040 10360 7104
rect 10424 7040 10440 7104
rect 10504 7040 10520 7104
rect 10584 7040 10600 7104
rect 10664 7040 10680 7104
rect 10744 7040 10752 7104
rect 10352 6016 10752 7040
rect 10352 5952 10360 6016
rect 10424 5952 10440 6016
rect 10504 5952 10520 6016
rect 10584 5952 10600 6016
rect 10664 5952 10680 6016
rect 10744 5952 10752 6016
rect 9995 5404 10061 5405
rect 9995 5340 9996 5404
rect 10060 5340 10061 5404
rect 9995 5339 10061 5340
rect 9811 5132 9877 5133
rect 9811 5068 9812 5132
rect 9876 5068 9877 5132
rect 9811 5067 9877 5068
rect 7352 4320 7360 4384
rect 7424 4320 7440 4384
rect 7504 4320 7520 4384
rect 7584 4320 7600 4384
rect 7664 4320 7680 4384
rect 7744 4320 7752 4384
rect 7352 3296 7752 4320
rect 9443 3908 9509 3909
rect 9443 3844 9444 3908
rect 9508 3844 9509 3908
rect 9443 3843 9509 3844
rect 9075 3364 9141 3365
rect 9075 3300 9076 3364
rect 9140 3300 9141 3364
rect 9075 3299 9141 3300
rect 7352 3232 7360 3296
rect 7424 3232 7440 3296
rect 7504 3232 7520 3296
rect 7584 3232 7600 3296
rect 7664 3232 7680 3296
rect 7744 3232 7752 3296
rect 7352 2208 7752 3232
rect 9078 2685 9138 3299
rect 9259 3092 9325 3093
rect 9259 3028 9260 3092
rect 9324 3028 9325 3092
rect 9259 3027 9325 3028
rect 9075 2684 9141 2685
rect 9075 2620 9076 2684
rect 9140 2620 9141 2684
rect 9075 2619 9141 2620
rect 9262 2413 9322 3027
rect 9259 2412 9325 2413
rect 9259 2348 9260 2412
rect 9324 2348 9325 2412
rect 9259 2347 9325 2348
rect 7352 2144 7360 2208
rect 7424 2144 7440 2208
rect 7504 2144 7520 2208
rect 7584 2144 7600 2208
rect 7664 2144 7680 2208
rect 7744 2144 7752 2208
rect 7352 1120 7752 2144
rect 9446 1733 9506 3843
rect 9811 3772 9877 3773
rect 9811 3708 9812 3772
rect 9876 3708 9877 3772
rect 9811 3707 9877 3708
rect 9814 2821 9874 3707
rect 9811 2820 9877 2821
rect 9811 2756 9812 2820
rect 9876 2756 9877 2820
rect 9811 2755 9877 2756
rect 9443 1732 9509 1733
rect 9443 1668 9444 1732
rect 9508 1668 9509 1732
rect 9443 1667 9509 1668
rect 7352 1056 7360 1120
rect 7424 1056 7440 1120
rect 7504 1056 7520 1120
rect 7584 1056 7600 1120
rect 7664 1056 7680 1120
rect 7744 1056 7752 1120
rect 7352 496 7752 1056
rect 9998 917 10058 5339
rect 10352 4928 10752 5952
rect 10352 4864 10360 4928
rect 10424 4864 10440 4928
rect 10504 4864 10520 4928
rect 10584 4864 10600 4928
rect 10664 4864 10680 4928
rect 10744 4864 10752 4928
rect 10352 3840 10752 4864
rect 10352 3776 10360 3840
rect 10424 3776 10440 3840
rect 10504 3776 10520 3840
rect 10584 3776 10600 3840
rect 10664 3776 10680 3840
rect 10744 3776 10752 3840
rect 10352 2752 10752 3776
rect 11102 3365 11162 9419
rect 11099 3364 11165 3365
rect 11099 3300 11100 3364
rect 11164 3300 11165 3364
rect 11099 3299 11165 3300
rect 10352 2688 10360 2752
rect 10424 2688 10440 2752
rect 10504 2688 10520 2752
rect 10584 2688 10600 2752
rect 10664 2688 10680 2752
rect 10744 2688 10752 2752
rect 10352 1664 10752 2688
rect 13126 2685 13186 13363
rect 13352 13088 13752 14112
rect 13352 13024 13360 13088
rect 13424 13024 13440 13088
rect 13504 13024 13520 13088
rect 13584 13024 13600 13088
rect 13664 13024 13680 13088
rect 13744 13024 13752 13088
rect 13352 12000 13752 13024
rect 16352 14720 16752 15280
rect 16352 14656 16360 14720
rect 16424 14656 16440 14720
rect 16504 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16752 14720
rect 16352 13632 16752 14656
rect 16352 13568 16360 13632
rect 16424 13568 16440 13632
rect 16504 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16752 13632
rect 15699 12884 15765 12885
rect 15699 12820 15700 12884
rect 15764 12820 15765 12884
rect 15699 12819 15765 12820
rect 14963 12612 15029 12613
rect 14963 12548 14964 12612
rect 15028 12548 15029 12612
rect 14963 12547 15029 12548
rect 13352 11936 13360 12000
rect 13424 11936 13440 12000
rect 13504 11936 13520 12000
rect 13584 11936 13600 12000
rect 13664 11936 13680 12000
rect 13744 11936 13752 12000
rect 13352 10912 13752 11936
rect 13352 10848 13360 10912
rect 13424 10848 13440 10912
rect 13504 10848 13520 10912
rect 13584 10848 13600 10912
rect 13664 10848 13680 10912
rect 13744 10848 13752 10912
rect 13352 9824 13752 10848
rect 13352 9760 13360 9824
rect 13424 9760 13440 9824
rect 13504 9760 13520 9824
rect 13584 9760 13600 9824
rect 13664 9760 13680 9824
rect 13744 9760 13752 9824
rect 13352 8736 13752 9760
rect 14779 9212 14845 9213
rect 14779 9148 14780 9212
rect 14844 9148 14845 9212
rect 14779 9147 14845 9148
rect 13352 8672 13360 8736
rect 13424 8672 13440 8736
rect 13504 8672 13520 8736
rect 13584 8672 13600 8736
rect 13664 8672 13680 8736
rect 13744 8672 13752 8736
rect 13352 7648 13752 8672
rect 13352 7584 13360 7648
rect 13424 7584 13440 7648
rect 13504 7584 13520 7648
rect 13584 7584 13600 7648
rect 13664 7584 13680 7648
rect 13744 7584 13752 7648
rect 13352 6560 13752 7584
rect 13352 6496 13360 6560
rect 13424 6496 13440 6560
rect 13504 6496 13520 6560
rect 13584 6496 13600 6560
rect 13664 6496 13680 6560
rect 13744 6496 13752 6560
rect 13352 5472 13752 6496
rect 14782 5813 14842 9147
rect 14779 5812 14845 5813
rect 14779 5748 14780 5812
rect 14844 5748 14845 5812
rect 14779 5747 14845 5748
rect 13352 5408 13360 5472
rect 13424 5408 13440 5472
rect 13504 5408 13520 5472
rect 13584 5408 13600 5472
rect 13664 5408 13680 5472
rect 13744 5408 13752 5472
rect 13352 4384 13752 5408
rect 13352 4320 13360 4384
rect 13424 4320 13440 4384
rect 13504 4320 13520 4384
rect 13584 4320 13600 4384
rect 13664 4320 13680 4384
rect 13744 4320 13752 4384
rect 13352 3296 13752 4320
rect 13352 3232 13360 3296
rect 13424 3232 13440 3296
rect 13504 3232 13520 3296
rect 13584 3232 13600 3296
rect 13664 3232 13680 3296
rect 13744 3232 13752 3296
rect 13123 2684 13189 2685
rect 13123 2620 13124 2684
rect 13188 2620 13189 2684
rect 13123 2619 13189 2620
rect 10352 1600 10360 1664
rect 10424 1600 10440 1664
rect 10504 1600 10520 1664
rect 10584 1600 10600 1664
rect 10664 1600 10680 1664
rect 10744 1600 10752 1664
rect 9995 916 10061 917
rect 9995 852 9996 916
rect 10060 852 10061 916
rect 9995 851 10061 852
rect 10352 576 10752 1600
rect 10352 512 10360 576
rect 10424 512 10440 576
rect 10504 512 10520 576
rect 10584 512 10600 576
rect 10664 512 10680 576
rect 10744 512 10752 576
rect 10352 496 10752 512
rect 13352 2208 13752 3232
rect 13352 2144 13360 2208
rect 13424 2144 13440 2208
rect 13504 2144 13520 2208
rect 13584 2144 13600 2208
rect 13664 2144 13680 2208
rect 13744 2144 13752 2208
rect 13352 1120 13752 2144
rect 14966 2141 15026 12547
rect 15147 10300 15213 10301
rect 15147 10236 15148 10300
rect 15212 10236 15213 10300
rect 15147 10235 15213 10236
rect 15150 5541 15210 10235
rect 15702 6901 15762 12819
rect 16352 12544 16752 13568
rect 16352 12480 16360 12544
rect 16424 12480 16440 12544
rect 16504 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16752 12544
rect 16352 11456 16752 12480
rect 16352 11392 16360 11456
rect 16424 11392 16440 11456
rect 16504 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16752 11456
rect 16352 10368 16752 11392
rect 16352 10304 16360 10368
rect 16424 10304 16440 10368
rect 16504 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16752 10368
rect 16352 9280 16752 10304
rect 16352 9216 16360 9280
rect 16424 9216 16440 9280
rect 16504 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16752 9280
rect 16352 8192 16752 9216
rect 16352 8128 16360 8192
rect 16424 8128 16440 8192
rect 16504 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16752 8192
rect 16352 7104 16752 8128
rect 16352 7040 16360 7104
rect 16424 7040 16440 7104
rect 16504 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16752 7104
rect 15699 6900 15765 6901
rect 15699 6836 15700 6900
rect 15764 6836 15765 6900
rect 15699 6835 15765 6836
rect 16352 6016 16752 7040
rect 16352 5952 16360 6016
rect 16424 5952 16440 6016
rect 16504 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16752 6016
rect 15147 5540 15213 5541
rect 15147 5476 15148 5540
rect 15212 5476 15213 5540
rect 15147 5475 15213 5476
rect 16067 5540 16133 5541
rect 16067 5476 16068 5540
rect 16132 5476 16133 5540
rect 16067 5475 16133 5476
rect 14963 2140 15029 2141
rect 14963 2076 14964 2140
rect 15028 2076 15029 2140
rect 14963 2075 15029 2076
rect 16070 1461 16130 5475
rect 16352 4928 16752 5952
rect 16352 4864 16360 4928
rect 16424 4864 16440 4928
rect 16504 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16752 4928
rect 16352 3840 16752 4864
rect 16352 3776 16360 3840
rect 16424 3776 16440 3840
rect 16504 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16752 3840
rect 16352 2752 16752 3776
rect 16352 2688 16360 2752
rect 16424 2688 16440 2752
rect 16504 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16752 2752
rect 16352 1664 16752 2688
rect 16352 1600 16360 1664
rect 16424 1600 16440 1664
rect 16504 1600 16520 1664
rect 16584 1600 16600 1664
rect 16664 1600 16680 1664
rect 16744 1600 16752 1664
rect 16067 1460 16133 1461
rect 16067 1396 16068 1460
rect 16132 1396 16133 1460
rect 16067 1395 16133 1396
rect 13352 1056 13360 1120
rect 13424 1056 13440 1120
rect 13504 1056 13520 1120
rect 13584 1056 13600 1120
rect 13664 1056 13680 1120
rect 13744 1056 13752 1120
rect 13352 496 13752 1056
rect 16352 576 16752 1600
rect 16352 512 16360 576
rect 16424 512 16440 576
rect 16504 512 16520 576
rect 16584 512 16600 576
rect 16664 512 16680 576
rect 16744 512 16752 576
rect 16352 496 16752 512
rect 19352 15264 19752 15280
rect 19352 15200 19360 15264
rect 19424 15200 19440 15264
rect 19504 15200 19520 15264
rect 19584 15200 19600 15264
rect 19664 15200 19680 15264
rect 19744 15200 19752 15264
rect 19352 14176 19752 15200
rect 19352 14112 19360 14176
rect 19424 14112 19440 14176
rect 19504 14112 19520 14176
rect 19584 14112 19600 14176
rect 19664 14112 19680 14176
rect 19744 14112 19752 14176
rect 19352 13088 19752 14112
rect 19352 13024 19360 13088
rect 19424 13024 19440 13088
rect 19504 13024 19520 13088
rect 19584 13024 19600 13088
rect 19664 13024 19680 13088
rect 19744 13024 19752 13088
rect 19352 12000 19752 13024
rect 19352 11936 19360 12000
rect 19424 11936 19440 12000
rect 19504 11936 19520 12000
rect 19584 11936 19600 12000
rect 19664 11936 19680 12000
rect 19744 11936 19752 12000
rect 19352 10912 19752 11936
rect 19352 10848 19360 10912
rect 19424 10848 19440 10912
rect 19504 10848 19520 10912
rect 19584 10848 19600 10912
rect 19664 10848 19680 10912
rect 19744 10848 19752 10912
rect 19352 9824 19752 10848
rect 19352 9760 19360 9824
rect 19424 9760 19440 9824
rect 19504 9760 19520 9824
rect 19584 9760 19600 9824
rect 19664 9760 19680 9824
rect 19744 9760 19752 9824
rect 19352 8736 19752 9760
rect 22352 14720 22752 15280
rect 22352 14656 22360 14720
rect 22424 14656 22440 14720
rect 22504 14656 22520 14720
rect 22584 14656 22600 14720
rect 22664 14656 22680 14720
rect 22744 14656 22752 14720
rect 22352 13632 22752 14656
rect 22352 13568 22360 13632
rect 22424 13568 22440 13632
rect 22504 13568 22520 13632
rect 22584 13568 22600 13632
rect 22664 13568 22680 13632
rect 22744 13568 22752 13632
rect 22352 12544 22752 13568
rect 22352 12480 22360 12544
rect 22424 12480 22440 12544
rect 22504 12480 22520 12544
rect 22584 12480 22600 12544
rect 22664 12480 22680 12544
rect 22744 12480 22752 12544
rect 22352 11456 22752 12480
rect 22352 11392 22360 11456
rect 22424 11392 22440 11456
rect 22504 11392 22520 11456
rect 22584 11392 22600 11456
rect 22664 11392 22680 11456
rect 22744 11392 22752 11456
rect 22352 10368 22752 11392
rect 22352 10304 22360 10368
rect 22424 10304 22440 10368
rect 22504 10304 22520 10368
rect 22584 10304 22600 10368
rect 22664 10304 22680 10368
rect 22744 10304 22752 10368
rect 22352 9280 22752 10304
rect 22352 9216 22360 9280
rect 22424 9216 22440 9280
rect 22504 9216 22520 9280
rect 22584 9216 22600 9280
rect 22664 9216 22680 9280
rect 22744 9216 22752 9280
rect 19931 9212 19997 9213
rect 19931 9148 19932 9212
rect 19996 9148 19997 9212
rect 19931 9147 19997 9148
rect 19352 8672 19360 8736
rect 19424 8672 19440 8736
rect 19504 8672 19520 8736
rect 19584 8672 19600 8736
rect 19664 8672 19680 8736
rect 19744 8672 19752 8736
rect 19352 7648 19752 8672
rect 19934 8261 19994 9147
rect 19931 8260 19997 8261
rect 19931 8196 19932 8260
rect 19996 8196 19997 8260
rect 19931 8195 19997 8196
rect 19352 7584 19360 7648
rect 19424 7584 19440 7648
rect 19504 7584 19520 7648
rect 19584 7584 19600 7648
rect 19664 7584 19680 7648
rect 19744 7584 19752 7648
rect 19352 6560 19752 7584
rect 19352 6496 19360 6560
rect 19424 6496 19440 6560
rect 19504 6496 19520 6560
rect 19584 6496 19600 6560
rect 19664 6496 19680 6560
rect 19744 6496 19752 6560
rect 19352 5472 19752 6496
rect 22352 8192 22752 9216
rect 22352 8128 22360 8192
rect 22424 8128 22440 8192
rect 22504 8128 22520 8192
rect 22584 8128 22600 8192
rect 22664 8128 22680 8192
rect 22744 8128 22752 8192
rect 22352 7104 22752 8128
rect 22352 7040 22360 7104
rect 22424 7040 22440 7104
rect 22504 7040 22520 7104
rect 22584 7040 22600 7104
rect 22664 7040 22680 7104
rect 22744 7040 22752 7104
rect 22352 6016 22752 7040
rect 22352 5952 22360 6016
rect 22424 5952 22440 6016
rect 22504 5952 22520 6016
rect 22584 5952 22600 6016
rect 22664 5952 22680 6016
rect 22744 5952 22752 6016
rect 20667 5676 20733 5677
rect 20667 5612 20668 5676
rect 20732 5612 20733 5676
rect 20667 5611 20733 5612
rect 19352 5408 19360 5472
rect 19424 5408 19440 5472
rect 19504 5408 19520 5472
rect 19584 5408 19600 5472
rect 19664 5408 19680 5472
rect 19744 5408 19752 5472
rect 19352 4384 19752 5408
rect 19352 4320 19360 4384
rect 19424 4320 19440 4384
rect 19504 4320 19520 4384
rect 19584 4320 19600 4384
rect 19664 4320 19680 4384
rect 19744 4320 19752 4384
rect 19352 3296 19752 4320
rect 19352 3232 19360 3296
rect 19424 3232 19440 3296
rect 19504 3232 19520 3296
rect 19584 3232 19600 3296
rect 19664 3232 19680 3296
rect 19744 3232 19752 3296
rect 19352 2208 19752 3232
rect 20670 2685 20730 5611
rect 22352 4928 22752 5952
rect 22352 4864 22360 4928
rect 22424 4864 22440 4928
rect 22504 4864 22520 4928
rect 22584 4864 22600 4928
rect 22664 4864 22680 4928
rect 22744 4864 22752 4928
rect 22352 3840 22752 4864
rect 22352 3776 22360 3840
rect 22424 3776 22440 3840
rect 22504 3776 22520 3840
rect 22584 3776 22600 3840
rect 22664 3776 22680 3840
rect 22744 3776 22752 3840
rect 22352 2752 22752 3776
rect 22352 2688 22360 2752
rect 22424 2688 22440 2752
rect 22504 2688 22520 2752
rect 22584 2688 22600 2752
rect 22664 2688 22680 2752
rect 22744 2688 22752 2752
rect 20667 2684 20733 2685
rect 20667 2620 20668 2684
rect 20732 2620 20733 2684
rect 20667 2619 20733 2620
rect 19352 2144 19360 2208
rect 19424 2144 19440 2208
rect 19504 2144 19520 2208
rect 19584 2144 19600 2208
rect 19664 2144 19680 2208
rect 19744 2144 19752 2208
rect 19352 1120 19752 2144
rect 19352 1056 19360 1120
rect 19424 1056 19440 1120
rect 19504 1056 19520 1120
rect 19584 1056 19600 1120
rect 19664 1056 19680 1120
rect 19744 1056 19752 1120
rect 19352 496 19752 1056
rect 22352 1664 22752 2688
rect 22352 1600 22360 1664
rect 22424 1600 22440 1664
rect 22504 1600 22520 1664
rect 22584 1600 22600 1664
rect 22664 1600 22680 1664
rect 22744 1600 22752 1664
rect 22352 576 22752 1600
rect 22352 512 22360 576
rect 22424 512 22440 576
rect 22504 512 22520 576
rect 22584 512 22600 576
rect 22664 512 22680 576
rect 22744 512 22752 576
rect 22352 496 22752 512
use sky130_fd_sc_hd__dlymetal6s2s_1  _0516_
timestamp 1713545776
transform 1 0 21712 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0517_
timestamp 1713545776
transform -1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0518_
timestamp 1713545776
transform -1 0 6624 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0519_
timestamp 1713545776
transform -1 0 21896 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0520_
timestamp 1713545776
transform -1 0 17664 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0521_
timestamp 1713545776
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0522_
timestamp 1713545776
transform 1 0 17388 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0523_
timestamp 1713545776
transform 1 0 16744 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0524_
timestamp 1713545776
transform -1 0 18032 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0525_
timestamp 1713545776
transform 1 0 17388 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0526_
timestamp 1713545776
transform -1 0 21896 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0527_
timestamp 1713545776
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0528_
timestamp 1713545776
transform 1 0 22172 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0529_
timestamp 1713545776
transform -1 0 21160 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0530_
timestamp 1713545776
transform 1 0 18032 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0531_
timestamp 1713545776
transform 1 0 16836 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1713545776
transform 1 0 21252 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0533_
timestamp 1713545776
transform 1 0 16652 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0534_
timestamp 1713545776
transform 1 0 16284 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0535_
timestamp 1713545776
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0536_
timestamp 1713545776
transform -1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0537_
timestamp 1713545776
transform 1 0 2208 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0538_
timestamp 1713545776
transform -1 0 6256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0539_
timestamp 1713545776
transform 1 0 4324 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0540_
timestamp 1713545776
transform -1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0541_
timestamp 1713545776
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0542_
timestamp 1713545776
transform -1 0 4140 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0543_
timestamp 1713545776
transform -1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0544_
timestamp 1713545776
transform 1 0 4968 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0545_
timestamp 1713545776
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0546_
timestamp 1713545776
transform 1 0 4784 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0547_
timestamp 1713545776
transform -1 0 5520 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0548_
timestamp 1713545776
transform 1 0 5796 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _0549_
timestamp 1713545776
transform -1 0 5704 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0550_
timestamp 1713545776
transform 1 0 5244 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0551_
timestamp 1713545776
transform 1 0 6532 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0552_
timestamp 1713545776
transform 1 0 7360 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0553_
timestamp 1713545776
transform 1 0 13524 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _0554_
timestamp 1713545776
transform -1 0 14076 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0555_
timestamp 1713545776
transform -1 0 12972 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0556_
timestamp 1713545776
transform -1 0 13248 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0557_
timestamp 1713545776
transform 1 0 2668 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0558_
timestamp 1713545776
transform 1 0 3680 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0559_
timestamp 1713545776
transform 1 0 12236 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0560_
timestamp 1713545776
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1713545776
transform -1 0 18768 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0562_
timestamp 1713545776
transform 1 0 18676 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1713545776
transform -1 0 18216 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0564_
timestamp 1713545776
transform 1 0 17296 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0565_
timestamp 1713545776
transform -1 0 17204 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1713545776
transform -1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0567_
timestamp 1713545776
transform -1 0 21804 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0568_
timestamp 1713545776
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0569_
timestamp 1713545776
transform -1 0 10856 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0570_
timestamp 1713545776
transform 1 0 10488 0 1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__o311a_1  _0571_
timestamp 1713545776
transform 1 0 16100 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0572_
timestamp 1713545776
transform 1 0 15364 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0573_
timestamp 1713545776
transform 1 0 2852 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0574_
timestamp 1713545776
transform -1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0575_
timestamp 1713545776
transform 1 0 4324 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0576_
timestamp 1713545776
transform -1 0 4692 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0577_
timestamp 1713545776
transform 1 0 3404 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0578_
timestamp 1713545776
transform 1 0 5244 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0579_
timestamp 1713545776
transform 1 0 5980 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _0580_
timestamp 1713545776
transform 1 0 5796 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _0581_
timestamp 1713545776
transform -1 0 15916 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0582_
timestamp 1713545776
transform 1 0 16100 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1713545776
transform -1 0 15456 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0584_
timestamp 1713545776
transform 1 0 15916 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0585_
timestamp 1713545776
transform -1 0 15180 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0586_
timestamp 1713545776
transform 1 0 15732 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0587_
timestamp 1713545776
transform -1 0 18584 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0588_
timestamp 1713545776
transform 1 0 13064 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0589_
timestamp 1713545776
transform 1 0 13064 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _0590_
timestamp 1713545776
transform 1 0 16100 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _0591_
timestamp 1713545776
transform -1 0 16376 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0592_
timestamp 1713545776
transform -1 0 20976 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0593_
timestamp 1713545776
transform -1 0 19136 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0594_
timestamp 1713545776
transform -1 0 17848 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0595_
timestamp 1713545776
transform 1 0 6624 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0596_
timestamp 1713545776
transform -1 0 17388 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0597_
timestamp 1713545776
transform 1 0 16192 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0598_
timestamp 1713545776
transform 1 0 15364 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0599_
timestamp 1713545776
transform 1 0 13524 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0600_
timestamp 1713545776
transform -1 0 14352 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0601_
timestamp 1713545776
transform -1 0 13892 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0602_
timestamp 1713545776
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0603_
timestamp 1713545776
transform -1 0 11592 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0604_
timestamp 1713545776
transform -1 0 22264 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _0605_
timestamp 1713545776
transform 1 0 21252 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0606_
timestamp 1713545776
transform -1 0 22540 0 1 544
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0607_
timestamp 1713545776
transform -1 0 19228 0 -1 1632
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _0608_
timestamp 1713545776
transform -1 0 17388 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0609_
timestamp 1713545776
transform -1 0 17664 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0610_
timestamp 1713545776
transform -1 0 22540 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0611_
timestamp 1713545776
transform -1 0 14444 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0612_
timestamp 1713545776
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0613_
timestamp 1713545776
transform 1 0 4968 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0614_
timestamp 1713545776
transform -1 0 6348 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0615_
timestamp 1713545776
transform -1 0 6992 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _0616_
timestamp 1713545776
transform -1 0 5704 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_1  _0617_
timestamp 1713545776
transform -1 0 14536 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0618_
timestamp 1713545776
transform 1 0 13524 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0619_
timestamp 1713545776
transform -1 0 21988 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0620_
timestamp 1713545776
transform 1 0 18216 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0621_
timestamp 1713545776
transform -1 0 15456 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0622_
timestamp 1713545776
transform -1 0 13340 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0623_
timestamp 1713545776
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0624_
timestamp 1713545776
transform -1 0 16744 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0625_
timestamp 1713545776
transform -1 0 18124 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0626_
timestamp 1713545776
transform 1 0 17388 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0627_
timestamp 1713545776
transform 1 0 15456 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0628_
timestamp 1713545776
transform 1 0 12972 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1713545776
transform 1 0 12236 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0630_
timestamp 1713545776
transform 1 0 4416 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0631_
timestamp 1713545776
transform 1 0 7636 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0632_
timestamp 1713545776
transform 1 0 13524 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0633_
timestamp 1713545776
transform -1 0 17112 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0634_
timestamp 1713545776
transform 1 0 17112 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0635_
timestamp 1713545776
transform 1 0 4140 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0636_
timestamp 1713545776
transform -1 0 6716 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _0637_
timestamp 1713545776
transform 1 0 6072 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _0638_
timestamp 1713545776
transform 1 0 10304 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0639_
timestamp 1713545776
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0640_
timestamp 1713545776
transform 1 0 16100 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0641_
timestamp 1713545776
transform 1 0 11592 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0642_
timestamp 1713545776
transform -1 0 19228 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0643_
timestamp 1713545776
transform 1 0 17848 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0644_
timestamp 1713545776
transform 1 0 3680 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0645_
timestamp 1713545776
transform 1 0 4784 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1713545776
transform -1 0 22264 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0647_
timestamp 1713545776
transform -1 0 21712 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0648_
timestamp 1713545776
transform 1 0 20700 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0649_
timestamp 1713545776
transform 1 0 6256 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0650_
timestamp 1713545776
transform -1 0 7452 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1713545776
transform -1 0 7176 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0652_
timestamp 1713545776
transform 1 0 9568 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0653_
timestamp 1713545776
transform 1 0 9016 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1713545776
transform 1 0 10212 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0655_
timestamp 1713545776
transform 1 0 10212 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0656_
timestamp 1713545776
transform 1 0 11040 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0657_
timestamp 1713545776
transform 1 0 4048 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0658_
timestamp 1713545776
transform -1 0 5704 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1713545776
transform 1 0 18216 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0660_
timestamp 1713545776
transform 1 0 3772 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0661_
timestamp 1713545776
transform -1 0 4784 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0662_
timestamp 1713545776
transform 1 0 4784 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0663_
timestamp 1713545776
transform 1 0 6532 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0664_
timestamp 1713545776
transform 1 0 7360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0665_
timestamp 1713545776
transform 1 0 7084 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0666_
timestamp 1713545776
transform 1 0 7728 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0667_
timestamp 1713545776
transform -1 0 16468 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0668_
timestamp 1713545776
transform 1 0 5336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0669_
timestamp 1713545776
transform -1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0670_
timestamp 1713545776
transform 1 0 5796 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__o221a_1  _0671_
timestamp 1713545776
transform 1 0 13524 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0672_
timestamp 1713545776
transform 1 0 13524 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0673_
timestamp 1713545776
transform -1 0 8280 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0674_
timestamp 1713545776
transform 1 0 16928 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0675_
timestamp 1713545776
transform 1 0 8372 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0676_
timestamp 1713545776
transform 1 0 7544 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0677_
timestamp 1713545776
transform 1 0 16560 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0678_
timestamp 1713545776
transform -1 0 16560 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0679_
timestamp 1713545776
transform 1 0 16192 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_2  _0680_
timestamp 1713545776
transform 1 0 5704 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _0681_
timestamp 1713545776
transform 1 0 9936 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0682_
timestamp 1713545776
transform 1 0 10948 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0683_
timestamp 1713545776
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0684_
timestamp 1713545776
transform -1 0 6164 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0685_
timestamp 1713545776
transform -1 0 9016 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0686_
timestamp 1713545776
transform 1 0 8924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0687_
timestamp 1713545776
transform 1 0 6716 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0688_
timestamp 1713545776
transform 1 0 7360 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1713545776
transform 1 0 5796 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1713545776
transform 1 0 4600 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0691_
timestamp 1713545776
transform -1 0 5520 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0692_
timestamp 1713545776
transform 1 0 7636 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0693_
timestamp 1713545776
transform 1 0 8372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0694_
timestamp 1713545776
transform -1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0695_
timestamp 1713545776
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0696_
timestamp 1713545776
transform 1 0 9936 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0697_
timestamp 1713545776
transform 1 0 9936 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0698_
timestamp 1713545776
transform -1 0 11592 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0699_
timestamp 1713545776
transform 1 0 10856 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0700_
timestamp 1713545776
transform 1 0 8372 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0701_
timestamp 1713545776
transform -1 0 9936 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1713545776
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0703_
timestamp 1713545776
transform 1 0 7360 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0704_
timestamp 1713545776
transform -1 0 8924 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0705_
timestamp 1713545776
transform 1 0 9016 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0706_
timestamp 1713545776
transform -1 0 9844 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0707_
timestamp 1713545776
transform 1 0 9476 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0708_
timestamp 1713545776
transform -1 0 10856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0709_
timestamp 1713545776
transform -1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0710_
timestamp 1713545776
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0711_
timestamp 1713545776
transform 1 0 5520 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__o221a_1  _0712_
timestamp 1713545776
transform -1 0 14260 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0713_
timestamp 1713545776
transform 1 0 12880 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0714_
timestamp 1713545776
transform -1 0 10580 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0715_
timestamp 1713545776
transform 1 0 17848 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0716_
timestamp 1713545776
transform 1 0 9016 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0717_
timestamp 1713545776
transform -1 0 9844 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0718_
timestamp 1713545776
transform -1 0 9108 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0719_
timestamp 1713545776
transform 1 0 7636 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1713545776
transform 1 0 8924 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0721_
timestamp 1713545776
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1713545776
transform 1 0 7820 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0723_
timestamp 1713545776
transform 1 0 8004 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1713545776
transform -1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0725_
timestamp 1713545776
transform -1 0 10120 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0726_
timestamp 1713545776
transform 1 0 9108 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0727_
timestamp 1713545776
transform 1 0 9292 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1713545776
transform 1 0 9384 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0729_
timestamp 1713545776
transform 1 0 9752 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0730_
timestamp 1713545776
transform 1 0 10396 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0731_
timestamp 1713545776
transform -1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0732_
timestamp 1713545776
transform -1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0733_
timestamp 1713545776
transform 1 0 5796 0 -1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_1  _0734_
timestamp 1713545776
transform -1 0 9568 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0735_
timestamp 1713545776
transform 1 0 14996 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0736_
timestamp 1713545776
transform 1 0 8740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0737_
timestamp 1713545776
transform 1 0 10396 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0738_
timestamp 1713545776
transform -1 0 14352 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0739_
timestamp 1713545776
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0740_
timestamp 1713545776
transform 1 0 10580 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0741_
timestamp 1713545776
transform 1 0 17480 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0742_
timestamp 1713545776
transform 1 0 9200 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0743_
timestamp 1713545776
transform -1 0 10856 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0744_
timestamp 1713545776
transform -1 0 8924 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0745_
timestamp 1713545776
transform 1 0 12788 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0746_
timestamp 1713545776
transform -1 0 14168 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0747_
timestamp 1713545776
transform 1 0 10028 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _0748_
timestamp 1713545776
transform 1 0 10948 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0749_
timestamp 1713545776
transform -1 0 11500 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1713545776
transform -1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0751_
timestamp 1713545776
transform -1 0 5152 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1713545776
transform 1 0 6348 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0753_
timestamp 1713545776
transform -1 0 5888 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0754_
timestamp 1713545776
transform -1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0755_
timestamp 1713545776
transform 1 0 5888 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0756_
timestamp 1713545776
transform 1 0 13432 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0757_
timestamp 1713545776
transform -1 0 9568 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0758_
timestamp 1713545776
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0759_
timestamp 1713545776
transform 1 0 12604 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0760_
timestamp 1713545776
transform 1 0 13064 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0761_
timestamp 1713545776
transform 1 0 16652 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_2  _0762_
timestamp 1713545776
transform -1 0 11776 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0763_
timestamp 1713545776
transform -1 0 14352 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0764_
timestamp 1713545776
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0765_
timestamp 1713545776
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0766_
timestamp 1713545776
transform -1 0 20332 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1713545776
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0768_
timestamp 1713545776
transform 1 0 15088 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0769_
timestamp 1713545776
transform -1 0 16284 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0770_
timestamp 1713545776
transform -1 0 14996 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0771_
timestamp 1713545776
transform 1 0 15364 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0772_
timestamp 1713545776
transform 1 0 14996 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0773_
timestamp 1713545776
transform -1 0 12696 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0774_
timestamp 1713545776
transform 1 0 12236 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0775_
timestamp 1713545776
transform -1 0 15824 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0776_
timestamp 1713545776
transform 1 0 15272 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0777_
timestamp 1713545776
transform 1 0 14352 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0778_
timestamp 1713545776
transform 1 0 5428 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0779_
timestamp 1713545776
transform -1 0 15456 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0780_
timestamp 1713545776
transform 1 0 13064 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0781_
timestamp 1713545776
transform -1 0 13432 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0782_
timestamp 1713545776
transform -1 0 14168 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0783_
timestamp 1713545776
transform 1 0 13524 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0784_
timestamp 1713545776
transform -1 0 4876 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0785_
timestamp 1713545776
transform 1 0 10580 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0786_
timestamp 1713545776
transform 1 0 13524 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0787_
timestamp 1713545776
transform 1 0 12328 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0788_
timestamp 1713545776
transform -1 0 12236 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0789_
timestamp 1713545776
transform -1 0 12696 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0790_
timestamp 1713545776
transform -1 0 15732 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0791_
timestamp 1713545776
transform 1 0 5520 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0792_
timestamp 1713545776
transform 1 0 6348 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0793_
timestamp 1713545776
transform 1 0 15364 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0794_
timestamp 1713545776
transform 1 0 14996 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0795_
timestamp 1713545776
transform -1 0 11132 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0796_
timestamp 1713545776
transform -1 0 11684 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0797_
timestamp 1713545776
transform -1 0 12144 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0798_
timestamp 1713545776
transform -1 0 12144 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0799_
timestamp 1713545776
transform -1 0 13432 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0800_
timestamp 1713545776
transform 1 0 16560 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0801_
timestamp 1713545776
transform 1 0 3772 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0802_
timestamp 1713545776
transform 1 0 2852 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0803_
timestamp 1713545776
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0804_
timestamp 1713545776
transform 1 0 10948 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0805_
timestamp 1713545776
transform -1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0806_
timestamp 1713545776
transform 1 0 11776 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0807_
timestamp 1713545776
transform -1 0 10856 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0808_
timestamp 1713545776
transform -1 0 13432 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0809_
timestamp 1713545776
transform 1 0 2484 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0810_
timestamp 1713545776
transform -1 0 3128 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0811_
timestamp 1713545776
transform 1 0 11684 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0812_
timestamp 1713545776
transform -1 0 11684 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0813_
timestamp 1713545776
transform 1 0 10856 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0814_
timestamp 1713545776
transform 1 0 9752 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0815_
timestamp 1713545776
transform 1 0 18124 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0816_
timestamp 1713545776
transform 1 0 3220 0 1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0817_
timestamp 1713545776
transform -1 0 10856 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0818_
timestamp 1713545776
transform -1 0 11684 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0819_
timestamp 1713545776
transform 1 0 11224 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0820_
timestamp 1713545776
transform 1 0 9476 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0821_
timestamp 1713545776
transform 1 0 3036 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__o2bb2a_1  _0822_
timestamp 1713545776
transform 1 0 14352 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0823_
timestamp 1713545776
transform 1 0 12696 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0824_
timestamp 1713545776
transform 1 0 12144 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0825_
timestamp 1713545776
transform 1 0 11224 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0826_
timestamp 1713545776
transform 1 0 15180 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1713545776
transform -1 0 16376 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1713545776
transform 1 0 14812 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0829_
timestamp 1713545776
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0830_
timestamp 1713545776
transform 1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0831_
timestamp 1713545776
transform 1 0 15180 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0832_
timestamp 1713545776
transform -1 0 16560 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0833_
timestamp 1713545776
transform 1 0 15916 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0834_
timestamp 1713545776
transform -1 0 16652 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0835_
timestamp 1713545776
transform 1 0 13708 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 1713545776
transform 1 0 12972 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0837_
timestamp 1713545776
transform -1 0 16008 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0838_
timestamp 1713545776
transform -1 0 14904 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0839_
timestamp 1713545776
transform 1 0 14168 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0840_
timestamp 1713545776
transform -1 0 16008 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0841_
timestamp 1713545776
transform 1 0 11592 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 1713545776
transform 1 0 11684 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1713545776
transform 1 0 12144 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0844_
timestamp 1713545776
transform -1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0845_
timestamp 1713545776
transform -1 0 12604 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0846_
timestamp 1713545776
transform 1 0 12696 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0847_
timestamp 1713545776
transform 1 0 13524 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0848_
timestamp 1713545776
transform -1 0 12696 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0849_
timestamp 1713545776
transform -1 0 17204 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1713545776
transform 1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0851_
timestamp 1713545776
transform 1 0 15732 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0852_
timestamp 1713545776
transform -1 0 15364 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _0853_
timestamp 1713545776
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0854_
timestamp 1713545776
transform -1 0 15088 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0855_
timestamp 1713545776
transform -1 0 15732 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0856_
timestamp 1713545776
transform -1 0 16652 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0857_
timestamp 1713545776
transform 1 0 14444 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0858_
timestamp 1713545776
transform 1 0 10580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0859_
timestamp 1713545776
transform 1 0 10396 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0860_
timestamp 1713545776
transform -1 0 15180 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _0861_
timestamp 1713545776
transform -1 0 11960 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0862_
timestamp 1713545776
transform -1 0 12144 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0863_
timestamp 1713545776
transform -1 0 12236 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0864_
timestamp 1713545776
transform -1 0 19228 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0865_
timestamp 1713545776
transform 1 0 14076 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1713545776
transform 1 0 14628 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0867_
timestamp 1713545776
transform 1 0 13800 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0868_
timestamp 1713545776
transform -1 0 15732 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0869_
timestamp 1713545776
transform -1 0 14996 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0870_
timestamp 1713545776
transform -1 0 18032 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1713545776
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0872_
timestamp 1713545776
transform 1 0 10120 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0873_
timestamp 1713545776
transform -1 0 11684 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0874_
timestamp 1713545776
transform 1 0 11040 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0875_
timestamp 1713545776
transform 1 0 10580 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0876_
timestamp 1713545776
transform 1 0 12880 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0877_
timestamp 1713545776
transform 1 0 13984 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0878_
timestamp 1713545776
transform -1 0 14720 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0879_
timestamp 1713545776
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0880_
timestamp 1713545776
transform 1 0 13432 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0881_
timestamp 1713545776
transform -1 0 14720 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1713545776
transform -1 0 2576 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1713545776
transform -1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0884_
timestamp 1713545776
transform 1 0 2760 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0885_
timestamp 1713545776
transform -1 0 3680 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0886_
timestamp 1713545776
transform 1 0 3496 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0887_
timestamp 1713545776
transform 1 0 3956 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0888_
timestamp 1713545776
transform -1 0 22172 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0889_
timestamp 1713545776
transform -1 0 19688 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0890_
timestamp 1713545776
transform 1 0 2484 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1713545776
transform -1 0 3772 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0892_
timestamp 1713545776
transform 1 0 2300 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0893_
timestamp 1713545776
transform -1 0 3312 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0894_
timestamp 1713545776
transform 1 0 3128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0895_
timestamp 1713545776
transform 1 0 4600 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0896_
timestamp 1713545776
transform 1 0 3220 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0897_
timestamp 1713545776
transform -1 0 3772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0898_
timestamp 1713545776
transform 1 0 1932 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0899_
timestamp 1713545776
transform -1 0 3772 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0900_
timestamp 1713545776
transform -1 0 3496 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0901_
timestamp 1713545776
transform 1 0 2300 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0902_
timestamp 1713545776
transform 1 0 1932 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0903_
timestamp 1713545776
transform 1 0 1840 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _0904_
timestamp 1713545776
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0905_
timestamp 1713545776
transform -1 0 2576 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0906_
timestamp 1713545776
transform 1 0 2760 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0907_
timestamp 1713545776
transform 1 0 4600 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _0908_
timestamp 1713545776
transform -1 0 4600 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0909_
timestamp 1713545776
transform 1 0 20056 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1713545776
transform -1 0 21160 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _0911_
timestamp 1713545776
transform 1 0 21344 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _0912_
timestamp 1713545776
transform 1 0 20700 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _0913_
timestamp 1713545776
transform 1 0 21896 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0914_
timestamp 1713545776
transform -1 0 22172 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _0915_
timestamp 1713545776
transform 1 0 21252 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0916_
timestamp 1713545776
transform -1 0 20976 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0917_
timestamp 1713545776
transform -1 0 19688 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 1713545776
transform 1 0 18860 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0919_
timestamp 1713545776
transform 1 0 18308 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0920_
timestamp 1713545776
transform -1 0 19136 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0921_
timestamp 1713545776
transform -1 0 20424 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0922_
timestamp 1713545776
transform 1 0 19320 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0923_
timestamp 1713545776
transform -1 0 21344 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0924_
timestamp 1713545776
transform -1 0 20424 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1713545776
transform -1 0 19872 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 1713545776
transform 1 0 18952 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0927_
timestamp 1713545776
transform -1 0 19872 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0928_
timestamp 1713545776
transform -1 0 19596 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0929_
timestamp 1713545776
transform 1 0 19320 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1713545776
transform -1 0 19964 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0931_
timestamp 1713545776
transform -1 0 12236 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1713545776
transform -1 0 7912 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0933_
timestamp 1713545776
transform -1 0 6992 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0934_
timestamp 1713545776
transform 1 0 3772 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0935_
timestamp 1713545776
transform 1 0 5980 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0936_
timestamp 1713545776
transform 1 0 6532 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0937_
timestamp 1713545776
transform 1 0 7820 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0938_
timestamp 1713545776
transform 1 0 7820 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0939_
timestamp 1713545776
transform 1 0 18676 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0940_
timestamp 1713545776
transform 1 0 8464 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0941_
timestamp 1713545776
transform -1 0 9016 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0942_
timestamp 1713545776
transform -1 0 5428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0943_
timestamp 1713545776
transform -1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0944_
timestamp 1713545776
transform 1 0 18676 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0945_
timestamp 1713545776
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0946_
timestamp 1713545776
transform -1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0947_
timestamp 1713545776
transform -1 0 8648 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0948_
timestamp 1713545776
transform 1 0 8372 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0949_
timestamp 1713545776
transform -1 0 8556 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1713545776
transform 1 0 7452 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0951_
timestamp 1713545776
transform -1 0 9292 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0952_
timestamp 1713545776
transform -1 0 8924 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0953_
timestamp 1713545776
transform -1 0 11684 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1713545776
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0955_
timestamp 1713545776
transform -1 0 3036 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1713545776
transform 1 0 1748 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0957_
timestamp 1713545776
transform 1 0 2300 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0958_
timestamp 1713545776
transform -1 0 19596 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0959_
timestamp 1713545776
transform 1 0 1656 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0960_
timestamp 1713545776
transform -1 0 2300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0961_
timestamp 1713545776
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0962_
timestamp 1713545776
transform -1 0 3036 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0963_
timestamp 1713545776
transform 1 0 4876 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0964_
timestamp 1713545776
transform -1 0 1656 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0965_
timestamp 1713545776
transform 1 0 1656 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1713545776
transform 1 0 2300 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0967_
timestamp 1713545776
transform 1 0 1840 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0968_
timestamp 1713545776
transform 1 0 1472 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0969_
timestamp 1713545776
transform -1 0 2576 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0970_
timestamp 1713545776
transform -1 0 2852 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0971_
timestamp 1713545776
transform -1 0 2116 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0972_
timestamp 1713545776
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0973_
timestamp 1713545776
transform -1 0 2576 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0974_
timestamp 1713545776
transform -1 0 2116 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0975_
timestamp 1713545776
transform -1 0 1840 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0976_
timestamp 1713545776
transform 1 0 1196 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1713545776
transform 1 0 1932 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1713545776
transform 1 0 1840 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1713545776
transform -1 0 2944 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0980_
timestamp 1713545776
transform 1 0 1656 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0981_
timestamp 1713545776
transform 1 0 2024 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0982_
timestamp 1713545776
transform 1 0 1472 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1713545776
transform -1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0984_
timestamp 1713545776
transform 1 0 3220 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0985_
timestamp 1713545776
transform 1 0 2668 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0986_
timestamp 1713545776
transform -1 0 3128 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0987_
timestamp 1713545776
transform 1 0 16192 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1713545776
transform -1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0989_
timestamp 1713545776
transform -1 0 19412 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 1713545776
transform 1 0 16100 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1713545776
transform 1 0 14536 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0992_
timestamp 1713545776
transform 1 0 16284 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1713545776
transform 1 0 6348 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp 1713545776
transform 1 0 16100 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1713545776
transform 1 0 6900 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 1713545776
transform -1 0 20148 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1713545776
transform 1 0 19872 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1713545776
transform 1 0 18032 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1713545776
transform -1 0 12328 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 1713545776
transform -1 0 19688 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1713545776
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp 1713545776
transform -1 0 18952 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1713545776
transform -1 0 20240 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1713545776
transform 1 0 19872 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1713545776
transform 1 0 20240 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1006_
timestamp 1713545776
transform -1 0 20424 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1007_
timestamp 1713545776
transform 1 0 19596 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1008_
timestamp 1713545776
transform -1 0 21344 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1009_
timestamp 1713545776
transform 1 0 19504 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1010_
timestamp 1713545776
transform -1 0 20608 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1011_
timestamp 1713545776
transform 1 0 18124 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1012_
timestamp 1713545776
transform -1 0 18952 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1713545776
transform 1 0 18952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1014_
timestamp 1713545776
transform -1 0 20148 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1015_
timestamp 1713545776
transform -1 0 19136 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1016_
timestamp 1713545776
transform 1 0 18308 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1017_
timestamp 1713545776
transform -1 0 17848 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1018_
timestamp 1713545776
transform -1 0 18308 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 1713545776
transform -1 0 18216 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1020_
timestamp 1713545776
transform 1 0 18676 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1021_
timestamp 1713545776
transform -1 0 19136 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1022_
timestamp 1713545776
transform 1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1023_
timestamp 1713545776
transform -1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1024_
timestamp 1713545776
transform 1 0 17296 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1025_
timestamp 1713545776
transform 1 0 17664 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1026_
timestamp 1713545776
transform -1 0 19320 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1027_
timestamp 1713545776
transform -1 0 18952 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1028_
timestamp 1713545776
transform 1 0 17940 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1029_
timestamp 1713545776
transform 1 0 18400 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1030_
timestamp 1713545776
transform -1 0 18952 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1713545776
transform 1 0 18676 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1032_
timestamp 1713545776
transform 1 0 18676 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1713545776
transform 1 0 20148 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1034_
timestamp 1713545776
transform -1 0 19688 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1035_
timestamp 1713545776
transform -1 0 18400 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1036_
timestamp 1713545776
transform 1 0 20700 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1713545776
transform -1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1038_
timestamp 1713545776
transform 1 0 19596 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1039_
timestamp 1713545776
transform -1 0 20700 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1713545776
transform -1 0 20976 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1041_
timestamp 1713545776
transform -1 0 17296 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _1042_
timestamp 1713545776
transform 1 0 16284 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__or4b_1  _1043_
timestamp 1713545776
transform 1 0 19688 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1044_
timestamp 1713545776
transform 1 0 20424 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1713545776
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1046_
timestamp 1713545776
transform 1 0 17020 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1047_
timestamp 1713545776
transform 1 0 22632 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1048_
timestamp 1713545776
transform -1 0 21528 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1049_
timestamp 1713545776
transform 1 0 20884 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1050_
timestamp 1713545776
transform -1 0 22356 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 1713545776
transform -1 0 22632 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1052_
timestamp 1713545776
transform 1 0 18032 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1053_
timestamp 1713545776
transform -1 0 21896 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1054_
timestamp 1713545776
transform 1 0 20608 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1713545776
transform 1 0 21160 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1056_
timestamp 1713545776
transform -1 0 22816 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1057_
timestamp 1713545776
transform 1 0 21528 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1058_
timestamp 1713545776
transform 1 0 21620 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1059_
timestamp 1713545776
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1713545776
transform 1 0 828 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1713545776
transform 1 0 21436 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1713545776
transform 1 0 19688 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1713545776
transform 1 0 2208 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1713545776
transform -1 0 5060 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1713545776
transform 1 0 5796 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1713545776
transform 1 0 8372 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1713545776
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1713545776
transform 1 0 7728 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1713545776
transform 1 0 920 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1713545776
transform 1 0 1104 0 -1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1713545776
transform 1 0 1380 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1713545776
transform 1 0 1288 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1713545776
transform 1 0 2300 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1713545776
transform 1 0 828 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1713545776
transform 1 0 1196 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1713545776
transform 1 0 2576 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1713545776
transform 1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1713545776
transform 1 0 3496 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1713545776
transform -1 0 17572 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1713545776
transform 1 0 13800 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1713545776
transform -1 0 6348 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1713545776
transform 1 0 4232 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1713545776
transform 1 0 19688 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1713545776
transform 1 0 12328 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1713545776
transform 1 0 21620 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1713545776
transform 1 0 20148 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1713545776
transform 1 0 21252 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1713545776
transform 1 0 21252 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1713545776
transform 1 0 19688 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1713545776
transform 1 0 21436 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1713545776
transform 1 0 8096 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1092_
timestamp 1713545776
transform 1 0 18952 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1713545776
transform -1 0 20148 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1713545776
transform 1 0 21252 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1713545776
transform 1 0 21160 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1713545776
transform 1 0 21344 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1713545776
transform 1 0 21620 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1713545776
transform 1 0 1656 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1099_
timestamp 1713545776
transform 1 0 1380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1100_
timestamp 1713545776
transform -1 0 9108 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1101_
timestamp 1713545776
transform 1 0 9568 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1713545776
transform -1 0 17480 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1103_
timestamp 1713545776
transform -1 0 15180 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1713545776
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1713545776
transform -1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1713545776
transform -1 0 13800 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1713545776
transform -1 0 7544 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1713545776
transform -1 0 7912 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1713545776
transform 1 0 17296 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1713545776
transform 1 0 17480 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3
timestamp 1713545776
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_8
timestamp 1713545776
transform 1 0 1288 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 1713545776
transform 1 0 2852 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_39
timestamp 1713545776
transform 1 0 4140 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_44
timestamp 1713545776
transform 1 0 4600 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_48
timestamp 1713545776
transform 1 0 4968 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1713545776
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57
timestamp 1713545776
transform 1 0 5796 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_62
timestamp 1713545776
transform 1 0 6256 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_74
timestamp 1713545776
transform 1 0 7360 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1713545776
transform 1 0 8096 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1713545776
transform 1 0 8740 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1713545776
transform 1 0 9108 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_101
timestamp 1713545776
transform 1 0 9844 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_107
timestamp 1713545776
transform 1 0 10396 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1713545776
transform 1 0 10764 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_119
timestamp 1713545776
transform 1 0 11500 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_134
timestamp 1713545776
transform 1 0 12880 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_145
timestamp 1713545776
transform 1 0 13892 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_152
timestamp 1713545776
transform 1 0 14536 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_164
timestamp 1713545776
transform 1 0 15640 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_179
timestamp 1713545776
transform 1 0 17020 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_183
timestamp 1713545776
transform 1 0 17388 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_188
timestamp 1713545776
transform 1 0 17848 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_209
timestamp 1713545776
transform 1 0 19780 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_215
timestamp 1713545776
transform 1 0 20332 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_219
timestamp 1713545776
transform 1 0 20700 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_225
timestamp 1713545776
transform 1 0 21252 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_243
timestamp 1713545776
transform 1 0 22908 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_9
timestamp 1713545776
transform 1 0 1380 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_17
timestamp 1713545776
transform 1 0 2116 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_44
timestamp 1713545776
transform 1 0 4600 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_53
timestamp 1713545776
transform 1 0 5428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1713545776
transform 1 0 5796 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 1713545776
transform 1 0 6164 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_67
timestamp 1713545776
transform 1 0 6716 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_75
timestamp 1713545776
transform 1 0 7452 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_91
timestamp 1713545776
transform 1 0 8924 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_98
timestamp 1713545776
transform 1 0 9568 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1713545776
transform 1 0 10948 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_122
timestamp 1713545776
transform 1 0 11776 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_132
timestamp 1713545776
transform 1 0 12696 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_203
timestamp 1713545776
transform 1 0 19228 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_207
timestamp 1713545776
transform 1 0 19596 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_242
timestamp 1713545776
transform 1 0 22816 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_3
timestamp 1713545776
transform 1 0 828 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1713545776
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1713545776
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_29
timestamp 1713545776
transform 1 0 3220 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_61
timestamp 1713545776
transform 1 0 6164 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_68
timestamp 1713545776
transform 1 0 6808 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_97
timestamp 1713545776
transform 1 0 9476 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_103
timestamp 1713545776
transform 1 0 10028 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_120
timestamp 1713545776
transform 1 0 11592 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_126
timestamp 1713545776
transform 1 0 12144 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_130
timestamp 1713545776
transform 1 0 12512 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_145
timestamp 1713545776
transform 1 0 13892 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_155
timestamp 1713545776
transform 1 0 14812 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_176
timestamp 1713545776
transform 1 0 16744 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_186
timestamp 1713545776
transform 1 0 17664 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1713545776
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_203
timestamp 1713545776
transform 1 0 19228 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_215
timestamp 1713545776
transform 1 0 20332 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_236
timestamp 1713545776
transform 1 0 22264 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_244
timestamp 1713545776
transform 1 0 23000 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_3
timestamp 1713545776
transform 1 0 828 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_23
timestamp 1713545776
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_38
timestamp 1713545776
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1713545776
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1713545776
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1713545776
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1713545776
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_93
timestamp 1713545776
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_101
timestamp 1713545776
transform 1 0 9844 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_108
timestamp 1713545776
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_130
timestamp 1713545776
transform 1 0 12512 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_134
timestamp 1713545776
transform 1 0 12880 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_138
timestamp 1713545776
transform 1 0 13248 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_150
timestamp 1713545776
transform 1 0 14352 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_162
timestamp 1713545776
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_177
timestamp 1713545776
transform 1 0 16836 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_189
timestamp 1713545776
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_195
timestamp 1713545776
transform 1 0 18492 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_211
timestamp 1713545776
transform 1 0 19964 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1713545776
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 1713545776
transform 1 0 21252 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_243
timestamp 1713545776
transform 1 0 22908 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3
timestamp 1713545776
transform 1 0 828 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_12
timestamp 1713545776
transform 1 0 1656 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_16
timestamp 1713545776
transform 1 0 2024 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1713545776
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_34
timestamp 1713545776
transform 1 0 3680 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_46
timestamp 1713545776
transform 1 0 4784 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_58
timestamp 1713545776
transform 1 0 5888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_62
timestamp 1713545776
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_70
timestamp 1713545776
transform 1 0 6992 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_74
timestamp 1713545776
transform 1 0 7360 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1713545776
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_85
timestamp 1713545776
transform 1 0 8372 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_101
timestamp 1713545776
transform 1 0 9844 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_107
timestamp 1713545776
transform 1 0 10396 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_118
timestamp 1713545776
transform 1 0 11408 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_130
timestamp 1713545776
transform 1 0 12512 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1713545776
transform 1 0 17204 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1713545776
transform 1 0 18308 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_202
timestamp 1713545776
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_216
timestamp 1713545776
transform 1 0 20424 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_222
timestamp 1713545776
transform 1 0 20976 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_226
timestamp 1713545776
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_238
timestamp 1713545776
transform 1 0 22448 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_244
timestamp 1713545776
transform 1 0 23000 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_3
timestamp 1713545776
transform 1 0 828 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_20
timestamp 1713545776
transform 1 0 2392 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_27
timestamp 1713545776
transform 1 0 3036 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1713545776
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_71
timestamp 1713545776
transform 1 0 7084 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1713545776
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_121
timestamp 1713545776
transform 1 0 11684 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_130
timestamp 1713545776
transform 1 0 12512 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_146
timestamp 1713545776
transform 1 0 13984 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 1713545776
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_172
timestamp 1713545776
transform 1 0 16376 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_180
timestamp 1713545776
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_185
timestamp 1713545776
transform 1 0 17572 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_198
timestamp 1713545776
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_205
timestamp 1713545776
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_215
timestamp 1713545776
transform 1 0 20332 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1713545776
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_241
timestamp 1713545776
transform 1 0 22724 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 1713545776
transform 1 0 828 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_11
timestamp 1713545776
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_17
timestamp 1713545776
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_24
timestamp 1713545776
transform 1 0 2760 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1713545776
transform 1 0 3220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_37
timestamp 1713545776
transform 1 0 3956 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_45
timestamp 1713545776
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_54
timestamp 1713545776
transform 1 0 5520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_66
timestamp 1713545776
transform 1 0 6624 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_74
timestamp 1713545776
transform 1 0 7360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1713545776
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_88
timestamp 1713545776
transform 1 0 8648 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_105
timestamp 1713545776
transform 1 0 10212 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_117
timestamp 1713545776
transform 1 0 11316 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_129
timestamp 1713545776
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_156
timestamp 1713545776
transform 1 0 14904 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_174
timestamp 1713545776
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_186
timestamp 1713545776
transform 1 0 17664 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_192
timestamp 1713545776
transform 1 0 18216 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_207
timestamp 1713545776
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_242
timestamp 1713545776
transform 1 0 22816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1713545776
transform 1 0 828 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_7
timestamp 1713545776
transform 1 0 1196 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_24
timestamp 1713545776
transform 1 0 2760 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_30
timestamp 1713545776
transform 1 0 3312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_49
timestamp 1713545776
transform 1 0 5060 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1713545776
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_60
timestamp 1713545776
transform 1 0 6072 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_66
timestamp 1713545776
transform 1 0 6624 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_79
timestamp 1713545776
transform 1 0 7820 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_91
timestamp 1713545776
transform 1 0 8924 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_103
timestamp 1713545776
transform 1 0 10028 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_113
timestamp 1713545776
transform 1 0 10948 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_124
timestamp 1713545776
transform 1 0 11960 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_132
timestamp 1713545776
transform 1 0 12696 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_139
timestamp 1713545776
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_151
timestamp 1713545776
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_178
timestamp 1713545776
transform 1 0 16928 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_196
timestamp 1713545776
transform 1 0 18584 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_202
timestamp 1713545776
transform 1 0 19136 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_210
timestamp 1713545776
transform 1 0 19872 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_216
timestamp 1713545776
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_241
timestamp 1713545776
transform 1 0 22724 0 -1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1713545776
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_22
timestamp 1713545776
transform 1 0 2576 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1713545776
transform 1 0 3220 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_47
timestamp 1713545776
transform 1 0 4876 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_73
timestamp 1713545776
transform 1 0 7268 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1713545776
transform 1 0 8004 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_91
timestamp 1713545776
transform 1 0 8924 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_103
timestamp 1713545776
transform 1 0 10028 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_127
timestamp 1713545776
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_136
timestamp 1713545776
transform 1 0 13064 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_151
timestamp 1713545776
transform 1 0 14444 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_172
timestamp 1713545776
transform 1 0 16376 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_184
timestamp 1713545776
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_189
timestamp 1713545776
transform 1 0 17940 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_200
timestamp 1713545776
transform 1 0 18952 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_212
timestamp 1713545776
transform 1 0 20056 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_220
timestamp 1713545776
transform 1 0 20792 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_235
timestamp 1713545776
transform 1 0 22172 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_243
timestamp 1713545776
transform 1 0 22908 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1713545776
transform 1 0 828 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_11
timestamp 1713545776
transform 1 0 1564 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_35
timestamp 1713545776
transform 1 0 3772 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1713545776
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_73
timestamp 1713545776
transform 1 0 7268 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_96
timestamp 1713545776
transform 1 0 9384 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_108
timestamp 1713545776
transform 1 0 10488 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_121
timestamp 1713545776
transform 1 0 11684 0 -1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_147
timestamp 1713545776
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1713545776
transform 1 0 15732 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 1713545776
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_183
timestamp 1713545776
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_203
timestamp 1713545776
transform 1 0 19228 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_207
timestamp 1713545776
transform 1 0 19596 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1713545776
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_239
timestamp 1713545776
transform 1 0 22540 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1713545776
transform 1 0 828 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_9
timestamp 1713545776
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1713545776
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1713545776
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1713545776
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_53
timestamp 1713545776
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_75
timestamp 1713545776
transform 1 0 7452 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1713545776
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_92
timestamp 1713545776
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_104
timestamp 1713545776
transform 1 0 10120 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_131
timestamp 1713545776
transform 1 0 12604 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1713545776
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_147
timestamp 1713545776
transform 1 0 14076 0 1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_173
timestamp 1713545776
transform 1 0 16468 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_185
timestamp 1713545776
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_192
timestamp 1713545776
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_204
timestamp 1713545776
transform 1 0 19320 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_216
timestamp 1713545776
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_220
timestamp 1713545776
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_243
timestamp 1713545776
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1713545776
transform 1 0 828 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_11
timestamp 1713545776
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_17
timestamp 1713545776
transform 1 0 2116 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_34
timestamp 1713545776
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_38
timestamp 1713545776
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1713545776
transform 1 0 4692 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1713545776
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp 1713545776
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_78
timestamp 1713545776
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_98
timestamp 1713545776
transform 1 0 9568 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_106
timestamp 1713545776
transform 1 0 10304 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_129
timestamp 1713545776
transform 1 0 12420 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_137
timestamp 1713545776
transform 1 0 13156 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_150
timestamp 1713545776
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_158
timestamp 1713545776
transform 1 0 15088 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1713545776
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_169
timestamp 1713545776
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_173
timestamp 1713545776
transform 1 0 16468 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_177
timestamp 1713545776
transform 1 0 16836 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_181
timestamp 1713545776
transform 1 0 17204 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_186
timestamp 1713545776
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_198
timestamp 1713545776
transform 1 0 18768 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_210
timestamp 1713545776
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_218
timestamp 1713545776
transform 1 0 20608 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_234
timestamp 1713545776
transform 1 0 22080 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_242
timestamp 1713545776
transform 1 0 22816 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1713545776
transform 1 0 828 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_12
timestamp 1713545776
transform 1 0 1656 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1713545776
transform 1 0 7544 0 1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1713545776
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_97
timestamp 1713545776
transform 1 0 9476 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_101
timestamp 1713545776
transform 1 0 9844 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_127
timestamp 1713545776
transform 1 0 12236 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_164
timestamp 1713545776
transform 1 0 15640 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_188
timestamp 1713545776
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_217
timestamp 1713545776
transform 1 0 20516 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_224
timestamp 1713545776
transform 1 0 21160 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_236
timestamp 1713545776
transform 1 0 22264 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_244
timestamp 1713545776
transform 1 0 23000 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_19
timestamp 1713545776
transform 1 0 2300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_23
timestamp 1713545776
transform 1 0 2668 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_35
timestamp 1713545776
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_39
timestamp 1713545776
transform 1 0 4140 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_47
timestamp 1713545776
transform 1 0 4876 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1713545776
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_75
timestamp 1713545776
transform 1 0 7452 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_87
timestamp 1713545776
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 1713545776
transform 1 0 9936 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1713545776
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1713545776
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1713545776
transform 1 0 15640 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_169
timestamp 1713545776
transform 1 0 16100 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_202
timestamp 1713545776
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_206
timestamp 1713545776
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp 1713545776
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_242
timestamp 1713545776
transform 1 0 22816 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1713545776
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_15
timestamp 1713545776
transform 1 0 1932 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_35
timestamp 1713545776
transform 1 0 3772 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_43
timestamp 1713545776
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_48
timestamp 1713545776
transform 1 0 4968 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 1713545776
transform 1 0 7360 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1713545776
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_98
timestamp 1713545776
transform 1 0 9568 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_110
timestamp 1713545776
transform 1 0 10672 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_129
timestamp 1713545776
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_133
timestamp 1713545776
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_141
timestamp 1713545776
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_186
timestamp 1713545776
transform 1 0 17664 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1713545776
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_202
timestamp 1713545776
transform 1 0 19136 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_208
timestamp 1713545776
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_222
timestamp 1713545776
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_243
timestamp 1713545776
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1713545776
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_30
timestamp 1713545776
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_42
timestamp 1713545776
transform 1 0 4416 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1713545776
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1713545776
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_62
timestamp 1713545776
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_74
timestamp 1713545776
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_86
timestamp 1713545776
transform 1 0 8464 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_107
timestamp 1713545776
transform 1 0 10396 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1713545776
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_152
timestamp 1713545776
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1713545776
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_173
timestamp 1713545776
transform 1 0 16468 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_191
timestamp 1713545776
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_196
timestamp 1713545776
transform 1 0 18584 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_204
timestamp 1713545776
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_216
timestamp 1713545776
transform 1 0 20424 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_235
timestamp 1713545776
transform 1 0 22172 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_243
timestamp 1713545776
transform 1 0 22908 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1713545776
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_15
timestamp 1713545776
transform 1 0 1932 0 1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_35
timestamp 1713545776
transform 1 0 3772 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_72
timestamp 1713545776
transform 1 0 7176 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_101
timestamp 1713545776
transform 1 0 9844 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_109
timestamp 1713545776
transform 1 0 10580 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_115
timestamp 1713545776
transform 1 0 11132 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1713545776
transform 1 0 13156 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_181
timestamp 1713545776
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1713545776
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_215
timestamp 1713545776
transform 1 0 20332 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_242
timestamp 1713545776
transform 1 0 22816 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_3
timestamp 1713545776
transform 1 0 828 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_32
timestamp 1713545776
transform 1 0 3496 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_47
timestamp 1713545776
transform 1 0 4876 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_51
timestamp 1713545776
transform 1 0 5244 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1713545776
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_57
timestamp 1713545776
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_80
timestamp 1713545776
transform 1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_95
timestamp 1713545776
transform 1 0 9292 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_103
timestamp 1713545776
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_121
timestamp 1713545776
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_133
timestamp 1713545776
transform 1 0 12788 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_143
timestamp 1713545776
transform 1 0 13708 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_151
timestamp 1713545776
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_156
timestamp 1713545776
transform 1 0 14904 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_169
timestamp 1713545776
transform 1 0 16100 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_183
timestamp 1713545776
transform 1 0 17388 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_208
timestamp 1713545776
transform 1 0 19688 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_219
timestamp 1713545776
transform 1 0 20700 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1713545776
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_240
timestamp 1713545776
transform 1 0 22632 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_244
timestamp 1713545776
transform 1 0 23000 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1713545776
transform 1 0 828 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_11
timestamp 1713545776
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_17
timestamp 1713545776
transform 1 0 2116 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_25
timestamp 1713545776
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 1713545776
transform 1 0 3220 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_33
timestamp 1713545776
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_52
timestamp 1713545776
transform 1 0 5336 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_70
timestamp 1713545776
transform 1 0 6992 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1713545776
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_98
timestamp 1713545776
transform 1 0 9568 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_110
timestamp 1713545776
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_127
timestamp 1713545776
transform 1 0 12236 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_178
timestamp 1713545776
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_186
timestamp 1713545776
transform 1 0 17664 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1713545776
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_197
timestamp 1713545776
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_216
timestamp 1713545776
transform 1 0 20424 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_236
timestamp 1713545776
transform 1 0 22264 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_244
timestamp 1713545776
transform 1 0 23000 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1713545776
transform 1 0 828 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_23
timestamp 1713545776
transform 1 0 2668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_32
timestamp 1713545776
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_47
timestamp 1713545776
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1713545776
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_75
timestamp 1713545776
transform 1 0 7452 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_79
timestamp 1713545776
transform 1 0 7820 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_91
timestamp 1713545776
transform 1 0 8924 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_98
timestamp 1713545776
transform 1 0 9568 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_106
timestamp 1713545776
transform 1 0 10304 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1713545776
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1713545776
transform 1 0 10948 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_130
timestamp 1713545776
transform 1 0 12512 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1713545776
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_172
timestamp 1713545776
transform 1 0 16376 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_186
timestamp 1713545776
transform 1 0 17664 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_200
timestamp 1713545776
transform 1 0 18952 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_208
timestamp 1713545776
transform 1 0 19688 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_241
timestamp 1713545776
transform 1 0 22724 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1713545776
transform 1 0 828 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_14
timestamp 1713545776
transform 1 0 1840 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_22
timestamp 1713545776
transform 1 0 2576 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_39
timestamp 1713545776
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_50
timestamp 1713545776
transform 1 0 5152 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_58
timestamp 1713545776
transform 1 0 5888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_63
timestamp 1713545776
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_69
timestamp 1713545776
transform 1 0 6900 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1713545776
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1713545776
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_97
timestamp 1713545776
transform 1 0 9476 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_103
timestamp 1713545776
transform 1 0 10028 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_123
timestamp 1713545776
transform 1 0 11868 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_135
timestamp 1713545776
transform 1 0 12972 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1713545776
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_154
timestamp 1713545776
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_162
timestamp 1713545776
transform 1 0 15456 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_166
timestamp 1713545776
transform 1 0 15824 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_179
timestamp 1713545776
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_185
timestamp 1713545776
transform 1 0 17572 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1713545776
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_205
timestamp 1713545776
transform 1 0 19412 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_217
timestamp 1713545776
transform 1 0 20516 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_223
timestamp 1713545776
transform 1 0 21068 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_240
timestamp 1713545776
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_244
timestamp 1713545776
transform 1 0 23000 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1713545776
transform 1 0 828 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_11
timestamp 1713545776
transform 1 0 1564 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_37
timestamp 1713545776
transform 1 0 3956 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_41
timestamp 1713545776
transform 1 0 4324 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_45
timestamp 1713545776
transform 1 0 4692 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_67
timestamp 1713545776
transform 1 0 6716 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_94
timestamp 1713545776
transform 1 0 9200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_103
timestamp 1713545776
transform 1 0 10028 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_120
timestamp 1713545776
transform 1 0 11592 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_147
timestamp 1713545776
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_159
timestamp 1713545776
transform 1 0 15180 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_185
timestamp 1713545776
transform 1 0 17572 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_193
timestamp 1713545776
transform 1 0 18308 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_213
timestamp 1713545776
transform 1 0 20148 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 1713545776
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1713545776
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_237
timestamp 1713545776
transform 1 0 22356 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 1713545776
transform 1 0 828 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_48
timestamp 1713545776
transform 1 0 4968 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1713545776
transform 1 0 8372 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_93
timestamp 1713545776
transform 1 0 9108 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_100
timestamp 1713545776
transform 1 0 9752 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_108
timestamp 1713545776
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_122
timestamp 1713545776
transform 1 0 11776 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_154
timestamp 1713545776
transform 1 0 14720 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_166
timestamp 1713545776
transform 1 0 15824 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_176
timestamp 1713545776
transform 1 0 16744 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_188
timestamp 1713545776
transform 1 0 17848 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_210
timestamp 1713545776
transform 1 0 19872 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_238
timestamp 1713545776
transform 1 0 22448 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1713545776
transform 1 0 828 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_11
timestamp 1713545776
transform 1 0 1564 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_35
timestamp 1713545776
transform 1 0 3772 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_47
timestamp 1713545776
transform 1 0 4876 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1713545776
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1713545776
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_66
timestamp 1713545776
transform 1 0 6624 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_74
timestamp 1713545776
transform 1 0 7360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_80
timestamp 1713545776
transform 1 0 7912 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_88
timestamp 1713545776
transform 1 0 8648 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_92
timestamp 1713545776
transform 1 0 9016 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_122
timestamp 1713545776
transform 1 0 11776 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_134
timestamp 1713545776
transform 1 0 12880 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_146
timestamp 1713545776
transform 1 0 13984 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_158
timestamp 1713545776
transform 1 0 15088 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1713545776
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_181
timestamp 1713545776
transform 1 0 17204 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_200
timestamp 1713545776
transform 1 0 18952 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_205
timestamp 1713545776
transform 1 0 19412 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_214
timestamp 1713545776
transform 1 0 20240 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1713545776
transform 1 0 20976 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1713545776
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 1713545776
transform 1 0 828 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_11
timestamp 1713545776
transform 1 0 1564 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_18
timestamp 1713545776
transform 1 0 2208 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_22
timestamp 1713545776
transform 1 0 2576 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1713545776
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1713545776
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_41
timestamp 1713545776
transform 1 0 4324 0 1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_67
timestamp 1713545776
transform 1 0 6716 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1713545776
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_94
timestamp 1713545776
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_101
timestamp 1713545776
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_122
timestamp 1713545776
transform 1 0 11776 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_134
timestamp 1713545776
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1713545776
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1713545776
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_147
timestamp 1713545776
transform 1 0 14076 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_151
timestamp 1713545776
transform 1 0 14444 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_155
timestamp 1713545776
transform 1 0 14812 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_186
timestamp 1713545776
transform 1 0 17664 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1713545776
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_202
timestamp 1713545776
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_213
timestamp 1713545776
transform 1 0 20148 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_217
timestamp 1713545776
transform 1 0 20516 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_222
timestamp 1713545776
transform 1 0 20976 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_234
timestamp 1713545776
transform 1 0 22080 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_242
timestamp 1713545776
transform 1 0 22816 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_38
timestamp 1713545776
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1713545776
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_72
timestamp 1713545776
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_88
timestamp 1713545776
transform 1 0 8648 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_94
timestamp 1713545776
transform 1 0 9200 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_119
timestamp 1713545776
transform 1 0 11500 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_160
timestamp 1713545776
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_225
timestamp 1713545776
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1713545776
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_15
timestamp 1713545776
transform 1 0 1932 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1713545776
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1713545776
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_41
timestamp 1713545776
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_47
timestamp 1713545776
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_55
timestamp 1713545776
transform 1 0 5612 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_57
timestamp 1713545776
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_63
timestamp 1713545776
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_71
timestamp 1713545776
transform 1 0 7084 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1713545776
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_95
timestamp 1713545776
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_103
timestamp 1713545776
transform 1 0 10028 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_111
timestamp 1713545776
transform 1 0 10764 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_119
timestamp 1713545776
transform 1 0 11500 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_131
timestamp 1713545776
transform 1 0 12604 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1713545776
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_151
timestamp 1713545776
transform 1 0 14444 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_163
timestamp 1713545776
transform 1 0 15548 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_167
timestamp 1713545776
transform 1 0 15916 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_178
timestamp 1713545776
transform 1 0 16928 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_186
timestamp 1713545776
transform 1 0 17664 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_190
timestamp 1713545776
transform 1 0 18032 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_200
timestamp 1713545776
transform 1 0 18952 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_206
timestamp 1713545776
transform 1 0 19504 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_216
timestamp 1713545776
transform 1 0 20424 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_222
timestamp 1713545776
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_234
timestamp 1713545776
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_238
timestamp 1713545776
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1713545776
transform 1 0 2300 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1713545776
transform -1 0 23092 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1713545776
transform -1 0 23092 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1713545776
transform -1 0 22448 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1713545776
transform -1 0 22080 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1713545776
transform -1 0 20976 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1713545776
transform 1 0 20148 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1713545776
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1713545776
transform -1 0 18952 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1713545776
transform -1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1713545776
transform -1 0 7084 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1713545776
transform -1 0 10028 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1713545776
transform -1 0 6256 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1713545776
transform -1 0 5428 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1713545776
transform -1 0 4600 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1713545776
transform -1 0 3588 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1713545776
transform -1 0 4140 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1713545776
transform -1 0 2116 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1713545776
transform -1 0 1288 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1713545776
transform -1 0 1380 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1713545776
transform -1 0 7820 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1713545776
transform -1 0 10764 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1713545776
transform -1 0 14536 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1713545776
transform 1 0 13524 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1713545776
transform -1 0 12880 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1713545776
transform 1 0 12144 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1713545776
transform 1 0 10948 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1713545776
transform 1 0 10028 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1713545776
transform 1 0 9200 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1713545776
transform -1 0 8740 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1713545776
transform -1 0 4876 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1713545776
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1713545776
transform -1 0 8924 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1713545776
transform -1 0 11500 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1713545776
transform 1 0 22448 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1713545776
transform 1 0 22540 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1713545776
transform 1 0 20792 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1713545776
transform 1 0 19964 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1713545776
transform 1 0 19228 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1713545776
transform 1 0 18216 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1713545776
transform 1 0 17480 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1713545776
transform 1 0 16652 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1713545776
transform -1 0 5612 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1713545776
transform 1 0 8924 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_27
timestamp 1713545776
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1713545776
transform -1 0 23368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_28
timestamp 1713545776
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1713545776
transform -1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_29
timestamp 1713545776
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1713545776
transform -1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_30
timestamp 1713545776
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1713545776
transform -1 0 23368 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_31
timestamp 1713545776
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1713545776
transform -1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_32
timestamp 1713545776
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1713545776
transform -1 0 23368 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_33
timestamp 1713545776
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1713545776
transform -1 0 23368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_34
timestamp 1713545776
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1713545776
transform -1 0 23368 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_35
timestamp 1713545776
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1713545776
transform -1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_36
timestamp 1713545776
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1713545776
transform -1 0 23368 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_37
timestamp 1713545776
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1713545776
transform -1 0 23368 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_38
timestamp 1713545776
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1713545776
transform -1 0 23368 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_39
timestamp 1713545776
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1713545776
transform -1 0 23368 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_40
timestamp 1713545776
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1713545776
transform -1 0 23368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_41
timestamp 1713545776
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1713545776
transform -1 0 23368 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_42
timestamp 1713545776
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1713545776
transform -1 0 23368 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_43
timestamp 1713545776
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1713545776
transform -1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_44
timestamp 1713545776
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1713545776
transform -1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_45
timestamp 1713545776
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1713545776
transform -1 0 23368 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_46
timestamp 1713545776
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1713545776
transform -1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_47
timestamp 1713545776
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1713545776
transform -1 0 23368 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_48
timestamp 1713545776
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1713545776
transform -1 0 23368 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_49
timestamp 1713545776
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1713545776
transform -1 0 23368 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_50
timestamp 1713545776
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1713545776
transform -1 0 23368 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_51
timestamp 1713545776
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1713545776
transform -1 0 23368 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_52
timestamp 1713545776
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1713545776
transform -1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_53
timestamp 1713545776
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1713545776
transform -1 0 23368 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_54
timestamp 1713545776
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_55
timestamp 1713545776
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 1713545776
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1713545776
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1713545776
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1713545776
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1713545776
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1713545776
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 1713545776
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp 1713545776
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 1713545776
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_65
timestamp 1713545776
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp 1713545776
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 1713545776
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_68
timestamp 1713545776
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_69
timestamp 1713545776
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 1713545776
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_71
timestamp 1713545776
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_72
timestamp 1713545776
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_73
timestamp 1713545776
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_74
timestamp 1713545776
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp 1713545776
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_76
timestamp 1713545776
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 1713545776
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp 1713545776
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp 1713545776
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp 1713545776
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp 1713545776
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_82
timestamp 1713545776
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp 1713545776
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp 1713545776
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp 1713545776
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp 1713545776
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_87
timestamp 1713545776
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp 1713545776
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_89
timestamp 1713545776
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp 1713545776
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp 1713545776
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp 1713545776
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp 1713545776
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp 1713545776
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp 1713545776
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp 1713545776
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp 1713545776
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_98
timestamp 1713545776
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_99
timestamp 1713545776
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_100
timestamp 1713545776
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp 1713545776
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_102
timestamp 1713545776
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_103
timestamp 1713545776
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_104
timestamp 1713545776
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_105
timestamp 1713545776
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_106
timestamp 1713545776
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_107
timestamp 1713545776
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_108
timestamp 1713545776
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_109
timestamp 1713545776
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_110
timestamp 1713545776
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_111
timestamp 1713545776
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_112
timestamp 1713545776
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_113
timestamp 1713545776
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_114
timestamp 1713545776
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_115
timestamp 1713545776
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_116
timestamp 1713545776
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_117
timestamp 1713545776
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_118
timestamp 1713545776
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_119
timestamp 1713545776
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_120
timestamp 1713545776
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_121
timestamp 1713545776
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_122
timestamp 1713545776
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_123
timestamp 1713545776
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_124
timestamp 1713545776
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_125
timestamp 1713545776
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_126
timestamp 1713545776
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_127
timestamp 1713545776
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_128
timestamp 1713545776
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_129
timestamp 1713545776
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_130
timestamp 1713545776
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_131
timestamp 1713545776
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_132
timestamp 1713545776
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_133
timestamp 1713545776
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_134
timestamp 1713545776
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_135
timestamp 1713545776
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_136
timestamp 1713545776
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_137
timestamp 1713545776
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_138
timestamp 1713545776
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_139
timestamp 1713545776
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_140
timestamp 1713545776
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_141
timestamp 1713545776
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_142
timestamp 1713545776
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_143
timestamp 1713545776
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_144
timestamp 1713545776
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_145
timestamp 1713545776
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_146
timestamp 1713545776
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_147
timestamp 1713545776
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_148
timestamp 1713545776
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_149
timestamp 1713545776
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_150
timestamp 1713545776
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_151
timestamp 1713545776
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_152
timestamp 1713545776
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_153
timestamp 1713545776
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_154
timestamp 1713545776
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_155
timestamp 1713545776
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_156
timestamp 1713545776
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_157
timestamp 1713545776
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_158
timestamp 1713545776
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_159
timestamp 1713545776
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_160
timestamp 1713545776
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_161
timestamp 1713545776
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_162
timestamp 1713545776
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_163
timestamp 1713545776
transform 1 0 5704 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_164
timestamp 1713545776
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_165
timestamp 1713545776
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_166
timestamp 1713545776
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_167
timestamp 1713545776
transform 1 0 16008 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_168
timestamp 1713545776
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_169
timestamp 1713545776
transform 1 0 21160 0 1 14688
box -38 -48 130 592
<< labels >>
rlabel metal1 s 11960 14688 11960 14688 4 VGND
rlabel metal1 s 11960 15232 11960 15232 4 VPWR
rlabel metal1 s 1513 14450 1513 14450 4 _0000_
rlabel metal1 s 21512 2550 21512 2550 4 _0001_
rlabel metal1 s 19954 1394 19954 1394 4 _0002_
rlabel metal1 s 3818 1496 3818 1496 4 _0003_
rlabel metal1 s 5673 3638 5673 3638 4 _0004_
rlabel metal1 s 5658 5338 5658 5338 4 _0005_
rlabel metal1 s 8592 9486 8592 9486 4 _0006_
rlabel metal1 s 7309 12682 7309 12682 4 _0007_
rlabel metal1 s 8644 11322 8644 11322 4 _0008_
rlabel metal1 s 1334 3162 1334 3162 4 _0009_
rlabel metal1 s 1605 2550 1605 2550 4 _0010_
rlabel metal1 s 1789 714 1789 714 4 _0011_
rlabel metal1 s 1973 4726 1973 4726 4 _0012_
rlabel metal1 s 2520 5746 2520 5746 4 _0013_
rlabel metal1 s 1288 7514 1288 7514 4 _0014_
rlabel metal2 s 1513 11186 1513 11186 4 _0015_
rlabel metal2 s 2898 14246 2898 14246 4 _0016_
rlabel metal2 s 2617 13430 2617 13430 4 _0017_
rlabel metal1 s 3798 12648 3798 12648 4 _0018_
rlabel metal1 s 16610 12342 16610 12342 4 _0019_
rlabel metal2 s 14582 14246 14582 14246 4 _0020_
rlabel metal1 s 6133 13770 6133 13770 4 _0021_
rlabel metal1 s 4917 14450 4917 14450 4 _0022_
rlabel metal2 s 20005 14450 20005 14450 4 _0023_
rlabel metal1 s 12466 14416 12466 14416 4 _0024_
rlabel metal1 s 21834 14518 21834 14518 4 _0025_
rlabel metal2 s 20465 12750 20465 12750 4 _0026_
rlabel metal1 s 21374 3638 21374 3638 4 _0027_
rlabel metal1 s 20654 3978 20654 3978 4 _0028_
rlabel metal1 s 19718 5814 19718 5814 4 _0029_
rlabel metal1 s 21298 6120 21298 6120 4 _0030_
rlabel metal3 s 17434 7429 17434 7429 4 _0031_
rlabel metal1 s 18890 7242 18890 7242 4 _0032_
rlabel metal2 s 18722 12070 18722 12070 4 _0033_
rlabel metal1 s 21466 11254 21466 11254 4 _0034_
rlabel metal2 s 20930 11186 20930 11186 4 _0035_
rlabel metal2 s 20838 7718 20838 7718 4 _0036_
rlabel metal1 s 21742 13430 21742 13430 4 _0037_
rlabel metal1 s 16790 10030 16790 10030 4 _0038_
rlabel metal1 s 21298 10030 21298 10030 4 _0039_
rlabel metal1 s 6578 10642 6578 10642 4 _0040_
rlabel metal1 s 20102 11118 20102 11118 4 _0041_
rlabel metal1 s 16744 9486 16744 9486 4 _0042_
rlabel metal1 s 8786 13328 8786 13328 4 _0043_
rlabel metal1 s 16790 9036 16790 9036 4 _0044_
rlabel metal1 s 14490 9044 14490 9044 4 _0045_
rlabel metal1 s 17250 9690 17250 9690 4 _0046_
rlabel metal1 s 17158 10642 17158 10642 4 _0047_
rlabel metal1 s 5842 4590 5842 4590 4 _0048_
rlabel metal2 s 17894 4828 17894 4828 4 _0049_
rlabel metal2 s 18262 2176 18262 2176 4 _0050_
rlabel metal1 s 20838 6426 20838 6426 4 _0051_
rlabel metal1 s 17434 8840 17434 8840 4 _0052_
rlabel metal2 s 17342 9316 17342 9316 4 _0053_
rlabel metal2 s 22770 9656 22770 9656 4 _0054_
rlabel metal1 s 16744 10234 16744 10234 4 _0055_
rlabel metal1 s 6118 11322 6118 11322 4 _0056_
rlabel metal3 s 2530 12291 2530 12291 4 _0057_
rlabel metal1 s 2484 8398 2484 8398 4 _0058_
rlabel metal2 s 5934 7582 5934 7582 4 _0059_
rlabel metal1 s 7682 13396 7682 13396 4 _0060_
rlabel metal1 s 2530 8942 2530 8942 4 _0061_
rlabel metal1 s 5474 9690 5474 9690 4 _0062_
rlabel metal1 s 3726 8058 3726 8058 4 _0063_
rlabel metal1 s 5014 7990 5014 7990 4 _0064_
rlabel metal1 s 5336 9146 5336 9146 4 _0065_
rlabel metal1 s 5152 12750 5152 12750 4 _0066_
rlabel metal2 s 5106 9486 5106 9486 4 _0067_
rlabel metal2 s 5474 10642 5474 10642 4 _0068_
rlabel metal1 s 12926 12172 12926 12172 4 _0069_
rlabel metal2 s 5750 11747 5750 11747 4 _0070_
rlabel metal1 s 18262 13498 18262 13498 4 _0071_
rlabel metal1 s 18492 14382 18492 14382 4 _0072_
rlabel metal1 s 14214 9011 14214 9011 4 _0073_
rlabel metal2 s 13570 7412 13570 7412 4 _0074_
rlabel metal1 s 13064 2278 13064 2278 4 _0075_
rlabel metal2 s 16606 3213 16606 3213 4 _0076_
rlabel metal3 s 14858 2907 14858 2907 4 _0077_
rlabel metal1 s 12052 3434 12052 3434 4 _0078_
rlabel metal1 s 21758 4046 21758 4046 4 _0079_
rlabel metal2 s 18630 3842 18630 3842 4 _0080_
rlabel metal2 s 18906 1700 18906 1700 4 _0081_
rlabel metal1 s 17296 3570 17296 3570 4 _0082_
rlabel metal1 s 16376 2414 16376 2414 4 _0083_
rlabel metal1 s 16652 2482 16652 2482 4 _0084_
rlabel metal1 s 11730 13872 11730 13872 4 _0085_
rlabel metal1 s 13110 13804 13110 13804 4 _0086_
rlabel metal1 s 10488 5746 10488 5746 4 _0087_
rlabel metal1 s 9154 1496 9154 1496 4 _0088_
rlabel metal1 s 10672 3026 10672 3026 4 _0089_
rlabel metal1 s 15778 1904 15778 1904 4 _0090_
rlabel metal3 s 15571 5508 15571 5508 4 _0091_
rlabel metal1 s 21482 1938 21482 1938 4 _0092_
rlabel metal1 s 3358 6766 3358 6766 4 _0093_
rlabel metal1 s 4002 1938 4002 1938 4 _0094_
rlabel metal1 s 3542 6834 3542 6834 4 _0095_
rlabel metal1 s 3174 8602 3174 8602 4 _0096_
rlabel metal1 s 5750 7718 5750 7718 4 _0097_
rlabel metal1 s 16422 14994 16422 14994 4 _0098_
rlabel metal2 s 7314 5661 7314 5661 4 _0099_
rlabel metal1 s 15502 9486 15502 9486 4 _0100_
rlabel metal1 s 15042 9690 15042 9690 4 _0101_
rlabel metal1 s 14950 11696 14950 11696 4 _0102_
rlabel metal1 s 16422 11526 16422 11526 4 _0103_
rlabel metal2 s 15042 8857 15042 8857 4 _0104_
rlabel metal1 s 14306 8602 14306 8602 4 _0105_
rlabel metal1 s 17940 4726 17940 4726 4 _0106_
rlabel metal1 s 13156 11186 13156 11186 4 _0107_
rlabel metal1 s 15226 4692 15226 4692 4 _0108_
rlabel metal2 s 16882 4896 16882 4896 4 _0109_
rlabel metal2 s 15778 4998 15778 4998 4 _0110_
rlabel metal1 s 19044 13838 19044 13838 4 _0111_
rlabel metal1 s 18078 13396 18078 13396 4 _0112_
rlabel metal2 s 17618 13056 17618 13056 4 _0113_
rlabel metal1 s 17112 13838 17112 13838 4 _0114_
rlabel metal1 s 16422 12716 16422 12716 4 _0115_
rlabel metal1 s 16790 12614 16790 12614 4 _0116_
rlabel metal1 s 14904 1802 14904 1802 4 _0117_
rlabel metal1 s 12880 10166 12880 10166 4 _0118_
rlabel metal1 s 9798 12750 9798 12750 4 _0119_
rlabel metal1 s 11914 12274 11914 12274 4 _0120_
rlabel metal2 s 14628 3026 14628 3026 4 _0121_
rlabel metal1 s 22494 4012 22494 4012 4 _0122_
rlabel metal1 s 21850 1870 21850 1870 4 _0123_
rlabel metal1 s 19419 1394 19419 1394 4 _0124_
rlabel metal1 s 18078 1802 18078 1802 4 _0125_
rlabel metal1 s 16698 1938 16698 1938 4 _0126_
rlabel metal1 s 16514 1836 16514 1836 4 _0127_
rlabel metal1 s 21896 3910 21896 3910 4 _0128_
rlabel metal1 s 14168 4046 14168 4046 4 _0129_
rlabel metal2 s 2254 9180 2254 9180 4 _0130_
rlabel metal2 s 7038 7548 7038 7548 4 _0131_
rlabel metal2 s 5658 7072 5658 7072 4 _0132_
rlabel metal1 s 6716 10778 6716 10778 4 _0133_
rlabel metal1 s 7222 7752 7222 7752 4 _0134_
rlabel metal2 s 13754 7854 13754 7854 4 _0135_
rlabel metal1 s 11086 5066 11086 5066 4 _0136_
rlabel metal1 s 21712 1938 21712 1938 4 _0137_
rlabel metal2 s 19412 2618 19412 2618 4 _0138_
rlabel metal2 s 15226 5338 15226 5338 4 _0139_
rlabel metal1 s 13432 4046 13432 4046 4 _0140_
rlabel metal1 s 16238 1836 16238 1836 4 _0141_
rlabel metal1 s 13432 1190 13432 1190 4 _0142_
rlabel metal1 s 17250 14246 17250 14246 4 _0143_
rlabel metal1 s 16882 14450 16882 14450 4 _0144_
rlabel metal2 s 15778 1836 15778 1836 4 _0145_
rlabel metal1 s 11178 1904 11178 1904 4 _0146_
rlabel metal2 s 12650 5185 12650 5185 4 _0147_
rlabel metal1 s 11408 5134 11408 5134 4 _0148_
rlabel metal1 s 11132 6834 11132 6834 4 _0149_
rlabel metal1 s 12926 5678 12926 5678 4 _0150_
rlabel metal1 s 17296 5542 17296 5542 4 _0151_
rlabel metal1 s 8234 6970 8234 6970 4 _0152_
rlabel metal1 s 6256 12750 6256 12750 4 _0153_
rlabel metal2 s 9430 5882 9430 5882 4 _0154_
rlabel metal1 s 10764 5134 10764 5134 4 _0155_
rlabel metal2 s 11454 2077 11454 2077 4 _0156_
rlabel metal1 s 17020 1394 17020 1394 4 _0157_
rlabel metal1 s 11546 2414 11546 2414 4 _0158_
rlabel metal1 s 18584 1802 18584 1802 4 _0159_
rlabel metal1 s 8602 1972 8602 1972 4 _0160_
rlabel metal1 s 4600 1326 4600 1326 4 _0161_
rlabel metal1 s 6394 1428 6394 1428 4 _0162_
rlabel metal1 s 21620 1734 21620 1734 4 _0163_
rlabel metal1 s 20930 1904 20930 1904 4 _0164_
rlabel metal1 s 18906 1938 18906 1938 4 _0165_
rlabel metal1 s 6808 1394 6808 1394 4 _0166_
rlabel metal1 s 7130 1360 7130 1360 4 _0167_
rlabel metal1 s 8510 1870 8510 1870 4 _0168_
rlabel metal1 s 10258 1870 10258 1870 4 _0169_
rlabel metal2 s 10074 2312 10074 2312 4 _0170_
rlabel metal1 s 10396 1938 10396 1938 4 _0171_
rlabel metal1 s 11684 1394 11684 1394 4 _0172_
rlabel metal1 s 5014 4012 5014 4012 4 _0173_
rlabel metal1 s 5244 1870 5244 1870 4 _0174_
rlabel metal1 s 18400 2278 18400 2278 4 _0175_
rlabel metal1 s 4554 1904 4554 1904 4 _0176_
rlabel metal1 s 4830 1938 4830 1938 4 _0177_
rlabel metal1 s 5934 1904 5934 1904 4 _0178_
rlabel metal1 s 8280 1326 8280 1326 4 _0179_
rlabel metal1 s 7682 1938 7682 1938 4 _0180_
rlabel metal1 s 7958 1972 7958 1972 4 _0181_
rlabel metal1 s 7820 1530 7820 1530 4 _0182_
rlabel metal1 s 13984 6222 13984 6222 4 _0183_
rlabel metal1 s 8372 5814 8372 5814 4 _0184_
rlabel metal1 s 13800 8942 13800 8942 4 _0185_
rlabel metal2 s 7314 7616 7314 7616 4 _0186_
rlabel metal1 s 13800 6222 13800 6222 4 _0187_
rlabel metal2 s 13018 5457 13018 5457 4 _0188_
rlabel metal2 s 8786 1462 8786 1462 4 _0189_
rlabel metal3 s 16261 1428 16261 1428 4 _0190_
rlabel metal1 s 8970 5644 8970 5644 4 _0191_
rlabel metal1 s 21574 9690 21574 9690 4 _0192_
rlabel metal1 s 16100 8602 16100 8602 4 _0193_
rlabel metal1 s 16514 7412 16514 7412 4 _0194_
rlabel metal2 s 9982 7922 9982 7922 4 _0195_
rlabel metal1 s 10994 6868 10994 6868 4 _0196_
rlabel metal2 s 11270 4250 11270 4250 4 _0197_
rlabel metal1 s 18446 12614 18446 12614 4 _0198_
rlabel metal1 s 8280 1938 8280 1938 4 _0199_
rlabel metal1 s 8832 2958 8832 2958 4 _0200_
rlabel metal1 s 9522 2482 9522 2482 4 _0201_
rlabel metal2 s 7682 4862 7682 4862 4 _0202_
rlabel metal1 s 7820 4114 7820 4114 4 _0203_
rlabel metal1 s 5106 4080 5106 4080 4 _0204_
rlabel metal1 s 5244 4046 5244 4046 4 _0205_
rlabel metal1 s 7866 4012 7866 4012 4 _0206_
rlabel metal1 s 8004 3570 8004 3570 4 _0207_
rlabel metal1 s 8142 3604 8142 3604 4 _0208_
rlabel metal1 s 8234 3536 8234 3536 4 _0209_
rlabel metal1 s 9890 2958 9890 2958 4 _0210_
rlabel metal1 s 10948 2482 10948 2482 4 _0211_
rlabel metal1 s 11362 2516 11362 2516 4 _0212_
rlabel metal2 s 11546 2074 11546 2074 4 _0213_
rlabel metal1 s 9292 8330 9292 8330 4 _0214_
rlabel metal1 s 9016 4046 9016 4046 4 _0215_
rlabel metal2 s 20010 6953 20010 6953 4 _0216_
rlabel metal1 s 8234 4794 8234 4794 4 _0217_
rlabel metal1 s 9246 4087 9246 4087 4 _0218_
rlabel metal1 s 10534 3978 10534 3978 4 _0219_
rlabel metal3 s 9798 2805 9798 2805 4 _0220_
rlabel metal1 s 9890 2618 9890 2618 4 _0221_
rlabel metal1 s 9890 3468 9890 3468 4 _0222_
rlabel metal2 s 13340 7820 13340 7820 4 _0223_
rlabel metal1 s 9246 10064 9246 10064 4 _0224_
rlabel metal1 s 11914 9078 11914 9078 4 _0225_
rlabel metal1 s 13110 8432 13110 8432 4 _0226_
rlabel metal1 s 10442 3570 10442 3570 4 _0227_
rlabel metal2 s 9430 1887 9430 1887 4 _0228_
rlabel metal1 s 9246 1428 9246 1428 4 _0229_
rlabel metal1 s 8602 3638 8602 3638 4 _0230_
rlabel metal1 s 10166 13328 10166 13328 4 _0231_
rlabel metal1 s 8648 13838 8648 13838 4 _0232_
rlabel metal1 s 8832 14042 8832 14042 4 _0233_
rlabel metal2 s 7866 14484 7866 14484 4 _0234_
rlabel metal1 s 8142 14450 8142 14450 4 _0235_
rlabel metal2 s 9338 14314 9338 14314 4 _0236_
rlabel metal1 s 20930 9486 20930 9486 4 _0237_
rlabel metal1 s 9338 8976 9338 8976 4 _0238_
rlabel metal1 s 9338 13770 9338 13770 4 _0239_
rlabel metal1 s 10626 14416 10626 14416 4 _0240_
rlabel metal1 s 9936 14042 9936 14042 4 _0241_
rlabel metal1 s 10350 14484 10350 14484 4 _0242_
rlabel metal2 s 10902 12988 10902 12988 4 _0243_
rlabel metal1 s 10764 12750 10764 12750 4 _0244_
rlabel metal1 s 7176 11322 7176 11322 4 _0245_
rlabel metal1 s 10626 10166 10626 10166 4 _0246_
rlabel metal1 s 8661 10574 8661 10574 4 _0247_
rlabel metal1 s 14720 10234 14720 10234 4 _0248_
rlabel metal1 s 9476 13158 9476 13158 4 _0249_
rlabel metal2 s 17986 11390 17986 11390 4 _0250_
rlabel metal1 s 11914 10608 11914 10608 4 _0251_
rlabel metal1 s 11546 10778 11546 10778 4 _0252_
rlabel metal1 s 10120 12818 10120 12818 4 _0253_
rlabel metal1 s 9430 12716 9430 12716 4 _0254_
rlabel metal1 s 10856 13838 10856 13838 4 _0255_
rlabel metal1 s 9936 13838 9936 13838 4 _0256_
rlabel metal1 s 13386 12274 13386 12274 4 _0257_
rlabel metal1 s 13340 12954 13340 12954 4 _0258_
rlabel metal1 s 10764 13974 10764 13974 4 _0259_
rlabel metal1 s 11178 14042 11178 14042 4 _0260_
rlabel metal2 s 11178 13668 11178 13668 4 _0261_
rlabel metal1 s 4370 10982 4370 10982 4 _0262_
rlabel metal2 s 4048 9010 4048 9010 4 _0263_
rlabel metal1 s 6394 12886 6394 12886 4 _0264_
rlabel metal1 s 6762 12682 6762 12682 4 _0265_
rlabel metal1 s 6394 12716 6394 12716 4 _0266_
rlabel metal2 s 5934 13090 5934 13090 4 _0267_
rlabel metal1 s 13432 10166 13432 10166 4 _0268_
rlabel metal1 s 13110 9078 13110 9078 4 _0269_
rlabel metal3 s 12558 9316 12558 9316 4 _0270_
rlabel metal1 s 13432 9146 13432 9146 4 _0271_
rlabel metal1 s 12926 9962 12926 9962 4 _0272_
rlabel metal2 s 14490 12954 14490 12954 4 _0273_
rlabel metal1 s 14030 1292 14030 1292 4 _0274_
rlabel metal1 s 21528 5338 21528 5338 4 _0275_
rlabel metal1 s 21206 4046 21206 4046 4 _0276_
rlabel metal1 s 20194 2856 20194 2856 4 _0277_
rlabel metal1 s 15824 11118 15824 11118 4 _0278_
rlabel metal1 s 15364 10438 15364 10438 4 _0279_
rlabel metal2 s 15318 8092 15318 8092 4 _0280_
rlabel metal1 s 12742 5168 12742 5168 4 _0281_
rlabel metal1 s 15916 10574 15916 10574 4 _0282_
rlabel metal2 s 15318 3927 15318 3927 4 _0283_
rlabel metal2 s 12466 9282 12466 9282 4 _0284_
rlabel metal1 s 13294 12138 13294 12138 4 _0285_
rlabel metal1 s 15778 3094 15778 3094 4 _0286_
rlabel metal1 s 15042 3162 15042 3162 4 _0287_
rlabel metal1 s 5750 5168 5750 5168 4 _0288_
rlabel metal2 s 13754 11645 13754 11645 4 _0289_
rlabel metal1 s 13018 3706 13018 3706 4 _0290_
rlabel metal2 s 13478 3026 13478 3026 4 _0291_
rlabel metal1 s 14030 1394 14030 1394 4 _0292_
rlabel metal1 s 11408 4658 11408 4658 4 _0293_
rlabel metal2 s 12006 4828 12006 4828 4 _0294_
rlabel metal1 s 13202 4794 13202 4794 4 _0295_
rlabel metal2 s 11730 5219 11730 5219 4 _0296_
rlabel metal2 s 12282 2077 12282 2077 4 _0297_
rlabel metal1 s 18998 6120 18998 6120 4 _0298_
rlabel metal1 s 6394 6086 6394 6086 4 _0299_
rlabel metal1 s 8878 5711 8878 5711 4 _0300_
rlabel metal1 s 10626 9894 10626 9894 4 _0301_
rlabel metal1 s 11178 5712 11178 5712 4 _0302_
rlabel metal1 s 10948 7310 10948 7310 4 _0303_
rlabel metal2 s 11638 6052 11638 6052 4 _0304_
rlabel metal1 s 11914 986 11914 986 4 _0305_
rlabel metal2 s 9522 2533 9522 2533 4 _0306_
rlabel metal1 s 15456 6698 15456 6698 4 _0307_
rlabel metal1 s 4048 7446 4048 7446 4 _0308_
rlabel metal2 s 1978 6052 1978 6052 4 _0309_
rlabel metal1 s 13110 10506 13110 10506 4 _0310_
rlabel metal2 s 11086 7820 11086 7820 4 _0311_
rlabel metal1 s 12098 6834 12098 6834 4 _0312_
rlabel metal1 s 10442 1428 10442 1428 4 _0313_
rlabel metal1 s 13110 7276 13110 7276 4 _0314_
rlabel metal1 s 2668 8602 2668 8602 4 _0315_
rlabel metal1 s 2415 6834 2415 6834 4 _0316_
rlabel metal1 s 11178 9044 11178 9044 4 _0317_
rlabel metal1 s 11408 6290 11408 6290 4 _0318_
rlabel metal2 s 10166 2295 10166 2295 4 _0319_
rlabel metal1 s 11638 11764 11638 11764 4 _0320_
rlabel metal1 s 3542 11628 3542 11628 4 _0321_
rlabel metal1 s 11178 10132 11178 10132 4 _0322_
rlabel metal1 s 11684 10234 11684 10234 4 _0323_
rlabel metal1 s 11086 11866 11086 11866 4 _0324_
rlabel metal1 s 3358 12308 3358 12308 4 _0325_
rlabel metal2 s 13202 10676 13202 10676 4 _0326_
rlabel metal1 s 12696 10778 12696 10778 4 _0327_
rlabel metal1 s 11914 12410 11914 12410 4 _0328_
rlabel metal1 s 16422 1326 16422 1326 4 _0329_
rlabel metal1 s 16238 3094 16238 3094 4 _0330_
rlabel metal1 s 16146 2924 16146 2924 4 _0331_
rlabel metal1 s 14996 8466 14996 8466 4 _0332_
rlabel metal1 s 14812 6630 14812 6630 4 _0333_
rlabel metal1 s 16284 4046 16284 4046 4 _0334_
rlabel metal1 s 16422 3060 16422 3060 4 _0335_
rlabel metal1 s 16146 986 16146 986 4 _0336_
rlabel metal2 s 14490 3196 14490 3196 4 _0337_
rlabel metal1 s 14214 2958 14214 2958 4 _0338_
rlabel metal1 s 14950 4046 14950 4046 4 _0339_
rlabel metal1 s 14766 3026 14766 3026 4 _0340_
rlabel metal1 s 14904 2822 14904 2822 4 _0341_
rlabel metal2 s 11822 7905 11822 7905 4 _0342_
rlabel metal1 s 12144 4794 12144 4794 4 _0343_
rlabel metal1 s 12512 5746 12512 5746 4 _0344_
rlabel metal1 s 11730 7956 11730 7956 4 _0345_
rlabel metal1 s 13294 6800 13294 6800 4 _0346_
rlabel metal1 s 13616 5746 13616 5746 4 _0347_
rlabel metal1 s 12190 5644 12190 5644 4 _0348_
rlabel metal2 s 16882 1394 16882 1394 4 _0349_
rlabel metal1 s 15410 6188 15410 6188 4 _0350_
rlabel metal1 s 15824 6222 15824 6222 4 _0351_
rlabel metal1 s 11224 10574 11224 10574 4 _0352_
rlabel metal1 s 14858 6902 14858 6902 4 _0353_
rlabel metal1 s 15180 6222 15180 6222 4 _0354_
rlabel metal2 s 16238 1887 16238 1887 4 _0355_
rlabel metal1 s 18124 1326 18124 1326 4 _0356_
rlabel metal1 s 10810 6698 10810 6698 4 _0357_
rlabel metal1 s 12006 7276 12006 7276 4 _0358_
rlabel metal1 s 14030 11254 14030 11254 4 _0359_
rlabel metal1 s 11546 8058 11546 8058 4 _0360_
rlabel metal2 s 11730 7786 11730 7786 4 _0361_
rlabel metal1 s 18216 986 18216 986 4 _0362_
rlabel metal1 s 14352 6630 14352 6630 4 _0363_
rlabel metal1 s 14950 7310 14950 7310 4 _0364_
rlabel metal1 s 15042 7854 15042 7854 4 _0365_
rlabel metal2 s 14490 7854 14490 7854 4 _0366_
rlabel metal1 s 17526 1394 17526 1394 4 _0367_
rlabel metal2 s 10856 11730 10856 11730 4 _0368_
rlabel metal1 s 10672 11662 10672 11662 4 _0369_
rlabel metal2 s 10902 10982 10902 10982 4 _0370_
rlabel metal2 s 11086 11407 11086 11407 4 _0371_
rlabel metal1 s 12604 12818 12604 12818 4 _0372_
rlabel metal2 s 14122 11492 14122 11492 4 _0373_
rlabel metal1 s 14260 11662 14260 11662 4 _0374_
rlabel metal1 s 13432 11866 13432 11866 4 _0375_
rlabel metal1 s 14168 12410 14168 12410 4 _0376_
rlabel metal1 s 2714 9520 2714 9520 4 _0377_
rlabel metal1 s 2576 9622 2576 9622 4 _0378_
rlabel metal1 s 3956 8806 3956 8806 4 _0379_
rlabel metal1 s 3956 9010 3956 9010 4 _0380_
rlabel metal1 s 3358 9010 3358 9010 4 _0381_
rlabel metal1 s 21412 9010 21412 9010 4 _0382_
rlabel metal1 s 3680 9894 3680 9894 4 _0383_
rlabel metal2 s 2622 9894 2622 9894 4 _0384_
rlabel metal1 s 3404 7786 3404 7786 4 _0385_
rlabel metal1 s 3082 9044 3082 9044 4 _0386_
rlabel metal1 s 2530 10030 2530 10030 4 _0387_
rlabel metal1 s 3450 6970 3450 6970 4 _0388_
rlabel metal1 s 3450 9452 3450 9452 4 _0389_
rlabel metal2 s 3726 7786 3726 7786 4 _0390_
rlabel metal1 s 3082 7514 3082 7514 4 _0391_
rlabel metal1 s 2254 9112 2254 9112 4 _0392_
rlabel metal2 s 3266 9928 3266 9928 4 _0393_
rlabel metal1 s 2990 9996 2990 9996 4 _0394_
rlabel metal1 s 2254 10234 2254 10234 4 _0395_
rlabel metal1 s 1610 9962 1610 9962 4 _0396_
rlabel metal1 s 4048 10574 4048 10574 4 _0397_
rlabel metal2 s 3082 5474 3082 5474 4 _0398_
rlabel metal1 s 3864 10778 3864 10778 4 _0399_
rlabel metal1 s 4554 10574 4554 10574 4 _0400_
rlabel metal2 s 3818 10013 3818 10013 4 _0401_
rlabel metal1 s 19964 9010 19964 9010 4 _0402_
rlabel metal1 s 20378 7922 20378 7922 4 _0403_
rlabel metal1 s 21942 9452 21942 9452 4 _0404_
rlabel metal1 s 20838 8500 20838 8500 4 _0405_
rlabel metal1 s 21804 6834 21804 6834 4 _0406_
rlabel metal1 s 21850 5338 21850 5338 4 _0407_
rlabel metal1 s 21114 8398 21114 8398 4 _0408_
rlabel metal1 s 19642 8432 19642 8432 4 _0409_
rlabel metal1 s 19688 2618 19688 2618 4 _0410_
rlabel metal1 s 18722 2414 18722 2414 4 _0411_
rlabel metal1 s 19090 4624 19090 4624 4 _0412_
rlabel metal2 s 18906 4029 18906 4029 4 _0413_
rlabel metal1 s 19872 2890 19872 2890 4 _0414_
rlabel metal1 s 20516 2958 20516 2958 4 _0415_
rlabel metal2 s 19826 8806 19826 8806 4 _0416_
rlabel metal1 s 19563 3706 19563 3706 4 _0417_
rlabel metal3 s 17917 2924 17917 2924 4 _0418_
rlabel metal1 s 19550 12852 19550 12852 4 _0419_
rlabel metal1 s 20148 2414 20148 2414 4 _0420_
rlabel metal1 s 19918 2516 19918 2516 4 _0421_
rlabel metal1 s 6854 2958 6854 2958 4 _0422_
rlabel metal1 s 7038 2822 7038 2822 4 _0423_
rlabel metal1 s 4600 2482 4600 2482 4 _0424_
rlabel metal1 s 6486 3502 6486 3502 4 _0425_
rlabel metal1 s 7866 6868 7866 6868 4 _0426_
rlabel metal2 s 8050 6494 8050 6494 4 _0427_
rlabel metal1 s 17020 11730 17020 11730 4 _0428_
rlabel metal1 s 8556 5882 8556 5882 4 _0429_
rlabel metal1 s 5198 5202 5198 5202 4 _0430_
rlabel metal2 s 8234 9486 8234 9486 4 _0431_
rlabel metal1 s 9016 10030 9016 10030 4 _0432_
rlabel metal1 s 8556 9418 8556 9418 4 _0433_
rlabel metal1 s 8326 11118 8326 11118 4 _0434_
rlabel metal2 s 8418 11016 8418 11016 4 _0435_
rlabel metal1 s 7912 11322 7912 11322 4 _0436_
rlabel metal1 s 8970 10778 8970 10778 4 _0437_
rlabel metal3 s 7636 2856 7636 2856 4 _0438_
rlabel metal1 s 1978 2924 1978 2924 4 _0439_
rlabel metal1 s 2070 4080 2070 4080 4 _0440_
rlabel metal1 s 19412 10574 19412 10574 4 _0441_
rlabel metal1 s 1840 10234 1840 10234 4 _0442_
rlabel metal1 s 1886 4046 1886 4046 4 _0443_
rlabel metal2 s 2622 6664 2622 6664 4 _0444_
rlabel metal1 s 2346 5576 2346 5576 4 _0445_
rlabel metal1 s 1748 9894 1748 9894 4 _0446_
rlabel metal1 s 2530 5168 2530 5168 4 _0447_
rlabel metal1 s 2116 6426 2116 6426 4 _0448_
rlabel metal1 s 2530 6188 2530 6188 4 _0449_
rlabel metal1 s 2024 7310 2024 7310 4 _0450_
rlabel metal1 s 1610 6970 1610 6970 4 _0451_
rlabel metal1 s 1978 12784 1978 12784 4 _0452_
rlabel metal1 s 1840 10778 1840 10778 4 _0453_
rlabel metal1 s 1702 12886 1702 12886 4 _0454_
rlabel metal1 s 2300 12954 2300 12954 4 _0455_
rlabel metal1 s 2484 13158 2484 13158 4 _0456_
rlabel metal2 s 1702 12835 1702 12835 4 _0457_
rlabel metal2 s 1710 12614 1710 12614 4 _0458_
rlabel metal1 s 1840 12954 1840 12954 4 _0459_
rlabel metal1 s 2576 12750 2576 12750 4 _0460_
rlabel metal2 s 18354 7565 18354 7565 4 _0461_
rlabel metal2 s 16238 12070 16238 12070 4 _0462_
rlabel metal2 s 19182 13702 19182 13702 4 _0463_
rlabel metal1 s 15456 13838 15456 13838 4 _0464_
rlabel metal1 s 16284 14042 16284 14042 4 _0465_
rlabel metal1 s 7130 14926 7130 14926 4 _0466_
rlabel metal2 s 20102 14484 20102 14484 4 _0467_
rlabel metal2 s 18078 14960 18078 14960 4 _0468_
rlabel metal1 s 21068 14450 21068 14450 4 _0469_
rlabel metal1 s 20010 13396 20010 13396 4 _0470_
rlabel metal2 s 19918 11050 19918 11050 4 _0471_
rlabel metal1 s 20240 9690 20240 9690 4 _0472_
rlabel metal1 s 20332 9146 20332 9146 4 _0473_
rlabel metal1 s 20424 3706 20424 3706 4 _0474_
rlabel metal1 s 20056 4046 20056 4046 4 _0475_
rlabel metal1 s 18860 5338 18860 5338 4 _0476_
rlabel metal1 s 18952 5746 18952 5746 4 _0477_
rlabel metal1 s 18814 5814 18814 5814 4 _0478_
rlabel metal1 s 19504 10506 19504 10506 4 _0479_
rlabel metal1 s 18584 10778 18584 10778 4 _0480_
rlabel metal1 s 17848 5882 17848 5882 4 _0481_
rlabel metal1 s 18400 8398 18400 8398 4 _0482_
rlabel metal1 s 18722 6188 18722 6188 4 _0483_
rlabel metal2 s 18722 8092 18722 8092 4 _0484_
rlabel metal1 s 17618 7242 17618 7242 4 _0485_
rlabel metal1 s 18032 6698 18032 6698 4 _0486_
rlabel metal1 s 19274 9044 19274 9044 4 _0487_
rlabel metal2 s 19090 8738 19090 8738 4 _0488_
rlabel metal1 s 17986 7344 17986 7344 4 _0489_
rlabel metal1 s 19090 11696 19090 11696 4 _0490_
rlabel metal1 s 19044 11322 19044 11322 4 _0491_
rlabel metal2 s 19895 9452 19895 9452 4 _0492_
rlabel metal1 s 19182 10608 19182 10608 4 _0493_
rlabel metal1 s 20010 11254 20010 11254 4 _0494_
rlabel metal3 s 19734 11101 19734 11101 4 _0495_
rlabel metal2 s 21114 11424 21114 11424 4 _0496_
rlabel metal1 s 20286 9622 20286 9622 4 _0497_
rlabel metal2 s 20746 10778 20746 10778 4 _0498_
rlabel metal1 s 17894 8058 17894 8058 4 _0499_
rlabel metal2 s 19274 9792 19274 9792 4 _0500_
rlabel metal1 s 20608 8058 20608 8058 4 _0501_
rlabel metal1 s 20654 7344 20654 7344 4 _0502_
rlabel metal1 s 21574 8840 21574 8840 4 _0503_
rlabel metal1 s 21666 9044 21666 9044 4 _0504_
rlabel metal1 s 21022 5338 21022 5338 4 _0505_
rlabel metal1 s 22448 10030 22448 10030 4 _0506_
rlabel metal1 s 22540 9690 22540 9690 4 _0507_
rlabel metal2 s 22218 11458 22218 11458 4 _0508_
rlabel metal1 s 19688 4794 19688 4794 4 _0509_
rlabel metal1 s 21804 9146 21804 9146 4 _0510_
rlabel metal1 s 21160 4794 21160 4794 4 _0511_
rlabel metal1 s 21850 8602 21850 8602 4 _0512_
rlabel metal1 s 22402 9656 22402 9656 4 _0513_
rlabel metal1 s 21896 12818 21896 12818 4 _0514_
rlabel metal1 s 21528 12954 21528 12954 4 _0515_
rlabel metal2 s 6670 15412 6670 15412 4 b6
rlabel metal2 s 9614 15412 9614 15412 4 b7
rlabel metal2 s 5842 500 5842 500 4 b[0]
rlabel metal2 s 5014 500 5014 500 4 b[1]
rlabel metal2 s 4186 500 4186 500 4 b[2]
rlabel metal2 s 3358 500 3358 500 4 b[3]
rlabel metal2 s 2530 534 2530 534 4 b[4]
rlabel metal2 s 1702 483 1702 483 4 b[5]
rlabel metal2 s 874 415 874 415 4 b[6]
rlabel metal2 s 46 772 46 772 4 b[7]
rlabel metal3 s 21858 13940 21858 13940 4 clk
rlabel metal1 s 17434 7990 17434 7990 4 clknet_0_clk
rlabel metal1 s 1196 2482 1196 2482 4 clknet_2_0__leaf_clk
rlabel metal1 s 7774 9554 7774 9554 4 clknet_2_1__leaf_clk
rlabel metal1 s 18998 7412 18998 7412 4 clknet_2_2__leaf_clk
rlabel metal1 s 19734 14484 19734 14484 4 clknet_2_3__leaf_clk
rlabel metal1 s 5658 13702 5658 13702 4 divider\[0\]
rlabel metal1 s 5888 14518 5888 14518 4 divider\[1\]
rlabel metal1 s 7452 15130 7452 15130 4 g6
rlabel metal1 s 10442 15130 10442 15130 4 g7
rlabel metal2 s 14122 415 14122 415 4 g[0]
rlabel metal2 s 13294 500 13294 500 4 g[1]
rlabel metal2 s 12466 415 12466 415 4 g[2]
rlabel metal2 s 11638 500 11638 500 4 g[3]
rlabel metal2 s 10810 415 10810 415 4 g[4]
rlabel metal2 s 9982 500 9982 500 4 g[5]
rlabel metal2 s 9154 500 9154 500 4 g[6]
rlabel metal2 s 8326 500 8326 500 4 g[7]
rlabel metal2 s 15410 14076 15410 14076 4 gate
rlabel metal2 s 4646 15419 4646 15419 4 hblank
rlabel metal2 s 6210 15419 6210 15419 4 hsync
rlabel metal1 s 21298 14586 21298 14586 4 mode\[0\]
rlabel metal1 s 13524 14246 13524 14246 4 mode\[1\]
rlabel metal1 s 23230 14586 23230 14586 4 mode\[2\]
rlabel metal2 s 22862 11050 22862 11050 4 net1
rlabel metal1 s 2162 1870 2162 1870 4 net10
rlabel metal2 s 8970 9316 8970 9316 4 net11
rlabel metal2 s 15410 1020 15410 1020 4 net12
rlabel metal1 s 13018 850 13018 850 4 net13
rlabel metal1 s 4554 850 4554 850 4 net14
rlabel metal1 s 4002 782 4002 782 4 net15
rlabel metal1 s 4002 680 4002 680 4 net16
rlabel metal1 s 1978 1496 1978 1496 4 net17
rlabel metal1 s 1150 782 1150 782 4 net18
rlabel metal1 s 1196 1394 1196 1394 4 net19
rlabel metal1 s 22310 15368 22310 15368 4 net2
rlabel metal1 s 8234 14858 8234 14858 4 net20
rlabel metal4 s 10051 5372 10051 5372 4 net21
rlabel metal1 s 14444 782 14444 782 4 net22
rlabel metal1 s 13708 782 13708 782 4 net23
rlabel metal1 s 12742 782 12742 782 4 net24
rlabel metal1 s 12144 782 12144 782 4 net25
rlabel metal1 s 10948 782 10948 782 4 net26
rlabel metal1 s 10074 816 10074 816 4 net27
rlabel metal1 s 9154 782 9154 782 4 net28
rlabel metal1 s 8694 748 8694 748 4 net29
rlabel metal1 s 22218 15028 22218 15028 4 net3
rlabel metal1 s 4830 14892 4830 14892 4 net30
rlabel metal1 s 2070 13872 2070 13872 4 net31
rlabel metal3 s 12926 12869 12926 12869 4 net32
rlabel metal4 s 14973 2108 14973 2108 4 net33
rlabel metal1 s 16698 646 16698 646 4 net34
rlabel metal1 s 20930 816 20930 816 4 net35
rlabel metal1 s 20838 816 20838 816 4 net36
rlabel metal1 s 19550 782 19550 782 4 net37
rlabel metal1 s 19274 714 19274 714 4 net38
rlabel metal1 s 18124 782 18124 782 4 net39
rlabel metal1 s 16882 13294 16882 13294 4 net4
rlabel metal1 s 17480 782 17480 782 4 net40
rlabel metal1 s 16698 816 16698 816 4 net41
rlabel metal1 s 6808 14450 6808 14450 4 net42
rlabel metal1 s 8188 14314 8188 14314 4 net43
rlabel metal2 s 2530 14620 2530 14620 4 net44
rlabel metal1 s 17664 14382 17664 14382 4 net5
rlabel metal1 s 19964 13838 19964 13838 4 net6
rlabel metal1 s 18860 14586 18860 14586 4 net7
rlabel metal2 s 18906 14637 18906 14637 4 net8
rlabel metal2 s 18538 14144 18538 14144 4 net9
rlabel metal2 s 8142 15412 8142 15412 4 r6
rlabel metal2 s 11086 15412 11086 15412 4 r7
rlabel metal2 s 22374 0 22430 400 4 r[0]
port 28 nsew
rlabel metal2 s 21574 500 21574 500 4 r[1]
rlabel metal2 s 20746 500 20746 500 4 r[2]
rlabel metal2 s 19918 500 19918 500 4 r[3]
rlabel metal2 s 19090 500 19090 500 4 r[4]
rlabel metal2 s 18262 415 18262 415 4 r[5]
rlabel metal2 s 17434 500 17434 500 4 r[6]
rlabel metal2 s 16578 0 16634 400 4 r[7]
port 35 nsew
rlabel metal1 s 20562 3570 20562 3570 4 rampc\[0\]
rlabel metal1 s 21758 1326 21758 1326 4 rampc\[1\]
rlabel metal1 s 3864 1938 3864 1938 4 rampc\[2\]
rlabel metal1 s 4232 4046 4232 4046 4 rampc\[3\]
rlabel metal2 s 7222 5100 7222 5100 4 rampc\[4\]
rlabel metal1 s 8786 9010 8786 9010 4 rampc\[5\]
rlabel metal1 s 8878 12614 8878 12614 4 rampc\[6\]
rlabel metal1 s 9522 11152 9522 11152 4 rampc\[7\]
rlabel metal1 s 16054 11662 16054 11662 4 registered
rlabel metal1 s 23046 12784 23046 12784 4 rst_n
rlabel metal1 s 22954 14926 22954 14926 4 ui_in[0]
rlabel metal1 s 22264 14926 22264 14926 4 ui_in[1]
rlabel metal1 s 22034 14892 22034 14892 4 ui_in[2]
rlabel metal1 s 20792 14926 20792 14926 4 ui_in[3]
rlabel metal1 s 20286 14926 20286 14926 4 ui_in[4]
rlabel metal1 s 19320 14926 19320 14926 4 ui_in[5]
rlabel metal1 s 18584 14926 18584 14926 4 ui_in[6]
rlabel metal1 s 17756 14926 17756 14926 4 ui_in[7]
rlabel metal2 s 5198 15412 5198 15412 4 vblank
rlabel metal2 s 2346 3876 2346 3876 4 vga_sync.hpos\[0\]
rlabel metal2 s 21482 1955 21482 1955 4 vga_sync.hpos\[1\]
rlabel metal1 s 4094 1326 4094 1326 4 vga_sync.hpos\[2\]
rlabel metal1 s 4094 7820 4094 7820 4 vga_sync.hpos\[3\]
rlabel metal1 s 7130 4590 7130 4590 4 vga_sync.hpos\[4\]
rlabel metal2 s 9706 8772 9706 8772 4 vga_sync.hpos\[5\]
rlabel metal1 s 3634 11118 3634 11118 4 vga_sync.hpos\[6\]
rlabel metal1 s 4370 12274 4370 12274 4 vga_sync.hpos\[7\]
rlabel metal1 s 4048 8942 4048 8942 4 vga_sync.hpos\[8\]
rlabel metal1 s 5060 12274 5060 12274 4 vga_sync.hpos\[9\]
rlabel metal2 s 2254 14756 2254 14756 4 vga_sync.hsync
rlabel metal1 s 21160 12614 21160 12614 4 vga_sync.mode
rlabel metal1 s 22126 5163 22126 5163 4 vga_sync.o_vpos\[0\]
rlabel metal1 s 22218 4046 22218 4046 4 vga_sync.o_vpos\[1\]
rlabel metal1 s 22218 5780 22218 5780 4 vga_sync.o_vpos\[2\]
rlabel metal2 s 21896 6426 21896 6426 4 vga_sync.o_vpos\[3\]
rlabel metal3 s 16606 8381 16606 8381 4 vga_sync.o_vpos\[4\]
rlabel metal1 s 17388 8398 17388 8398 4 vga_sync.o_vpos\[5\]
rlabel metal1 s 17986 11594 17986 11594 4 vga_sync.o_vpos\[6\]
rlabel metal1 s 22218 10506 22218 10506 4 vga_sync.o_vpos\[7\]
rlabel metal1 s 22218 10608 22218 10608 4 vga_sync.o_vpos\[8\]
rlabel metal1 s 22862 8364 22862 8364 4 vga_sync.o_vpos\[9\]
rlabel metal1 s 23230 13158 23230 13158 4 vga_sync.vsync
rlabel metal2 s 9154 15419 9154 15419 4 vsync
flabel metal4 s 22352 496 22752 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 16352 496 16752 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 10352 496 10752 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4352 496 4752 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 19352 496 19752 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 13352 496 13752 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7352 496 7752 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1352 496 1752 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 6642 15600 6698 16000 0 FreeSans 280 90 0 0 b6
port 3 nsew
flabel metal2 s 9586 15600 9642 16000 0 FreeSans 280 90 0 0 b7
port 4 nsew
flabel metal2 s 5814 0 5870 400 0 FreeSans 280 90 0 0 b[0]
port 5 nsew
flabel metal2 s 4986 0 5042 400 0 FreeSans 280 90 0 0 b[1]
port 6 nsew
flabel metal2 s 4158 0 4214 400 0 FreeSans 280 90 0 0 b[2]
port 7 nsew
flabel metal2 s 3330 0 3386 400 0 FreeSans 280 90 0 0 b[3]
port 8 nsew
flabel metal2 s 2502 0 2558 400 0 FreeSans 280 90 0 0 b[4]
port 9 nsew
flabel metal2 s 1674 0 1730 400 0 FreeSans 280 90 0 0 b[5]
port 10 nsew
flabel metal2 s 846 0 902 400 0 FreeSans 280 90 0 0 b[6]
port 11 nsew
flabel metal2 s 18 0 74 400 0 FreeSans 280 90 0 0 b[7]
port 12 nsew
flabel metal3 s 23600 13880 24000 14000 0 FreeSans 600 0 0 0 clk
port 13 nsew
flabel metal2 s 7378 15600 7434 16000 0 FreeSans 280 90 0 0 g6
port 14 nsew
flabel metal2 s 10322 15600 10378 16000 0 FreeSans 280 90 0 0 g7
port 15 nsew
flabel metal2 s 14094 0 14150 400 0 FreeSans 280 90 0 0 g[0]
port 16 nsew
flabel metal2 s 13266 0 13322 400 0 FreeSans 280 90 0 0 g[1]
port 17 nsew
flabel metal2 s 12438 0 12494 400 0 FreeSans 280 90 0 0 g[2]
port 18 nsew
flabel metal2 s 11610 0 11666 400 0 FreeSans 280 90 0 0 g[3]
port 19 nsew
flabel metal2 s 10782 0 10838 400 0 FreeSans 280 90 0 0 g[4]
port 20 nsew
flabel metal2 s 9954 0 10010 400 0 FreeSans 280 90 0 0 g[5]
port 21 nsew
flabel metal2 s 9126 0 9182 400 0 FreeSans 280 90 0 0 g[6]
port 22 nsew
flabel metal2 s 8298 0 8354 400 0 FreeSans 280 90 0 0 g[7]
port 23 nsew
flabel metal2 s 4434 15600 4490 16000 0 FreeSans 280 90 0 0 hblank
port 24 nsew
flabel metal2 s 5906 15600 5962 16000 0 FreeSans 280 90 0 0 hsync
port 25 nsew
flabel metal2 s 8114 15600 8170 16000 0 FreeSans 280 90 0 0 r6
port 26 nsew
flabel metal2 s 11058 15600 11114 16000 0 FreeSans 280 90 0 0 r7
port 27 nsew
flabel metal2 s 22402 200 22402 200 0 FreeSans 280 90 0 0 r[0]
flabel metal2 s 21546 0 21602 400 0 FreeSans 280 90 0 0 r[1]
port 29 nsew
flabel metal2 s 20718 0 20774 400 0 FreeSans 280 90 0 0 r[2]
port 30 nsew
flabel metal2 s 19890 0 19946 400 0 FreeSans 280 90 0 0 r[3]
port 31 nsew
flabel metal2 s 19062 0 19118 400 0 FreeSans 280 90 0 0 r[4]
port 32 nsew
flabel metal2 s 18234 0 18290 400 0 FreeSans 280 90 0 0 r[5]
port 33 nsew
flabel metal2 s 17406 0 17462 400 0 FreeSans 280 90 0 0 r[6]
port 34 nsew
flabel metal2 s 16606 200 16606 200 0 FreeSans 280 90 0 0 r[7]
flabel metal3 s 23600 12792 24000 12912 0 FreeSans 600 0 0 0 rst_n
port 36 nsew
flabel metal2 s 22834 15600 22890 16000 0 FreeSans 280 90 0 0 ui_in[0]
port 37 nsew
flabel metal2 s 22098 15600 22154 16000 0 FreeSans 280 90 0 0 ui_in[1]
port 38 nsew
flabel metal2 s 21362 15600 21418 16000 0 FreeSans 280 90 0 0 ui_in[2]
port 39 nsew
flabel metal2 s 20626 15600 20682 16000 0 FreeSans 280 90 0 0 ui_in[3]
port 40 nsew
flabel metal2 s 19890 15600 19946 16000 0 FreeSans 280 90 0 0 ui_in[4]
port 41 nsew
flabel metal2 s 19154 15600 19210 16000 0 FreeSans 280 90 0 0 ui_in[5]
port 42 nsew
flabel metal2 s 18418 15600 18474 16000 0 FreeSans 280 90 0 0 ui_in[6]
port 43 nsew
flabel metal2 s 17682 15600 17738 16000 0 FreeSans 280 90 0 0 ui_in[7]
port 44 nsew
flabel metal2 s 5170 15600 5226 16000 0 FreeSans 280 90 0 0 vblank
port 45 nsew
flabel metal2 s 8850 15600 8906 16000 0 FreeSans 280 90 0 0 vsync
port 46 nsew
<< properties >>
string FIXED_BBOX 0 0 24000 16000
string GDS_END 2009418
string GDS_FILE controller.gds
string GDS_START 417510
<< end >>
