magic
tech sky130A
magscale 1 2
timestamp 1713524504
<< metal1 >>
rect 6686 26488 6742 26494
rect 7514 26488 7570 26494
rect 8342 26488 8398 26494
rect 9170 26488 9226 26494
rect 9998 26488 10054 26494
rect 10826 26488 10882 26494
rect 11654 26488 11710 26494
rect 12482 26488 12538 26494
rect 14966 26488 15022 26494
rect 15794 26488 15850 26494
rect 16622 26488 16678 26494
rect 17450 26488 17506 26494
rect 18278 26488 18334 26494
rect 19106 26488 19162 26494
rect 23246 26488 23302 26494
rect 24074 26488 24130 26494
rect 24902 26488 24958 26494
rect 25730 26488 25786 26494
rect 6742 26432 7048 26488
rect 6686 26426 6742 26432
rect 6992 25992 7048 26432
rect 7570 26432 7848 26488
rect 7514 26426 7570 26432
rect 7792 25992 7848 26432
rect 8398 26432 8648 26488
rect 8342 26426 8398 26432
rect 8592 25992 8648 26432
rect 9226 26432 9448 26488
rect 9170 26426 9226 26432
rect 9392 26032 9448 26432
rect 10054 26432 10248 26488
rect 9998 26426 10054 26432
rect 10192 25992 10248 26432
rect 10882 26432 11048 26488
rect 10826 26426 10882 26432
rect 10992 26032 11048 26432
rect 11710 26432 11848 26488
rect 11654 26426 11710 26432
rect 11792 26032 11848 26432
rect 12538 26432 12648 26488
rect 12482 26426 12538 26432
rect 12592 25972 12648 26432
rect 15022 26432 15248 26488
rect 14966 26426 15022 26432
rect 15192 26032 15248 26432
rect 15850 26432 16048 26488
rect 15794 26426 15850 26432
rect 15992 26012 16048 26432
rect 16678 26432 16848 26488
rect 16622 26426 16678 26432
rect 16792 26032 16848 26432
rect 17506 26432 17648 26488
rect 17450 26426 17506 26432
rect 17592 26032 17648 26432
rect 18334 26432 18448 26488
rect 18278 26426 18334 26432
rect 18392 25992 18448 26432
rect 19162 26432 19268 26488
rect 19928 26432 19934 26488
rect 19990 26432 20068 26488
rect 20756 26432 20762 26488
rect 20818 26432 20824 26488
rect 23302 26432 23448 26488
rect 19106 26426 19162 26432
rect 19212 25972 19268 26432
rect 20012 25992 20068 26432
rect 20762 25992 20818 26432
rect 23246 26426 23302 26432
rect 23392 26052 23448 26432
rect 24130 26432 24248 26488
rect 24074 26426 24130 26432
rect 24192 26032 24248 26432
rect 24958 26432 25048 26488
rect 24902 26426 24958 26432
rect 24992 26012 25048 26432
rect 25786 26432 25900 26488
rect 26552 26432 26558 26488
rect 26614 26432 26620 26488
rect 27380 26432 27386 26488
rect 27442 26432 27448 26488
rect 28208 26432 28214 26488
rect 28270 26432 28276 26488
rect 28976 26440 29042 26496
rect 29098 26440 29104 26496
rect 25730 26426 25786 26432
rect 25844 26052 25900 26432
rect 26558 26032 26614 26432
rect 27386 26032 27442 26432
rect 28214 25992 28270 26432
rect 28976 25970 29032 26440
<< via1 >>
rect 6686 26432 6742 26488
rect 7514 26432 7570 26488
rect 8342 26432 8398 26488
rect 9170 26432 9226 26488
rect 9998 26432 10054 26488
rect 10826 26432 10882 26488
rect 11654 26432 11710 26488
rect 12482 26432 12538 26488
rect 14966 26432 15022 26488
rect 15794 26432 15850 26488
rect 16622 26432 16678 26488
rect 17450 26432 17506 26488
rect 18278 26432 18334 26488
rect 19106 26432 19162 26488
rect 19934 26432 19990 26488
rect 20762 26432 20818 26488
rect 23246 26432 23302 26488
rect 24074 26432 24130 26488
rect 24902 26432 24958 26488
rect 25730 26432 25786 26488
rect 26558 26432 26614 26488
rect 27386 26432 27442 26488
rect 28214 26432 28270 26488
rect 29042 26440 29098 26496
<< metal2 >>
rect 11102 44264 11162 44266
rect 11838 44264 11898 44266
rect 12574 44264 12634 44266
rect 13310 44264 13370 44266
rect 14046 44264 14106 44266
rect 14782 44264 14842 44266
rect 15518 44264 15578 44266
rect 16254 44264 16314 44266
rect 16990 44264 17050 44266
rect 17726 44264 17786 44266
rect 24350 44264 24410 44266
rect 25086 44264 25146 44266
rect 25822 44264 25882 44266
rect 26558 44264 26618 44266
rect 27294 44264 27354 44266
rect 28030 44264 28090 44266
rect 28766 44264 28826 44266
rect 29502 44264 29562 44266
rect 11095 44208 11104 44264
rect 11160 44208 11169 44264
rect 11831 44208 11840 44264
rect 11896 44208 11905 44264
rect 12567 44208 12576 44264
rect 12632 44208 12641 44264
rect 13303 44208 13312 44264
rect 13368 44208 13377 44264
rect 14039 44208 14048 44264
rect 14104 44208 14113 44264
rect 14775 44208 14784 44264
rect 14840 44208 14849 44264
rect 15511 44208 15520 44264
rect 15576 44208 15585 44264
rect 16247 44208 16256 44264
rect 16312 44208 16321 44264
rect 16983 44208 16992 44264
rect 17048 44208 17057 44264
rect 17719 44208 17728 44264
rect 17784 44208 17793 44264
rect 24343 44208 24352 44264
rect 24408 44208 24417 44264
rect 25079 44208 25088 44264
rect 25144 44208 25153 44264
rect 25815 44208 25824 44264
rect 25880 44208 25889 44264
rect 26551 44208 26560 44264
rect 26616 44208 26625 44264
rect 27287 44208 27296 44264
rect 27352 44208 27361 44264
rect 28023 44208 28032 44264
rect 28088 44208 28097 44264
rect 28759 44208 28768 44264
rect 28824 44208 28833 44264
rect 29495 44208 29504 44264
rect 29560 44208 29569 44264
rect 11102 43388 11162 44208
rect 11838 43388 11898 44208
rect 12574 43388 12634 44208
rect 13310 43388 13370 44208
rect 14046 43388 14106 44208
rect 14782 43388 14842 44208
rect 15518 43388 15578 44208
rect 16254 43388 16314 44208
rect 16990 43388 17050 44208
rect 17726 43388 17786 44208
rect 24350 43388 24410 44208
rect 25086 43388 25146 44208
rect 25822 43388 25882 44208
rect 26558 43388 26618 44208
rect 27294 43388 27354 44208
rect 28030 43388 28090 44208
rect 28766 43388 28826 44208
rect 29502 43388 29562 44208
rect 6686 26488 6742 27794
rect 7514 26488 7570 27794
rect 8342 26488 8398 27794
rect 9170 26488 9226 27794
rect 9998 26488 10054 27808
rect 10826 26488 10882 27794
rect 11654 26488 11710 27794
rect 12482 26488 12538 27794
rect 14966 26488 15022 27794
rect 15794 26488 15850 27794
rect 16622 26488 16678 27794
rect 17450 26488 17506 27794
rect 18278 26488 18334 27794
rect 19106 26488 19162 27794
rect 19934 26488 19990 27794
rect 6680 26432 6686 26488
rect 6742 26432 6748 26488
rect 7508 26432 7514 26488
rect 7570 26432 7576 26488
rect 8336 26432 8342 26488
rect 8398 26432 8404 26488
rect 9164 26432 9170 26488
rect 9226 26432 9232 26488
rect 9992 26432 9998 26488
rect 10054 26432 10060 26488
rect 10820 26432 10826 26488
rect 10882 26432 10888 26488
rect 11648 26432 11654 26488
rect 11710 26432 11716 26488
rect 12476 26432 12482 26488
rect 12538 26432 12544 26488
rect 14960 26432 14966 26488
rect 15022 26432 15028 26488
rect 15788 26432 15794 26488
rect 15850 26432 15856 26488
rect 16616 26432 16622 26488
rect 16678 26432 16684 26488
rect 17444 26432 17450 26488
rect 17506 26432 17512 26488
rect 18272 26432 18278 26488
rect 18334 26432 18340 26488
rect 19100 26432 19106 26488
rect 19162 26432 19168 26488
rect 19934 26426 19990 26432
rect 20762 26488 20818 27794
rect 23246 26488 23302 27794
rect 24074 26488 24130 27794
rect 24902 26488 24958 27794
rect 25730 26488 25786 27794
rect 26558 26488 26614 27794
rect 23240 26432 23246 26488
rect 23302 26432 23308 26488
rect 24068 26432 24074 26488
rect 24130 26432 24136 26488
rect 24896 26432 24902 26488
rect 24958 26432 24964 26488
rect 25724 26432 25730 26488
rect 25786 26432 25792 26488
rect 20762 26426 20818 26432
rect 26558 26426 26614 26432
rect 27386 26488 27442 27794
rect 27386 26426 27442 26432
rect 28214 26488 28270 27794
rect 29042 26496 29098 27794
rect 29042 26434 29098 26440
rect 28214 26426 28270 26432
<< via2 >>
rect 11104 44208 11160 44264
rect 11840 44208 11896 44264
rect 12576 44208 12632 44264
rect 13312 44208 13368 44264
rect 14048 44208 14104 44264
rect 14784 44208 14840 44264
rect 15520 44208 15576 44264
rect 16256 44208 16312 44264
rect 16992 44208 17048 44264
rect 17728 44208 17784 44264
rect 24352 44208 24408 44264
rect 25088 44208 25144 44264
rect 25824 44208 25880 44264
rect 26560 44208 26616 44264
rect 27296 44208 27352 44264
rect 28032 44208 28088 44264
rect 28768 44208 28824 44264
rect 29504 44208 29560 44264
<< metal3 >>
rect 11094 44554 11100 44618
rect 11164 44554 11170 44618
rect 11830 44554 11836 44618
rect 11900 44554 11906 44618
rect 12566 44554 12572 44618
rect 12636 44554 12642 44618
rect 13302 44554 13308 44618
rect 13372 44554 13378 44618
rect 14038 44554 14044 44618
rect 14108 44554 14114 44618
rect 14774 44554 14780 44618
rect 14844 44554 14850 44618
rect 15510 44554 15516 44618
rect 15580 44554 15586 44618
rect 16246 44554 16252 44618
rect 16316 44554 16322 44618
rect 16982 44554 16988 44618
rect 17052 44554 17058 44618
rect 17718 44554 17724 44618
rect 17788 44554 17794 44618
rect 24342 44554 24348 44618
rect 24412 44554 24418 44618
rect 25078 44554 25084 44618
rect 25148 44554 25154 44618
rect 25814 44554 25820 44618
rect 25884 44554 25890 44618
rect 26550 44554 26556 44618
rect 26620 44554 26626 44618
rect 27286 44554 27292 44618
rect 27356 44554 27362 44618
rect 28022 44554 28028 44618
rect 28092 44554 28098 44618
rect 28758 44554 28764 44618
rect 28828 44554 28834 44618
rect 29494 44554 29500 44618
rect 29564 44554 29570 44618
rect 11102 44269 11162 44554
rect 11838 44269 11898 44554
rect 12574 44269 12634 44554
rect 13310 44269 13370 44554
rect 14046 44269 14106 44554
rect 14782 44269 14842 44554
rect 15518 44269 15578 44554
rect 16254 44269 16314 44554
rect 16990 44269 17050 44554
rect 17726 44269 17786 44554
rect 24350 44269 24410 44554
rect 25086 44269 25146 44554
rect 25822 44269 25882 44554
rect 26558 44269 26618 44554
rect 27294 44269 27354 44554
rect 28030 44269 28090 44554
rect 28766 44269 28826 44554
rect 29502 44269 29562 44554
rect 11099 44264 11165 44269
rect 11099 44208 11104 44264
rect 11160 44208 11165 44264
rect 11099 44203 11165 44208
rect 11835 44264 11901 44269
rect 11835 44208 11840 44264
rect 11896 44208 11901 44264
rect 11835 44203 11901 44208
rect 12571 44264 12637 44269
rect 12571 44208 12576 44264
rect 12632 44208 12637 44264
rect 12571 44203 12637 44208
rect 13307 44264 13373 44269
rect 13307 44208 13312 44264
rect 13368 44208 13373 44264
rect 13307 44203 13373 44208
rect 14043 44264 14109 44269
rect 14043 44208 14048 44264
rect 14104 44208 14109 44264
rect 14043 44203 14109 44208
rect 14779 44264 14845 44269
rect 14779 44208 14784 44264
rect 14840 44208 14845 44264
rect 14779 44203 14845 44208
rect 15515 44264 15581 44269
rect 15515 44208 15520 44264
rect 15576 44208 15581 44264
rect 15515 44203 15581 44208
rect 16251 44264 16317 44269
rect 16251 44208 16256 44264
rect 16312 44208 16317 44264
rect 16251 44203 16317 44208
rect 16987 44264 17053 44269
rect 16987 44208 16992 44264
rect 17048 44208 17053 44264
rect 16987 44203 17053 44208
rect 17723 44264 17789 44269
rect 17723 44208 17728 44264
rect 17784 44208 17789 44264
rect 17723 44203 17789 44208
rect 24347 44264 24413 44269
rect 24347 44208 24352 44264
rect 24408 44208 24413 44264
rect 24347 44203 24413 44208
rect 25083 44264 25149 44269
rect 25083 44208 25088 44264
rect 25144 44208 25149 44264
rect 25083 44203 25149 44208
rect 25819 44264 25885 44269
rect 25819 44208 25824 44264
rect 25880 44208 25885 44264
rect 25819 44203 25885 44208
rect 26555 44264 26621 44269
rect 26555 44208 26560 44264
rect 26616 44208 26621 44264
rect 26555 44203 26621 44208
rect 27291 44264 27357 44269
rect 27291 44208 27296 44264
rect 27352 44208 27357 44264
rect 27291 44203 27357 44208
rect 28027 44264 28093 44269
rect 28027 44208 28032 44264
rect 28088 44208 28093 44264
rect 28027 44203 28093 44208
rect 28763 44264 28829 44269
rect 28763 44208 28768 44264
rect 28824 44208 28829 44264
rect 28763 44203 28829 44208
rect 29499 44264 29565 44269
rect 29499 44208 29504 44264
rect 29560 44208 29565 44264
rect 29499 44203 29565 44208
rect 30964 42339 31044 42340
rect 30959 42261 30965 42339
rect 31043 42261 31049 42339
rect 30964 41722 31044 42261
rect 30304 41642 31044 41722
rect 30804 41201 30876 41202
rect 30799 41131 30805 41201
rect 30875 41131 30881 41201
rect 30804 40620 30876 41131
rect 30294 40548 30876 40620
<< via3 >>
rect 11100 44554 11164 44618
rect 11836 44554 11900 44618
rect 12572 44554 12636 44618
rect 13308 44554 13372 44618
rect 14044 44554 14108 44618
rect 14780 44554 14844 44618
rect 15516 44554 15580 44618
rect 16252 44554 16316 44618
rect 16988 44554 17052 44618
rect 17724 44554 17788 44618
rect 24348 44554 24412 44618
rect 25084 44554 25148 44618
rect 25820 44554 25884 44618
rect 26556 44554 26620 44618
rect 27292 44554 27356 44618
rect 28028 44554 28092 44618
rect 28764 44554 28828 44618
rect 29500 44554 29564 44618
rect 30965 42261 31043 42339
rect 30805 41131 30875 41201
<< metal4 >>
rect 798 44438 858 45152
rect 1534 44438 1594 45152
rect 2270 44438 2330 45152
rect 3006 44438 3066 45152
rect 3742 44438 3802 45152
rect 4478 44438 4538 45152
rect 5214 44438 5274 45152
rect 5950 44438 6010 45152
rect 6686 44438 6746 45152
rect 7422 44438 7482 45152
rect 8158 44438 8218 45152
rect 8894 44438 8954 45152
rect 9630 44438 9690 45152
rect 10366 44438 10426 45152
rect 11102 44619 11162 45152
rect 11838 44619 11898 45152
rect 12574 44619 12634 45152
rect 13310 44619 13370 45152
rect 14046 44619 14106 45152
rect 14782 44619 14842 45152
rect 15518 44619 15578 45152
rect 16254 44619 16314 45152
rect 16990 44619 17050 45152
rect 17726 44619 17786 45152
rect 18462 44854 18522 45152
rect 19198 44854 19258 45152
rect 19934 44854 19994 45152
rect 20670 44854 20730 45152
rect 21406 44854 21466 45152
rect 22142 44854 22202 45152
rect 22878 44854 22938 45152
rect 23614 44854 23674 45152
rect 24350 44619 24410 45152
rect 25086 44619 25146 45152
rect 25822 44619 25882 45152
rect 26558 44619 26618 45152
rect 27294 44619 27354 45152
rect 28030 44619 28090 45152
rect 28766 44619 28826 45152
rect 29502 44619 29562 45152
rect 11099 44618 11165 44619
rect 11099 44554 11100 44618
rect 11164 44554 11165 44618
rect 11099 44553 11165 44554
rect 11835 44618 11901 44619
rect 11835 44554 11836 44618
rect 11900 44554 11901 44618
rect 11835 44553 11901 44554
rect 12571 44618 12637 44619
rect 12571 44554 12572 44618
rect 12636 44554 12637 44618
rect 12571 44553 12637 44554
rect 13307 44618 13373 44619
rect 13307 44554 13308 44618
rect 13372 44554 13373 44618
rect 13307 44553 13373 44554
rect 14043 44618 14109 44619
rect 14043 44554 14044 44618
rect 14108 44554 14109 44618
rect 14043 44553 14109 44554
rect 14779 44618 14845 44619
rect 14779 44554 14780 44618
rect 14844 44554 14845 44618
rect 14779 44553 14845 44554
rect 15515 44618 15581 44619
rect 15515 44554 15516 44618
rect 15580 44554 15581 44618
rect 15515 44553 15581 44554
rect 16251 44618 16317 44619
rect 16251 44554 16252 44618
rect 16316 44554 16317 44618
rect 16251 44553 16317 44554
rect 16987 44618 17053 44619
rect 16987 44554 16988 44618
rect 17052 44554 17053 44618
rect 16987 44553 17053 44554
rect 17723 44618 17789 44619
rect 17723 44554 17724 44618
rect 17788 44554 17789 44618
rect 17723 44553 17789 44554
rect 24347 44618 24413 44619
rect 24347 44554 24348 44618
rect 24412 44554 24413 44618
rect 24347 44553 24413 44554
rect 25083 44618 25149 44619
rect 25083 44554 25084 44618
rect 25148 44554 25149 44618
rect 25083 44553 25149 44554
rect 25819 44618 25885 44619
rect 25819 44554 25820 44618
rect 25884 44554 25885 44618
rect 25819 44553 25885 44554
rect 26555 44618 26621 44619
rect 26555 44554 26556 44618
rect 26620 44554 26621 44618
rect 26555 44553 26621 44554
rect 27291 44618 27357 44619
rect 27291 44554 27292 44618
rect 27356 44554 27357 44618
rect 27291 44553 27357 44554
rect 28027 44618 28093 44619
rect 28027 44554 28028 44618
rect 28092 44554 28093 44618
rect 28027 44553 28093 44554
rect 28763 44618 28829 44619
rect 28763 44554 28764 44618
rect 28828 44554 28829 44618
rect 28763 44553 28829 44554
rect 29499 44618 29565 44619
rect 29499 44554 29500 44618
rect 29564 44554 29565 44618
rect 29499 44553 29565 44554
rect 11102 44438 11162 44553
rect 11838 44438 11898 44553
rect 12574 44438 12634 44553
rect 13310 44438 13370 44553
rect 14046 44438 14106 44553
rect 14782 44438 14842 44553
rect 15518 44438 15578 44553
rect 16254 44438 16314 44553
rect 16990 44438 17050 44553
rect 200 6137 500 44152
rect 2100 43926 5800 44438
rect 30238 44256 30298 45152
rect 30238 44196 30600 44256
rect 1083 6137 1285 6138
rect 200 5937 1285 6137
rect 200 1000 500 5937
rect 1083 5936 1285 5937
rect 3800 1000 4100 43926
rect 30540 42024 30600 44196
rect 30974 42340 31034 45152
rect 31710 44952 31770 45152
rect 30964 42339 31044 42340
rect 30964 42261 30965 42339
rect 31043 42261 31044 42339
rect 30964 42260 31044 42261
rect 30540 41964 30870 42024
rect 30810 41202 30870 41964
rect 30804 41201 30876 41202
rect 30804 41131 30805 41201
rect 30875 41131 30876 41201
rect 30804 41130 30876 41131
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 488
rect 31312 0 31432 488
use controller  controller_0
timestamp 1713497815
transform 1 0 6668 0 1 27738
box 14 0 24000 16000
use inverter  inverter_0
timestamp 1712241802
transform 1 0 6274 0 1 2809
box -410 547 1220 2810
use r2r  r2r_0
timestamp 1713380768
transform 0 1 28786 -1 0 25766
box -400 -5786 14766 800
use r2r  r2r_blue
timestamp 1713380768
transform 0 1 12386 -1 0 25766
box -400 -5786 14766 800
use r2r  r2r_green
timestamp 1713380768
transform 0 1 20586 -1 0 25766
box -400 -5786 14766 800
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 3800 1000 4100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
