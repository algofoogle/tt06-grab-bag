magic
tech sky130A
magscale 1 2
timestamp 1713487838
<< metal2 >>
rect 24398 43377 24482 43382
rect 24394 43303 24403 43377
rect 24477 43303 24486 43377
rect 23658 43078 23743 43083
rect 22760 43055 22840 43060
rect 22756 42985 22765 43055
rect 22835 42985 22844 43055
rect 23654 43003 23663 43078
rect 23738 43003 23747 43078
rect 22053 42932 22147 42936
rect 21408 42927 22152 42932
rect 21408 42833 22053 42927
rect 22147 42833 22152 42927
rect 21408 42828 22152 42833
rect 21408 41948 21512 42828
rect 22053 42824 22147 42828
rect 22760 42780 22840 42985
rect 23658 42783 23743 43003
rect 22240 42700 22840 42780
rect 22240 41960 22320 42700
rect 23078 42698 23743 42783
rect 24398 42782 24482 43303
rect 25304 42921 25376 42925
rect 27193 42923 27288 42928
rect 23898 42698 24482 42782
rect 24719 42916 25381 42921
rect 24719 42844 25304 42916
rect 25376 42844 25381 42916
rect 25561 42915 25640 42920
rect 25557 42846 25566 42915
rect 25635 42846 25644 42915
rect 26382 42914 26459 42919
rect 26378 42847 26387 42914
rect 26454 42847 26463 42914
rect 24719 42839 25381 42844
rect 23078 41958 23163 42698
rect 23898 41958 23982 42698
rect 24719 41939 24801 42839
rect 25304 42835 25376 42839
rect 25561 41941 25640 42846
rect 26382 41942 26459 42847
rect 27189 42838 27198 42923
rect 27283 42838 27292 42923
rect 28854 42921 28946 42926
rect 28041 42915 28120 42920
rect 28037 42846 28046 42915
rect 28115 42846 28124 42915
rect 27193 41953 27288 42838
rect 28041 41941 28120 42846
rect 28850 42839 28859 42921
rect 28941 42839 28950 42921
rect 29697 42918 29783 42923
rect 30514 42921 30606 42926
rect 29693 42842 29702 42918
rect 29778 42842 29787 42918
rect 28854 41934 28946 42839
rect 29697 41937 29783 42842
rect 30510 42839 30519 42921
rect 30601 42839 30610 42921
rect 30514 41954 30606 42839
<< via2 >>
rect 24403 43303 24477 43377
rect 22765 42985 22835 43055
rect 23663 43003 23738 43078
rect 22053 42833 22147 42927
rect 25304 42844 25376 42916
rect 25566 42846 25635 42915
rect 26387 42847 26454 42914
rect 27198 42838 27283 42923
rect 28046 42846 28115 42915
rect 28859 42839 28941 42921
rect 29702 42842 29778 42918
rect 30519 42839 30601 42921
<< metal3 >>
rect 25561 44299 25640 44300
rect 25556 44222 25562 44299
rect 25639 44222 25645 44299
rect 25075 43382 25157 43387
rect 24398 43381 25158 43382
rect 24398 43377 25075 43381
rect 24398 43303 24403 43377
rect 24477 43303 25075 43377
rect 24398 43299 25075 43303
rect 25157 43299 25158 43381
rect 25299 43380 25381 43381
rect 25294 43300 25300 43380
rect 25380 43300 25386 43380
rect 24398 43298 25158 43299
rect 25075 43293 25157 43298
rect 24099 43083 24182 43088
rect 23658 43082 24183 43083
rect 23658 43078 24099 43082
rect 22049 43072 22151 43077
rect 22048 43071 22152 43072
rect 22048 42969 22049 43071
rect 22151 42969 22152 43071
rect 23321 43060 23399 43065
rect 22760 43059 23400 43060
rect 22760 43055 23321 43059
rect 22760 42985 22765 43055
rect 22835 42985 23321 43055
rect 22760 42981 23321 42985
rect 23399 42981 23400 43059
rect 23658 43003 23663 43078
rect 23738 43003 24099 43078
rect 23658 42999 24099 43003
rect 24182 42999 24183 43082
rect 23658 42998 24183 42999
rect 24099 42993 24182 42998
rect 22760 42980 23400 42981
rect 23321 42975 23399 42980
rect 22048 42927 22152 42969
rect 22048 42833 22053 42927
rect 22147 42833 22152 42927
rect 25299 42916 25381 43300
rect 25299 42844 25304 42916
rect 25376 42844 25381 42916
rect 25299 42839 25381 42844
rect 25561 42915 25640 44222
rect 26382 44098 26459 44099
rect 26377 44023 26383 44098
rect 26458 44023 26464 44098
rect 25561 42846 25566 42915
rect 25635 42846 25640 42915
rect 25561 42841 25640 42846
rect 26382 42914 26459 44023
rect 26382 42847 26387 42914
rect 26454 42847 26459 42914
rect 26382 42842 26459 42847
rect 27193 43852 27288 43868
rect 27193 43788 27208 43852
rect 27272 43788 27288 43852
rect 27193 42923 27288 43788
rect 28041 43599 28120 43600
rect 28036 43522 28042 43599
rect 28119 43522 28125 43599
rect 27193 42838 27198 42923
rect 27283 42838 27288 42923
rect 28041 42915 28120 43522
rect 28854 43365 28946 43366
rect 28849 43275 28855 43365
rect 28945 43275 28951 43365
rect 28041 42846 28046 42915
rect 28115 42846 28120 42915
rect 28041 42841 28120 42846
rect 28854 42921 28946 43275
rect 30514 43125 30606 43126
rect 29697 43122 29783 43123
rect 29692 43038 29698 43122
rect 29782 43038 29788 43122
rect 27193 42833 27288 42838
rect 28854 42839 28859 42921
rect 28941 42839 28946 42921
rect 28854 42834 28946 42839
rect 29697 42918 29783 43038
rect 30509 43035 30515 43125
rect 30605 43035 30611 43125
rect 29697 42842 29702 42918
rect 29778 42842 29783 42918
rect 29697 42837 29783 42842
rect 30514 42921 30606 43035
rect 30514 42839 30519 42921
rect 30601 42839 30606 42921
rect 30514 42834 30606 42839
rect 22048 42828 22152 42833
<< via3 >>
rect 25562 44222 25639 44299
rect 25075 43299 25157 43381
rect 25300 43300 25380 43380
rect 22049 42969 22151 43071
rect 23321 42981 23399 43059
rect 24099 42999 24182 43082
rect 26383 44023 26458 44098
rect 27208 43788 27272 43852
rect 28042 43522 28119 43599
rect 28855 43275 28945 43365
rect 29698 43038 29782 43122
rect 30515 43035 30605 43125
<< metal4 >>
rect 798 44438 858 45152
rect 1534 44438 1594 45152
rect 2270 44438 2330 45152
rect 3006 44438 3066 45152
rect 3742 44438 3802 45152
rect 4478 44438 4538 45152
rect 5214 44438 5274 45152
rect 5950 44438 6010 45152
rect 6686 44438 6746 45152
rect 7422 44438 7482 45152
rect 8158 44438 8218 45152
rect 8894 44438 8954 45152
rect 9630 44438 9690 45152
rect 10366 44438 10426 45152
rect 11102 44438 11162 45152
rect 11838 44438 11898 45152
rect 12574 44438 12634 45152
rect 13310 44438 13370 45152
rect 14046 44438 14106 45152
rect 14782 44438 14842 45152
rect 15518 44438 15578 45152
rect 16254 44438 16314 45152
rect 16990 44438 17050 45152
rect 17726 44688 17786 45152
rect 18462 44688 18522 45152
rect 19198 44688 19258 45152
rect 19934 44688 19994 45152
rect 20670 44688 20730 45152
rect 21406 44688 21466 45152
rect 22142 44688 22202 45152
rect 200 6137 500 44152
rect 2100 43926 5800 44438
rect 1083 6137 1285 6138
rect 200 5937 1285 6137
rect 200 1000 500 5937
rect 1083 5936 1285 5937
rect 3800 1000 4100 43926
rect 22878 43310 22938 45152
rect 23614 43310 23674 45152
rect 24350 43630 24410 45152
rect 22530 43250 22938 43310
rect 23330 43250 23674 43310
rect 24110 43570 24410 43630
rect 22048 43071 22152 43072
rect 22048 42969 22049 43071
rect 22151 43050 22152 43071
rect 22530 43050 22590 43250
rect 23330 43060 23390 43250
rect 24110 43083 24170 43570
rect 25086 43382 25146 45152
rect 25822 44490 25882 45152
rect 25310 44430 25882 44490
rect 25074 43381 25158 43382
rect 25310 43381 25370 44430
rect 25561 44299 25640 44300
rect 25561 44222 25562 44299
rect 25639 44290 25640 44299
rect 26558 44290 26618 45152
rect 25639 44230 26618 44290
rect 25639 44222 25640 44230
rect 25561 44221 25640 44222
rect 26382 44098 26459 44099
rect 26382 44023 26383 44098
rect 26458 44090 26459 44098
rect 27294 44090 27354 45152
rect 26458 44030 27354 44090
rect 26458 44023 26459 44030
rect 26382 44022 26459 44023
rect 27207 43852 27273 43853
rect 27207 43788 27208 43852
rect 27272 43850 27273 43852
rect 28030 43850 28090 45152
rect 27272 43790 28090 43850
rect 27272 43788 27273 43790
rect 27207 43787 27273 43788
rect 28041 43599 28120 43600
rect 28041 43522 28042 43599
rect 28119 43590 28120 43599
rect 28766 43590 28826 45152
rect 29502 44817 29562 45152
rect 28119 43530 28826 43590
rect 28119 43522 28120 43530
rect 28041 43521 28120 43522
rect 25074 43299 25075 43381
rect 25157 43299 25158 43381
rect 25299 43380 25381 43381
rect 25299 43300 25300 43380
rect 25380 43300 25381 43380
rect 25299 43299 25381 43300
rect 28854 43365 28946 43366
rect 25074 43298 25158 43299
rect 28854 43275 28855 43365
rect 28945 43353 28946 43365
rect 29499 43353 29565 44817
rect 28945 43287 29565 43353
rect 28945 43275 28946 43287
rect 28854 43274 28946 43275
rect 29697 43122 29783 43123
rect 24098 43082 24183 43083
rect 22151 42990 22590 43050
rect 23320 43059 23400 43060
rect 22151 42969 22152 42990
rect 23320 42981 23321 43059
rect 23399 42981 23400 43059
rect 24098 42999 24099 43082
rect 24182 42999 24183 43082
rect 29697 43038 29698 43122
rect 29782 43110 29783 43122
rect 30238 43110 30298 45152
rect 29782 43050 30298 43110
rect 30514 43125 30606 43126
rect 29782 43038 29783 43050
rect 29697 43037 29783 43038
rect 30514 43035 30515 43125
rect 30605 43110 30606 43125
rect 30974 43110 31034 45152
rect 31710 44952 31770 45152
rect 30605 43050 31034 43110
rect 30605 43035 30606 43050
rect 30514 43034 30606 43035
rect 24098 42998 24183 42999
rect 23320 42980 23400 42981
rect 22048 42968 22152 42969
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 488
rect 31312 0 31432 488
use controller  controller_0
timestamp 1713486661
transform 1 0 13590 0 1 24046
box 514 0 17724 18245
use inverter  inverter_0
timestamp 1712241802
transform 1 0 6274 0 1 2809
box -410 547 1220 2810
use r2r  r2r_blue
timestamp 1713380768
transform 0 1 15786 -1 0 20766
box -400 -5786 14766 800
use r2r  r2r_green
timestamp 1713380768
transform 0 1 23186 -1 0 20766
box -400 -5786 14766 800
use r2r  r2r_red
timestamp 1713380768
transform 0 1 30586 -1 0 20766
box -400 -5786 14766 800
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 3800 1000 4100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
