MACRO tt_um_algofoogle_tt06_grab_bag
  CLASS BLOCK ;
  FOREIGN tt_um_algofoogle_tt06_grab_bag ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 19.000 5.000 20.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 70.520 205.855 156.460 207.460 ;
      LAYER pwell ;
        RECT 70.715 204.655 72.085 205.465 ;
        RECT 72.095 204.655 73.465 205.465 ;
        RECT 73.485 204.655 76.225 205.335 ;
        RECT 76.235 204.655 77.605 205.435 ;
        RECT 77.615 205.335 78.960 205.565 ;
        RECT 79.455 205.335 80.385 205.565 ;
        RECT 77.615 204.655 79.445 205.335 ;
        RECT 79.455 204.655 83.355 205.335 ;
        RECT 83.605 204.740 84.035 205.525 ;
        RECT 84.150 205.335 85.070 205.565 ;
        RECT 87.735 205.335 89.080 205.565 ;
        RECT 84.150 204.655 87.615 205.335 ;
        RECT 87.735 204.655 89.565 205.335 ;
        RECT 89.575 204.655 90.945 205.465 ;
        RECT 90.955 205.335 92.300 205.565 ;
        RECT 90.955 204.655 92.785 205.335 ;
        RECT 92.795 204.655 95.535 205.335 ;
        RECT 96.485 204.740 96.915 205.525 ;
        RECT 96.945 204.655 99.685 205.335 ;
        RECT 100.630 204.655 102.445 205.565 ;
        RECT 103.860 205.335 105.205 205.565 ;
        RECT 105.700 205.335 107.045 205.565 ;
        RECT 108.000 205.335 109.345 205.565 ;
        RECT 103.375 204.655 105.205 205.335 ;
        RECT 105.215 204.655 107.045 205.335 ;
        RECT 107.515 204.655 109.345 205.335 ;
        RECT 109.365 204.740 109.795 205.525 ;
        RECT 109.825 204.655 111.175 205.565 ;
        RECT 111.655 205.335 113.000 205.565 ;
        RECT 111.655 204.655 113.485 205.335 ;
        RECT 113.495 204.655 114.865 205.435 ;
        RECT 115.795 204.655 117.165 205.435 ;
        RECT 117.175 204.655 118.545 205.435 ;
        RECT 118.650 205.335 119.570 205.565 ;
        RECT 118.650 204.655 122.115 205.335 ;
        RECT 122.245 204.740 122.675 205.525 ;
        RECT 123.155 205.335 124.085 205.565 ;
        RECT 127.295 205.335 128.225 205.565 ;
        RECT 131.530 205.335 132.450 205.565 ;
        RECT 123.155 204.655 127.055 205.335 ;
        RECT 127.295 204.655 131.195 205.335 ;
        RECT 131.530 204.655 134.995 205.335 ;
        RECT 135.125 204.740 135.555 205.525 ;
        RECT 135.575 204.655 136.945 205.435 ;
        RECT 136.955 204.655 138.325 205.435 ;
        RECT 138.335 204.655 139.705 205.435 ;
        RECT 144.150 205.335 145.060 205.555 ;
        RECT 146.595 205.335 147.945 205.565 ;
        RECT 140.635 204.655 147.945 205.335 ;
        RECT 148.005 204.740 148.435 205.525 ;
        RECT 149.575 205.335 153.505 205.565 ;
        RECT 149.090 204.655 153.505 205.335 ;
        RECT 153.515 204.655 154.885 205.465 ;
        RECT 154.895 204.655 156.265 205.465 ;
        RECT 70.855 204.445 71.025 204.655 ;
        RECT 72.235 204.465 72.405 204.655 ;
        RECT 73.155 204.445 73.325 204.635 ;
        RECT 75.915 204.465 76.085 204.655 ;
        RECT 77.295 204.465 77.465 204.655 ;
        RECT 79.135 204.465 79.305 204.655 ;
        RECT 79.870 204.465 80.040 204.655 ;
        RECT 80.515 204.445 80.685 204.635 ;
        RECT 83.270 204.445 83.440 204.635 ;
        RECT 83.735 204.445 83.905 204.635 ;
        RECT 87.415 204.465 87.585 204.655 ;
        RECT 89.255 204.465 89.425 204.655 ;
        RECT 89.715 204.465 89.885 204.655 ;
        RECT 92.015 204.445 92.185 204.635 ;
        RECT 92.475 204.465 92.645 204.655 ;
        RECT 92.935 204.465 93.105 204.655 ;
        RECT 93.405 204.445 93.575 204.635 ;
        RECT 95.695 204.445 95.865 204.635 ;
        RECT 96.150 204.495 96.270 204.605 ;
        RECT 97.075 204.445 97.245 204.635 ;
        RECT 99.375 204.465 99.545 204.655 ;
        RECT 99.845 204.500 100.005 204.610 ;
        RECT 100.290 204.495 100.410 204.605 ;
        RECT 100.755 204.465 100.925 204.655 ;
        RECT 103.515 204.635 103.685 204.655 ;
        RECT 102.605 204.500 102.765 204.610 ;
        RECT 103.510 204.465 103.685 204.635 ;
        RECT 103.985 204.490 104.145 204.600 ;
        RECT 70.715 203.635 72.085 204.445 ;
        RECT 73.015 203.765 80.325 204.445 ;
        RECT 76.530 203.545 77.440 203.765 ;
        RECT 78.975 203.535 80.325 203.765 ;
        RECT 80.375 203.635 82.205 204.445 ;
        RECT 82.235 203.535 83.585 204.445 ;
        RECT 83.595 203.765 90.905 204.445 ;
        RECT 87.110 203.545 88.020 203.765 ;
        RECT 89.555 203.535 90.905 203.765 ;
        RECT 90.955 203.665 92.325 204.445 ;
        RECT 93.255 203.665 94.625 204.445 ;
        RECT 94.635 203.665 96.005 204.445 ;
        RECT 96.485 203.575 96.915 204.360 ;
        RECT 97.035 203.535 100.145 204.445 ;
        RECT 100.615 204.415 101.550 204.445 ;
        RECT 103.510 204.415 103.680 204.465 ;
        RECT 105.170 204.445 105.340 204.635 ;
        RECT 105.355 204.465 105.525 204.655 ;
        RECT 107.190 204.495 107.310 204.605 ;
        RECT 107.655 204.465 107.825 204.655 ;
        RECT 110.875 204.465 111.045 204.655 ;
        RECT 111.330 204.495 111.450 204.605 ;
        RECT 113.175 204.465 113.345 204.655 ;
        RECT 113.635 204.465 113.805 204.655 ;
        RECT 115.025 204.500 115.185 204.610 ;
        RECT 115.935 204.445 116.105 204.635 ;
        RECT 116.855 204.465 117.025 204.655 ;
        RECT 117.315 204.445 117.485 204.655 ;
        RECT 118.050 204.445 118.220 204.635 ;
        RECT 121.915 204.605 122.085 204.655 ;
        RECT 122.835 204.605 123.005 204.635 ;
        RECT 121.910 204.495 122.085 204.605 ;
        RECT 122.830 204.495 123.005 204.605 ;
        RECT 121.915 204.465 122.085 204.495 ;
        RECT 122.835 204.445 123.005 204.495 ;
        RECT 123.570 204.465 123.740 204.655 ;
        RECT 124.215 204.445 124.385 204.635 ;
        RECT 125.595 204.445 125.765 204.635 ;
        RECT 127.710 204.465 127.880 204.655 ;
        RECT 132.950 204.495 133.070 204.605 ;
        RECT 134.325 204.445 134.495 204.635 ;
        RECT 134.795 204.465 134.965 204.655 ;
        RECT 135.715 204.445 135.885 204.635 ;
        RECT 136.635 204.465 136.805 204.655 ;
        RECT 137.095 204.445 137.265 204.635 ;
        RECT 138.015 204.465 138.185 204.655 ;
        RECT 139.395 204.465 139.565 204.655 ;
        RECT 139.865 204.500 140.025 204.610 ;
        RECT 140.775 204.465 140.945 204.655 ;
        RECT 149.090 204.635 149.200 204.655 ;
        RECT 153.655 204.635 153.825 204.655 ;
        RECT 145.375 204.445 145.545 204.635 ;
        RECT 146.755 204.445 146.925 204.635 ;
        RECT 147.225 204.490 147.385 204.600 ;
        RECT 148.590 204.495 148.710 204.605 ;
        RECT 148.870 204.465 149.200 204.635 ;
        RECT 153.645 204.465 153.825 204.635 ;
        RECT 154.125 204.490 154.285 204.600 ;
        RECT 148.870 204.445 149.040 204.465 ;
        RECT 153.645 204.445 153.815 204.465 ;
        RECT 155.955 204.445 156.125 204.655 ;
        RECT 100.615 204.215 103.680 204.415 ;
        RECT 100.615 203.735 103.825 204.215 ;
        RECT 100.615 203.535 101.565 203.735 ;
        RECT 102.895 203.535 103.825 203.735 ;
        RECT 104.755 203.765 108.655 204.445 ;
        RECT 108.935 203.765 116.245 204.445 ;
        RECT 104.755 203.535 105.685 203.765 ;
        RECT 108.935 203.535 110.285 203.765 ;
        RECT 111.820 203.545 112.730 203.765 ;
        RECT 116.255 203.665 117.625 204.445 ;
        RECT 117.635 203.765 121.535 204.445 ;
        RECT 117.635 203.535 118.565 203.765 ;
        RECT 122.245 203.575 122.675 204.360 ;
        RECT 122.695 203.635 124.065 204.445 ;
        RECT 124.075 203.665 125.445 204.445 ;
        RECT 125.455 203.765 132.765 204.445 ;
        RECT 128.970 203.545 129.880 203.765 ;
        RECT 131.415 203.535 132.765 203.765 ;
        RECT 133.275 203.665 134.645 204.445 ;
        RECT 135.575 203.665 136.945 204.445 ;
        RECT 136.955 203.765 144.265 204.445 ;
        RECT 140.470 203.545 141.380 203.765 ;
        RECT 142.915 203.535 144.265 203.765 ;
        RECT 144.315 203.665 145.685 204.445 ;
        RECT 145.695 203.665 147.065 204.445 ;
        RECT 148.005 203.575 148.435 204.360 ;
        RECT 148.455 203.765 152.355 204.445 ;
        RECT 148.455 203.535 149.385 203.765 ;
        RECT 152.595 203.665 153.965 204.445 ;
        RECT 154.895 203.635 156.265 204.445 ;
      LAYER nwell ;
        RECT 70.520 200.415 156.460 203.245 ;
      LAYER pwell ;
        RECT 70.715 199.215 72.085 200.025 ;
        RECT 72.095 199.215 73.925 200.025 ;
        RECT 77.450 199.895 78.360 200.115 ;
        RECT 79.895 199.895 81.245 200.125 ;
        RECT 73.935 199.215 81.245 199.895 ;
        RECT 82.215 199.215 83.585 199.995 ;
        RECT 83.605 199.300 84.035 200.085 ;
        RECT 84.095 199.895 85.445 200.125 ;
        RECT 86.980 199.895 87.890 200.115 ;
        RECT 95.390 199.895 96.300 200.115 ;
        RECT 97.835 199.895 99.185 200.125 ;
        RECT 102.435 199.895 103.365 200.125 ;
        RECT 84.095 199.215 91.405 199.895 ;
        RECT 91.875 199.215 99.185 199.895 ;
        RECT 99.465 199.215 103.365 199.895 ;
        RECT 104.495 200.035 105.445 200.125 ;
        RECT 104.495 199.215 106.425 200.035 ;
        RECT 106.615 199.215 107.965 200.125 ;
        RECT 107.985 199.215 109.335 200.125 ;
        RECT 109.365 199.300 109.795 200.085 ;
        RECT 110.735 199.215 113.485 200.125 ;
        RECT 117.930 199.895 118.840 200.115 ;
        RECT 120.375 199.895 121.725 200.125 ;
        RECT 114.415 199.215 121.725 199.895 ;
        RECT 121.775 199.215 124.525 200.125 ;
        RECT 128.195 199.895 129.125 200.125 ;
        RECT 125.225 199.215 129.125 199.895 ;
        RECT 129.135 199.215 131.885 200.125 ;
        RECT 132.355 199.215 135.105 200.125 ;
        RECT 135.125 199.300 135.555 200.085 ;
        RECT 135.575 199.895 136.505 200.125 ;
        RECT 145.215 199.895 146.145 200.125 ;
        RECT 149.670 199.895 150.580 200.115 ;
        RECT 152.115 199.895 153.465 200.125 ;
        RECT 135.575 199.215 139.475 199.895 ;
        RECT 139.715 199.215 141.545 199.895 ;
        RECT 142.245 199.215 146.145 199.895 ;
        RECT 146.155 199.215 153.465 199.895 ;
        RECT 153.515 199.215 154.885 200.025 ;
        RECT 154.895 199.215 156.265 200.025 ;
        RECT 70.855 199.005 71.025 199.215 ;
        RECT 72.235 199.005 72.405 199.215 ;
        RECT 74.075 199.025 74.245 199.215 ;
        RECT 74.995 199.005 75.165 199.195 ;
        RECT 80.055 199.025 80.225 199.195 ;
        RECT 80.055 199.005 80.075 199.025 ;
        RECT 70.715 198.195 72.085 199.005 ;
        RECT 72.095 198.195 74.845 199.005 ;
        RECT 74.855 198.095 77.605 199.005 ;
        RECT 77.625 198.325 80.075 199.005 ;
        RECT 80.520 198.975 80.690 199.195 ;
        RECT 81.445 199.060 81.605 199.170 ;
        RECT 82.355 199.025 82.525 199.215 ;
        RECT 83.745 199.005 83.915 199.195 ;
        RECT 85.125 199.050 85.285 199.160 ;
        RECT 86.945 199.005 87.115 199.195 ;
        RECT 88.325 199.005 88.495 199.195 ;
        RECT 89.705 199.005 89.875 199.195 ;
        RECT 91.095 199.025 91.265 199.215 ;
        RECT 92.015 199.195 92.185 199.215 ;
        RECT 91.555 199.165 91.725 199.195 ;
        RECT 91.550 199.055 91.725 199.165 ;
        RECT 91.555 199.005 91.725 199.055 ;
        RECT 92.015 199.025 92.190 199.195 ;
        RECT 92.020 199.005 92.190 199.025 ;
        RECT 95.245 199.005 95.415 199.195 ;
        RECT 97.085 199.005 97.255 199.195 ;
        RECT 98.450 199.005 98.620 199.195 ;
        RECT 99.835 199.005 100.005 199.195 ;
        RECT 101.670 199.055 101.790 199.165 ;
        RECT 102.780 199.025 102.950 199.215 ;
        RECT 106.275 199.195 106.425 199.215 ;
        RECT 103.525 199.060 103.685 199.170 ;
        RECT 104.435 199.005 104.605 199.195 ;
        RECT 106.275 199.025 106.445 199.195 ;
        RECT 107.650 199.025 107.820 199.215 ;
        RECT 108.115 199.195 108.285 199.215 ;
        RECT 108.110 199.025 108.285 199.195 ;
        RECT 108.110 199.005 108.280 199.025 ;
        RECT 108.575 199.005 108.745 199.195 ;
        RECT 109.965 199.060 110.125 199.170 ;
        RECT 110.875 199.025 111.045 199.215 ;
        RECT 112.265 199.050 112.425 199.160 ;
        RECT 113.645 199.060 113.805 199.170 ;
        RECT 114.085 199.005 114.255 199.195 ;
        RECT 114.555 199.165 114.725 199.215 ;
        RECT 114.550 199.055 114.725 199.165 ;
        RECT 114.555 199.025 114.725 199.055 ;
        RECT 115.025 199.005 115.195 199.195 ;
        RECT 116.395 199.005 116.565 199.195 ;
        RECT 119.155 199.005 119.325 199.195 ;
        RECT 121.915 199.165 122.085 199.215 ;
        RECT 121.910 199.055 122.085 199.165 ;
        RECT 121.915 199.025 122.085 199.055 ;
        RECT 122.835 199.005 123.005 199.195 ;
        RECT 124.670 199.055 124.790 199.165 ;
        RECT 125.605 199.050 125.765 199.160 ;
        RECT 127.430 199.005 127.600 199.195 ;
        RECT 128.540 199.025 128.710 199.215 ;
        RECT 129.275 199.025 129.445 199.215 ;
        RECT 132.495 199.195 132.665 199.215 ;
        RECT 132.060 199.165 132.230 199.195 ;
        RECT 132.030 199.055 132.230 199.165 ;
        RECT 132.060 199.025 132.230 199.055 ;
        RECT 132.490 199.025 132.665 199.195 ;
        RECT 132.060 199.005 132.170 199.025 ;
        RECT 82.650 198.975 83.585 199.005 ;
        RECT 80.520 198.775 83.585 198.975 ;
        RECT 77.625 198.095 79.585 198.325 ;
        RECT 80.375 198.295 83.585 198.775 ;
        RECT 80.375 198.095 81.305 198.295 ;
        RECT 82.635 198.095 83.585 198.295 ;
        RECT 83.595 198.225 84.965 199.005 ;
        RECT 85.895 198.225 87.265 199.005 ;
        RECT 87.275 198.225 88.645 199.005 ;
        RECT 88.655 198.225 90.025 199.005 ;
        RECT 90.035 198.325 91.865 199.005 ;
        RECT 91.875 198.095 94.795 199.005 ;
        RECT 95.095 198.225 96.465 199.005 ;
        RECT 96.485 198.135 96.915 198.920 ;
        RECT 96.935 198.225 98.305 199.005 ;
        RECT 98.335 198.095 99.685 199.005 ;
        RECT 99.695 198.195 101.525 199.005 ;
        RECT 101.995 198.095 104.745 199.005 ;
        RECT 104.950 198.095 108.425 199.005 ;
        RECT 108.435 198.195 112.105 199.005 ;
        RECT 113.035 198.225 114.405 199.005 ;
        RECT 114.875 198.225 116.245 199.005 ;
        RECT 116.255 198.095 119.005 199.005 ;
        RECT 119.015 198.195 121.765 199.005 ;
        RECT 122.245 198.135 122.675 198.920 ;
        RECT 122.695 198.095 125.445 199.005 ;
        RECT 126.395 198.095 127.745 199.005 ;
        RECT 127.755 198.325 132.170 199.005 ;
        RECT 132.490 198.975 132.660 199.025 ;
        RECT 135.715 199.005 135.885 199.195 ;
        RECT 135.990 199.025 136.160 199.215 ;
        RECT 136.170 199.055 136.290 199.165 ;
        RECT 136.635 199.005 136.805 199.195 ;
        RECT 139.395 199.005 139.565 199.195 ;
        RECT 141.235 199.025 141.405 199.215 ;
        RECT 141.690 199.055 141.810 199.165 ;
        RECT 142.165 199.005 142.335 199.195 ;
        RECT 143.535 199.005 143.705 199.195 ;
        RECT 145.375 199.005 145.545 199.195 ;
        RECT 145.560 199.025 145.730 199.215 ;
        RECT 146.295 199.025 146.465 199.215 ;
        RECT 147.675 199.005 147.845 199.195 ;
        RECT 148.595 199.005 148.765 199.195 ;
        RECT 151.350 199.055 151.470 199.165 ;
        RECT 152.735 199.005 152.905 199.195 ;
        RECT 153.655 199.025 153.825 199.215 ;
        RECT 154.105 199.005 154.275 199.195 ;
        RECT 154.570 199.055 154.690 199.165 ;
        RECT 155.955 199.005 156.125 199.215 ;
        RECT 133.690 198.975 134.645 199.005 ;
        RECT 127.755 198.095 131.685 198.325 ;
        RECT 132.365 198.295 134.645 198.975 ;
        RECT 133.690 198.095 134.645 198.295 ;
        RECT 134.655 198.225 136.025 199.005 ;
        RECT 136.495 198.095 139.245 199.005 ;
        RECT 139.255 198.095 142.005 199.005 ;
        RECT 142.015 198.225 143.385 199.005 ;
        RECT 143.395 198.195 145.225 199.005 ;
        RECT 145.235 198.225 146.605 199.005 ;
        RECT 146.615 198.225 147.985 199.005 ;
        RECT 148.005 198.135 148.435 198.920 ;
        RECT 148.455 198.195 151.205 199.005 ;
        RECT 151.685 198.095 153.035 199.005 ;
        RECT 153.055 198.225 154.425 199.005 ;
        RECT 154.895 198.195 156.265 199.005 ;
      LAYER nwell ;
        RECT 70.520 194.975 156.460 197.805 ;
      LAYER pwell ;
        RECT 70.715 193.775 72.085 194.585 ;
        RECT 75.610 194.455 76.520 194.675 ;
        RECT 78.055 194.455 79.405 194.685 ;
        RECT 72.095 193.775 79.405 194.455 ;
        RECT 79.455 193.775 81.285 194.585 ;
        RECT 81.295 194.455 82.215 194.685 ;
        RECT 81.295 193.775 83.585 194.455 ;
        RECT 83.605 193.860 84.035 194.645 ;
        RECT 84.055 193.775 86.975 194.685 ;
        RECT 87.355 193.775 90.355 194.685 ;
        RECT 93.695 194.455 94.625 194.685 ;
        RECT 90.955 193.775 94.625 194.455 ;
        RECT 94.635 194.455 95.565 194.685 ;
        RECT 101.430 194.455 102.350 194.685 ;
        RECT 104.990 194.455 106.125 194.685 ;
        RECT 94.635 193.775 98.305 194.455 ;
        RECT 98.885 193.775 102.350 194.455 ;
        RECT 102.915 193.775 106.125 194.455 ;
        RECT 106.135 194.485 107.065 194.685 ;
        RECT 108.400 194.485 109.345 194.685 ;
        RECT 106.135 194.005 109.345 194.485 ;
        RECT 106.275 193.805 109.345 194.005 ;
        RECT 109.365 193.860 109.795 194.645 ;
        RECT 111.150 194.485 112.105 194.685 ;
        RECT 109.825 193.805 112.105 194.485 ;
        RECT 70.855 193.565 71.025 193.775 ;
        RECT 72.235 193.565 72.405 193.775 ;
        RECT 75.000 193.565 75.170 193.755 ;
        RECT 76.835 193.565 77.005 193.755 ;
        RECT 78.675 193.565 78.845 193.755 ;
        RECT 79.595 193.585 79.765 193.775 ;
        RECT 80.060 193.565 80.230 193.755 ;
        RECT 83.275 193.585 83.445 193.775 ;
        RECT 84.200 193.585 84.370 193.775 ;
        RECT 87.415 193.755 87.585 193.775 ;
        RECT 87.415 193.585 87.610 193.755 ;
        RECT 87.870 193.615 87.990 193.725 ;
        RECT 87.440 193.565 87.550 193.585 ;
        RECT 88.335 193.565 88.505 193.755 ;
        RECT 90.630 193.615 90.750 193.725 ;
        RECT 91.095 193.585 91.265 193.775 ;
        RECT 97.995 193.585 98.165 193.775 ;
        RECT 98.450 193.615 98.570 193.725 ;
        RECT 98.915 193.585 99.085 193.775 ;
        RECT 101.215 193.565 101.385 193.755 ;
        RECT 101.670 193.615 101.790 193.725 ;
        RECT 70.715 192.755 72.085 193.565 ;
        RECT 72.095 192.755 74.845 193.565 ;
        RECT 74.855 192.655 76.685 193.565 ;
        RECT 76.710 192.655 78.525 193.565 ;
        RECT 78.535 192.755 79.905 193.565 ;
        RECT 79.915 192.655 82.835 193.565 ;
        RECT 83.135 192.885 87.550 193.565 ;
        RECT 88.195 192.885 96.465 193.565 ;
        RECT 96.945 193.525 97.865 193.565 ;
        RECT 83.135 192.655 87.065 192.885 ;
        RECT 95.015 192.655 96.465 192.885 ;
        RECT 96.485 192.695 96.915 193.480 ;
        RECT 96.935 193.335 97.865 193.525 ;
        RECT 99.955 193.335 101.525 193.565 ;
        RECT 102.135 193.335 102.305 193.755 ;
        RECT 102.590 193.615 102.710 193.725 ;
        RECT 103.055 193.585 103.225 193.775 ;
        RECT 106.275 193.565 106.445 193.805 ;
        RECT 108.400 193.775 109.345 193.805 ;
        RECT 109.950 193.585 110.120 193.805 ;
        RECT 111.150 193.775 112.105 193.805 ;
        RECT 112.115 193.775 117.625 194.585 ;
        RECT 117.635 193.775 123.145 194.585 ;
        RECT 125.495 194.455 126.845 194.685 ;
        RECT 128.380 194.455 129.290 194.675 ;
        RECT 123.615 193.775 125.445 194.455 ;
        RECT 125.495 193.775 132.805 194.455 ;
        RECT 132.815 193.775 134.185 194.555 ;
        RECT 135.125 193.860 135.555 194.645 ;
        RECT 135.575 193.775 136.945 194.555 ;
        RECT 136.955 193.775 138.325 194.555 ;
        RECT 139.255 194.485 140.185 194.685 ;
        RECT 141.515 194.485 142.465 194.685 ;
        RECT 139.255 194.005 142.465 194.485 ;
        RECT 139.400 193.805 142.465 194.005 ;
        RECT 112.255 193.585 112.425 193.775 ;
        RECT 114.550 193.615 114.670 193.725 ;
        RECT 115.015 193.565 115.185 193.755 ;
        RECT 116.855 193.565 117.025 193.755 ;
        RECT 117.775 193.585 117.945 193.775 ;
        RECT 103.415 193.335 106.125 193.565 ;
        RECT 96.935 192.975 101.525 193.335 ;
        RECT 96.945 192.885 101.525 192.975 ;
        RECT 102.030 192.885 106.125 193.335 ;
        RECT 106.135 192.885 114.405 193.565 ;
        RECT 114.875 192.885 116.705 193.565 ;
        RECT 96.945 192.655 99.945 192.885 ;
        RECT 102.030 192.655 103.405 192.885 ;
        RECT 105.175 192.655 106.125 192.885 ;
        RECT 112.955 192.655 114.405 192.885 ;
        RECT 116.715 192.755 118.545 193.565 ;
        RECT 118.555 193.535 119.500 193.565 ;
        RECT 120.990 193.535 121.160 193.755 ;
        RECT 121.465 193.610 121.625 193.720 ;
        RECT 122.845 193.565 123.015 193.755 ;
        RECT 123.290 193.615 123.410 193.725 ;
        RECT 124.215 193.565 124.385 193.755 ;
        RECT 125.135 193.585 125.305 193.775 ;
        RECT 126.050 193.615 126.170 193.725 ;
        RECT 128.355 193.585 128.525 193.755 ;
        RECT 128.355 193.565 128.505 193.585 ;
        RECT 118.555 192.855 121.305 193.535 ;
        RECT 118.555 192.655 119.500 192.855 ;
        RECT 122.245 192.695 122.675 193.480 ;
        RECT 122.695 192.785 124.065 193.565 ;
        RECT 124.075 192.755 125.905 193.565 ;
        RECT 126.575 192.745 128.505 193.565 ;
        RECT 128.820 193.535 128.990 193.755 ;
        RECT 132.045 193.565 132.215 193.755 ;
        RECT 132.495 193.585 132.665 193.775 ;
        RECT 133.415 193.565 133.585 193.755 ;
        RECT 133.865 193.585 134.035 193.775 ;
        RECT 134.345 193.620 134.505 193.730 ;
        RECT 135.725 193.585 135.895 193.775 ;
        RECT 136.170 193.615 136.290 193.725 ;
        RECT 136.635 193.565 136.805 193.755 ;
        RECT 137.105 193.585 137.275 193.775 ;
        RECT 139.400 193.755 139.570 193.805 ;
        RECT 141.530 193.775 142.465 193.805 ;
        RECT 142.475 193.775 145.225 194.585 ;
        RECT 145.235 193.775 146.605 194.555 ;
        RECT 150.590 194.455 151.500 194.675 ;
        RECT 153.035 194.455 154.385 194.685 ;
        RECT 147.075 193.775 154.385 194.455 ;
        RECT 154.895 193.775 156.265 194.585 ;
        RECT 138.485 193.610 138.645 193.730 ;
        RECT 139.395 193.585 139.570 193.755 ;
        RECT 142.615 193.585 142.785 193.775 ;
        RECT 145.375 193.585 145.545 193.775 ;
        RECT 146.750 193.615 146.870 193.725 ;
        RECT 147.215 193.585 147.385 193.775 ;
        RECT 139.395 193.565 139.565 193.585 ;
        RECT 147.665 193.565 147.835 193.755 ;
        RECT 148.595 193.565 148.765 193.755 ;
        RECT 154.125 193.610 154.285 193.720 ;
        RECT 154.570 193.615 154.690 193.725 ;
        RECT 155.955 193.565 156.125 193.775 ;
        RECT 130.950 193.535 131.885 193.565 ;
        RECT 128.820 193.335 131.885 193.535 ;
        RECT 128.675 192.855 131.885 193.335 ;
        RECT 126.575 192.655 127.525 192.745 ;
        RECT 128.675 192.655 129.605 192.855 ;
        RECT 130.935 192.655 131.885 192.855 ;
        RECT 131.895 192.785 133.265 193.565 ;
        RECT 133.275 192.755 136.025 193.565 ;
        RECT 136.510 192.655 138.325 193.565 ;
        RECT 139.255 192.885 146.565 193.565 ;
        RECT 142.770 192.665 143.680 192.885 ;
        RECT 145.215 192.655 146.565 192.885 ;
        RECT 146.615 192.785 147.985 193.565 ;
        RECT 148.005 192.695 148.435 193.480 ;
        RECT 148.455 192.755 153.965 193.565 ;
        RECT 154.895 192.755 156.265 193.565 ;
      LAYER nwell ;
        RECT 70.520 189.535 156.460 192.365 ;
      LAYER pwell ;
        RECT 81.035 189.155 81.985 189.245 ;
        RECT 70.715 188.335 72.085 189.145 ;
        RECT 72.095 188.335 77.605 189.145 ;
        RECT 77.615 188.335 80.365 189.145 ;
        RECT 81.035 188.335 82.965 189.155 ;
        RECT 83.605 188.420 84.035 189.205 ;
        RECT 84.055 188.335 85.425 189.115 ;
        RECT 85.455 188.335 86.805 189.245 ;
        RECT 86.815 188.335 89.735 189.245 ;
        RECT 90.035 188.335 91.405 189.115 ;
        RECT 91.415 188.335 96.925 189.245 ;
        RECT 96.935 188.335 98.305 189.145 ;
        RECT 98.350 189.015 99.725 189.245 ;
        RECT 101.495 189.015 102.445 189.245 ;
        RECT 98.350 188.565 102.445 189.015 ;
        RECT 70.855 188.125 71.025 188.335 ;
        RECT 72.235 188.285 72.405 188.335 ;
        RECT 72.230 188.175 72.405 188.285 ;
        RECT 72.235 188.145 72.405 188.175 ;
        RECT 72.695 188.125 72.865 188.315 ;
        RECT 77.755 188.145 77.925 188.335 ;
        RECT 82.815 188.315 82.965 188.335 ;
        RECT 80.510 188.175 80.630 188.285 ;
        RECT 80.965 188.125 81.135 188.315 ;
        RECT 82.815 188.145 82.985 188.315 ;
        RECT 83.275 188.285 83.445 188.315 ;
        RECT 83.270 188.175 83.445 188.285 ;
        RECT 83.275 188.125 83.445 188.175 ;
        RECT 83.745 188.125 83.915 188.315 ;
        RECT 84.205 188.145 84.375 188.335 ;
        RECT 85.125 188.125 85.295 188.315 ;
        RECT 86.490 188.280 86.660 188.335 ;
        RECT 86.490 188.170 86.665 188.280 ;
        RECT 86.490 188.145 86.660 188.170 ;
        RECT 86.960 188.145 87.130 188.335 ;
        RECT 89.255 188.145 89.425 188.315 ;
        RECT 89.725 188.170 89.885 188.280 ;
        RECT 90.185 188.145 90.355 188.335 ;
        RECT 89.255 188.125 89.420 188.145 ;
        RECT 90.645 188.125 90.815 188.315 ;
        RECT 91.555 188.145 91.725 188.335 ;
        RECT 96.180 188.145 96.350 188.315 ;
        RECT 97.075 188.145 97.245 188.335 ;
        RECT 96.180 188.125 96.290 188.145 ;
        RECT 97.985 188.125 98.155 188.315 ;
        RECT 98.455 188.125 98.625 188.565 ;
        RECT 99.735 188.335 102.445 188.565 ;
        RECT 102.455 188.335 103.825 189.115 ;
        RECT 103.835 189.015 104.785 189.245 ;
        RECT 106.555 189.015 107.930 189.245 ;
        RECT 103.835 188.565 107.930 189.015 ;
        RECT 103.835 188.335 106.545 188.565 ;
        RECT 99.835 188.125 100.005 188.315 ;
        RECT 102.605 188.145 102.775 188.335 ;
        RECT 107.655 188.145 107.825 188.565 ;
        RECT 107.975 188.335 109.345 189.145 ;
        RECT 109.365 188.420 109.795 189.205 ;
        RECT 109.815 188.335 111.185 189.115 ;
        RECT 112.115 188.335 113.485 189.115 ;
        RECT 120.775 189.015 122.225 189.245 ;
        RECT 113.955 188.335 122.225 189.015 ;
        RECT 122.235 189.015 123.155 189.245 ;
        RECT 130.715 189.155 131.665 189.245 ;
        RECT 122.235 188.335 124.525 189.015 ;
        RECT 124.535 188.335 126.365 189.015 ;
        RECT 126.375 188.335 127.745 189.115 ;
        RECT 127.755 188.335 129.125 189.115 ;
        RECT 129.135 188.335 130.505 189.115 ;
        RECT 130.715 188.335 132.645 189.155 ;
        RECT 132.815 188.335 134.185 189.115 ;
        RECT 135.125 188.420 135.555 189.205 ;
        RECT 135.575 188.335 137.405 189.245 ;
        RECT 137.725 189.015 138.655 189.245 ;
        RECT 143.230 189.015 144.140 189.235 ;
        RECT 145.675 189.015 147.025 189.245 ;
        RECT 137.725 188.335 139.560 189.015 ;
        RECT 139.715 188.335 147.025 189.015 ;
        RECT 147.115 188.335 150.285 189.245 ;
        RECT 151.215 188.335 152.585 189.115 ;
        RECT 152.595 188.335 153.965 189.115 ;
        RECT 154.895 188.335 156.265 189.145 ;
        RECT 108.115 188.125 108.285 188.335 ;
        RECT 110.865 188.145 111.035 188.335 ;
        RECT 111.345 188.180 111.505 188.290 ;
        RECT 112.265 188.145 112.435 188.335 ;
        RECT 113.630 188.175 113.750 188.285 ;
        RECT 114.095 188.145 114.265 188.335 ;
        RECT 117.305 188.125 117.475 188.315 ;
        RECT 70.715 187.315 72.085 188.125 ;
        RECT 72.555 187.445 79.865 188.125 ;
        RECT 76.070 187.225 76.980 187.445 ;
        RECT 78.515 187.215 79.865 187.445 ;
        RECT 79.915 187.345 81.285 188.125 ;
        RECT 81.295 187.445 83.585 188.125 ;
        RECT 81.295 187.215 82.215 187.445 ;
        RECT 83.595 187.345 84.965 188.125 ;
        RECT 84.975 187.345 86.345 188.125 ;
        RECT 87.585 187.445 89.420 188.125 ;
        RECT 87.585 187.215 88.515 187.445 ;
        RECT 90.495 187.345 91.865 188.125 ;
        RECT 91.875 187.445 96.290 188.125 ;
        RECT 91.875 187.215 95.805 187.445 ;
        RECT 96.485 187.255 96.915 188.040 ;
        RECT 96.935 187.345 98.305 188.125 ;
        RECT 98.315 187.315 99.685 188.125 ;
        RECT 99.695 187.445 107.965 188.125 ;
        RECT 107.975 187.445 116.245 188.125 ;
        RECT 106.515 187.215 107.965 187.445 ;
        RECT 114.795 187.215 116.245 187.445 ;
        RECT 116.255 187.345 117.625 188.125 ;
        RECT 117.775 187.895 117.945 188.315 ;
        RECT 121.910 188.175 122.030 188.285 ;
        RECT 123.745 188.125 123.915 188.315 ;
        RECT 124.215 188.285 124.385 188.335 ;
        RECT 124.210 188.175 124.385 188.285 ;
        RECT 124.215 188.145 124.385 188.175 ;
        RECT 124.675 188.125 124.845 188.335 ;
        RECT 127.425 188.145 127.595 188.335 ;
        RECT 128.805 188.145 128.975 188.335 ;
        RECT 129.285 188.145 129.455 188.335 ;
        RECT 132.495 188.315 132.645 188.335 ;
        RECT 133.865 188.315 134.035 188.335 ;
        RECT 132.495 188.145 132.665 188.315 ;
        RECT 133.865 188.145 134.045 188.315 ;
        RECT 134.345 188.180 134.505 188.290 ;
        RECT 137.090 188.145 137.260 188.335 ;
        RECT 139.395 188.315 139.560 188.335 ;
        RECT 139.395 188.145 139.565 188.315 ;
        RECT 139.855 188.145 140.025 188.335 ;
        RECT 142.130 188.145 142.300 188.315 ;
        RECT 147.215 188.145 147.385 188.335 ;
        RECT 133.875 188.125 134.045 188.145 ;
        RECT 142.190 188.125 142.300 188.145 ;
        RECT 147.675 188.125 147.845 188.315 ;
        RECT 150.435 188.145 150.605 188.315 ;
        RECT 150.435 188.125 150.585 188.145 ;
        RECT 151.805 188.125 151.975 188.315 ;
        RECT 152.265 188.145 152.435 188.335 ;
        RECT 153.185 188.125 153.355 188.315 ;
        RECT 153.645 188.145 153.815 188.335 ;
        RECT 154.125 188.180 154.285 188.290 ;
        RECT 154.575 188.125 154.745 188.315 ;
        RECT 155.955 188.125 156.125 188.335 ;
        RECT 119.055 187.895 121.765 188.125 ;
        RECT 117.670 187.445 121.765 187.895 ;
        RECT 117.670 187.215 119.045 187.445 ;
        RECT 120.815 187.215 121.765 187.445 ;
        RECT 122.245 187.255 122.675 188.040 ;
        RECT 122.695 187.345 124.065 188.125 ;
        RECT 124.535 187.445 133.640 188.125 ;
        RECT 133.735 187.445 142.005 188.125 ;
        RECT 142.190 187.445 146.605 188.125 ;
        RECT 140.555 187.215 142.005 187.445 ;
        RECT 142.675 187.215 146.605 187.445 ;
        RECT 146.615 187.345 147.985 188.125 ;
        RECT 148.005 187.255 148.435 188.040 ;
        RECT 148.655 187.305 150.585 188.125 ;
        RECT 150.755 187.345 152.125 188.125 ;
        RECT 152.135 187.345 153.505 188.125 ;
        RECT 153.515 187.345 154.885 188.125 ;
        RECT 154.895 187.315 156.265 188.125 ;
        RECT 148.655 187.215 149.605 187.305 ;
      LAYER nwell ;
        RECT 70.520 184.095 156.460 186.925 ;
      LAYER pwell ;
        RECT 70.715 182.895 72.085 183.705 ;
        RECT 72.095 182.895 73.925 183.705 ;
        RECT 74.395 182.895 75.745 183.805 ;
        RECT 75.775 182.895 77.605 183.805 ;
        RECT 77.615 182.895 80.365 183.705 ;
        RECT 80.375 183.605 81.305 183.805 ;
        RECT 82.635 183.605 83.585 183.805 ;
        RECT 80.375 183.125 83.585 183.605 ;
        RECT 80.520 182.925 83.585 183.125 ;
        RECT 83.605 182.980 84.035 183.765 ;
        RECT 87.570 183.575 88.480 183.795 ;
        RECT 90.015 183.575 91.365 183.805 ;
        RECT 70.855 182.685 71.025 182.895 ;
        RECT 72.235 182.685 72.405 182.895 ;
        RECT 74.070 182.735 74.190 182.845 ;
        RECT 74.540 182.705 74.710 182.895 ;
        RECT 77.290 182.705 77.460 182.895 ;
        RECT 77.755 182.705 77.925 182.895 ;
        RECT 79.595 182.685 79.765 182.875 ;
        RECT 80.520 182.705 80.690 182.925 ;
        RECT 82.650 182.895 83.585 182.925 ;
        RECT 84.055 182.895 91.365 183.575 ;
        RECT 92.335 182.895 93.705 183.675 ;
        RECT 94.375 183.575 98.305 183.805 ;
        RECT 93.890 182.895 98.305 183.575 ;
        RECT 98.315 183.575 99.245 183.805 ;
        RECT 98.315 182.895 102.215 183.575 ;
        RECT 102.455 182.895 103.825 183.675 ;
        RECT 103.835 182.895 109.345 183.705 ;
        RECT 109.365 182.980 109.795 183.765 ;
        RECT 109.815 182.895 111.645 183.575 ;
        RECT 111.655 182.895 115.325 183.705 ;
        RECT 115.335 182.895 116.705 183.675 ;
        RECT 123.535 183.575 124.985 183.805 ;
        RECT 116.715 182.895 124.985 183.575 ;
        RECT 124.995 182.895 126.365 183.705 ;
        RECT 126.375 182.895 127.745 183.675 ;
        RECT 127.755 182.895 129.125 183.675 ;
        RECT 130.055 182.895 132.975 183.805 ;
        RECT 133.275 182.895 135.105 183.705 ;
        RECT 135.125 182.980 135.555 183.765 ;
        RECT 135.575 182.895 136.945 183.675 ;
        RECT 137.615 183.575 141.545 183.805 ;
        RECT 142.675 183.575 146.605 183.805 ;
        RECT 150.590 183.575 151.500 183.795 ;
        RECT 153.035 183.575 154.385 183.805 ;
        RECT 137.130 182.895 141.545 183.575 ;
        RECT 142.190 182.895 146.605 183.575 ;
        RECT 147.075 182.895 154.385 183.575 ;
        RECT 154.895 182.895 156.265 183.705 ;
        RECT 82.350 182.735 82.470 182.845 ;
        RECT 82.815 182.685 82.985 182.875 ;
        RECT 84.195 182.845 84.365 182.895 ;
        RECT 84.190 182.735 84.365 182.845 ;
        RECT 84.195 182.705 84.365 182.735 ;
        RECT 85.575 182.685 85.745 182.875 ;
        RECT 86.945 182.685 87.115 182.875 ;
        RECT 91.580 182.850 91.750 182.875 ;
        RECT 91.565 182.740 91.750 182.850 ;
        RECT 91.580 182.705 91.750 182.740 ;
        RECT 91.990 182.705 92.160 182.875 ;
        RECT 93.385 182.705 93.555 182.895 ;
        RECT 93.890 182.875 94.000 182.895 ;
        RECT 93.830 182.705 94.000 182.875 ;
        RECT 98.730 182.705 98.900 182.895 ;
        RECT 98.915 182.705 99.085 182.875 ;
        RECT 99.350 182.705 99.520 182.875 ;
        RECT 102.605 182.705 102.775 182.895 ;
        RECT 103.975 182.875 104.145 182.895 ;
        RECT 103.975 182.705 104.150 182.875 ;
        RECT 91.580 182.685 91.690 182.705 ;
        RECT 70.715 181.875 72.085 182.685 ;
        RECT 72.095 182.005 79.405 182.685 ;
        RECT 75.610 181.785 76.520 182.005 ;
        RECT 78.055 181.775 79.405 182.005 ;
        RECT 79.455 181.875 82.205 182.685 ;
        RECT 82.675 181.905 84.045 182.685 ;
        RECT 84.525 181.775 85.875 182.685 ;
        RECT 85.895 181.905 87.265 182.685 ;
        RECT 87.275 182.005 91.690 182.685 ;
        RECT 92.050 182.685 92.160 182.705 ;
        RECT 98.915 182.685 99.065 182.705 ;
        RECT 92.050 182.005 96.465 182.685 ;
        RECT 87.275 181.775 91.205 182.005 ;
        RECT 92.535 181.775 96.465 182.005 ;
        RECT 96.485 181.815 96.915 182.600 ;
        RECT 97.135 181.865 99.065 182.685 ;
        RECT 99.410 182.685 99.520 182.705 ;
        RECT 103.980 182.685 104.150 182.705 ;
        RECT 109.495 182.705 109.665 182.875 ;
        RECT 109.495 182.685 109.645 182.705 ;
        RECT 110.865 182.685 111.035 182.875 ;
        RECT 111.335 182.685 111.505 182.895 ;
        RECT 111.795 182.705 111.965 182.895 ;
        RECT 116.385 182.705 116.555 182.895 ;
        RECT 116.855 182.685 117.025 182.895 ;
        RECT 122.835 182.685 123.005 182.875 ;
        RECT 124.670 182.735 124.790 182.845 ;
        RECT 125.135 182.685 125.305 182.895 ;
        RECT 126.525 182.705 126.695 182.895 ;
        RECT 128.805 182.705 128.975 182.895 ;
        RECT 129.285 182.740 129.445 182.850 ;
        RECT 130.200 182.705 130.370 182.895 ;
        RECT 132.495 182.685 132.665 182.875 ;
        RECT 133.415 182.705 133.585 182.895 ;
        RECT 136.170 182.735 136.290 182.845 ;
        RECT 136.625 182.705 136.795 182.895 ;
        RECT 137.130 182.875 137.240 182.895 ;
        RECT 142.190 182.875 142.300 182.895 ;
        RECT 137.070 182.705 137.240 182.875 ;
        RECT 137.550 182.685 137.720 182.875 ;
        RECT 138.015 182.685 138.185 182.875 ;
        RECT 140.775 182.685 140.945 182.875 ;
        RECT 141.690 182.735 141.810 182.845 ;
        RECT 142.130 182.705 142.300 182.875 ;
        RECT 146.750 182.735 146.870 182.845 ;
        RECT 147.215 182.705 147.385 182.895 ;
        RECT 148.605 182.730 148.765 182.840 ;
        RECT 152.275 182.685 152.445 182.875 ;
        RECT 154.575 182.845 154.745 182.875 ;
        RECT 154.570 182.735 154.745 182.845 ;
        RECT 154.575 182.705 154.745 182.735 ;
        RECT 154.575 182.685 154.725 182.705 ;
        RECT 155.955 182.685 156.125 182.895 ;
        RECT 99.410 182.005 103.825 182.685 ;
        RECT 97.135 181.775 98.085 181.865 ;
        RECT 99.895 181.775 103.825 182.005 ;
        RECT 103.835 181.775 107.505 182.685 ;
        RECT 107.715 181.865 109.645 182.685 ;
        RECT 109.815 181.905 111.185 182.685 ;
        RECT 111.195 181.875 116.705 182.685 ;
        RECT 116.715 181.875 122.225 182.685 ;
        RECT 107.715 181.775 108.665 181.865 ;
        RECT 122.245 181.815 122.675 182.600 ;
        RECT 122.695 181.875 124.525 182.685 ;
        RECT 124.995 182.005 132.305 182.685 ;
        RECT 128.510 181.785 129.420 182.005 ;
        RECT 130.955 181.775 132.305 182.005 ;
        RECT 132.355 181.875 136.025 182.685 ;
        RECT 136.515 181.775 137.865 182.685 ;
        RECT 137.875 182.005 140.625 182.685 ;
        RECT 140.635 182.005 147.945 182.685 ;
        RECT 139.695 181.775 140.625 182.005 ;
        RECT 144.150 181.785 145.060 182.005 ;
        RECT 146.595 181.775 147.945 182.005 ;
        RECT 148.005 181.815 148.435 182.600 ;
        RECT 149.375 181.775 152.545 182.685 ;
        RECT 152.795 181.865 154.725 182.685 ;
        RECT 154.895 181.875 156.265 182.685 ;
        RECT 152.795 181.775 153.745 181.865 ;
      LAYER nwell ;
        RECT 70.520 178.655 156.460 181.485 ;
      LAYER pwell ;
        RECT 70.715 177.455 72.085 178.265 ;
        RECT 72.095 177.455 74.845 178.265 ;
        RECT 74.855 177.455 76.205 178.365 ;
        RECT 76.695 178.135 77.615 178.365 ;
        RECT 76.695 177.455 78.985 178.135 ;
        RECT 78.995 177.455 80.825 178.365 ;
        RECT 80.835 177.455 83.585 178.265 ;
        RECT 83.605 177.540 84.035 178.325 ;
        RECT 84.055 177.455 85.885 178.265 ;
        RECT 86.355 177.455 87.725 178.235 ;
        RECT 87.735 177.455 90.945 178.365 ;
        RECT 91.040 177.455 100.145 178.135 ;
        RECT 100.155 177.455 103.825 178.265 ;
        RECT 104.755 177.455 108.415 178.365 ;
        RECT 109.365 177.540 109.795 178.325 ;
        RECT 110.735 178.165 111.680 178.365 ;
        RECT 113.495 178.165 114.440 178.365 ;
        RECT 110.735 177.485 113.485 178.165 ;
        RECT 113.495 177.485 116.245 178.165 ;
        RECT 110.735 177.455 111.680 177.485 ;
        RECT 70.855 177.245 71.025 177.455 ;
        RECT 72.235 177.245 72.405 177.455 ;
        RECT 75.000 177.265 75.170 177.455 ;
        RECT 78.675 177.435 78.845 177.455 ;
        RECT 75.910 177.295 76.030 177.405 ;
        RECT 76.370 177.295 76.490 177.405 ;
        RECT 78.215 177.265 78.385 177.435 ;
        RECT 78.675 177.265 78.850 177.435 ;
        RECT 80.510 177.265 80.680 177.455 ;
        RECT 78.215 177.245 78.365 177.265 ;
        RECT 78.680 177.245 78.850 177.265 ;
        RECT 80.975 177.245 81.145 177.455 ;
        RECT 84.195 177.265 84.365 177.455 ;
        RECT 86.030 177.295 86.150 177.405 ;
        RECT 87.405 177.265 87.575 177.455 ;
        RECT 88.335 177.245 88.505 177.435 ;
        RECT 90.635 177.265 90.805 177.455 ;
        RECT 91.555 177.245 91.725 177.435 ;
        RECT 94.325 177.245 94.495 177.435 ;
        RECT 95.705 177.290 95.865 177.400 ;
        RECT 97.085 177.245 97.255 177.435 ;
        RECT 98.455 177.245 98.625 177.435 ;
        RECT 99.835 177.265 100.005 177.455 ;
        RECT 100.295 177.265 100.465 177.455 ;
        RECT 101.210 177.295 101.330 177.405 ;
        RECT 101.675 177.245 101.845 177.435 ;
        RECT 103.985 177.300 104.145 177.410 ;
        RECT 106.735 177.245 106.905 177.435 ;
        RECT 107.190 177.245 107.360 177.435 ;
        RECT 108.120 177.265 108.290 177.455 ;
        RECT 108.575 177.245 108.745 177.435 ;
        RECT 109.965 177.300 110.125 177.410 ;
        RECT 113.170 177.265 113.340 177.485 ;
        RECT 113.495 177.455 114.440 177.485 ;
        RECT 115.930 177.435 116.100 177.485 ;
        RECT 116.265 177.455 118.995 178.365 ;
        RECT 119.165 177.455 124.985 178.365 ;
        RECT 124.995 177.455 126.365 178.235 ;
        RECT 126.395 177.455 127.745 178.365 ;
        RECT 127.755 177.455 129.585 178.365 ;
        RECT 130.515 177.455 131.885 178.235 ;
        RECT 131.895 178.135 132.815 178.365 ;
        RECT 131.895 177.455 134.185 178.135 ;
        RECT 135.125 177.540 135.555 178.325 ;
        RECT 135.575 178.165 136.505 178.365 ;
        RECT 137.835 178.165 138.785 178.365 ;
        RECT 135.575 177.685 138.785 178.165 ;
        RECT 135.720 177.485 138.785 177.685 ;
        RECT 70.715 176.435 72.085 177.245 ;
        RECT 72.095 176.435 75.765 177.245 ;
        RECT 76.435 176.425 78.365 177.245 ;
        RECT 76.435 176.335 77.385 176.425 ;
        RECT 78.535 176.335 80.365 177.245 ;
        RECT 80.835 176.565 88.145 177.245 ;
        RECT 88.195 176.565 91.405 177.245 ;
        RECT 91.555 177.015 94.165 177.245 ;
        RECT 84.350 176.345 85.260 176.565 ;
        RECT 86.795 176.335 88.145 176.565 ;
        RECT 90.270 176.335 91.405 176.565 ;
        RECT 91.415 176.335 94.165 177.015 ;
        RECT 94.175 176.465 95.545 177.245 ;
        RECT 96.485 176.375 96.915 177.160 ;
        RECT 96.935 176.465 98.305 177.245 ;
        RECT 98.315 176.435 101.065 177.245 ;
        RECT 101.545 176.335 102.895 177.245 ;
        RECT 102.985 176.335 107.045 177.245 ;
        RECT 107.075 176.335 108.425 177.245 ;
        RECT 108.435 176.435 111.185 177.245 ;
        RECT 111.195 177.215 112.140 177.245 ;
        RECT 113.630 177.215 113.800 177.435 ;
        RECT 115.930 177.265 116.110 177.435 ;
        RECT 113.955 177.215 114.910 177.245 ;
        RECT 115.940 177.215 116.110 177.265 ;
        RECT 116.395 177.245 116.565 177.455 ;
        RECT 121.915 177.265 122.085 177.435 ;
        RECT 121.915 177.245 122.065 177.265 ;
        RECT 122.835 177.245 123.005 177.435 ;
        RECT 124.215 177.245 124.385 177.435 ;
        RECT 124.675 177.265 124.845 177.455 ;
        RECT 126.045 177.265 126.215 177.455 ;
        RECT 127.430 177.265 127.600 177.455 ;
        RECT 129.270 177.265 129.440 177.455 ;
        RECT 129.745 177.300 129.905 177.410 ;
        RECT 130.195 177.245 130.365 177.435 ;
        RECT 131.565 177.265 131.735 177.455 ;
        RECT 133.875 177.265 134.045 177.455 ;
        RECT 134.345 177.300 134.505 177.410 ;
        RECT 135.720 177.265 135.890 177.485 ;
        RECT 137.850 177.455 138.785 177.485 ;
        RECT 138.795 178.135 139.715 178.365 ;
        RECT 142.145 178.135 143.075 178.365 ;
        RECT 147.830 178.135 148.740 178.355 ;
        RECT 150.275 178.135 151.625 178.365 ;
        RECT 138.795 177.455 141.085 178.135 ;
        RECT 141.240 177.455 143.075 178.135 ;
        RECT 144.315 177.455 151.625 178.135 ;
        RECT 151.675 177.455 154.425 178.265 ;
        RECT 154.895 177.455 156.265 178.265 ;
        RECT 139.395 177.245 139.565 177.435 ;
        RECT 140.775 177.265 140.945 177.455 ;
        RECT 141.240 177.435 141.405 177.455 ;
        RECT 141.235 177.405 141.405 177.435 ;
        RECT 141.230 177.295 141.405 177.405 ;
        RECT 143.545 177.300 143.705 177.410 ;
        RECT 141.235 177.265 141.405 177.295 ;
        RECT 144.455 177.265 144.625 177.455 ;
        RECT 145.860 177.265 146.030 177.435 ;
        RECT 145.860 177.245 145.970 177.265 ;
        RECT 147.670 177.245 147.840 177.435 ;
        RECT 149.515 177.245 149.685 177.435 ;
        RECT 149.970 177.295 150.090 177.405 ;
        RECT 151.815 177.265 151.985 177.455 ;
        RECT 152.735 177.245 152.905 177.435 ;
        RECT 153.195 177.245 153.365 177.435 ;
        RECT 154.570 177.295 154.690 177.405 ;
        RECT 155.955 177.245 156.125 177.455 ;
        RECT 111.195 176.535 113.945 177.215 ;
        RECT 113.955 176.535 116.235 177.215 ;
        RECT 111.195 176.335 112.140 176.535 ;
        RECT 113.955 176.335 114.910 176.535 ;
        RECT 116.255 176.435 119.925 177.245 ;
        RECT 120.135 176.425 122.065 177.245 ;
        RECT 120.135 176.335 121.085 176.425 ;
        RECT 122.245 176.375 122.675 177.160 ;
        RECT 122.695 176.435 124.065 177.245 ;
        RECT 124.075 176.335 129.915 177.245 ;
        RECT 130.055 176.565 139.160 177.245 ;
        RECT 139.255 176.435 141.085 177.245 ;
        RECT 141.555 176.565 145.970 177.245 ;
        RECT 141.555 176.335 145.485 176.565 ;
        RECT 146.155 176.335 147.985 177.245 ;
        RECT 148.005 176.375 148.435 177.160 ;
        RECT 148.455 176.465 149.825 177.245 ;
        RECT 150.305 176.335 153.035 177.245 ;
        RECT 153.055 176.435 154.885 177.245 ;
        RECT 154.895 176.435 156.265 177.245 ;
      LAYER nwell ;
        RECT 70.520 173.215 156.460 176.045 ;
      LAYER pwell ;
        RECT 70.715 172.015 72.085 172.825 ;
        RECT 72.095 172.015 74.845 172.825 ;
        RECT 75.315 172.015 76.665 172.925 ;
        RECT 76.695 172.015 82.205 172.825 ;
        RECT 82.215 172.015 83.585 172.825 ;
        RECT 83.605 172.100 84.035 172.885 ;
        RECT 84.055 172.015 85.425 172.825 ;
        RECT 85.435 172.695 89.365 172.925 ;
        RECT 90.495 172.725 91.445 172.925 ;
        RECT 85.435 172.015 89.850 172.695 ;
        RECT 90.495 172.045 94.165 172.725 ;
        RECT 97.170 172.695 98.305 172.925 ;
        RECT 90.495 172.015 91.445 172.045 ;
        RECT 70.855 171.805 71.025 172.015 ;
        RECT 72.235 171.805 72.405 172.015 ;
        RECT 74.990 171.855 75.110 171.965 ;
        RECT 75.460 171.825 75.630 172.015 ;
        RECT 76.835 171.825 77.005 172.015 ;
        RECT 79.595 171.805 79.765 171.995 ;
        RECT 82.355 171.825 82.525 172.015 ;
        RECT 84.195 171.825 84.365 172.015 ;
        RECT 89.740 171.995 89.850 172.015 ;
        RECT 86.960 171.805 87.130 171.995 ;
        RECT 89.740 171.825 89.910 171.995 ;
        RECT 90.170 171.855 90.290 171.965 ;
        RECT 70.715 170.995 72.085 171.805 ;
        RECT 72.095 171.125 79.405 171.805 ;
        RECT 79.455 171.125 86.765 171.805 ;
        RECT 75.610 170.905 76.520 171.125 ;
        RECT 78.055 170.895 79.405 171.125 ;
        RECT 82.970 170.905 83.880 171.125 ;
        RECT 85.415 170.895 86.765 171.125 ;
        RECT 86.815 170.895 90.485 171.805 ;
        RECT 90.630 171.775 90.800 171.995 ;
        RECT 92.930 171.855 93.050 171.965 ;
        RECT 93.395 171.805 93.565 171.995 ;
        RECT 93.850 171.825 94.020 172.045 ;
        RECT 95.095 172.015 98.305 172.695 ;
        RECT 98.315 172.015 101.985 172.925 ;
        RECT 102.915 172.015 106.125 172.925 ;
        RECT 106.135 172.015 107.505 172.795 ;
        RECT 107.515 172.015 109.345 172.825 ;
        RECT 109.365 172.100 109.795 172.885 ;
        RECT 131.175 172.835 132.125 172.925 ;
        RECT 110.360 172.015 119.465 172.695 ;
        RECT 119.475 172.015 124.985 172.825 ;
        RECT 124.995 172.015 130.505 172.825 ;
        RECT 131.175 172.015 133.105 172.835 ;
        RECT 133.275 172.015 134.625 172.925 ;
        RECT 135.125 172.100 135.555 172.885 ;
        RECT 135.775 172.835 136.725 172.925 ;
        RECT 135.775 172.015 137.705 172.835 ;
        RECT 137.875 172.015 139.705 172.825 ;
        RECT 139.715 172.725 140.645 172.925 ;
        RECT 141.975 172.725 142.925 172.925 ;
        RECT 139.715 172.245 142.925 172.725 ;
        RECT 143.985 172.695 144.915 172.925 ;
        RECT 139.860 172.045 142.925 172.245 ;
        RECT 94.325 171.860 94.485 171.970 ;
        RECT 95.235 171.825 95.405 172.015 ;
        RECT 97.075 171.805 97.245 171.995 ;
        RECT 98.460 171.825 98.630 172.015 ;
        RECT 99.375 171.805 99.545 171.995 ;
        RECT 102.145 171.860 102.305 171.970 ;
        RECT 104.435 171.825 104.605 171.995 ;
        RECT 104.435 171.805 104.600 171.825 ;
        RECT 104.890 171.805 105.060 171.995 ;
        RECT 105.815 171.825 105.985 172.015 ;
        RECT 106.285 171.995 106.455 172.015 ;
        RECT 106.275 171.825 106.455 171.995 ;
        RECT 107.655 171.995 107.825 172.015 ;
        RECT 107.655 171.825 107.830 171.995 ;
        RECT 109.950 171.855 110.070 171.965 ;
        RECT 111.330 171.855 111.450 171.965 ;
        RECT 106.275 171.805 106.445 171.825 ;
        RECT 107.660 171.805 107.830 171.825 ;
        RECT 91.830 171.775 92.785 171.805 ;
        RECT 90.505 171.095 92.785 171.775 ;
        RECT 93.255 171.125 96.465 171.805 ;
        RECT 91.830 170.895 92.785 171.095 ;
        RECT 95.330 170.895 96.465 171.125 ;
        RECT 96.485 170.935 96.915 171.720 ;
        RECT 96.935 171.125 99.225 171.805 ;
        RECT 98.305 170.895 99.225 171.125 ;
        RECT 99.335 170.895 102.445 171.805 ;
        RECT 102.765 171.125 104.600 171.805 ;
        RECT 102.765 170.895 103.695 171.125 ;
        RECT 104.775 170.895 106.125 171.805 ;
        RECT 106.135 170.995 107.505 171.805 ;
        RECT 107.515 170.895 111.185 171.805 ;
        RECT 111.655 171.775 112.600 171.805 ;
        RECT 114.090 171.775 114.260 171.995 ;
        RECT 115.465 171.805 115.635 171.995 ;
        RECT 116.855 171.805 117.025 171.995 ;
        RECT 117.325 171.850 117.485 171.960 ;
        RECT 118.235 171.805 118.405 171.995 ;
        RECT 119.155 171.825 119.325 172.015 ;
        RECT 119.615 171.825 119.785 172.015 ;
        RECT 120.070 171.855 120.190 171.965 ;
        RECT 120.530 171.805 120.700 171.995 ;
        RECT 121.910 171.855 122.030 171.965 ;
        RECT 122.835 171.805 123.005 171.995 ;
        RECT 125.135 171.825 125.305 172.015 ;
        RECT 132.955 171.995 133.105 172.015 ;
        RECT 130.650 171.855 130.770 171.965 ;
        RECT 131.105 171.805 131.275 171.995 ;
        RECT 132.485 171.805 132.655 171.995 ;
        RECT 132.955 171.805 133.125 171.995 ;
        RECT 133.420 171.825 133.590 172.015 ;
        RECT 137.555 171.995 137.705 172.015 ;
        RECT 134.790 171.855 134.910 171.965 ;
        RECT 135.265 171.805 135.435 171.995 ;
        RECT 136.635 171.805 136.805 171.995 ;
        RECT 137.555 171.825 137.725 171.995 ;
        RECT 138.015 171.825 138.185 172.015 ;
        RECT 139.860 171.825 140.030 172.045 ;
        RECT 141.990 172.015 142.925 172.045 ;
        RECT 143.080 172.015 144.915 172.695 ;
        RECT 145.235 172.015 146.605 172.795 ;
        RECT 146.615 172.015 149.365 172.825 ;
        RECT 149.475 172.015 152.585 172.925 ;
        RECT 152.595 172.015 154.425 172.825 ;
        RECT 154.895 172.015 156.265 172.825 ;
        RECT 143.080 171.995 143.245 172.015 ;
        RECT 138.035 171.805 138.185 171.825 ;
        RECT 140.315 171.805 140.485 171.995 ;
        RECT 143.075 171.825 143.245 171.995 ;
        RECT 144.915 171.805 145.085 171.995 ;
        RECT 145.375 171.805 145.545 171.995 ;
        RECT 146.285 171.825 146.455 172.015 ;
        RECT 146.755 171.825 146.925 172.015 ;
        RECT 148.595 171.805 148.765 171.995 ;
        RECT 149.515 171.825 149.685 172.015 ;
        RECT 152.735 171.995 152.905 172.015 ;
        RECT 152.730 171.825 152.905 171.995 ;
        RECT 152.730 171.805 152.900 171.825 ;
        RECT 153.195 171.805 153.365 171.995 ;
        RECT 154.570 171.855 154.690 171.965 ;
        RECT 155.955 171.805 156.125 172.015 ;
        RECT 111.655 171.095 114.405 171.775 ;
        RECT 111.655 170.895 112.600 171.095 ;
        RECT 114.415 171.025 115.785 171.805 ;
        RECT 115.805 170.895 117.155 171.805 ;
        RECT 118.110 170.895 119.925 171.805 ;
        RECT 120.415 170.895 121.765 171.805 ;
        RECT 122.245 170.935 122.675 171.720 ;
        RECT 122.695 171.125 130.005 171.805 ;
        RECT 126.210 170.905 127.120 171.125 ;
        RECT 128.655 170.895 130.005 171.125 ;
        RECT 130.055 171.025 131.425 171.805 ;
        RECT 131.435 171.025 132.805 171.805 ;
        RECT 132.815 170.995 134.645 171.805 ;
        RECT 135.115 171.025 136.485 171.805 ;
        RECT 136.495 170.995 137.865 171.805 ;
        RECT 138.035 170.985 139.965 171.805 ;
        RECT 140.175 170.995 143.845 171.805 ;
        RECT 139.015 170.895 139.965 170.985 ;
        RECT 143.865 170.895 145.215 171.805 ;
        RECT 145.245 170.895 147.975 171.805 ;
        RECT 148.005 170.935 148.435 171.720 ;
        RECT 148.555 170.895 151.665 171.805 ;
        RECT 151.695 170.895 153.045 171.805 ;
        RECT 153.065 170.895 154.415 171.805 ;
        RECT 154.895 170.995 156.265 171.805 ;
      LAYER nwell ;
        RECT 70.520 167.775 156.460 170.605 ;
      LAYER pwell ;
        RECT 70.715 166.575 72.085 167.385 ;
        RECT 75.610 167.255 76.520 167.475 ;
        RECT 78.055 167.255 79.405 167.485 ;
        RECT 72.095 166.575 79.405 167.255 ;
        RECT 79.455 166.575 80.825 167.355 ;
        RECT 80.845 166.575 82.195 167.485 ;
        RECT 82.215 166.575 83.585 167.385 ;
        RECT 83.605 166.660 84.035 167.445 ;
        RECT 84.055 166.575 86.805 167.385 ;
        RECT 86.815 166.575 88.185 167.355 ;
        RECT 88.215 166.575 89.565 167.485 ;
        RECT 90.120 166.575 99.225 167.255 ;
        RECT 99.235 166.575 102.905 167.485 ;
        RECT 102.915 166.575 108.425 167.385 ;
        RECT 109.365 166.660 109.795 167.445 ;
        RECT 109.815 166.575 113.485 167.385 ;
        RECT 113.495 166.575 114.865 167.355 ;
        RECT 114.875 166.575 116.705 167.385 ;
        RECT 116.715 166.575 120.385 167.485 ;
        RECT 123.910 167.255 124.820 167.475 ;
        RECT 126.355 167.255 128.125 167.485 ;
        RECT 120.395 166.575 128.125 167.255 ;
        RECT 128.215 167.285 129.160 167.485 ;
        RECT 128.215 166.605 130.965 167.285 ;
        RECT 128.215 166.575 129.160 166.605 ;
        RECT 70.855 166.365 71.025 166.575 ;
        RECT 72.235 166.365 72.405 166.575 ;
        RECT 75.925 166.410 76.085 166.520 ;
        RECT 76.835 166.365 77.005 166.555 ;
        RECT 79.605 166.385 79.775 166.575 ;
        RECT 80.975 166.385 81.145 166.575 ;
        RECT 82.355 166.385 82.525 166.575 ;
        RECT 84.195 166.385 84.365 166.575 ;
        RECT 86.965 166.385 87.135 166.575 ;
        RECT 89.250 166.385 89.420 166.575 ;
        RECT 89.710 166.415 89.830 166.525 ;
        RECT 91.095 166.365 91.265 166.555 ;
        RECT 91.530 166.385 91.700 166.555 ;
        RECT 96.150 166.415 96.270 166.525 ;
        RECT 97.070 166.415 97.190 166.525 ;
        RECT 91.590 166.365 91.700 166.385 ;
        RECT 98.450 166.365 98.620 166.555 ;
        RECT 98.915 166.385 99.085 166.575 ;
        RECT 99.380 166.385 99.550 166.575 ;
        RECT 100.755 166.385 100.925 166.555 ;
        RECT 100.755 166.365 100.920 166.385 ;
        RECT 101.220 166.365 101.390 166.555 ;
        RECT 103.055 166.385 103.225 166.575 ;
        RECT 104.895 166.365 105.065 166.555 ;
        RECT 106.275 166.365 106.445 166.555 ;
        RECT 108.090 166.385 108.260 166.555 ;
        RECT 108.585 166.420 108.745 166.530 ;
        RECT 109.955 166.385 110.125 166.575 ;
        RECT 108.150 166.365 108.260 166.385 ;
        RECT 112.720 166.365 112.890 166.555 ;
        RECT 113.645 166.385 113.815 166.575 ;
        RECT 115.015 166.385 115.185 166.575 ;
        RECT 116.395 166.365 116.565 166.555 ;
        RECT 118.230 166.415 118.350 166.525 ;
        RECT 118.695 166.365 118.865 166.555 ;
        RECT 120.070 166.385 120.240 166.575 ;
        RECT 120.535 166.385 120.705 166.575 ;
        RECT 121.910 166.415 122.030 166.525 ;
        RECT 124.675 166.385 124.845 166.555 ;
        RECT 124.675 166.365 124.840 166.385 ;
        RECT 126.975 166.365 127.145 166.555 ;
        RECT 127.435 166.365 127.605 166.555 ;
        RECT 129.270 166.415 129.390 166.525 ;
        RECT 130.650 166.365 130.820 166.605 ;
        RECT 130.975 166.575 132.345 167.355 ;
        RECT 132.355 166.575 133.725 167.385 ;
        RECT 133.735 166.575 135.105 167.355 ;
        RECT 135.125 166.660 135.555 167.445 ;
        RECT 136.625 167.255 137.555 167.485 ;
        RECT 135.720 166.575 137.555 167.255 ;
        RECT 138.530 166.575 142.005 167.485 ;
        RECT 145.530 167.255 146.440 167.475 ;
        RECT 147.975 167.255 149.325 167.485 ;
        RECT 150.955 167.255 154.885 167.485 ;
        RECT 142.015 166.575 149.325 167.255 ;
        RECT 150.470 166.575 154.885 167.255 ;
        RECT 154.895 166.575 156.265 167.385 ;
        RECT 131.125 166.555 131.295 166.575 ;
        RECT 132.495 166.555 132.665 166.575 ;
        RECT 131.115 166.385 131.295 166.555 ;
        RECT 132.470 166.385 132.665 166.555 ;
        RECT 134.785 166.385 134.955 166.575 ;
        RECT 135.720 166.555 135.885 166.575 ;
        RECT 141.690 166.555 141.860 166.575 ;
        RECT 135.715 166.385 135.885 166.555 ;
        RECT 137.070 166.385 137.240 166.555 ;
        RECT 138.010 166.415 138.130 166.525 ;
        RECT 141.690 166.385 141.875 166.555 ;
        RECT 142.155 166.385 142.325 166.575 ;
        RECT 150.470 166.555 150.580 166.575 ;
        RECT 131.115 166.365 131.285 166.385 ;
        RECT 132.530 166.365 132.640 166.385 ;
        RECT 137.130 166.365 137.240 166.385 ;
        RECT 141.705 166.365 141.875 166.385 ;
        RECT 143.995 166.365 144.165 166.555 ;
        RECT 144.455 166.365 144.625 166.555 ;
        RECT 146.290 166.415 146.410 166.525 ;
        RECT 147.675 166.365 147.845 166.555 ;
        RECT 149.525 166.420 149.685 166.530 ;
        RECT 150.410 166.385 150.580 166.555 ;
        RECT 152.760 166.385 152.930 166.555 ;
        RECT 152.760 166.365 152.870 166.385 ;
        RECT 153.205 166.365 153.375 166.555 ;
        RECT 154.570 166.415 154.690 166.525 ;
        RECT 155.955 166.365 156.125 166.575 ;
        RECT 70.715 165.555 72.085 166.365 ;
        RECT 72.095 165.555 75.765 166.365 ;
        RECT 76.695 165.685 84.005 166.365 ;
        RECT 80.210 165.465 81.120 165.685 ;
        RECT 82.655 165.455 84.005 165.685 ;
        RECT 84.095 165.685 91.405 166.365 ;
        RECT 91.590 165.685 96.005 166.365 ;
        RECT 84.095 165.455 85.445 165.685 ;
        RECT 86.980 165.465 87.890 165.685 ;
        RECT 92.075 165.455 96.005 165.685 ;
        RECT 96.485 165.495 96.915 166.280 ;
        RECT 97.415 165.455 98.765 166.365 ;
        RECT 99.085 165.685 100.920 166.365 ;
        RECT 99.085 165.455 100.015 165.685 ;
        RECT 101.075 165.455 104.745 166.365 ;
        RECT 104.765 165.455 106.115 166.365 ;
        RECT 106.135 165.555 107.965 166.365 ;
        RECT 108.150 165.685 112.565 166.365 ;
        RECT 108.635 165.455 112.565 165.685 ;
        RECT 112.575 165.455 116.050 166.365 ;
        RECT 116.255 165.555 118.085 166.365 ;
        RECT 118.555 165.455 121.765 166.365 ;
        RECT 122.245 165.495 122.675 166.280 ;
        RECT 123.005 165.685 124.840 166.365 ;
        RECT 124.995 165.685 127.285 166.365 ;
        RECT 123.005 165.455 123.935 165.685 ;
        RECT 124.995 165.455 125.915 165.685 ;
        RECT 127.295 165.555 129.125 166.365 ;
        RECT 129.615 165.455 130.965 166.365 ;
        RECT 130.975 165.555 132.345 166.365 ;
        RECT 132.530 165.685 136.945 166.365 ;
        RECT 137.130 165.685 141.545 166.365 ;
        RECT 133.015 165.455 136.945 165.685 ;
        RECT 137.615 165.455 141.545 165.685 ;
        RECT 141.555 165.585 142.925 166.365 ;
        RECT 142.945 165.455 144.295 166.365 ;
        RECT 144.315 165.555 146.145 166.365 ;
        RECT 146.625 165.455 147.975 166.365 ;
        RECT 148.005 165.495 148.435 166.280 ;
        RECT 148.455 165.685 152.870 166.365 ;
        RECT 148.455 165.455 152.385 165.685 ;
        RECT 153.055 165.585 154.425 166.365 ;
        RECT 154.895 165.555 156.265 166.365 ;
      LAYER nwell ;
        RECT 70.520 162.335 156.460 165.165 ;
      LAYER pwell ;
        RECT 70.715 161.135 72.085 161.945 ;
        RECT 72.135 161.815 73.485 162.045 ;
        RECT 75.020 161.815 75.930 162.035 ;
        RECT 72.135 161.135 79.445 161.815 ;
        RECT 79.455 161.135 83.125 161.945 ;
        RECT 83.605 161.220 84.035 162.005 ;
        RECT 84.055 161.135 86.805 161.945 ;
        RECT 86.965 161.135 92.785 162.045 ;
        RECT 92.830 161.815 94.205 162.045 ;
        RECT 95.975 161.815 96.925 162.045 ;
        RECT 92.830 161.365 96.925 161.815 ;
        RECT 70.855 160.925 71.025 161.135 ;
        RECT 72.235 160.925 72.405 161.115 ;
        RECT 75.920 160.925 76.090 161.115 ;
        RECT 77.755 160.925 77.925 161.115 ;
        RECT 79.135 160.945 79.305 161.135 ;
        RECT 79.595 160.945 79.765 161.135 ;
        RECT 82.815 160.945 82.985 161.115 ;
        RECT 83.285 161.085 83.455 161.115 ;
        RECT 83.270 160.975 83.455 161.085 ;
        RECT 82.815 160.925 82.980 160.945 ;
        RECT 83.285 160.925 83.455 160.975 ;
        RECT 84.195 160.945 84.365 161.135 ;
        RECT 84.655 160.925 84.825 161.115 ;
        RECT 88.345 160.925 88.515 161.115 ;
        RECT 89.725 160.925 89.895 161.115 ;
        RECT 70.715 160.115 72.085 160.925 ;
        RECT 72.095 160.115 75.765 160.925 ;
        RECT 75.775 160.015 77.605 160.925 ;
        RECT 77.715 160.015 80.825 160.925 ;
        RECT 81.145 160.245 82.980 160.925 ;
        RECT 81.145 160.015 82.075 160.245 ;
        RECT 83.135 160.145 84.505 160.925 ;
        RECT 84.515 160.115 88.185 160.925 ;
        RECT 88.195 160.145 89.565 160.925 ;
        RECT 89.575 160.145 90.945 160.925 ;
        RECT 91.100 160.895 91.270 161.115 ;
        RECT 92.475 160.945 92.645 161.135 ;
        RECT 92.935 160.945 93.105 161.365 ;
        RECT 94.215 161.135 96.925 161.365 ;
        RECT 96.935 161.135 100.145 162.045 ;
        RECT 100.155 161.815 101.085 162.045 ;
        RECT 100.155 161.135 102.905 161.815 ;
        RECT 102.925 161.135 104.275 162.045 ;
        RECT 104.295 161.135 105.645 162.045 ;
        RECT 106.145 161.135 108.875 162.045 ;
        RECT 109.365 161.220 109.795 162.005 ;
        RECT 110.935 161.815 114.865 162.045 ;
        RECT 110.450 161.135 114.865 161.815 ;
        RECT 114.875 161.135 116.225 162.045 ;
        RECT 116.715 161.135 120.385 162.045 ;
        RECT 120.395 161.135 123.145 161.945 ;
        RECT 123.465 161.815 124.395 162.045 ;
        RECT 123.465 161.135 125.300 161.815 ;
        RECT 125.455 161.135 126.825 161.915 ;
        RECT 126.835 161.135 132.345 161.945 ;
        RECT 132.355 161.135 135.105 161.945 ;
        RECT 135.125 161.220 135.555 162.005 ;
        RECT 135.725 161.135 139.380 162.045 ;
        RECT 139.715 161.135 145.225 161.945 ;
        RECT 145.235 161.135 147.065 161.945 ;
        RECT 151.050 161.815 151.960 162.035 ;
        RECT 153.495 161.815 154.845 162.045 ;
        RECT 147.535 161.135 154.845 161.815 ;
        RECT 154.895 161.135 156.265 161.945 ;
        RECT 94.785 160.925 94.955 161.115 ;
        RECT 97.075 161.085 97.245 161.135 ;
        RECT 96.150 160.975 96.270 161.085 ;
        RECT 97.070 160.975 97.245 161.085 ;
        RECT 97.075 160.945 97.245 160.975 ;
        RECT 97.535 160.925 97.705 161.115 ;
        RECT 99.835 160.925 100.005 161.115 ;
        RECT 102.135 160.925 102.305 161.115 ;
        RECT 102.595 160.945 102.765 161.135 ;
        RECT 103.055 160.945 103.225 161.135 ;
        RECT 104.440 160.945 104.610 161.135 ;
        RECT 105.810 160.975 105.930 161.085 ;
        RECT 106.275 160.945 106.445 161.135 ;
        RECT 110.450 161.115 110.560 161.135 ;
        RECT 115.940 161.115 116.110 161.135 ;
        RECT 109.980 161.085 110.150 161.115 ;
        RECT 109.030 160.975 109.150 161.085 ;
        RECT 109.950 160.975 110.150 161.085 ;
        RECT 109.980 160.945 110.150 160.975 ;
        RECT 110.390 160.945 110.585 161.115 ;
        RECT 109.980 160.925 110.090 160.945 ;
        RECT 110.415 160.925 110.585 160.945 ;
        RECT 115.935 160.945 116.110 161.115 ;
        RECT 116.390 160.975 116.510 161.085 ;
        RECT 116.860 160.945 117.030 161.135 ;
        RECT 115.935 160.925 116.105 160.945 ;
        RECT 119.610 160.925 119.780 161.115 ;
        RECT 120.535 160.945 120.705 161.135 ;
        RECT 125.135 161.115 125.300 161.135 ;
        RECT 121.905 160.925 122.075 161.115 ;
        RECT 122.845 160.970 123.005 161.080 ;
        RECT 125.135 160.945 125.305 161.115 ;
        RECT 126.055 160.925 126.225 161.115 ;
        RECT 126.505 160.945 126.675 161.135 ;
        RECT 126.975 160.945 127.145 161.135 ;
        RECT 130.195 160.945 130.365 161.115 ;
        RECT 130.195 160.925 130.355 160.945 ;
        RECT 130.665 160.925 130.835 161.115 ;
        RECT 132.035 160.925 132.205 161.115 ;
        RECT 132.495 160.945 132.665 161.135 ;
        RECT 135.725 161.115 135.885 161.135 ;
        RECT 134.790 160.975 134.910 161.085 ;
        RECT 135.255 160.945 135.425 161.115 ;
        RECT 135.715 160.945 135.885 161.115 ;
        RECT 139.395 160.945 139.565 161.115 ;
        RECT 139.855 160.945 140.025 161.135 ;
        RECT 143.530 160.975 143.650 161.085 ;
        RECT 135.265 160.925 135.425 160.945 ;
        RECT 139.405 160.925 139.565 160.945 ;
        RECT 144.920 160.925 145.090 161.115 ;
        RECT 145.375 160.945 145.545 161.135 ;
        RECT 147.675 161.085 147.845 161.135 ;
        RECT 147.210 160.975 147.330 161.085 ;
        RECT 147.670 160.975 147.845 161.085 ;
        RECT 147.675 160.945 147.845 160.975 ;
        RECT 145.380 160.925 145.545 160.945 ;
        RECT 148.595 160.925 148.765 161.115 ;
        RECT 151.815 160.925 151.985 161.115 ;
        RECT 152.275 160.925 152.445 161.115 ;
        RECT 155.955 160.925 156.125 161.135 ;
        RECT 93.675 160.895 94.625 160.925 ;
        RECT 90.955 160.215 94.625 160.895 ;
        RECT 93.675 160.015 94.625 160.215 ;
        RECT 94.635 160.145 96.005 160.925 ;
        RECT 96.485 160.055 96.915 160.840 ;
        RECT 97.395 160.245 99.685 160.925 ;
        RECT 99.695 160.245 101.985 160.925 ;
        RECT 98.765 160.015 99.685 160.245 ;
        RECT 101.065 160.015 101.985 160.245 ;
        RECT 101.995 160.115 105.665 160.925 ;
        RECT 105.675 160.245 110.090 160.925 ;
        RECT 105.675 160.015 109.605 160.245 ;
        RECT 110.275 160.115 115.785 160.925 ;
        RECT 115.795 160.115 119.465 160.925 ;
        RECT 119.495 160.015 120.845 160.925 ;
        RECT 120.855 160.145 122.225 160.925 ;
        RECT 122.245 160.055 122.675 160.840 ;
        RECT 123.615 160.015 126.365 160.925 ;
        RECT 126.700 160.015 130.355 160.925 ;
        RECT 130.515 160.145 131.885 160.925 ;
        RECT 131.895 160.115 134.645 160.925 ;
        RECT 135.265 160.015 138.920 160.925 ;
        RECT 139.405 160.015 143.060 160.925 ;
        RECT 143.855 160.015 145.205 160.925 ;
        RECT 145.380 160.245 147.215 160.925 ;
        RECT 146.285 160.015 147.215 160.245 ;
        RECT 148.005 160.055 148.435 160.840 ;
        RECT 148.455 160.245 150.745 160.925 ;
        RECT 149.825 160.015 150.745 160.245 ;
        RECT 150.755 160.145 152.125 160.925 ;
        RECT 152.135 160.115 154.885 160.925 ;
        RECT 154.895 160.115 156.265 160.925 ;
      LAYER nwell ;
        RECT 70.520 156.895 156.460 159.725 ;
      LAYER pwell ;
        RECT 70.715 155.695 72.085 156.505 ;
        RECT 72.095 155.695 77.605 156.505 ;
        RECT 77.615 155.695 78.965 156.605 ;
        RECT 78.995 155.695 80.345 156.605 ;
        RECT 81.515 156.515 82.465 156.605 ;
        RECT 80.535 155.695 82.465 156.515 ;
        RECT 83.605 155.780 84.035 156.565 ;
        RECT 84.055 155.695 85.885 156.505 ;
        RECT 86.355 155.695 89.105 156.605 ;
        RECT 89.175 155.695 90.945 156.605 ;
        RECT 90.955 155.695 92.305 156.605 ;
        RECT 92.795 155.695 94.165 156.475 ;
        RECT 94.635 155.695 96.005 156.475 ;
        RECT 96.015 155.695 97.385 156.475 ;
        RECT 97.395 155.695 98.765 156.475 ;
        RECT 99.695 155.695 101.065 156.475 ;
        RECT 101.075 155.695 106.585 156.505 ;
        RECT 106.595 155.695 109.345 156.505 ;
        RECT 109.365 155.780 109.795 156.565 ;
        RECT 110.140 155.695 113.795 156.605 ;
        RECT 113.955 155.695 116.705 156.605 ;
        RECT 117.635 155.695 119.005 156.475 ;
        RECT 119.035 155.695 120.385 156.605 ;
        RECT 120.395 155.695 121.765 156.475 ;
        RECT 121.775 155.695 123.145 156.505 ;
        RECT 123.155 155.695 126.075 156.605 ;
        RECT 126.375 155.695 128.205 156.505 ;
        RECT 128.215 155.695 129.585 156.475 ;
        RECT 129.595 155.695 130.965 156.475 ;
        RECT 130.975 155.695 134.645 156.505 ;
        RECT 135.125 155.780 135.555 156.565 ;
        RECT 135.575 155.695 137.405 156.505 ;
        RECT 137.415 155.695 140.165 156.605 ;
        RECT 140.175 155.695 142.925 156.605 ;
        RECT 142.935 155.695 145.685 156.605 ;
        RECT 145.695 155.695 151.205 156.505 ;
        RECT 151.235 155.695 152.585 156.605 ;
        RECT 152.595 155.695 154.425 156.505 ;
        RECT 154.895 155.695 156.265 156.505 ;
        RECT 70.855 155.485 71.025 155.695 ;
        RECT 72.235 155.485 72.405 155.695 ;
        RECT 78.680 155.505 78.850 155.695 ;
        RECT 79.595 155.485 79.765 155.675 ;
        RECT 80.060 155.505 80.230 155.695 ;
        RECT 80.535 155.675 80.685 155.695 ;
        RECT 80.515 155.505 80.685 155.675 ;
        RECT 81.445 155.485 81.615 155.675 ;
        RECT 82.815 155.485 82.985 155.675 ;
        RECT 84.195 155.505 84.365 155.695 ;
        RECT 88.795 155.675 88.965 155.695 ;
        RECT 85.570 155.535 85.690 155.645 ;
        RECT 86.030 155.535 86.150 155.645 ;
        RECT 88.795 155.505 88.970 155.675 ;
        RECT 88.800 155.485 88.970 155.505 ;
        RECT 70.715 154.675 72.085 155.485 ;
        RECT 72.095 154.805 79.405 155.485 ;
        RECT 75.610 154.585 76.520 154.805 ;
        RECT 78.055 154.575 79.405 154.805 ;
        RECT 79.455 154.675 81.285 155.485 ;
        RECT 81.295 154.705 82.665 155.485 ;
        RECT 82.675 154.675 85.425 155.485 ;
        RECT 85.895 154.575 89.095 155.485 ;
        RECT 89.250 155.455 89.420 155.675 ;
        RECT 90.630 155.505 90.800 155.695 ;
        RECT 91.100 155.505 91.270 155.695 ;
        RECT 92.945 155.675 93.115 155.695 ;
        RECT 91.560 155.485 91.730 155.675 ;
        RECT 92.470 155.535 92.590 155.645 ;
        RECT 92.935 155.505 93.115 155.675 ;
        RECT 94.310 155.535 94.430 155.645 ;
        RECT 94.785 155.505 94.955 155.695 ;
        RECT 96.165 155.505 96.335 155.695 ;
        RECT 92.935 155.485 93.105 155.505 ;
        RECT 97.075 155.485 97.245 155.675 ;
        RECT 97.545 155.505 97.715 155.695 ;
        RECT 98.925 155.540 99.085 155.650 ;
        RECT 99.845 155.505 100.015 155.695 ;
        RECT 101.215 155.505 101.385 155.695 ;
        RECT 105.350 155.485 105.520 155.675 ;
        RECT 105.815 155.485 105.985 155.675 ;
        RECT 106.735 155.505 106.905 155.695 ;
        RECT 113.635 155.675 113.795 155.695 ;
        RECT 116.395 155.675 116.565 155.695 ;
        RECT 107.195 155.505 107.365 155.675 ;
        RECT 111.345 155.530 111.505 155.640 ;
        RECT 113.635 155.505 113.805 155.675 ;
        RECT 116.395 155.505 116.590 155.675 ;
        RECT 107.205 155.485 107.365 155.505 ;
        RECT 116.420 155.485 116.530 155.505 ;
        RECT 116.865 155.485 117.035 155.675 ;
        RECT 117.785 155.505 117.955 155.695 ;
        RECT 119.150 155.675 119.320 155.695 ;
        RECT 118.245 155.530 118.405 155.640 ;
        RECT 119.150 155.505 119.330 155.675 ;
        RECT 120.545 155.505 120.715 155.695 ;
        RECT 121.915 155.505 122.085 155.695 ;
        RECT 123.300 155.505 123.470 155.695 ;
        RECT 126.515 155.505 126.685 155.695 ;
        RECT 119.160 155.485 119.330 155.505 ;
        RECT 126.515 155.485 126.675 155.505 ;
        RECT 126.975 155.485 127.145 155.675 ;
        RECT 129.265 155.505 129.435 155.695 ;
        RECT 130.645 155.505 130.815 155.695 ;
        RECT 131.115 155.505 131.285 155.695 ;
        RECT 132.495 155.485 132.665 155.675 ;
        RECT 134.790 155.535 134.910 155.645 ;
        RECT 135.715 155.505 135.885 155.695 ;
        RECT 136.185 155.530 136.345 155.640 ;
        RECT 137.105 155.485 137.275 155.675 ;
        RECT 138.475 155.485 138.645 155.675 ;
        RECT 139.855 155.505 140.025 155.695 ;
        RECT 142.615 155.505 142.785 155.695 ;
        RECT 143.075 155.505 143.245 155.695 ;
        RECT 143.995 155.485 144.165 155.675 ;
        RECT 145.835 155.505 146.005 155.695 ;
        RECT 151.350 155.675 151.520 155.695 ;
        RECT 147.670 155.535 147.790 155.645 ;
        RECT 148.590 155.535 148.710 155.645 ;
        RECT 150.895 155.505 151.065 155.675 ;
        RECT 151.350 155.505 151.525 155.675 ;
        RECT 152.735 155.505 152.905 155.695 ;
        RECT 154.570 155.535 154.690 155.645 ;
        RECT 150.895 155.485 151.060 155.505 ;
        RECT 151.355 155.485 151.525 155.505 ;
        RECT 155.955 155.485 156.125 155.695 ;
        RECT 90.450 155.455 91.405 155.485 ;
        RECT 89.125 154.775 91.405 155.455 ;
        RECT 90.450 154.575 91.405 154.775 ;
        RECT 91.415 154.575 92.765 155.485 ;
        RECT 92.795 154.675 96.465 155.485 ;
        RECT 96.485 154.615 96.915 155.400 ;
        RECT 96.935 154.675 102.445 155.485 ;
        RECT 102.745 154.575 105.665 155.485 ;
        RECT 105.675 154.675 107.045 155.485 ;
        RECT 107.205 154.575 110.860 155.485 ;
        RECT 112.115 154.805 116.530 155.485 ;
        RECT 112.115 154.575 116.045 154.805 ;
        RECT 116.715 154.705 118.085 155.485 ;
        RECT 119.015 154.575 121.935 155.485 ;
        RECT 122.245 154.615 122.675 155.400 ;
        RECT 123.020 154.575 126.675 155.485 ;
        RECT 126.835 154.675 132.345 155.485 ;
        RECT 132.355 154.675 136.025 155.485 ;
        RECT 136.955 154.705 138.325 155.485 ;
        RECT 138.335 154.675 143.845 155.485 ;
        RECT 143.855 154.675 147.525 155.485 ;
        RECT 148.005 154.615 148.435 155.400 ;
        RECT 149.225 154.805 151.060 155.485 ;
        RECT 149.225 154.575 150.155 154.805 ;
        RECT 151.215 154.675 154.885 155.485 ;
        RECT 154.895 154.675 156.265 155.485 ;
      LAYER nwell ;
        RECT 70.520 151.455 156.460 154.285 ;
      LAYER pwell ;
        RECT 70.715 150.255 72.085 151.065 ;
        RECT 72.095 150.255 77.605 151.065 ;
        RECT 77.615 150.255 80.365 151.065 ;
        RECT 80.835 150.255 82.205 151.035 ;
        RECT 82.215 150.255 83.585 151.065 ;
        RECT 83.605 150.340 84.035 151.125 ;
        RECT 84.055 150.255 89.565 151.065 ;
        RECT 89.575 150.255 95.085 151.065 ;
        RECT 95.095 150.255 96.925 151.065 ;
        RECT 96.935 150.255 98.305 151.035 ;
        RECT 98.975 150.935 102.905 151.165 ;
        RECT 98.490 150.255 102.905 150.935 ;
        RECT 103.240 150.255 106.895 151.165 ;
        RECT 107.055 150.255 108.425 151.035 ;
        RECT 109.365 150.340 109.795 151.125 ;
        RECT 109.815 150.255 112.565 151.165 ;
        RECT 112.575 150.255 113.945 151.035 ;
        RECT 113.955 150.255 119.465 151.065 ;
        RECT 119.475 150.255 123.145 151.065 ;
        RECT 123.155 150.255 125.905 151.165 ;
        RECT 125.915 150.255 127.285 151.065 ;
        RECT 127.295 150.255 128.665 151.035 ;
        RECT 128.675 150.255 130.505 151.065 ;
        RECT 130.975 150.255 132.345 151.035 ;
        RECT 132.355 150.255 135.105 151.065 ;
        RECT 135.125 150.340 135.555 151.125 ;
        RECT 135.725 150.255 139.380 151.165 ;
        RECT 139.715 150.255 142.465 151.165 ;
        RECT 144.055 150.935 147.985 151.165 ;
        RECT 143.570 150.255 147.985 150.935 ;
        RECT 148.015 150.255 149.365 151.165 ;
        RECT 149.375 150.255 150.725 151.165 ;
        RECT 150.765 150.255 152.115 151.165 ;
        RECT 152.135 150.255 153.505 151.035 ;
        RECT 153.515 150.255 154.885 151.065 ;
        RECT 154.895 150.255 156.265 151.065 ;
        RECT 70.855 150.045 71.025 150.255 ;
        RECT 72.235 150.045 72.405 150.255 ;
        RECT 77.755 150.065 77.925 150.255 ;
        RECT 79.605 150.090 79.765 150.200 ;
        RECT 80.510 150.095 80.630 150.205 ;
        RECT 81.430 150.045 81.600 150.235 ;
        RECT 81.885 150.065 82.055 150.255 ;
        RECT 82.355 150.065 82.525 150.255 ;
        RECT 83.275 150.045 83.445 150.235 ;
        RECT 83.730 150.095 83.850 150.205 ;
        RECT 84.195 150.065 84.365 150.255 ;
        RECT 86.035 150.065 86.205 150.235 ;
        RECT 86.035 150.045 86.185 150.065 ;
        RECT 87.870 150.045 88.040 150.235 ;
        RECT 88.310 150.065 88.480 150.235 ;
        RECT 89.715 150.065 89.885 150.255 ;
        RECT 88.370 150.045 88.480 150.065 ;
        RECT 92.935 150.045 93.105 150.235 ;
        RECT 95.235 150.065 95.405 150.255 ;
        RECT 97.985 150.065 98.155 150.255 ;
        RECT 98.490 150.235 98.600 150.255 ;
        RECT 106.735 150.235 106.895 150.255 ;
        RECT 98.430 150.065 98.600 150.235 ;
        RECT 100.755 150.065 100.925 150.235 ;
        RECT 100.755 150.045 100.915 150.065 ;
        RECT 101.215 150.045 101.385 150.235 ;
        RECT 102.595 150.045 102.765 150.235 ;
        RECT 105.355 150.045 105.525 150.235 ;
        RECT 106.735 150.065 106.905 150.235 ;
        RECT 108.105 150.065 108.275 150.255 ;
        RECT 108.585 150.100 108.745 150.210 ;
        RECT 109.955 150.065 110.125 150.255 ;
        RECT 110.875 150.045 111.045 150.235 ;
        RECT 112.725 150.065 112.895 150.255 ;
        RECT 114.095 150.065 114.265 150.255 ;
        RECT 119.615 150.235 119.785 150.255 ;
        RECT 115.935 150.045 116.105 150.235 ;
        RECT 118.235 150.065 118.405 150.235 ;
        RECT 119.605 150.065 119.785 150.235 ;
        RECT 118.235 150.045 118.400 150.065 ;
        RECT 119.605 150.045 119.775 150.065 ;
        RECT 120.075 150.045 120.245 150.235 ;
        RECT 121.910 150.095 122.030 150.205 ;
        RECT 122.835 150.045 123.005 150.235 ;
        RECT 123.295 150.065 123.465 150.255 ;
        RECT 126.055 150.065 126.225 150.255 ;
        RECT 126.515 150.045 126.685 150.235 ;
        RECT 127.445 150.065 127.615 150.255 ;
        RECT 128.815 150.065 128.985 150.255 ;
        RECT 130.650 150.095 130.770 150.205 ;
        RECT 131.110 150.045 131.280 150.235 ;
        RECT 131.575 150.045 131.745 150.235 ;
        RECT 132.025 150.065 132.195 150.255 ;
        RECT 132.495 150.065 132.665 150.255 ;
        RECT 135.725 150.235 135.885 150.255 ;
        RECT 142.155 150.235 142.325 150.255 ;
        RECT 143.570 150.235 143.680 150.255 ;
        RECT 134.795 150.045 134.965 150.235 ;
        RECT 135.715 150.065 135.885 150.235 ;
        RECT 138.015 150.045 138.185 150.235 ;
        RECT 140.770 150.095 140.890 150.205 ;
        RECT 142.145 150.065 142.325 150.235 ;
        RECT 142.625 150.100 142.785 150.210 ;
        RECT 143.510 150.065 143.695 150.235 ;
        RECT 142.145 150.045 142.315 150.065 ;
        RECT 143.525 150.045 143.695 150.065 ;
        RECT 147.675 150.065 147.845 150.235 ;
        RECT 148.130 150.065 148.300 150.255 ;
        RECT 147.675 150.045 147.835 150.065 ;
        RECT 149.515 150.045 149.685 150.235 ;
        RECT 149.970 150.095 150.090 150.205 ;
        RECT 150.440 150.045 150.610 150.255 ;
        RECT 150.895 150.065 151.065 150.255 ;
        RECT 152.740 150.045 152.910 150.235 ;
        RECT 153.185 150.065 153.355 150.255 ;
        RECT 153.655 150.065 153.825 150.255 ;
        RECT 154.125 150.090 154.285 150.200 ;
        RECT 155.955 150.045 156.125 150.255 ;
        RECT 70.715 149.235 72.085 150.045 ;
        RECT 72.095 149.365 79.405 150.045 ;
        RECT 75.610 149.145 76.520 149.365 ;
        RECT 78.055 149.135 79.405 149.365 ;
        RECT 80.395 149.135 81.745 150.045 ;
        RECT 81.755 149.135 83.570 150.045 ;
        RECT 84.255 149.225 86.185 150.045 ;
        RECT 84.255 149.135 85.205 149.225 ;
        RECT 86.355 149.135 88.185 150.045 ;
        RECT 88.370 149.365 92.785 150.045 ;
        RECT 88.855 149.135 92.785 149.365 ;
        RECT 92.795 149.235 96.465 150.045 ;
        RECT 96.485 149.175 96.915 149.960 ;
        RECT 97.260 149.135 100.915 150.045 ;
        RECT 101.075 149.235 102.445 150.045 ;
        RECT 102.455 149.135 105.205 150.045 ;
        RECT 105.215 149.235 110.725 150.045 ;
        RECT 110.735 149.235 113.485 150.045 ;
        RECT 113.495 149.135 116.245 150.045 ;
        RECT 116.565 149.365 118.400 150.045 ;
        RECT 116.565 149.135 117.495 149.365 ;
        RECT 118.555 149.265 119.925 150.045 ;
        RECT 119.935 149.235 121.765 150.045 ;
        RECT 122.245 149.175 122.675 149.960 ;
        RECT 122.695 149.235 126.365 150.045 ;
        RECT 126.375 149.235 127.745 150.045 ;
        RECT 127.950 149.135 131.425 150.045 ;
        RECT 131.435 149.135 134.645 150.045 ;
        RECT 134.655 149.135 137.865 150.045 ;
        RECT 137.875 149.235 140.625 150.045 ;
        RECT 141.095 149.265 142.465 150.045 ;
        RECT 142.475 149.265 143.845 150.045 ;
        RECT 144.180 149.135 147.835 150.045 ;
        RECT 148.005 149.175 148.435 149.960 ;
        RECT 148.465 149.135 149.815 150.045 ;
        RECT 150.295 149.135 152.505 150.045 ;
        RECT 152.595 149.135 153.945 150.045 ;
        RECT 154.895 149.235 156.265 150.045 ;
      LAYER nwell ;
        RECT 70.520 146.015 156.460 148.845 ;
      LAYER pwell ;
        RECT 70.715 144.815 72.085 145.625 ;
        RECT 72.115 144.815 73.465 145.725 ;
        RECT 73.485 144.815 74.835 145.725 ;
        RECT 75.905 145.495 76.835 145.725 ;
        RECT 75.000 144.815 76.835 145.495 ;
        RECT 77.155 145.495 78.075 145.725 ;
        RECT 77.155 144.815 79.445 145.495 ;
        RECT 79.455 144.815 81.285 145.725 ;
        RECT 81.295 145.495 82.215 145.725 ;
        RECT 81.295 144.815 83.585 145.495 ;
        RECT 83.605 144.900 84.035 145.685 ;
        RECT 84.975 144.815 87.895 145.725 ;
        RECT 88.195 144.815 89.565 145.595 ;
        RECT 89.575 144.815 92.325 145.625 ;
        RECT 92.485 144.815 96.140 145.725 ;
        RECT 96.475 144.815 98.305 145.625 ;
        RECT 99.435 145.495 103.365 145.725 ;
        RECT 98.950 144.815 103.365 145.495 ;
        RECT 103.375 144.815 106.585 145.725 ;
        RECT 106.595 144.815 109.345 145.625 ;
        RECT 109.365 144.900 109.795 145.685 ;
        RECT 109.815 144.815 113.025 145.725 ;
        RECT 113.035 144.815 114.405 145.595 ;
        RECT 114.415 144.815 117.625 145.725 ;
        RECT 118.880 144.815 122.535 145.725 ;
        RECT 122.695 144.815 125.445 145.725 ;
        RECT 125.455 144.815 127.285 145.625 ;
        RECT 127.445 144.815 131.100 145.725 ;
        RECT 131.435 144.815 132.805 145.595 ;
        RECT 132.815 144.815 134.645 145.625 ;
        RECT 135.125 144.900 135.555 145.685 ;
        RECT 135.575 144.815 138.785 145.725 ;
        RECT 138.795 144.815 144.305 145.625 ;
        RECT 144.315 144.815 149.825 145.625 ;
        RECT 149.835 144.815 153.505 145.625 ;
        RECT 153.515 144.815 154.885 145.625 ;
        RECT 154.895 144.815 156.265 145.625 ;
        RECT 70.855 144.605 71.025 144.815 ;
        RECT 72.230 144.795 72.400 144.815 ;
        RECT 72.230 144.625 72.405 144.795 ;
        RECT 74.535 144.625 74.705 144.815 ;
        RECT 75.000 144.795 75.165 144.815 ;
        RECT 72.235 144.605 72.405 144.625 ;
        RECT 74.995 144.605 75.165 144.795 ;
        RECT 75.450 144.655 75.570 144.765 ;
        RECT 77.295 144.605 77.465 144.795 ;
        RECT 77.755 144.605 77.925 144.795 ;
        RECT 79.135 144.625 79.305 144.815 ;
        RECT 79.600 144.625 79.770 144.815 ;
        RECT 83.275 144.625 83.445 144.815 ;
        RECT 85.120 144.795 85.290 144.815 ;
        RECT 84.205 144.660 84.365 144.770 ;
        RECT 84.650 144.605 84.820 144.795 ;
        RECT 85.115 144.625 85.290 144.795 ;
        RECT 85.115 144.605 85.285 144.625 ;
        RECT 86.495 144.605 86.665 144.795 ;
        RECT 88.345 144.625 88.515 144.815 ;
        RECT 89.715 144.625 89.885 144.815 ;
        RECT 92.485 144.795 92.645 144.815 ;
        RECT 92.010 144.655 92.130 144.765 ;
        RECT 92.475 144.625 92.645 144.795 ;
        RECT 96.615 144.625 96.785 144.815 ;
        RECT 98.950 144.795 99.060 144.815 ;
        RECT 97.075 144.625 97.245 144.795 ;
        RECT 98.450 144.655 98.570 144.765 ;
        RECT 98.890 144.625 99.060 144.795 ;
        RECT 92.485 144.605 92.645 144.625 ;
        RECT 97.085 144.605 97.245 144.625 ;
        RECT 101.215 144.605 101.385 144.795 ;
        RECT 103.515 144.625 103.685 144.815 ;
        RECT 104.895 144.605 105.065 144.795 ;
        RECT 106.735 144.625 106.905 144.815 ;
        RECT 109.035 144.625 109.205 144.795 ;
        RECT 109.035 144.605 109.195 144.625 ;
        RECT 109.495 144.605 109.665 144.795 ;
        RECT 109.955 144.625 110.125 144.815 ;
        RECT 113.185 144.625 113.355 144.815 ;
        RECT 117.315 144.625 117.485 144.815 ;
        RECT 122.375 144.795 122.535 144.815 ;
        RECT 117.785 144.660 117.945 144.770 ;
        RECT 118.695 144.625 118.865 144.795 ;
        RECT 118.695 144.605 118.855 144.625 ;
        RECT 119.155 144.605 119.325 144.795 ;
        RECT 121.910 144.655 122.030 144.765 ;
        RECT 122.375 144.625 122.545 144.795 ;
        RECT 122.835 144.605 123.005 144.815 ;
        RECT 125.595 144.795 125.765 144.815 ;
        RECT 127.445 144.795 127.605 144.815 ;
        RECT 125.585 144.625 125.765 144.795 ;
        RECT 126.055 144.625 126.225 144.795 ;
        RECT 127.435 144.625 127.605 144.795 ;
        RECT 128.330 144.625 128.500 144.795 ;
        RECT 132.485 144.625 132.655 144.815 ;
        RECT 125.585 144.605 125.755 144.625 ;
        RECT 126.060 144.605 126.225 144.625 ;
        RECT 128.390 144.605 128.500 144.625 ;
        RECT 132.955 144.605 133.125 144.815 ;
        RECT 134.790 144.655 134.910 144.765 ;
        RECT 135.710 144.655 135.830 144.765 ;
        RECT 138.475 144.625 138.645 144.815 ;
        RECT 138.935 144.795 139.105 144.815 ;
        RECT 138.930 144.625 139.105 144.795 ;
        RECT 139.405 144.650 139.565 144.760 ;
        RECT 142.155 144.625 142.325 144.795 ;
        RECT 138.930 144.605 139.100 144.625 ;
        RECT 142.155 144.605 142.320 144.625 ;
        RECT 143.540 144.605 143.710 144.795 ;
        RECT 143.995 144.605 144.165 144.795 ;
        RECT 144.455 144.625 144.625 144.815 ;
        RECT 147.670 144.655 147.790 144.765 ;
        RECT 148.590 144.655 148.710 144.765 ;
        RECT 149.975 144.625 150.145 144.815 ;
        RECT 151.815 144.605 151.985 144.795 ;
        RECT 152.275 144.605 152.445 144.795 ;
        RECT 153.655 144.625 153.825 144.815 ;
        RECT 155.955 144.605 156.125 144.815 ;
        RECT 70.715 143.795 72.085 144.605 ;
        RECT 72.095 143.795 73.925 144.605 ;
        RECT 73.935 143.825 75.305 144.605 ;
        RECT 75.775 143.925 77.605 144.605 ;
        RECT 77.615 143.795 83.125 144.605 ;
        RECT 83.135 143.695 84.965 144.605 ;
        RECT 84.975 143.825 86.345 144.605 ;
        RECT 86.355 143.795 91.865 144.605 ;
        RECT 92.485 143.695 96.140 144.605 ;
        RECT 96.485 143.735 96.915 144.520 ;
        RECT 97.085 143.695 100.740 144.605 ;
        RECT 101.075 143.795 102.445 144.605 ;
        RECT 102.455 143.695 105.205 144.605 ;
        RECT 105.540 143.695 109.195 144.605 ;
        RECT 109.355 143.795 114.865 144.605 ;
        RECT 115.200 143.695 118.855 144.605 ;
        RECT 119.015 143.795 121.765 144.605 ;
        RECT 122.245 143.735 122.675 144.520 ;
        RECT 122.695 143.795 124.525 144.605 ;
        RECT 124.535 143.825 125.905 144.605 ;
        RECT 126.060 143.925 127.895 144.605 ;
        RECT 128.390 143.925 132.805 144.605 ;
        RECT 126.965 143.695 127.895 143.925 ;
        RECT 128.875 143.695 132.805 143.925 ;
        RECT 132.815 143.795 135.565 144.605 ;
        RECT 136.325 143.695 139.245 144.605 ;
        RECT 140.485 143.925 142.320 144.605 ;
        RECT 140.485 143.695 141.415 143.925 ;
        RECT 142.475 143.695 143.825 144.605 ;
        RECT 143.855 143.795 147.525 144.605 ;
        RECT 148.005 143.735 148.435 144.520 ;
        RECT 148.915 143.695 152.085 144.605 ;
        RECT 152.135 143.795 154.885 144.605 ;
        RECT 154.895 143.795 156.265 144.605 ;
      LAYER nwell ;
        RECT 70.520 140.575 156.460 143.405 ;
      LAYER pwell ;
        RECT 70.715 139.375 72.085 140.185 ;
        RECT 75.610 140.055 76.520 140.275 ;
        RECT 78.055 140.055 79.405 140.285 ;
        RECT 72.095 139.375 79.405 140.055 ;
        RECT 79.655 140.195 80.605 140.285 ;
        RECT 79.655 139.375 81.585 140.195 ;
        RECT 81.755 139.375 83.585 140.055 ;
        RECT 83.605 139.460 84.035 140.245 ;
        RECT 87.570 140.055 88.480 140.275 ;
        RECT 90.015 140.055 91.365 140.285 ;
        RECT 84.055 139.375 91.365 140.055 ;
        RECT 91.415 139.375 94.165 140.185 ;
        RECT 94.635 139.375 98.110 140.285 ;
        RECT 98.315 139.375 101.065 140.285 ;
        RECT 101.075 139.375 103.825 140.185 ;
        RECT 103.835 139.375 106.585 140.285 ;
        RECT 106.595 139.375 109.345 140.185 ;
        RECT 109.365 139.460 109.795 140.245 ;
        RECT 109.815 139.375 115.325 140.185 ;
        RECT 115.815 139.375 117.165 140.285 ;
        RECT 117.175 139.375 119.925 140.185 ;
        RECT 120.395 140.055 124.325 140.285 ;
        RECT 120.395 139.375 124.810 140.055 ;
        RECT 124.995 139.375 126.365 140.155 ;
        RECT 126.835 140.055 130.765 140.285 ;
        RECT 126.835 139.375 131.250 140.055 ;
        RECT 132.185 139.375 135.105 140.285 ;
        RECT 135.125 139.460 135.555 140.245 ;
        RECT 135.575 139.375 139.050 140.285 ;
        RECT 139.255 139.375 142.175 140.285 ;
        RECT 143.395 140.055 144.315 140.285 ;
        RECT 143.395 139.375 146.980 140.055 ;
        RECT 147.155 139.375 150.155 140.285 ;
        RECT 150.295 139.375 151.665 140.185 ;
        RECT 151.685 139.375 154.885 140.285 ;
        RECT 154.895 139.375 156.265 140.185 ;
        RECT 70.855 139.165 71.025 139.375 ;
        RECT 72.235 139.165 72.405 139.375 ;
        RECT 81.435 139.355 81.585 139.375 ;
        RECT 75.915 139.165 76.085 139.355 ;
        RECT 77.295 139.165 77.465 139.355 ;
        RECT 80.060 139.165 80.230 139.355 ;
        RECT 81.435 139.185 81.605 139.355 ;
        RECT 81.895 139.185 82.065 139.375 ;
        RECT 82.355 139.165 82.525 139.355 ;
        RECT 84.195 139.185 84.365 139.375 ;
        RECT 86.980 139.185 87.150 139.355 ;
        RECT 86.980 139.165 87.090 139.185 ;
        RECT 87.415 139.165 87.585 139.355 ;
        RECT 91.555 139.185 91.725 139.375 ;
        RECT 92.935 139.165 93.105 139.355 ;
        RECT 94.315 139.325 94.485 139.355 ;
        RECT 94.310 139.215 94.485 139.325 ;
        RECT 94.315 139.185 94.485 139.215 ;
        RECT 94.780 139.185 94.950 139.375 ;
        RECT 97.070 139.215 97.190 139.325 ;
        RECT 99.375 139.185 99.545 139.355 ;
        RECT 94.320 139.165 94.485 139.185 ;
        RECT 99.375 139.165 99.540 139.185 ;
        RECT 99.845 139.165 100.015 139.355 ;
        RECT 100.755 139.185 100.925 139.375 ;
        RECT 101.215 139.165 101.385 139.375 ;
        RECT 103.975 139.185 104.145 139.375 ;
        RECT 104.905 139.210 105.065 139.320 ;
        RECT 105.820 139.165 105.990 139.355 ;
        RECT 106.735 139.185 106.905 139.375 ;
        RECT 109.495 139.165 109.665 139.355 ;
        RECT 109.955 139.185 110.125 139.375 ;
        RECT 112.250 139.215 112.370 139.325 ;
        RECT 112.715 139.185 112.885 139.355 ;
        RECT 115.480 139.325 115.650 139.355 ;
        RECT 115.010 139.215 115.130 139.325 ;
        RECT 115.470 139.215 115.650 139.325 ;
        RECT 112.720 139.165 112.885 139.185 ;
        RECT 115.480 139.165 115.650 139.215 ;
        RECT 115.930 139.185 116.100 139.375 ;
        RECT 117.315 139.185 117.485 139.375 ;
        RECT 124.700 139.355 124.810 139.375 ;
        RECT 120.070 139.215 120.190 139.325 ;
        RECT 121.910 139.165 122.080 139.355 ;
        RECT 122.835 139.165 123.005 139.355 ;
        RECT 124.700 139.185 124.870 139.355 ;
        RECT 125.590 139.215 125.710 139.325 ;
        RECT 126.045 139.185 126.215 139.375 ;
        RECT 131.140 139.355 131.250 139.375 ;
        RECT 126.510 139.215 126.630 139.325 ;
        RECT 128.355 139.165 128.525 139.355 ;
        RECT 128.825 139.165 128.995 139.355 ;
        RECT 131.120 139.185 131.310 139.355 ;
        RECT 131.575 139.325 131.745 139.355 ;
        RECT 131.570 139.215 131.745 139.325 ;
        RECT 131.120 139.165 131.290 139.185 ;
        RECT 131.575 139.165 131.745 139.215 ;
        RECT 134.790 139.185 134.960 139.375 ;
        RECT 135.720 139.185 135.890 139.375 ;
        RECT 136.630 139.165 136.800 139.355 ;
        RECT 138.020 139.165 138.190 139.355 ;
        RECT 139.400 139.185 139.570 139.375 ;
        RECT 141.230 139.165 141.400 139.355 ;
        RECT 141.670 139.185 141.840 139.355 ;
        RECT 142.625 139.220 142.785 139.330 ;
        RECT 143.540 139.185 143.710 139.375 ;
        RECT 141.730 139.165 141.840 139.185 ;
        RECT 146.295 139.165 146.465 139.355 ;
        RECT 147.215 139.185 147.385 139.375 ;
        RECT 150.435 139.185 150.605 139.375 ;
        RECT 151.810 139.355 151.980 139.375 ;
        RECT 151.355 139.165 151.525 139.355 ;
        RECT 151.810 139.185 151.990 139.355 ;
        RECT 154.570 139.215 154.690 139.325 ;
        RECT 70.715 138.355 72.085 139.165 ;
        RECT 72.095 138.355 75.765 139.165 ;
        RECT 75.775 138.355 77.145 139.165 ;
        RECT 77.165 138.255 79.895 139.165 ;
        RECT 79.915 138.255 81.265 139.165 ;
        RECT 81.305 138.255 82.655 139.165 ;
        RECT 82.675 138.485 87.090 139.165 ;
        RECT 82.675 138.255 86.605 138.485 ;
        RECT 87.275 138.355 92.785 139.165 ;
        RECT 92.795 138.355 94.165 139.165 ;
        RECT 94.320 138.485 96.155 139.165 ;
        RECT 95.225 138.255 96.155 138.485 ;
        RECT 96.485 138.295 96.915 139.080 ;
        RECT 97.705 138.485 99.540 139.165 ;
        RECT 97.705 138.255 98.635 138.485 ;
        RECT 99.695 138.385 101.065 139.165 ;
        RECT 101.075 138.355 104.745 139.165 ;
        RECT 105.675 138.255 109.150 139.165 ;
        RECT 109.355 138.355 112.105 139.165 ;
        RECT 112.720 138.485 114.555 139.165 ;
        RECT 113.625 138.255 114.555 138.485 ;
        RECT 115.335 138.255 118.810 139.165 ;
        RECT 119.305 138.255 122.225 139.165 ;
        RECT 122.245 138.295 122.675 139.080 ;
        RECT 122.695 138.355 125.445 139.165 ;
        RECT 125.915 138.485 128.665 139.165 ;
        RECT 125.915 138.255 126.845 138.485 ;
        RECT 128.675 138.385 130.045 139.165 ;
        RECT 130.055 138.255 131.405 139.165 ;
        RECT 131.435 138.355 133.265 139.165 ;
        RECT 133.470 138.255 136.945 139.165 ;
        RECT 136.955 138.255 138.305 139.165 ;
        RECT 138.625 138.255 141.545 139.165 ;
        RECT 141.730 138.485 146.145 139.165 ;
        RECT 142.215 138.255 146.145 138.485 ;
        RECT 146.155 138.355 147.985 139.165 ;
        RECT 148.005 138.295 148.435 139.080 ;
        RECT 148.455 138.255 151.625 139.165 ;
        RECT 151.820 139.135 151.990 139.185 ;
        RECT 155.955 139.165 156.125 139.375 ;
        RECT 153.480 139.135 154.425 139.165 ;
        RECT 151.675 138.455 154.425 139.135 ;
        RECT 153.480 138.255 154.425 138.455 ;
        RECT 154.895 138.355 156.265 139.165 ;
      LAYER nwell ;
        RECT 70.520 135.135 156.460 137.965 ;
      LAYER pwell ;
        RECT 70.715 133.935 72.085 134.745 ;
        RECT 72.095 133.935 74.845 134.745 ;
        RECT 75.415 133.935 78.525 134.845 ;
        RECT 78.535 133.935 79.885 134.845 ;
        RECT 79.915 133.935 83.585 134.745 ;
        RECT 83.605 134.020 84.035 134.805 ;
        RECT 84.055 133.935 85.885 134.745 ;
        RECT 86.375 133.935 87.725 134.845 ;
        RECT 88.875 134.755 89.825 134.845 ;
        RECT 87.895 133.935 89.825 134.755 ;
        RECT 90.235 134.755 91.185 134.845 ;
        RECT 90.235 133.935 92.165 134.755 ;
        RECT 92.335 133.935 94.165 134.745 ;
        RECT 94.195 133.935 95.545 134.845 ;
        RECT 95.555 133.935 99.225 134.845 ;
        RECT 99.525 133.935 102.445 134.845 ;
        RECT 102.915 133.935 104.285 134.715 ;
        RECT 104.295 133.935 105.665 134.715 ;
        RECT 105.965 133.935 108.885 134.845 ;
        RECT 109.365 134.020 109.795 134.805 ;
        RECT 109.815 133.935 113.485 134.745 ;
        RECT 113.495 133.935 114.865 134.745 ;
        RECT 114.875 133.935 117.795 134.845 ;
        RECT 118.095 133.935 123.605 134.745 ;
        RECT 123.615 133.935 126.365 134.745 ;
        RECT 126.835 133.935 130.045 134.845 ;
        RECT 130.055 133.935 133.725 134.745 ;
        RECT 133.735 133.935 135.105 134.715 ;
        RECT 135.125 134.020 135.555 134.805 ;
        RECT 135.575 133.935 138.495 134.845 ;
        RECT 139.105 134.615 140.035 134.845 ;
        RECT 139.105 133.935 140.940 134.615 ;
        RECT 141.095 133.935 143.845 134.745 ;
        RECT 144.975 134.615 148.905 134.845 ;
        RECT 150.320 134.615 151.665 134.845 ;
        RECT 144.490 133.935 148.905 134.615 ;
        RECT 149.835 133.935 151.665 134.615 ;
        RECT 151.675 133.935 153.505 134.845 ;
        RECT 153.535 133.935 154.885 134.845 ;
        RECT 154.895 133.935 156.265 134.745 ;
        RECT 70.855 133.725 71.025 133.935 ;
        RECT 72.235 133.725 72.405 133.935 ;
        RECT 74.990 133.775 75.110 133.885 ;
        RECT 75.455 133.725 75.625 133.935 ;
        RECT 78.680 133.745 78.850 133.935 ;
        RECT 80.055 133.745 80.225 133.935 ;
        RECT 80.975 133.725 81.145 133.915 ;
        RECT 82.810 133.775 82.930 133.885 ;
        RECT 83.280 133.725 83.450 133.915 ;
        RECT 84.195 133.745 84.365 133.935 ;
        RECT 85.575 133.725 85.745 133.915 ;
        RECT 86.030 133.775 86.150 133.885 ;
        RECT 87.410 133.745 87.580 133.935 ;
        RECT 87.895 133.915 88.045 133.935 ;
        RECT 92.015 133.915 92.165 133.935 ;
        RECT 87.875 133.745 88.045 133.915 ;
        RECT 88.340 133.725 88.510 133.915 ;
        RECT 89.715 133.725 89.885 133.915 ;
        RECT 92.015 133.745 92.185 133.915 ;
        RECT 92.475 133.745 92.645 133.935 ;
        RECT 94.310 133.745 94.480 133.935 ;
        RECT 95.235 133.725 95.405 133.915 ;
        RECT 95.700 133.745 95.870 133.935 ;
        RECT 97.075 133.725 97.245 133.915 ;
        RECT 100.745 133.725 100.915 133.915 ;
        RECT 101.215 133.725 101.385 133.915 ;
        RECT 102.130 133.745 102.300 133.935 ;
        RECT 102.590 133.775 102.710 133.885 ;
        RECT 103.065 133.745 103.235 133.935 ;
        RECT 103.970 133.775 104.090 133.885 ;
        RECT 104.445 133.745 104.615 133.935 ;
        RECT 106.275 133.745 106.445 133.915 ;
        RECT 106.275 133.725 106.440 133.745 ;
        RECT 106.735 133.725 106.905 133.915 ;
        RECT 108.570 133.745 108.740 133.935 ;
        RECT 109.030 133.775 109.150 133.885 ;
        RECT 109.955 133.745 110.125 133.935 ;
        RECT 112.245 133.725 112.415 133.915 ;
        RECT 113.635 133.745 113.805 133.935 ;
        RECT 115.020 133.745 115.190 133.935 ;
        RECT 115.475 133.725 115.645 133.915 ;
        RECT 118.235 133.745 118.405 133.935 ;
        RECT 120.995 133.725 121.165 133.915 ;
        RECT 122.835 133.725 123.005 133.915 ;
        RECT 123.755 133.745 123.925 133.935 ;
        RECT 124.685 133.725 124.855 133.915 ;
        RECT 126.055 133.725 126.225 133.915 ;
        RECT 126.510 133.775 126.630 133.885 ;
        RECT 126.965 133.745 127.135 133.935 ;
        RECT 130.195 133.915 130.365 133.935 ;
        RECT 128.810 133.775 128.930 133.885 ;
        RECT 130.185 133.745 130.365 133.915 ;
        RECT 130.185 133.725 130.355 133.745 ;
        RECT 130.655 133.725 130.825 133.915 ;
        RECT 132.045 133.725 132.215 133.915 ;
        RECT 133.415 133.725 133.585 133.915 ;
        RECT 133.885 133.745 134.055 133.935 ;
        RECT 135.720 133.745 135.890 133.935 ;
        RECT 140.775 133.915 140.940 133.935 ;
        RECT 137.095 133.725 137.265 133.915 ;
        RECT 138.480 133.725 138.650 133.915 ;
        RECT 140.775 133.745 140.945 133.915 ;
        RECT 141.235 133.745 141.405 133.935 ;
        RECT 144.490 133.915 144.600 133.935 ;
        RECT 142.620 133.725 142.790 133.915 ;
        RECT 143.070 133.775 143.190 133.885 ;
        RECT 143.990 133.775 144.110 133.885 ;
        RECT 144.430 133.745 144.620 133.915 ;
        RECT 144.450 133.725 144.620 133.745 ;
        RECT 144.920 133.725 145.090 133.915 ;
        RECT 146.295 133.725 146.465 133.915 ;
        RECT 148.595 133.725 148.765 133.915 ;
        RECT 149.065 133.780 149.225 133.890 ;
        RECT 149.975 133.745 150.145 133.935 ;
        RECT 150.890 133.775 151.010 133.885 ;
        RECT 151.820 133.745 151.990 133.935 ;
        RECT 153.195 133.745 153.365 133.915 ;
        RECT 153.650 133.745 153.820 133.935 ;
        RECT 153.195 133.725 153.360 133.745 ;
        RECT 154.580 133.725 154.750 133.915 ;
        RECT 155.955 133.725 156.125 133.935 ;
        RECT 70.715 132.915 72.085 133.725 ;
        RECT 72.195 132.815 75.305 133.725 ;
        RECT 75.315 132.915 80.825 133.725 ;
        RECT 80.835 132.915 82.665 133.725 ;
        RECT 83.135 132.815 85.425 133.725 ;
        RECT 85.435 132.915 88.185 133.725 ;
        RECT 88.195 132.815 89.545 133.725 ;
        RECT 89.575 132.915 95.085 133.725 ;
        RECT 95.095 132.915 96.465 133.725 ;
        RECT 96.485 132.855 96.915 133.640 ;
        RECT 96.935 132.815 99.685 133.725 ;
        RECT 99.695 132.945 101.065 133.725 ;
        RECT 101.075 132.915 103.825 133.725 ;
        RECT 104.605 133.045 106.440 133.725 ;
        RECT 104.605 132.815 105.535 133.045 ;
        RECT 106.595 132.915 112.105 133.725 ;
        RECT 112.115 132.815 115.325 133.725 ;
        RECT 115.335 132.915 120.845 133.725 ;
        RECT 120.855 132.915 122.225 133.725 ;
        RECT 122.245 132.855 122.675 133.640 ;
        RECT 122.695 133.045 124.525 133.725 ;
        RECT 124.535 132.945 125.905 133.725 ;
        RECT 125.915 132.915 128.665 133.725 ;
        RECT 129.135 132.945 130.505 133.725 ;
        RECT 130.515 132.945 131.885 133.725 ;
        RECT 131.895 132.945 133.265 133.725 ;
        RECT 133.275 132.915 136.945 133.725 ;
        RECT 136.955 132.915 138.325 133.725 ;
        RECT 138.335 132.815 141.255 133.725 ;
        RECT 141.555 132.815 142.905 133.725 ;
        RECT 143.415 132.815 144.765 133.725 ;
        RECT 144.775 132.815 146.125 133.725 ;
        RECT 146.155 133.045 147.985 133.725 ;
        RECT 146.640 132.815 147.985 133.045 ;
        RECT 148.005 132.855 148.435 133.640 ;
        RECT 148.455 133.045 150.745 133.725 ;
        RECT 149.825 132.815 150.745 133.045 ;
        RECT 151.525 133.045 153.360 133.725 ;
        RECT 151.525 132.815 152.455 133.045 ;
        RECT 153.515 132.815 154.865 133.725 ;
        RECT 154.895 132.915 156.265 133.725 ;
      LAYER nwell ;
        RECT 70.520 129.695 156.460 132.525 ;
      LAYER pwell ;
        RECT 70.715 128.495 72.085 129.305 ;
        RECT 72.095 128.495 73.925 129.305 ;
        RECT 74.035 128.495 77.145 129.405 ;
        RECT 77.635 128.495 78.985 129.405 ;
        RECT 79.005 128.495 81.735 129.405 ;
        RECT 81.775 128.495 83.125 129.405 ;
        RECT 83.605 128.580 84.035 129.365 ;
        RECT 85.425 129.175 86.345 129.405 ;
        RECT 84.055 128.495 86.345 129.175 ;
        RECT 86.355 128.495 89.565 129.405 ;
        RECT 91.650 129.175 92.785 129.405 ;
        RECT 89.575 128.495 92.785 129.175 ;
        RECT 92.875 128.495 95.875 129.405 ;
        RECT 96.015 128.495 97.845 129.305 ;
        RECT 98.395 128.495 101.395 129.405 ;
        RECT 101.825 128.495 104.745 129.405 ;
        RECT 105.415 129.175 109.345 129.405 ;
        RECT 104.930 128.495 109.345 129.175 ;
        RECT 109.365 128.580 109.795 129.365 ;
        RECT 111.395 129.315 112.345 129.405 ;
        RECT 109.815 128.495 111.185 129.275 ;
        RECT 111.395 128.495 113.325 129.315 ;
        RECT 113.495 128.495 116.245 129.405 ;
        RECT 116.265 128.495 118.995 129.405 ;
        RECT 119.015 128.495 120.385 129.275 ;
        RECT 120.395 128.495 121.765 129.275 ;
        RECT 121.775 128.495 123.145 129.275 ;
        RECT 123.615 128.495 124.985 129.275 ;
        RECT 124.995 129.175 128.925 129.405 ;
        RECT 124.995 128.495 129.410 129.175 ;
        RECT 129.595 128.495 130.965 129.275 ;
        RECT 130.975 128.495 134.450 129.405 ;
        RECT 135.125 128.580 135.555 129.365 ;
        RECT 135.865 128.495 138.785 129.405 ;
        RECT 138.805 128.495 140.155 129.405 ;
        RECT 140.195 128.495 141.545 129.405 ;
        RECT 141.555 129.175 142.900 129.405 ;
        RECT 144.535 129.315 145.485 129.405 ;
        RECT 141.555 128.495 143.385 129.175 ;
        RECT 143.555 128.495 145.485 129.315 ;
        RECT 145.695 128.495 149.825 129.405 ;
        RECT 149.835 129.205 150.785 129.405 ;
        RECT 149.835 128.525 153.505 129.205 ;
        RECT 149.835 128.495 150.785 128.525 ;
        RECT 70.855 128.285 71.025 128.495 ;
        RECT 72.235 128.285 72.405 128.495 ;
        RECT 74.075 128.305 74.245 128.495 ;
        RECT 74.535 128.285 74.705 128.475 ;
        RECT 74.990 128.335 75.110 128.445 ;
        RECT 76.375 128.285 76.545 128.475 ;
        RECT 76.835 128.285 77.005 128.475 ;
        RECT 77.290 128.335 77.410 128.445 ;
        RECT 77.750 128.305 77.920 128.495 ;
        RECT 78.215 128.305 78.385 128.475 ;
        RECT 80.510 128.335 80.630 128.445 ;
        RECT 78.220 128.285 78.385 128.305 ;
        RECT 80.975 128.285 81.145 128.475 ;
        RECT 81.435 128.305 81.605 128.495 ;
        RECT 81.890 128.305 82.060 128.495 ;
        RECT 83.270 128.335 83.390 128.445 ;
        RECT 84.195 128.305 84.365 128.495 ;
        RECT 86.490 128.285 86.660 128.475 ;
        RECT 86.960 128.285 87.130 128.475 ;
        RECT 89.265 128.305 89.435 128.495 ;
        RECT 89.715 128.475 89.885 128.495 ;
        RECT 89.715 128.305 89.890 128.475 ;
        RECT 90.185 128.330 90.345 128.440 ;
        RECT 89.720 128.285 89.890 128.305 ;
        RECT 91.095 128.285 91.265 128.475 ;
        RECT 92.935 128.305 93.105 128.495 ;
        RECT 94.310 128.335 94.430 128.445 ;
        RECT 95.695 128.285 95.865 128.475 ;
        RECT 96.155 128.445 96.325 128.495 ;
        RECT 96.150 128.335 96.325 128.445 ;
        RECT 96.155 128.305 96.325 128.335 ;
        RECT 97.075 128.285 97.245 128.475 ;
        RECT 97.990 128.335 98.110 128.445 ;
        RECT 98.455 128.305 98.625 128.495 ;
        RECT 104.430 128.475 104.600 128.495 ;
        RECT 104.930 128.475 105.040 128.495 ;
        RECT 109.965 128.475 110.135 128.495 ;
        RECT 113.175 128.475 113.325 128.495 ;
        RECT 100.295 128.285 100.465 128.475 ;
        RECT 102.595 128.285 102.765 128.475 ;
        RECT 103.980 128.285 104.150 128.475 ;
        RECT 104.430 128.305 104.605 128.475 ;
        RECT 104.870 128.305 105.040 128.475 ;
        RECT 104.435 128.285 104.605 128.305 ;
        RECT 109.495 128.285 109.665 128.475 ;
        RECT 109.955 128.305 110.135 128.475 ;
        RECT 111.790 128.335 111.910 128.445 ;
        RECT 109.955 128.285 110.125 128.305 ;
        RECT 112.255 128.285 112.425 128.475 ;
        RECT 113.175 128.305 113.345 128.475 ;
        RECT 113.635 128.305 113.805 128.495 ;
        RECT 115.020 128.285 115.190 128.475 ;
        RECT 118.695 128.285 118.865 128.495 ;
        RECT 120.065 128.305 120.235 128.495 ;
        RECT 121.445 128.305 121.615 128.495 ;
        RECT 121.910 128.335 122.030 128.445 ;
        RECT 122.825 128.305 122.995 128.495 ;
        RECT 123.290 128.335 123.410 128.445 ;
        RECT 124.665 128.305 124.835 128.495 ;
        RECT 129.300 128.475 129.410 128.495 ;
        RECT 125.135 128.285 125.305 128.475 ;
        RECT 127.895 128.285 128.065 128.475 ;
        RECT 129.300 128.305 129.470 128.475 ;
        RECT 129.735 128.305 129.905 128.495 ;
        RECT 131.120 128.475 131.290 128.495 ;
        RECT 130.655 128.285 130.825 128.475 ;
        RECT 131.115 128.305 131.290 128.475 ;
        RECT 131.115 128.285 131.285 128.305 ;
        RECT 133.875 128.285 134.045 128.475 ;
        RECT 134.790 128.335 134.910 128.445 ;
        RECT 136.635 128.285 136.805 128.475 ;
        RECT 138.470 128.305 138.640 128.495 ;
        RECT 139.855 128.305 140.025 128.495 ;
        RECT 141.230 128.305 141.400 128.495 ;
        RECT 141.695 128.285 141.865 128.475 ;
        RECT 142.155 128.285 142.325 128.475 ;
        RECT 143.075 128.305 143.245 128.495 ;
        RECT 143.555 128.475 143.705 128.495 ;
        RECT 143.535 128.305 143.705 128.475 ;
        RECT 143.995 128.285 144.165 128.475 ;
        RECT 145.840 128.305 146.010 128.495 ;
        RECT 153.190 128.475 153.360 128.525 ;
        RECT 153.515 128.495 154.865 129.405 ;
        RECT 154.895 128.495 156.265 129.305 ;
        RECT 153.660 128.475 153.830 128.495 ;
        RECT 147.225 128.330 147.385 128.440 ;
        RECT 148.595 128.285 148.765 128.475 ;
        RECT 153.190 128.305 153.365 128.475 ;
        RECT 153.655 128.305 153.830 128.475 ;
        RECT 153.195 128.285 153.360 128.305 ;
        RECT 153.655 128.285 153.825 128.305 ;
        RECT 155.955 128.285 156.125 128.495 ;
        RECT 70.715 127.475 72.085 128.285 ;
        RECT 72.095 127.475 73.465 128.285 ;
        RECT 73.475 127.505 74.845 128.285 ;
        RECT 75.315 127.505 76.685 128.285 ;
        RECT 76.695 127.475 78.065 128.285 ;
        RECT 78.220 127.605 80.055 128.285 ;
        RECT 80.835 127.605 83.125 128.285 ;
        RECT 79.125 127.375 80.055 127.605 ;
        RECT 82.205 127.375 83.125 127.605 ;
        RECT 83.885 127.375 86.805 128.285 ;
        RECT 86.815 127.375 88.645 128.285 ;
        RECT 88.655 127.375 90.005 128.285 ;
        RECT 90.995 127.375 94.165 128.285 ;
        RECT 94.635 127.505 96.005 128.285 ;
        RECT 96.485 127.415 96.915 128.200 ;
        RECT 97.015 127.375 100.015 128.285 ;
        RECT 100.155 127.505 101.525 128.285 ;
        RECT 101.535 127.505 102.905 128.285 ;
        RECT 102.915 127.375 104.265 128.285 ;
        RECT 104.295 127.375 107.045 128.285 ;
        RECT 107.055 127.375 109.805 128.285 ;
        RECT 109.815 127.475 111.645 128.285 ;
        RECT 112.115 127.375 114.865 128.285 ;
        RECT 114.875 127.375 118.350 128.285 ;
        RECT 118.635 127.375 121.635 128.285 ;
        RECT 122.245 127.415 122.675 128.200 ;
        RECT 122.695 127.375 125.445 128.285 ;
        RECT 125.465 127.605 128.205 128.285 ;
        RECT 128.215 127.375 130.965 128.285 ;
        RECT 130.975 127.375 133.725 128.285 ;
        RECT 133.735 127.375 136.485 128.285 ;
        RECT 136.495 127.375 139.245 128.285 ;
        RECT 139.255 127.375 142.005 128.285 ;
        RECT 142.015 127.605 143.845 128.285 ;
        RECT 142.500 127.375 143.845 127.605 ;
        RECT 143.955 127.375 147.065 128.285 ;
        RECT 148.005 127.415 148.435 128.200 ;
        RECT 148.455 127.605 151.195 128.285 ;
        RECT 151.525 127.605 153.360 128.285 ;
        RECT 151.525 127.375 152.455 127.605 ;
        RECT 153.515 127.475 154.885 128.285 ;
        RECT 154.895 127.475 156.265 128.285 ;
      LAYER nwell ;
        RECT 70.520 124.255 156.460 127.085 ;
      LAYER pwell ;
        RECT 70.715 123.055 72.085 123.865 ;
        RECT 72.095 123.735 73.440 123.965 ;
        RECT 72.095 123.055 73.925 123.735 ;
        RECT 73.945 123.055 76.685 123.735 ;
        RECT 76.695 123.055 78.525 123.865 ;
        RECT 78.995 123.055 80.825 123.965 ;
        RECT 80.835 123.735 82.180 123.965 ;
        RECT 80.835 123.055 82.665 123.735 ;
        RECT 83.605 123.140 84.035 123.925 ;
        RECT 84.055 123.735 85.400 123.965 ;
        RECT 85.895 123.735 87.240 123.965 ;
        RECT 84.055 123.055 85.885 123.735 ;
        RECT 85.895 123.055 87.725 123.735 ;
        RECT 87.735 123.055 89.565 123.865 ;
        RECT 89.575 123.735 90.920 123.965 ;
        RECT 89.575 123.055 91.405 123.735 ;
        RECT 91.415 123.055 93.245 123.865 ;
        RECT 93.255 123.735 94.600 123.965 ;
        RECT 93.255 123.055 95.085 123.735 ;
        RECT 95.095 123.055 96.465 123.865 ;
        RECT 96.485 123.140 96.915 123.925 ;
        RECT 96.935 123.735 98.280 123.965 ;
        RECT 96.935 123.055 98.765 123.735 ;
        RECT 98.775 123.055 100.605 123.865 ;
        RECT 100.615 123.735 101.960 123.965 ;
        RECT 100.615 123.055 102.445 123.735 ;
        RECT 102.455 123.055 104.285 123.865 ;
        RECT 104.780 123.735 106.125 123.965 ;
        RECT 104.295 123.055 106.125 123.735 ;
        RECT 106.135 123.055 107.505 123.865 ;
        RECT 107.515 123.735 108.860 123.965 ;
        RECT 107.515 123.055 109.345 123.735 ;
        RECT 109.365 123.140 109.795 123.925 ;
        RECT 109.815 123.055 112.555 123.735 ;
        RECT 112.575 123.055 113.945 123.865 ;
        RECT 113.965 123.055 116.705 123.735 ;
        RECT 116.715 123.055 119.465 123.965 ;
        RECT 119.475 123.055 122.215 123.735 ;
        RECT 122.245 123.140 122.675 123.925 ;
        RECT 122.695 123.055 125.445 123.965 ;
        RECT 126.115 123.875 127.065 123.965 ;
        RECT 126.115 123.055 128.045 123.875 ;
        RECT 128.225 123.055 130.965 123.735 ;
        RECT 131.435 123.055 134.185 123.965 ;
        RECT 135.125 123.140 135.555 123.925 ;
        RECT 135.575 123.055 138.315 123.735 ;
        RECT 139.255 123.055 142.005 123.965 ;
        RECT 142.015 123.055 144.765 123.965 ;
        RECT 144.775 123.055 147.515 123.735 ;
        RECT 148.005 123.140 148.435 123.925 ;
        RECT 152.355 123.875 153.305 123.965 ;
        RECT 148.455 123.055 151.195 123.735 ;
        RECT 151.375 123.055 153.305 123.875 ;
        RECT 153.515 123.055 154.885 123.865 ;
        RECT 154.895 123.055 156.265 123.865 ;
        RECT 70.855 122.865 71.025 123.055 ;
        RECT 73.615 122.865 73.785 123.055 ;
        RECT 76.375 122.865 76.545 123.055 ;
        RECT 76.835 122.865 77.005 123.055 ;
        RECT 78.670 122.895 78.790 123.005 ;
        RECT 79.140 122.865 79.310 123.055 ;
        RECT 82.355 122.865 82.525 123.055 ;
        RECT 82.825 122.900 82.985 123.010 ;
        RECT 85.575 122.865 85.745 123.055 ;
        RECT 87.415 122.865 87.585 123.055 ;
        RECT 87.875 122.865 88.045 123.055 ;
        RECT 91.095 122.865 91.265 123.055 ;
        RECT 91.555 122.865 91.725 123.055 ;
        RECT 94.775 122.865 94.945 123.055 ;
        RECT 95.235 122.865 95.405 123.055 ;
        RECT 98.455 122.865 98.625 123.055 ;
        RECT 98.915 122.865 99.085 123.055 ;
        RECT 102.135 122.865 102.305 123.055 ;
        RECT 102.595 122.865 102.765 123.055 ;
        RECT 104.435 122.865 104.605 123.055 ;
        RECT 106.275 122.865 106.445 123.055 ;
        RECT 109.035 122.865 109.205 123.055 ;
        RECT 109.955 122.865 110.125 123.055 ;
        RECT 112.715 122.865 112.885 123.055 ;
        RECT 116.395 122.865 116.565 123.055 ;
        RECT 119.155 122.865 119.325 123.055 ;
        RECT 119.615 122.865 119.785 123.055 ;
        RECT 125.135 122.865 125.305 123.055 ;
        RECT 127.895 123.035 128.045 123.055 ;
        RECT 125.590 122.895 125.710 123.005 ;
        RECT 127.895 122.865 128.065 123.035 ;
        RECT 130.655 122.865 130.825 123.055 ;
        RECT 131.110 122.895 131.230 123.005 ;
        RECT 131.575 122.865 131.745 123.055 ;
        RECT 134.345 122.900 134.505 123.010 ;
        RECT 135.715 122.865 135.885 123.055 ;
        RECT 138.485 122.900 138.645 123.010 ;
        RECT 141.695 122.865 141.865 123.055 ;
        RECT 144.455 122.865 144.625 123.055 ;
        RECT 144.915 122.865 145.085 123.055 ;
        RECT 147.670 122.895 147.790 123.005 ;
        RECT 148.595 122.865 148.765 123.055 ;
        RECT 151.375 123.035 151.525 123.055 ;
        RECT 151.355 122.865 151.525 123.035 ;
        RECT 153.655 122.865 153.825 123.055 ;
        RECT 155.955 122.865 156.125 123.055 ;
        RECT 50.930 58.110 53.280 103.830 ;
        RECT 54.930 58.110 57.280 103.830 ;
        RECT 58.930 58.110 61.280 103.830 ;
        RECT 62.930 58.110 65.280 103.830 ;
        RECT 66.930 58.110 69.280 103.830 ;
        RECT 70.930 58.110 73.280 103.830 ;
        RECT 74.930 58.110 77.280 103.830 ;
        RECT 78.930 58.110 81.280 103.830 ;
        RECT 87.930 58.110 90.280 103.830 ;
        RECT 91.930 58.110 94.280 103.830 ;
        RECT 95.930 58.110 98.280 103.830 ;
        RECT 99.930 58.110 102.280 103.830 ;
        RECT 103.930 58.110 106.280 103.830 ;
        RECT 107.930 58.110 110.280 103.830 ;
        RECT 111.930 58.110 114.280 103.830 ;
        RECT 115.930 58.110 118.280 103.830 ;
        RECT 124.930 58.110 127.280 103.830 ;
        RECT 128.930 58.110 131.280 103.830 ;
        RECT 132.930 58.110 135.280 103.830 ;
        RECT 136.930 58.110 139.280 103.830 ;
        RECT 140.930 58.110 143.280 103.830 ;
        RECT 144.930 58.110 147.280 103.830 ;
        RECT 148.930 58.110 151.280 103.830 ;
        RECT 152.930 58.110 155.280 103.830 ;
        RECT 50.930 30.460 53.280 55.830 ;
        RECT 54.930 30.460 57.280 55.830 ;
        RECT 58.930 30.460 61.280 55.830 ;
        RECT 62.930 30.460 65.280 55.830 ;
        RECT 66.930 30.460 69.280 55.830 ;
        RECT 70.930 30.460 73.280 55.830 ;
        RECT 74.930 30.460 77.280 55.830 ;
        RECT 78.930 30.460 81.280 55.830 ;
        RECT 87.930 30.460 90.280 55.830 ;
        RECT 91.930 30.460 94.280 55.830 ;
        RECT 95.930 30.460 98.280 55.830 ;
        RECT 99.930 30.460 102.280 55.830 ;
        RECT 103.930 30.460 106.280 55.830 ;
        RECT 107.930 30.460 110.280 55.830 ;
        RECT 111.930 30.460 114.280 55.830 ;
        RECT 115.930 30.460 118.280 55.830 ;
        RECT 124.930 30.460 127.280 55.830 ;
        RECT 128.930 30.460 131.280 55.830 ;
        RECT 132.930 30.460 135.280 55.830 ;
        RECT 136.930 30.460 139.280 55.830 ;
        RECT 140.930 30.460 143.280 55.830 ;
        RECT 144.930 30.460 147.280 55.830 ;
        RECT 148.930 30.460 151.280 55.830 ;
        RECT 152.930 30.460 155.280 55.830 ;
      LAYER nwell ;
        RECT 31.105 16.780 33.215 26.970 ;
      LAYER pwell ;
        RECT 33.920 18.845 36.030 24.945 ;
      LAYER li1 ;
        RECT 70.710 207.185 156.270 207.355 ;
        RECT 70.795 206.095 72.005 207.185 ;
        RECT 72.175 206.095 73.385 207.185 ;
        RECT 73.610 206.315 73.895 207.185 ;
        RECT 74.065 206.555 74.325 207.015 ;
        RECT 74.500 206.725 74.755 207.185 ;
        RECT 74.925 206.555 75.185 207.015 ;
        RECT 74.065 206.385 75.185 206.555 ;
        RECT 75.355 206.385 75.665 207.185 ;
        RECT 74.065 206.135 74.325 206.385 ;
        RECT 75.835 206.215 76.145 207.015 ;
        RECT 70.795 205.385 71.315 205.925 ;
        RECT 71.485 205.555 72.005 206.095 ;
        RECT 72.175 205.385 72.695 205.925 ;
        RECT 72.865 205.555 73.385 206.095 ;
        RECT 73.570 205.965 74.325 206.135 ;
        RECT 75.115 206.045 76.145 206.215 ;
        RECT 73.570 205.455 73.975 205.965 ;
        RECT 75.115 205.795 75.285 206.045 ;
        RECT 74.145 205.625 75.285 205.795 ;
        RECT 70.795 204.635 72.005 205.385 ;
        RECT 72.175 204.635 73.385 205.385 ;
        RECT 73.570 205.285 75.220 205.455 ;
        RECT 75.455 205.305 75.805 205.875 ;
        RECT 73.615 204.635 73.895 205.115 ;
        RECT 74.065 204.895 74.325 205.285 ;
        RECT 74.500 204.635 74.755 205.115 ;
        RECT 74.925 204.895 75.220 205.285 ;
        RECT 75.975 205.135 76.145 206.045 ;
        RECT 75.400 204.635 75.675 205.115 ;
        RECT 75.845 204.805 76.145 205.135 ;
        RECT 76.315 206.110 76.585 207.015 ;
        RECT 76.755 206.425 77.085 207.185 ;
        RECT 77.265 206.255 77.435 207.015 ;
        RECT 76.315 205.310 76.485 206.110 ;
        RECT 76.770 206.085 77.435 206.255 ;
        RECT 76.770 205.940 76.940 206.085 ;
        RECT 77.700 206.035 77.960 207.185 ;
        RECT 78.135 206.110 78.390 207.015 ;
        RECT 78.560 206.425 78.890 207.185 ;
        RECT 79.105 206.255 79.275 207.015 ;
        RECT 76.655 205.610 76.940 205.940 ;
        RECT 76.770 205.355 76.940 205.610 ;
        RECT 77.175 205.535 77.505 205.905 ;
        RECT 76.315 204.805 76.575 205.310 ;
        RECT 76.770 205.185 77.435 205.355 ;
        RECT 76.755 204.635 77.085 205.015 ;
        RECT 77.265 204.805 77.435 205.185 ;
        RECT 77.700 204.635 77.960 205.475 ;
        RECT 78.135 205.380 78.305 206.110 ;
        RECT 78.560 206.085 79.275 206.255 ;
        RECT 78.560 205.875 78.730 206.085 ;
        RECT 79.540 206.045 79.875 207.015 ;
        RECT 80.045 206.045 80.215 207.185 ;
        RECT 80.385 206.845 82.415 207.015 ;
        RECT 78.475 205.545 78.730 205.875 ;
        RECT 78.135 204.805 78.390 205.380 ;
        RECT 78.560 205.355 78.730 205.545 ;
        RECT 79.010 205.535 79.365 205.905 ;
        RECT 79.540 205.375 79.710 206.045 ;
        RECT 80.385 205.875 80.555 206.845 ;
        RECT 79.880 205.545 80.135 205.875 ;
        RECT 80.360 205.545 80.555 205.875 ;
        RECT 80.725 206.505 81.850 206.675 ;
        RECT 79.965 205.375 80.135 205.545 ;
        RECT 80.725 205.375 80.895 206.505 ;
        RECT 78.560 205.185 79.275 205.355 ;
        RECT 78.560 204.635 78.890 205.015 ;
        RECT 79.105 204.805 79.275 205.185 ;
        RECT 79.540 204.805 79.795 205.375 ;
        RECT 79.965 205.205 80.895 205.375 ;
        RECT 81.065 206.165 82.075 206.335 ;
        RECT 81.065 205.365 81.235 206.165 ;
        RECT 81.440 205.485 81.715 205.965 ;
        RECT 81.435 205.315 81.715 205.485 ;
        RECT 80.720 205.170 80.895 205.205 ;
        RECT 79.965 204.635 80.295 205.035 ;
        RECT 80.720 204.805 81.250 205.170 ;
        RECT 81.440 204.805 81.715 205.315 ;
        RECT 81.885 204.805 82.075 206.165 ;
        RECT 82.245 206.180 82.415 206.845 ;
        RECT 82.585 206.425 82.755 207.185 ;
        RECT 82.990 206.425 83.505 206.835 ;
        RECT 82.245 205.990 82.995 206.180 ;
        RECT 83.165 205.615 83.505 206.425 ;
        RECT 83.675 206.020 83.965 207.185 ;
        RECT 84.135 206.045 84.520 207.015 ;
        RECT 84.690 206.725 85.015 207.185 ;
        RECT 85.535 206.555 85.815 207.015 ;
        RECT 84.690 206.335 85.815 206.555 ;
        RECT 82.275 205.445 83.505 205.615 ;
        RECT 82.255 204.635 82.765 205.170 ;
        RECT 82.985 204.840 83.230 205.445 ;
        RECT 84.135 205.375 84.415 206.045 ;
        RECT 84.690 205.875 85.140 206.335 ;
        RECT 86.005 206.165 86.405 207.015 ;
        RECT 86.805 206.725 87.075 207.185 ;
        RECT 87.245 206.555 87.530 207.015 ;
        RECT 84.585 205.545 85.140 205.875 ;
        RECT 85.310 205.605 86.405 206.165 ;
        RECT 84.690 205.435 85.140 205.545 ;
        RECT 83.675 204.635 83.965 205.360 ;
        RECT 84.135 204.805 84.520 205.375 ;
        RECT 84.690 205.265 85.815 205.435 ;
        RECT 84.690 204.635 85.015 205.095 ;
        RECT 85.535 204.805 85.815 205.265 ;
        RECT 86.005 204.805 86.405 205.605 ;
        RECT 86.575 206.335 87.530 206.555 ;
        RECT 86.575 205.435 86.785 206.335 ;
        RECT 86.955 205.605 87.645 206.165 ;
        RECT 87.820 206.035 88.080 207.185 ;
        RECT 88.255 206.110 88.510 207.015 ;
        RECT 88.680 206.425 89.010 207.185 ;
        RECT 89.225 206.255 89.395 207.015 ;
        RECT 86.575 205.265 87.530 205.435 ;
        RECT 86.805 204.635 87.075 205.095 ;
        RECT 87.245 204.805 87.530 205.265 ;
        RECT 87.820 204.635 88.080 205.475 ;
        RECT 88.255 205.380 88.425 206.110 ;
        RECT 88.680 206.085 89.395 206.255 ;
        RECT 89.655 206.095 90.865 207.185 ;
        RECT 88.680 205.875 88.850 206.085 ;
        RECT 88.595 205.545 88.850 205.875 ;
        RECT 88.255 204.805 88.510 205.380 ;
        RECT 88.680 205.355 88.850 205.545 ;
        RECT 89.130 205.535 89.485 205.905 ;
        RECT 89.655 205.385 90.175 205.925 ;
        RECT 90.345 205.555 90.865 206.095 ;
        RECT 91.040 206.035 91.300 207.185 ;
        RECT 91.475 206.110 91.730 207.015 ;
        RECT 91.900 206.425 92.230 207.185 ;
        RECT 92.445 206.255 92.615 207.015 ;
        RECT 88.680 205.185 89.395 205.355 ;
        RECT 88.680 204.635 89.010 205.015 ;
        RECT 89.225 204.805 89.395 205.185 ;
        RECT 89.655 204.635 90.865 205.385 ;
        RECT 91.040 204.635 91.300 205.475 ;
        RECT 91.475 205.380 91.645 206.110 ;
        RECT 91.900 206.085 92.615 206.255 ;
        RECT 92.875 206.215 93.185 207.015 ;
        RECT 93.355 206.385 93.665 207.185 ;
        RECT 93.835 206.555 94.095 207.015 ;
        RECT 94.265 206.725 94.520 207.185 ;
        RECT 94.695 206.555 94.955 207.015 ;
        RECT 93.835 206.385 94.955 206.555 ;
        RECT 94.315 206.335 94.485 206.385 ;
        RECT 91.900 205.875 92.070 206.085 ;
        RECT 92.875 206.045 93.905 206.215 ;
        RECT 91.815 205.545 92.070 205.875 ;
        RECT 91.475 204.805 91.730 205.380 ;
        RECT 91.900 205.355 92.070 205.545 ;
        RECT 92.350 205.535 92.705 205.905 ;
        RECT 91.900 205.185 92.615 205.355 ;
        RECT 91.900 204.635 92.230 205.015 ;
        RECT 92.445 204.805 92.615 205.185 ;
        RECT 92.875 205.135 93.045 206.045 ;
        RECT 93.215 205.305 93.565 205.875 ;
        RECT 93.735 205.795 93.905 206.045 ;
        RECT 94.695 206.135 94.955 206.385 ;
        RECT 95.125 206.315 95.410 207.185 ;
        RECT 94.695 205.965 95.450 206.135 ;
        RECT 96.555 206.020 96.845 207.185 ;
        RECT 97.070 206.315 97.355 207.185 ;
        RECT 97.525 206.555 97.785 207.015 ;
        RECT 97.960 206.725 98.215 207.185 ;
        RECT 98.385 206.555 98.645 207.015 ;
        RECT 97.525 206.385 98.645 206.555 ;
        RECT 98.815 206.385 99.125 207.185 ;
        RECT 97.525 206.135 97.785 206.385 ;
        RECT 99.295 206.215 99.605 207.015 ;
        RECT 93.735 205.625 94.875 205.795 ;
        RECT 95.045 205.455 95.450 205.965 ;
        RECT 93.800 205.285 95.450 205.455 ;
        RECT 97.030 205.965 97.785 206.135 ;
        RECT 98.575 206.045 99.605 206.215 ;
        RECT 100.705 206.235 100.980 207.005 ;
        RECT 101.150 206.575 101.480 207.005 ;
        RECT 101.650 206.745 101.845 207.185 ;
        RECT 102.025 206.575 102.355 207.005 ;
        RECT 101.150 206.405 102.355 206.575 ;
        RECT 100.705 206.045 101.290 206.235 ;
        RECT 101.460 206.075 102.355 206.405 ;
        RECT 103.545 206.255 103.715 207.015 ;
        RECT 103.930 206.425 104.260 207.185 ;
        RECT 103.545 206.085 104.260 206.255 ;
        RECT 104.430 206.110 104.685 207.015 ;
        RECT 97.030 205.455 97.435 205.965 ;
        RECT 98.575 205.795 98.745 206.045 ;
        RECT 97.605 205.625 98.745 205.795 ;
        RECT 92.875 204.805 93.175 205.135 ;
        RECT 93.345 204.635 93.620 205.115 ;
        RECT 93.800 204.895 94.095 205.285 ;
        RECT 94.265 204.635 94.520 205.115 ;
        RECT 94.695 204.895 94.955 205.285 ;
        RECT 95.125 204.635 95.405 205.115 ;
        RECT 96.555 204.635 96.845 205.360 ;
        RECT 97.030 205.285 98.680 205.455 ;
        RECT 98.915 205.305 99.265 205.875 ;
        RECT 97.075 204.635 97.355 205.115 ;
        RECT 97.525 204.895 97.785 205.285 ;
        RECT 97.960 204.635 98.215 205.115 ;
        RECT 98.385 204.895 98.680 205.285 ;
        RECT 99.435 205.135 99.605 206.045 ;
        RECT 100.705 205.225 100.945 205.875 ;
        RECT 101.115 205.375 101.290 206.045 ;
        RECT 101.460 205.545 101.875 205.875 ;
        RECT 102.055 205.545 102.350 205.875 ;
        RECT 101.115 205.195 101.445 205.375 ;
        RECT 98.860 204.635 99.135 205.115 ;
        RECT 99.305 204.805 99.605 205.135 ;
        RECT 100.720 204.635 101.050 205.025 ;
        RECT 101.220 204.815 101.445 205.195 ;
        RECT 101.645 204.925 101.875 205.545 ;
        RECT 103.455 205.535 103.810 205.905 ;
        RECT 104.090 205.875 104.260 206.085 ;
        RECT 104.090 205.545 104.345 205.875 ;
        RECT 102.055 204.635 102.355 205.365 ;
        RECT 104.090 205.355 104.260 205.545 ;
        RECT 104.515 205.380 104.685 206.110 ;
        RECT 104.860 206.035 105.120 207.185 ;
        RECT 105.385 206.255 105.555 207.015 ;
        RECT 105.770 206.425 106.100 207.185 ;
        RECT 105.385 206.085 106.100 206.255 ;
        RECT 106.270 206.110 106.525 207.015 ;
        RECT 105.295 205.535 105.650 205.905 ;
        RECT 105.930 205.875 106.100 206.085 ;
        RECT 105.930 205.545 106.185 205.875 ;
        RECT 103.545 205.185 104.260 205.355 ;
        RECT 103.545 204.805 103.715 205.185 ;
        RECT 103.930 204.635 104.260 205.015 ;
        RECT 104.430 204.805 104.685 205.380 ;
        RECT 104.860 204.635 105.120 205.475 ;
        RECT 105.930 205.355 106.100 205.545 ;
        RECT 106.355 205.380 106.525 206.110 ;
        RECT 106.700 206.035 106.960 207.185 ;
        RECT 107.685 206.255 107.855 207.015 ;
        RECT 108.070 206.425 108.400 207.185 ;
        RECT 107.685 206.085 108.400 206.255 ;
        RECT 108.570 206.110 108.825 207.015 ;
        RECT 107.595 205.535 107.950 205.905 ;
        RECT 108.230 205.875 108.400 206.085 ;
        RECT 108.230 205.545 108.485 205.875 ;
        RECT 105.385 205.185 106.100 205.355 ;
        RECT 105.385 204.805 105.555 205.185 ;
        RECT 105.770 204.635 106.100 205.015 ;
        RECT 106.270 204.805 106.525 205.380 ;
        RECT 106.700 204.635 106.960 205.475 ;
        RECT 108.230 205.355 108.400 205.545 ;
        RECT 108.655 205.380 108.825 206.110 ;
        RECT 109.000 206.035 109.260 207.185 ;
        RECT 109.435 206.020 109.725 207.185 ;
        RECT 109.955 206.045 110.165 207.185 ;
        RECT 110.335 206.035 110.665 207.015 ;
        RECT 110.835 206.045 111.065 207.185 ;
        RECT 111.740 206.035 112.000 207.185 ;
        RECT 112.175 206.110 112.430 207.015 ;
        RECT 112.600 206.425 112.930 207.185 ;
        RECT 113.145 206.255 113.315 207.015 ;
        RECT 107.685 205.185 108.400 205.355 ;
        RECT 107.685 204.805 107.855 205.185 ;
        RECT 108.070 204.635 108.400 205.015 ;
        RECT 108.570 204.805 108.825 205.380 ;
        RECT 109.000 204.635 109.260 205.475 ;
        RECT 109.435 204.635 109.725 205.360 ;
        RECT 109.955 204.635 110.165 205.455 ;
        RECT 110.335 205.435 110.585 206.035 ;
        RECT 110.755 205.625 111.085 205.875 ;
        RECT 110.335 204.805 110.665 205.435 ;
        RECT 110.835 204.635 111.065 205.455 ;
        RECT 111.740 204.635 112.000 205.475 ;
        RECT 112.175 205.380 112.345 206.110 ;
        RECT 112.600 206.085 113.315 206.255 ;
        RECT 113.665 206.255 113.835 207.015 ;
        RECT 114.015 206.425 114.345 207.185 ;
        RECT 113.665 206.085 114.330 206.255 ;
        RECT 114.515 206.110 114.785 207.015 ;
        RECT 112.600 205.875 112.770 206.085 ;
        RECT 114.160 205.940 114.330 206.085 ;
        RECT 112.515 205.545 112.770 205.875 ;
        RECT 112.175 204.805 112.430 205.380 ;
        RECT 112.600 205.355 112.770 205.545 ;
        RECT 113.050 205.535 113.405 205.905 ;
        RECT 113.595 205.535 113.925 205.905 ;
        RECT 114.160 205.610 114.445 205.940 ;
        RECT 114.160 205.355 114.330 205.610 ;
        RECT 112.600 205.185 113.315 205.355 ;
        RECT 112.600 204.635 112.930 205.015 ;
        RECT 113.145 204.805 113.315 205.185 ;
        RECT 113.665 205.185 114.330 205.355 ;
        RECT 114.615 205.310 114.785 206.110 ;
        RECT 113.665 204.805 113.835 205.185 ;
        RECT 114.015 204.635 114.345 205.015 ;
        RECT 114.525 204.805 114.785 205.310 ;
        RECT 115.875 206.110 116.145 207.015 ;
        RECT 116.315 206.425 116.645 207.185 ;
        RECT 116.825 206.255 116.995 207.015 ;
        RECT 115.875 205.310 116.045 206.110 ;
        RECT 116.330 206.085 116.995 206.255 ;
        RECT 117.345 206.255 117.515 207.015 ;
        RECT 117.695 206.425 118.025 207.185 ;
        RECT 117.345 206.085 118.010 206.255 ;
        RECT 118.195 206.110 118.465 207.015 ;
        RECT 116.330 205.940 116.500 206.085 ;
        RECT 116.215 205.610 116.500 205.940 ;
        RECT 117.840 205.940 118.010 206.085 ;
        RECT 116.330 205.355 116.500 205.610 ;
        RECT 116.735 205.535 117.065 205.905 ;
        RECT 117.275 205.535 117.605 205.905 ;
        RECT 117.840 205.610 118.125 205.940 ;
        RECT 117.840 205.355 118.010 205.610 ;
        RECT 115.875 204.805 116.135 205.310 ;
        RECT 116.330 205.185 116.995 205.355 ;
        RECT 116.315 204.635 116.645 205.015 ;
        RECT 116.825 204.805 116.995 205.185 ;
        RECT 117.345 205.185 118.010 205.355 ;
        RECT 118.295 205.310 118.465 206.110 ;
        RECT 117.345 204.805 117.515 205.185 ;
        RECT 117.695 204.635 118.025 205.015 ;
        RECT 118.205 204.805 118.465 205.310 ;
        RECT 118.635 206.045 119.020 207.015 ;
        RECT 119.190 206.725 119.515 207.185 ;
        RECT 120.035 206.555 120.315 207.015 ;
        RECT 119.190 206.335 120.315 206.555 ;
        RECT 118.635 205.375 118.915 206.045 ;
        RECT 119.190 205.875 119.640 206.335 ;
        RECT 120.505 206.165 120.905 207.015 ;
        RECT 121.305 206.725 121.575 207.185 ;
        RECT 121.745 206.555 122.030 207.015 ;
        RECT 119.085 205.545 119.640 205.875 ;
        RECT 119.810 205.605 120.905 206.165 ;
        RECT 119.190 205.435 119.640 205.545 ;
        RECT 118.635 204.805 119.020 205.375 ;
        RECT 119.190 205.265 120.315 205.435 ;
        RECT 119.190 204.635 119.515 205.095 ;
        RECT 120.035 204.805 120.315 205.265 ;
        RECT 120.505 204.805 120.905 205.605 ;
        RECT 121.075 206.335 122.030 206.555 ;
        RECT 121.075 205.435 121.285 206.335 ;
        RECT 121.455 205.605 122.145 206.165 ;
        RECT 122.315 206.020 122.605 207.185 ;
        RECT 123.240 206.045 123.575 207.015 ;
        RECT 123.745 206.045 123.915 207.185 ;
        RECT 124.085 206.845 126.115 207.015 ;
        RECT 121.075 205.265 122.030 205.435 ;
        RECT 123.240 205.375 123.410 206.045 ;
        RECT 124.085 205.875 124.255 206.845 ;
        RECT 123.580 205.545 123.835 205.875 ;
        RECT 124.060 205.545 124.255 205.875 ;
        RECT 124.425 206.505 125.550 206.675 ;
        RECT 123.665 205.375 123.835 205.545 ;
        RECT 124.425 205.375 124.595 206.505 ;
        RECT 121.305 204.635 121.575 205.095 ;
        RECT 121.745 204.805 122.030 205.265 ;
        RECT 122.315 204.635 122.605 205.360 ;
        RECT 123.240 204.805 123.495 205.375 ;
        RECT 123.665 205.205 124.595 205.375 ;
        RECT 124.765 206.165 125.775 206.335 ;
        RECT 124.765 205.365 124.935 206.165 ;
        RECT 125.140 205.825 125.415 205.965 ;
        RECT 125.135 205.655 125.415 205.825 ;
        RECT 124.420 205.170 124.595 205.205 ;
        RECT 123.665 204.635 123.995 205.035 ;
        RECT 124.420 204.805 124.950 205.170 ;
        RECT 125.140 204.805 125.415 205.655 ;
        RECT 125.585 204.805 125.775 206.165 ;
        RECT 125.945 206.180 126.115 206.845 ;
        RECT 126.285 206.425 126.455 207.185 ;
        RECT 126.690 206.425 127.205 206.835 ;
        RECT 125.945 205.990 126.695 206.180 ;
        RECT 126.865 205.615 127.205 206.425 ;
        RECT 125.975 205.445 127.205 205.615 ;
        RECT 127.380 206.045 127.715 207.015 ;
        RECT 127.885 206.045 128.055 207.185 ;
        RECT 128.225 206.845 130.255 207.015 ;
        RECT 125.955 204.635 126.465 205.170 ;
        RECT 126.685 204.840 126.930 205.445 ;
        RECT 127.380 205.375 127.550 206.045 ;
        RECT 128.225 205.875 128.395 206.845 ;
        RECT 127.720 205.545 127.975 205.875 ;
        RECT 128.200 205.545 128.395 205.875 ;
        RECT 128.565 206.505 129.690 206.675 ;
        RECT 127.805 205.375 127.975 205.545 ;
        RECT 128.565 205.375 128.735 206.505 ;
        RECT 127.380 204.805 127.635 205.375 ;
        RECT 127.805 205.205 128.735 205.375 ;
        RECT 128.905 206.165 129.915 206.335 ;
        RECT 128.905 205.365 129.075 206.165 ;
        RECT 129.280 205.485 129.555 205.965 ;
        RECT 129.275 205.315 129.555 205.485 ;
        RECT 128.560 205.170 128.735 205.205 ;
        RECT 127.805 204.635 128.135 205.035 ;
        RECT 128.560 204.805 129.090 205.170 ;
        RECT 129.280 204.805 129.555 205.315 ;
        RECT 129.725 204.805 129.915 206.165 ;
        RECT 130.085 206.180 130.255 206.845 ;
        RECT 130.425 206.425 130.595 207.185 ;
        RECT 130.830 206.425 131.345 206.835 ;
        RECT 130.085 205.990 130.835 206.180 ;
        RECT 131.005 205.615 131.345 206.425 ;
        RECT 130.115 205.445 131.345 205.615 ;
        RECT 131.515 206.045 131.900 207.015 ;
        RECT 132.070 206.725 132.395 207.185 ;
        RECT 132.915 206.555 133.195 207.015 ;
        RECT 132.070 206.335 133.195 206.555 ;
        RECT 130.095 204.635 130.605 205.170 ;
        RECT 130.825 204.840 131.070 205.445 ;
        RECT 131.515 205.375 131.795 206.045 ;
        RECT 132.070 205.875 132.520 206.335 ;
        RECT 133.385 206.165 133.785 207.015 ;
        RECT 134.185 206.725 134.455 207.185 ;
        RECT 134.625 206.555 134.910 207.015 ;
        RECT 131.965 205.545 132.520 205.875 ;
        RECT 132.690 205.605 133.785 206.165 ;
        RECT 132.070 205.435 132.520 205.545 ;
        RECT 131.515 204.805 131.900 205.375 ;
        RECT 132.070 205.265 133.195 205.435 ;
        RECT 132.070 204.635 132.395 205.095 ;
        RECT 132.915 204.805 133.195 205.265 ;
        RECT 133.385 204.805 133.785 205.605 ;
        RECT 133.955 206.335 134.910 206.555 ;
        RECT 133.955 205.435 134.165 206.335 ;
        RECT 134.335 205.605 135.025 206.165 ;
        RECT 135.195 206.020 135.485 207.185 ;
        RECT 135.655 206.110 135.925 207.015 ;
        RECT 136.095 206.425 136.425 207.185 ;
        RECT 136.605 206.255 136.775 207.015 ;
        RECT 133.955 205.265 134.910 205.435 ;
        RECT 134.185 204.635 134.455 205.095 ;
        RECT 134.625 204.805 134.910 205.265 ;
        RECT 135.195 204.635 135.485 205.360 ;
        RECT 135.655 205.310 135.825 206.110 ;
        RECT 136.110 206.085 136.775 206.255 ;
        RECT 137.035 206.110 137.305 207.015 ;
        RECT 137.475 206.425 137.805 207.185 ;
        RECT 137.985 206.255 138.155 207.015 ;
        RECT 136.110 205.940 136.280 206.085 ;
        RECT 135.995 205.610 136.280 205.940 ;
        RECT 136.110 205.355 136.280 205.610 ;
        RECT 136.515 205.535 136.845 205.905 ;
        RECT 135.655 204.805 135.915 205.310 ;
        RECT 136.110 205.185 136.775 205.355 ;
        RECT 136.095 204.635 136.425 205.015 ;
        RECT 136.605 204.805 136.775 205.185 ;
        RECT 137.035 205.310 137.205 206.110 ;
        RECT 137.490 206.085 138.155 206.255 ;
        RECT 138.415 206.110 138.685 207.015 ;
        RECT 138.855 206.425 139.185 207.185 ;
        RECT 139.365 206.255 139.535 207.015 ;
        RECT 140.805 206.515 140.975 207.015 ;
        RECT 141.145 206.685 141.475 207.185 ;
        RECT 140.805 206.345 141.470 206.515 ;
        RECT 137.490 205.940 137.660 206.085 ;
        RECT 137.375 205.610 137.660 205.940 ;
        RECT 137.490 205.355 137.660 205.610 ;
        RECT 137.895 205.535 138.225 205.905 ;
        RECT 137.035 204.805 137.295 205.310 ;
        RECT 137.490 205.185 138.155 205.355 ;
        RECT 137.475 204.635 137.805 205.015 ;
        RECT 137.985 204.805 138.155 205.185 ;
        RECT 138.415 205.310 138.585 206.110 ;
        RECT 138.870 206.085 139.535 206.255 ;
        RECT 138.870 205.940 139.040 206.085 ;
        RECT 138.755 205.610 139.040 205.940 ;
        RECT 138.870 205.355 139.040 205.610 ;
        RECT 139.275 205.535 139.605 205.905 ;
        RECT 140.720 205.525 141.070 206.175 ;
        RECT 141.240 205.355 141.470 206.345 ;
        RECT 138.415 204.805 138.675 205.310 ;
        RECT 138.870 205.185 139.535 205.355 ;
        RECT 138.855 204.635 139.185 205.015 ;
        RECT 139.365 204.805 139.535 205.185 ;
        RECT 140.805 205.185 141.470 205.355 ;
        RECT 140.805 204.895 140.975 205.185 ;
        RECT 141.145 204.635 141.475 205.015 ;
        RECT 141.645 204.895 141.830 207.015 ;
        RECT 142.070 206.725 142.335 207.185 ;
        RECT 142.505 206.590 142.755 207.015 ;
        RECT 142.965 206.740 144.070 206.910 ;
        RECT 142.450 206.460 142.755 206.590 ;
        RECT 142.000 205.265 142.280 206.215 ;
        RECT 142.450 205.355 142.620 206.460 ;
        RECT 142.790 205.675 143.030 206.270 ;
        RECT 143.200 206.205 143.730 206.570 ;
        RECT 143.200 205.505 143.370 206.205 ;
        RECT 143.900 206.125 144.070 206.740 ;
        RECT 144.240 206.385 144.410 207.185 ;
        RECT 144.580 206.685 144.830 207.015 ;
        RECT 145.055 206.715 145.940 206.885 ;
        RECT 143.900 206.035 144.410 206.125 ;
        RECT 142.450 205.225 142.675 205.355 ;
        RECT 142.845 205.285 143.370 205.505 ;
        RECT 143.540 205.865 144.410 206.035 ;
        RECT 142.085 204.635 142.335 205.095 ;
        RECT 142.505 205.085 142.675 205.225 ;
        RECT 143.540 205.085 143.710 205.865 ;
        RECT 144.240 205.795 144.410 205.865 ;
        RECT 143.920 205.615 144.120 205.645 ;
        RECT 144.580 205.615 144.750 206.685 ;
        RECT 144.920 205.795 145.110 206.515 ;
        RECT 143.920 205.315 144.750 205.615 ;
        RECT 145.280 205.585 145.600 206.545 ;
        RECT 142.505 204.915 142.840 205.085 ;
        RECT 143.035 204.915 143.710 205.085 ;
        RECT 144.030 204.635 144.400 205.135 ;
        RECT 144.580 205.085 144.750 205.315 ;
        RECT 145.135 205.255 145.600 205.585 ;
        RECT 145.770 205.875 145.940 206.715 ;
        RECT 146.120 206.685 146.435 207.185 ;
        RECT 146.665 206.455 147.005 207.015 ;
        RECT 146.110 206.080 147.005 206.455 ;
        RECT 147.175 206.175 147.345 207.185 ;
        RECT 146.815 205.875 147.005 206.080 ;
        RECT 147.515 206.125 147.845 206.970 ;
        RECT 147.515 206.045 147.905 206.125 ;
        RECT 147.690 205.995 147.905 206.045 ;
        RECT 148.075 206.020 148.365 207.185 ;
        RECT 148.995 206.590 149.430 207.015 ;
        RECT 149.600 206.760 149.985 207.185 ;
        RECT 148.995 206.420 149.985 206.590 ;
        RECT 145.770 205.545 146.645 205.875 ;
        RECT 146.815 205.545 147.565 205.875 ;
        RECT 145.770 205.085 145.940 205.545 ;
        RECT 146.815 205.375 147.015 205.545 ;
        RECT 147.735 205.415 147.905 205.995 ;
        RECT 148.995 205.545 149.480 206.250 ;
        RECT 149.650 205.875 149.985 206.420 ;
        RECT 150.155 206.225 150.580 207.015 ;
        RECT 150.750 206.590 151.025 207.015 ;
        RECT 151.195 206.760 151.580 207.185 ;
        RECT 150.750 206.395 151.580 206.590 ;
        RECT 150.155 206.045 151.060 206.225 ;
        RECT 149.650 205.545 150.060 205.875 ;
        RECT 150.230 205.545 151.060 206.045 ;
        RECT 151.230 205.875 151.580 206.395 ;
        RECT 151.750 206.225 151.995 207.015 ;
        RECT 152.185 206.590 152.440 207.015 ;
        RECT 152.610 206.760 152.995 207.185 ;
        RECT 152.185 206.395 152.995 206.590 ;
        RECT 151.750 206.045 152.475 206.225 ;
        RECT 151.230 205.545 151.655 205.875 ;
        RECT 151.825 205.545 152.475 206.045 ;
        RECT 152.645 205.875 152.995 206.395 ;
        RECT 153.165 206.045 153.425 207.015 ;
        RECT 153.595 206.095 154.805 207.185 ;
        RECT 152.645 205.545 153.070 205.875 ;
        RECT 147.680 205.375 147.905 205.415 ;
        RECT 149.650 205.375 149.985 205.545 ;
        RECT 150.230 205.375 150.580 205.545 ;
        RECT 151.230 205.375 151.580 205.545 ;
        RECT 151.825 205.375 151.995 205.545 ;
        RECT 152.645 205.375 152.995 205.545 ;
        RECT 153.240 205.375 153.425 206.045 ;
        RECT 144.580 204.915 144.985 205.085 ;
        RECT 145.155 204.915 145.940 205.085 ;
        RECT 146.215 204.635 146.425 205.165 ;
        RECT 146.685 204.850 147.015 205.375 ;
        RECT 147.525 205.290 147.905 205.375 ;
        RECT 147.185 204.635 147.355 205.245 ;
        RECT 147.525 204.855 147.855 205.290 ;
        RECT 148.075 204.635 148.365 205.360 ;
        RECT 148.995 205.205 149.985 205.375 ;
        RECT 148.995 204.805 149.430 205.205 ;
        RECT 149.600 204.635 149.985 205.035 ;
        RECT 150.155 204.805 150.580 205.375 ;
        RECT 150.770 205.205 151.580 205.375 ;
        RECT 150.770 204.805 151.025 205.205 ;
        RECT 151.195 204.635 151.580 205.035 ;
        RECT 151.750 204.805 151.995 205.375 ;
        RECT 152.185 205.205 152.995 205.375 ;
        RECT 152.185 204.805 152.440 205.205 ;
        RECT 152.610 204.635 152.995 205.035 ;
        RECT 153.165 204.805 153.425 205.375 ;
        RECT 153.595 205.385 154.115 205.925 ;
        RECT 154.285 205.555 154.805 206.095 ;
        RECT 154.975 206.095 156.185 207.185 ;
        RECT 154.975 205.555 155.495 206.095 ;
        RECT 155.665 205.385 156.185 205.925 ;
        RECT 153.595 204.635 154.805 205.385 ;
        RECT 154.975 204.635 156.185 205.385 ;
        RECT 70.710 204.465 156.270 204.635 ;
        RECT 70.795 203.715 72.005 204.465 ;
        RECT 73.185 203.915 73.355 204.205 ;
        RECT 73.525 204.085 73.855 204.465 ;
        RECT 73.185 203.745 73.850 203.915 ;
        RECT 70.795 203.175 71.315 203.715 ;
        RECT 71.485 203.005 72.005 203.545 ;
        RECT 70.795 201.915 72.005 203.005 ;
        RECT 73.100 202.925 73.450 203.575 ;
        RECT 73.620 202.755 73.850 203.745 ;
        RECT 73.185 202.585 73.850 202.755 ;
        RECT 73.185 202.085 73.355 202.585 ;
        RECT 73.525 201.915 73.855 202.415 ;
        RECT 74.025 202.085 74.210 204.205 ;
        RECT 74.465 204.005 74.715 204.465 ;
        RECT 74.885 204.015 75.220 204.185 ;
        RECT 75.415 204.015 76.090 204.185 ;
        RECT 74.885 203.875 75.055 204.015 ;
        RECT 74.380 202.885 74.660 203.835 ;
        RECT 74.830 203.745 75.055 203.875 ;
        RECT 74.830 202.640 75.000 203.745 ;
        RECT 75.225 203.595 75.750 203.815 ;
        RECT 75.170 202.830 75.410 203.425 ;
        RECT 75.580 202.895 75.750 203.595 ;
        RECT 75.920 203.235 76.090 204.015 ;
        RECT 76.410 203.965 76.780 204.465 ;
        RECT 76.960 204.015 77.365 204.185 ;
        RECT 77.535 204.015 78.320 204.185 ;
        RECT 76.960 203.785 77.130 204.015 ;
        RECT 76.300 203.485 77.130 203.785 ;
        RECT 77.515 203.515 77.980 203.845 ;
        RECT 76.300 203.455 76.500 203.485 ;
        RECT 76.620 203.235 76.790 203.305 ;
        RECT 75.920 203.065 76.790 203.235 ;
        RECT 76.280 202.975 76.790 203.065 ;
        RECT 74.830 202.510 75.135 202.640 ;
        RECT 75.580 202.530 76.110 202.895 ;
        RECT 74.450 201.915 74.715 202.375 ;
        RECT 74.885 202.085 75.135 202.510 ;
        RECT 76.280 202.360 76.450 202.975 ;
        RECT 75.345 202.190 76.450 202.360 ;
        RECT 76.620 201.915 76.790 202.715 ;
        RECT 76.960 202.415 77.130 203.485 ;
        RECT 77.300 202.585 77.490 203.305 ;
        RECT 77.660 202.555 77.980 203.515 ;
        RECT 78.150 203.555 78.320 204.015 ;
        RECT 78.595 203.935 78.805 204.465 ;
        RECT 79.065 203.725 79.395 204.250 ;
        RECT 79.565 203.855 79.735 204.465 ;
        RECT 79.905 203.810 80.235 204.245 ;
        RECT 79.905 203.725 80.285 203.810 ;
        RECT 79.195 203.555 79.395 203.725 ;
        RECT 80.060 203.685 80.285 203.725 ;
        RECT 78.150 203.225 79.025 203.555 ;
        RECT 79.195 203.225 79.945 203.555 ;
        RECT 76.960 202.085 77.210 202.415 ;
        RECT 78.150 202.385 78.320 203.225 ;
        RECT 79.195 203.020 79.385 203.225 ;
        RECT 80.115 203.105 80.285 203.685 ;
        RECT 80.455 203.695 82.125 204.465 ;
        RECT 80.455 203.175 81.205 203.695 ;
        RECT 82.305 203.655 82.575 204.465 ;
        RECT 82.745 203.655 83.075 204.295 ;
        RECT 83.245 203.655 83.485 204.465 ;
        RECT 83.765 203.915 83.935 204.205 ;
        RECT 84.105 204.085 84.435 204.465 ;
        RECT 83.765 203.745 84.430 203.915 ;
        RECT 80.070 203.055 80.285 203.105 ;
        RECT 78.490 202.645 79.385 203.020 ;
        RECT 79.895 202.975 80.285 203.055 ;
        RECT 81.375 203.005 82.125 203.525 ;
        RECT 82.295 203.225 82.645 203.475 ;
        RECT 82.815 203.055 82.985 203.655 ;
        RECT 83.155 203.225 83.505 203.475 ;
        RECT 77.435 202.215 78.320 202.385 ;
        RECT 78.500 201.915 78.815 202.415 ;
        RECT 79.045 202.085 79.385 202.645 ;
        RECT 79.555 201.915 79.725 202.925 ;
        RECT 79.895 202.130 80.225 202.975 ;
        RECT 80.455 201.915 82.125 203.005 ;
        RECT 82.305 201.915 82.635 203.055 ;
        RECT 82.815 202.885 83.495 203.055 ;
        RECT 83.680 202.925 84.030 203.575 ;
        RECT 83.165 202.100 83.495 202.885 ;
        RECT 84.200 202.755 84.430 203.745 ;
        RECT 83.765 202.585 84.430 202.755 ;
        RECT 83.765 202.085 83.935 202.585 ;
        RECT 84.105 201.915 84.435 202.415 ;
        RECT 84.605 202.085 84.790 204.205 ;
        RECT 85.045 204.005 85.295 204.465 ;
        RECT 85.465 204.015 85.800 204.185 ;
        RECT 85.995 204.015 86.670 204.185 ;
        RECT 85.465 203.875 85.635 204.015 ;
        RECT 84.960 202.885 85.240 203.835 ;
        RECT 85.410 203.745 85.635 203.875 ;
        RECT 85.410 202.640 85.580 203.745 ;
        RECT 85.805 203.595 86.330 203.815 ;
        RECT 85.750 202.830 85.990 203.425 ;
        RECT 86.160 202.895 86.330 203.595 ;
        RECT 86.500 203.235 86.670 204.015 ;
        RECT 86.990 203.965 87.360 204.465 ;
        RECT 87.540 204.015 87.945 204.185 ;
        RECT 88.115 204.015 88.900 204.185 ;
        RECT 87.540 203.785 87.710 204.015 ;
        RECT 86.880 203.485 87.710 203.785 ;
        RECT 88.095 203.515 88.560 203.845 ;
        RECT 86.880 203.455 87.080 203.485 ;
        RECT 87.200 203.235 87.370 203.305 ;
        RECT 86.500 203.065 87.370 203.235 ;
        RECT 86.860 202.975 87.370 203.065 ;
        RECT 85.410 202.510 85.715 202.640 ;
        RECT 86.160 202.530 86.690 202.895 ;
        RECT 85.030 201.915 85.295 202.375 ;
        RECT 85.465 202.085 85.715 202.510 ;
        RECT 86.860 202.360 87.030 202.975 ;
        RECT 85.925 202.190 87.030 202.360 ;
        RECT 87.200 201.915 87.370 202.715 ;
        RECT 87.540 202.415 87.710 203.485 ;
        RECT 87.880 202.585 88.070 203.305 ;
        RECT 88.240 202.555 88.560 203.515 ;
        RECT 88.730 203.555 88.900 204.015 ;
        RECT 89.175 203.935 89.385 204.465 ;
        RECT 89.645 203.725 89.975 204.250 ;
        RECT 90.145 203.855 90.315 204.465 ;
        RECT 90.485 203.810 90.815 204.245 ;
        RECT 90.485 203.725 90.865 203.810 ;
        RECT 89.775 203.555 89.975 203.725 ;
        RECT 90.640 203.685 90.865 203.725 ;
        RECT 88.730 203.225 89.605 203.555 ;
        RECT 89.775 203.225 90.525 203.555 ;
        RECT 87.540 202.085 87.790 202.415 ;
        RECT 88.730 202.385 88.900 203.225 ;
        RECT 89.775 203.020 89.965 203.225 ;
        RECT 90.695 203.105 90.865 203.685 ;
        RECT 90.650 203.055 90.865 203.105 ;
        RECT 89.070 202.645 89.965 203.020 ;
        RECT 90.475 202.975 90.865 203.055 ;
        RECT 91.035 203.790 91.295 204.295 ;
        RECT 91.475 204.085 91.805 204.465 ;
        RECT 91.985 203.915 92.155 204.295 ;
        RECT 91.035 202.990 91.205 203.790 ;
        RECT 91.490 203.745 92.155 203.915 ;
        RECT 93.425 203.915 93.595 204.295 ;
        RECT 93.775 204.085 94.105 204.465 ;
        RECT 93.425 203.745 94.090 203.915 ;
        RECT 94.285 203.790 94.545 204.295 ;
        RECT 91.490 203.490 91.660 203.745 ;
        RECT 91.375 203.160 91.660 203.490 ;
        RECT 91.895 203.195 92.225 203.565 ;
        RECT 93.355 203.195 93.695 203.565 ;
        RECT 93.920 203.490 94.090 203.745 ;
        RECT 91.490 203.015 91.660 203.160 ;
        RECT 93.920 203.160 94.195 203.490 ;
        RECT 93.920 203.015 94.090 203.160 ;
        RECT 88.015 202.215 88.900 202.385 ;
        RECT 89.080 201.915 89.395 202.415 ;
        RECT 89.625 202.085 89.965 202.645 ;
        RECT 90.135 201.915 90.305 202.925 ;
        RECT 90.475 202.130 90.805 202.975 ;
        RECT 91.035 202.085 91.305 202.990 ;
        RECT 91.490 202.845 92.155 203.015 ;
        RECT 91.475 201.915 91.805 202.675 ;
        RECT 91.985 202.085 92.155 202.845 ;
        RECT 93.415 202.845 94.090 203.015 ;
        RECT 94.365 202.990 94.545 203.790 ;
        RECT 93.415 202.085 93.595 202.845 ;
        RECT 93.775 201.915 94.105 202.675 ;
        RECT 94.275 202.085 94.545 202.990 ;
        RECT 94.715 203.790 94.975 204.295 ;
        RECT 95.155 204.085 95.485 204.465 ;
        RECT 95.665 203.915 95.835 204.295 ;
        RECT 94.715 202.990 94.885 203.790 ;
        RECT 95.170 203.745 95.835 203.915 ;
        RECT 95.170 203.490 95.340 203.745 ;
        RECT 96.555 203.740 96.845 204.465 ;
        RECT 97.015 203.725 97.480 204.270 ;
        RECT 95.055 203.160 95.340 203.490 ;
        RECT 95.575 203.195 95.905 203.565 ;
        RECT 95.170 203.015 95.340 203.160 ;
        RECT 94.715 202.085 94.985 202.990 ;
        RECT 95.170 202.845 95.835 203.015 ;
        RECT 95.155 201.915 95.485 202.675 ;
        RECT 95.665 202.085 95.835 202.845 ;
        RECT 96.555 201.915 96.845 203.080 ;
        RECT 97.015 202.765 97.185 203.725 ;
        RECT 97.985 203.645 98.155 204.465 ;
        RECT 98.325 203.815 98.655 204.295 ;
        RECT 98.825 204.075 99.175 204.465 ;
        RECT 99.345 203.895 99.575 204.295 ;
        RECT 99.065 203.815 99.575 203.895 ;
        RECT 98.325 203.725 99.575 203.815 ;
        RECT 99.745 203.725 100.065 204.205 ;
        RECT 98.325 203.645 99.235 203.725 ;
        RECT 97.355 203.105 97.600 203.555 ;
        RECT 97.860 203.275 98.555 203.475 ;
        RECT 98.725 203.305 99.325 203.475 ;
        RECT 98.725 203.105 98.895 203.305 ;
        RECT 99.555 203.135 99.725 203.555 ;
        RECT 97.355 202.935 98.895 203.105 ;
        RECT 99.065 202.965 99.725 203.135 ;
        RECT 99.065 202.765 99.235 202.965 ;
        RECT 99.895 202.795 100.065 203.725 ;
        RECT 97.015 202.595 99.235 202.765 ;
        RECT 99.405 202.595 100.065 202.795 ;
        RECT 100.695 203.815 100.955 204.295 ;
        RECT 101.125 204.005 101.455 204.465 ;
        RECT 101.645 203.825 101.845 204.245 ;
        RECT 100.695 202.785 100.865 203.815 ;
        RECT 101.035 203.125 101.265 203.555 ;
        RECT 101.435 203.305 101.845 203.825 ;
        RECT 102.015 203.980 102.805 204.245 ;
        RECT 102.015 203.125 102.270 203.980 ;
        RECT 102.985 203.645 103.315 204.065 ;
        RECT 103.485 203.645 103.745 204.465 ;
        RECT 104.840 203.725 105.095 204.295 ;
        RECT 105.265 204.065 105.595 204.465 ;
        RECT 106.020 203.930 106.550 204.295 ;
        RECT 106.020 203.895 106.195 203.930 ;
        RECT 105.265 203.725 106.195 203.895 ;
        RECT 106.740 203.785 107.015 204.295 ;
        RECT 102.985 203.555 103.235 203.645 ;
        RECT 102.440 203.305 103.235 203.555 ;
        RECT 101.035 202.955 102.825 203.125 ;
        RECT 97.015 201.915 97.315 202.425 ;
        RECT 97.485 202.085 97.815 202.595 ;
        RECT 99.405 202.425 99.575 202.595 ;
        RECT 97.985 201.915 98.615 202.425 ;
        RECT 99.195 202.255 99.575 202.425 ;
        RECT 99.745 201.915 100.045 202.425 ;
        RECT 100.695 202.085 100.970 202.785 ;
        RECT 101.140 202.660 101.855 202.955 ;
        RECT 102.075 202.595 102.405 202.785 ;
        RECT 101.180 201.915 101.395 202.460 ;
        RECT 101.565 202.085 102.040 202.425 ;
        RECT 102.210 202.420 102.405 202.595 ;
        RECT 102.575 202.590 102.825 202.955 ;
        RECT 102.210 201.915 102.825 202.420 ;
        RECT 103.065 202.085 103.235 203.305 ;
        RECT 103.405 202.595 103.745 203.475 ;
        RECT 104.840 203.055 105.010 203.725 ;
        RECT 105.265 203.555 105.435 203.725 ;
        RECT 105.180 203.225 105.435 203.555 ;
        RECT 105.660 203.225 105.855 203.555 ;
        RECT 103.485 201.915 103.745 202.425 ;
        RECT 104.840 202.085 105.175 203.055 ;
        RECT 105.345 201.915 105.515 203.055 ;
        RECT 105.685 202.255 105.855 203.225 ;
        RECT 106.025 202.595 106.195 203.725 ;
        RECT 106.365 202.935 106.535 203.735 ;
        RECT 106.735 203.615 107.015 203.785 ;
        RECT 106.740 203.135 107.015 203.615 ;
        RECT 107.185 202.935 107.375 204.295 ;
        RECT 107.555 203.930 108.065 204.465 ;
        RECT 108.285 203.655 108.530 204.260 ;
        RECT 109.025 203.810 109.355 204.245 ;
        RECT 109.525 203.855 109.695 204.465 ;
        RECT 108.975 203.725 109.355 203.810 ;
        RECT 109.865 203.725 110.195 204.250 ;
        RECT 110.455 203.935 110.665 204.465 ;
        RECT 110.940 204.015 111.725 204.185 ;
        RECT 111.895 204.015 112.300 204.185 ;
        RECT 108.975 203.685 109.200 203.725 ;
        RECT 107.575 203.485 108.805 203.655 ;
        RECT 106.365 202.765 107.375 202.935 ;
        RECT 107.545 202.920 108.295 203.110 ;
        RECT 106.025 202.425 107.150 202.595 ;
        RECT 107.545 202.255 107.715 202.920 ;
        RECT 108.465 202.675 108.805 203.485 ;
        RECT 108.975 203.105 109.145 203.685 ;
        RECT 109.865 203.555 110.065 203.725 ;
        RECT 110.940 203.555 111.110 204.015 ;
        RECT 109.315 203.225 110.065 203.555 ;
        RECT 110.235 203.225 111.110 203.555 ;
        RECT 108.975 203.055 109.190 203.105 ;
        RECT 108.975 202.975 109.365 203.055 ;
        RECT 105.685 202.085 107.715 202.255 ;
        RECT 107.885 201.915 108.055 202.675 ;
        RECT 108.290 202.265 108.805 202.675 ;
        RECT 109.035 202.130 109.365 202.975 ;
        RECT 109.875 203.020 110.065 203.225 ;
        RECT 109.535 201.915 109.705 202.925 ;
        RECT 109.875 202.645 110.770 203.020 ;
        RECT 109.875 202.085 110.215 202.645 ;
        RECT 110.445 201.915 110.760 202.415 ;
        RECT 110.940 202.385 111.110 203.225 ;
        RECT 111.280 203.515 111.745 203.845 ;
        RECT 112.130 203.785 112.300 204.015 ;
        RECT 112.480 203.965 112.850 204.465 ;
        RECT 113.170 204.015 113.845 204.185 ;
        RECT 114.040 204.015 114.375 204.185 ;
        RECT 111.280 202.555 111.600 203.515 ;
        RECT 112.130 203.485 112.960 203.785 ;
        RECT 111.770 202.585 111.960 203.305 ;
        RECT 112.130 202.415 112.300 203.485 ;
        RECT 112.760 203.455 112.960 203.485 ;
        RECT 112.470 203.235 112.640 203.305 ;
        RECT 113.170 203.235 113.340 204.015 ;
        RECT 114.205 203.875 114.375 204.015 ;
        RECT 114.545 204.005 114.795 204.465 ;
        RECT 112.470 203.065 113.340 203.235 ;
        RECT 113.510 203.595 114.035 203.815 ;
        RECT 114.205 203.745 114.430 203.875 ;
        RECT 112.470 202.975 112.980 203.065 ;
        RECT 110.940 202.215 111.825 202.385 ;
        RECT 112.050 202.085 112.300 202.415 ;
        RECT 112.470 201.915 112.640 202.715 ;
        RECT 112.810 202.360 112.980 202.975 ;
        RECT 113.510 202.895 113.680 203.595 ;
        RECT 113.150 202.530 113.680 202.895 ;
        RECT 113.850 202.830 114.090 203.425 ;
        RECT 114.260 202.640 114.430 203.745 ;
        RECT 114.600 202.885 114.880 203.835 ;
        RECT 114.125 202.510 114.430 202.640 ;
        RECT 112.810 202.190 113.915 202.360 ;
        RECT 114.125 202.085 114.375 202.510 ;
        RECT 114.545 201.915 114.810 202.375 ;
        RECT 115.050 202.085 115.235 204.205 ;
        RECT 115.405 204.085 115.735 204.465 ;
        RECT 115.905 203.915 116.075 204.205 ;
        RECT 115.410 203.745 116.075 203.915 ;
        RECT 116.335 203.790 116.595 204.295 ;
        RECT 116.775 204.085 117.105 204.465 ;
        RECT 117.285 203.915 117.455 204.295 ;
        RECT 115.410 202.755 115.640 203.745 ;
        RECT 115.810 202.925 116.160 203.575 ;
        RECT 116.335 202.990 116.505 203.790 ;
        RECT 116.790 203.745 117.455 203.915 ;
        RECT 116.790 203.490 116.960 203.745 ;
        RECT 117.720 203.725 117.975 204.295 ;
        RECT 118.145 204.065 118.475 204.465 ;
        RECT 118.900 203.930 119.430 204.295 ;
        RECT 118.900 203.895 119.075 203.930 ;
        RECT 118.145 203.725 119.075 203.895 ;
        RECT 116.675 203.160 116.960 203.490 ;
        RECT 117.195 203.195 117.525 203.565 ;
        RECT 116.790 203.015 116.960 203.160 ;
        RECT 117.720 203.055 117.890 203.725 ;
        RECT 118.145 203.555 118.315 203.725 ;
        RECT 118.060 203.225 118.315 203.555 ;
        RECT 118.540 203.225 118.735 203.555 ;
        RECT 115.410 202.585 116.075 202.755 ;
        RECT 115.405 201.915 115.735 202.415 ;
        RECT 115.905 202.085 116.075 202.585 ;
        RECT 116.335 202.085 116.605 202.990 ;
        RECT 116.790 202.845 117.455 203.015 ;
        RECT 116.775 201.915 117.105 202.675 ;
        RECT 117.285 202.085 117.455 202.845 ;
        RECT 117.720 202.085 118.055 203.055 ;
        RECT 118.225 201.915 118.395 203.055 ;
        RECT 118.565 202.255 118.735 203.225 ;
        RECT 118.905 202.595 119.075 203.725 ;
        RECT 119.245 202.935 119.415 203.735 ;
        RECT 119.620 203.445 119.895 204.295 ;
        RECT 119.615 203.275 119.895 203.445 ;
        RECT 119.620 203.135 119.895 203.275 ;
        RECT 120.065 202.935 120.255 204.295 ;
        RECT 120.435 203.930 120.945 204.465 ;
        RECT 121.165 203.655 121.410 204.260 ;
        RECT 122.315 203.740 122.605 204.465 ;
        RECT 122.775 203.715 123.985 204.465 ;
        RECT 124.245 203.915 124.415 204.295 ;
        RECT 124.595 204.085 124.925 204.465 ;
        RECT 124.245 203.745 124.910 203.915 ;
        RECT 125.105 203.790 125.365 204.295 ;
        RECT 120.455 203.485 121.685 203.655 ;
        RECT 119.245 202.765 120.255 202.935 ;
        RECT 120.425 202.920 121.175 203.110 ;
        RECT 118.905 202.425 120.030 202.595 ;
        RECT 120.425 202.255 120.595 202.920 ;
        RECT 121.345 202.675 121.685 203.485 ;
        RECT 122.775 203.175 123.295 203.715 ;
        RECT 118.565 202.085 120.595 202.255 ;
        RECT 120.765 201.915 120.935 202.675 ;
        RECT 121.170 202.265 121.685 202.675 ;
        RECT 122.315 201.915 122.605 203.080 ;
        RECT 123.465 203.005 123.985 203.545 ;
        RECT 124.175 203.195 124.505 203.565 ;
        RECT 124.740 203.490 124.910 203.745 ;
        RECT 124.740 203.160 125.025 203.490 ;
        RECT 124.740 203.015 124.910 203.160 ;
        RECT 122.775 201.915 123.985 203.005 ;
        RECT 124.245 202.845 124.910 203.015 ;
        RECT 125.195 202.990 125.365 203.790 ;
        RECT 125.625 203.915 125.795 204.205 ;
        RECT 125.965 204.085 126.295 204.465 ;
        RECT 125.625 203.745 126.290 203.915 ;
        RECT 124.245 202.085 124.415 202.845 ;
        RECT 124.595 201.915 124.925 202.675 ;
        RECT 125.095 202.085 125.365 202.990 ;
        RECT 125.540 202.925 125.890 203.575 ;
        RECT 126.060 202.755 126.290 203.745 ;
        RECT 125.625 202.585 126.290 202.755 ;
        RECT 125.625 202.085 125.795 202.585 ;
        RECT 125.965 201.915 126.295 202.415 ;
        RECT 126.465 202.085 126.650 204.205 ;
        RECT 126.905 204.005 127.155 204.465 ;
        RECT 127.325 204.015 127.660 204.185 ;
        RECT 127.855 204.015 128.530 204.185 ;
        RECT 127.325 203.875 127.495 204.015 ;
        RECT 126.820 202.885 127.100 203.835 ;
        RECT 127.270 203.745 127.495 203.875 ;
        RECT 127.270 202.640 127.440 203.745 ;
        RECT 127.665 203.595 128.190 203.815 ;
        RECT 127.610 202.830 127.850 203.425 ;
        RECT 128.020 202.895 128.190 203.595 ;
        RECT 128.360 203.235 128.530 204.015 ;
        RECT 128.850 203.965 129.220 204.465 ;
        RECT 129.400 204.015 129.805 204.185 ;
        RECT 129.975 204.015 130.760 204.185 ;
        RECT 129.400 203.785 129.570 204.015 ;
        RECT 128.740 203.485 129.570 203.785 ;
        RECT 129.955 203.515 130.420 203.845 ;
        RECT 128.740 203.455 128.940 203.485 ;
        RECT 129.060 203.235 129.230 203.305 ;
        RECT 128.360 203.065 129.230 203.235 ;
        RECT 128.720 202.975 129.230 203.065 ;
        RECT 127.270 202.510 127.575 202.640 ;
        RECT 128.020 202.530 128.550 202.895 ;
        RECT 126.890 201.915 127.155 202.375 ;
        RECT 127.325 202.085 127.575 202.510 ;
        RECT 128.720 202.360 128.890 202.975 ;
        RECT 127.785 202.190 128.890 202.360 ;
        RECT 129.060 201.915 129.230 202.715 ;
        RECT 129.400 202.415 129.570 203.485 ;
        RECT 129.740 202.585 129.930 203.305 ;
        RECT 130.100 202.555 130.420 203.515 ;
        RECT 130.590 203.555 130.760 204.015 ;
        RECT 131.035 203.935 131.245 204.465 ;
        RECT 131.505 203.725 131.835 204.250 ;
        RECT 132.005 203.855 132.175 204.465 ;
        RECT 132.345 203.810 132.675 204.245 ;
        RECT 132.345 203.725 132.725 203.810 ;
        RECT 131.635 203.555 131.835 203.725 ;
        RECT 132.500 203.685 132.725 203.725 ;
        RECT 130.590 203.225 131.465 203.555 ;
        RECT 131.635 203.225 132.385 203.555 ;
        RECT 129.400 202.085 129.650 202.415 ;
        RECT 130.590 202.385 130.760 203.225 ;
        RECT 131.635 203.020 131.825 203.225 ;
        RECT 132.555 203.105 132.725 203.685 ;
        RECT 132.510 203.055 132.725 203.105 ;
        RECT 130.930 202.645 131.825 203.020 ;
        RECT 132.335 202.975 132.725 203.055 ;
        RECT 133.355 203.790 133.615 204.295 ;
        RECT 133.795 204.085 134.125 204.465 ;
        RECT 134.305 203.915 134.475 204.295 ;
        RECT 133.355 202.990 133.535 203.790 ;
        RECT 133.810 203.745 134.475 203.915 ;
        RECT 135.745 203.915 135.915 204.295 ;
        RECT 136.095 204.085 136.425 204.465 ;
        RECT 135.745 203.745 136.410 203.915 ;
        RECT 136.605 203.790 136.865 204.295 ;
        RECT 133.810 203.490 133.980 203.745 ;
        RECT 133.705 203.160 133.980 203.490 ;
        RECT 134.205 203.195 134.545 203.565 ;
        RECT 135.675 203.195 136.005 203.565 ;
        RECT 136.240 203.490 136.410 203.745 ;
        RECT 133.810 203.015 133.980 203.160 ;
        RECT 136.240 203.160 136.525 203.490 ;
        RECT 136.240 203.015 136.410 203.160 ;
        RECT 129.875 202.215 130.760 202.385 ;
        RECT 130.940 201.915 131.255 202.415 ;
        RECT 131.485 202.085 131.825 202.645 ;
        RECT 131.995 201.915 132.165 202.925 ;
        RECT 132.335 202.130 132.665 202.975 ;
        RECT 133.355 202.085 133.625 202.990 ;
        RECT 133.810 202.845 134.485 203.015 ;
        RECT 133.795 201.915 134.125 202.675 ;
        RECT 134.305 202.085 134.485 202.845 ;
        RECT 135.745 202.845 136.410 203.015 ;
        RECT 136.695 202.990 136.865 203.790 ;
        RECT 137.125 203.915 137.295 204.205 ;
        RECT 137.465 204.085 137.795 204.465 ;
        RECT 137.125 203.745 137.790 203.915 ;
        RECT 135.745 202.085 135.915 202.845 ;
        RECT 136.095 201.915 136.425 202.675 ;
        RECT 136.595 202.085 136.865 202.990 ;
        RECT 137.040 202.925 137.390 203.575 ;
        RECT 137.560 202.755 137.790 203.745 ;
        RECT 137.125 202.585 137.790 202.755 ;
        RECT 137.125 202.085 137.295 202.585 ;
        RECT 137.465 201.915 137.795 202.415 ;
        RECT 137.965 202.085 138.150 204.205 ;
        RECT 138.405 204.005 138.655 204.465 ;
        RECT 138.825 204.015 139.160 204.185 ;
        RECT 139.355 204.015 140.030 204.185 ;
        RECT 138.825 203.875 138.995 204.015 ;
        RECT 138.320 202.885 138.600 203.835 ;
        RECT 138.770 203.745 138.995 203.875 ;
        RECT 138.770 202.640 138.940 203.745 ;
        RECT 139.165 203.595 139.690 203.815 ;
        RECT 139.110 202.830 139.350 203.425 ;
        RECT 139.520 202.895 139.690 203.595 ;
        RECT 139.860 203.235 140.030 204.015 ;
        RECT 140.350 203.965 140.720 204.465 ;
        RECT 140.900 204.015 141.305 204.185 ;
        RECT 141.475 204.015 142.260 204.185 ;
        RECT 140.900 203.785 141.070 204.015 ;
        RECT 140.240 203.485 141.070 203.785 ;
        RECT 141.455 203.515 141.920 203.845 ;
        RECT 140.240 203.455 140.440 203.485 ;
        RECT 140.560 203.235 140.730 203.305 ;
        RECT 139.860 203.065 140.730 203.235 ;
        RECT 140.220 202.975 140.730 203.065 ;
        RECT 138.770 202.510 139.075 202.640 ;
        RECT 139.520 202.530 140.050 202.895 ;
        RECT 138.390 201.915 138.655 202.375 ;
        RECT 138.825 202.085 139.075 202.510 ;
        RECT 140.220 202.360 140.390 202.975 ;
        RECT 139.285 202.190 140.390 202.360 ;
        RECT 140.560 201.915 140.730 202.715 ;
        RECT 140.900 202.415 141.070 203.485 ;
        RECT 141.240 202.585 141.430 203.305 ;
        RECT 141.600 202.555 141.920 203.515 ;
        RECT 142.090 203.555 142.260 204.015 ;
        RECT 142.535 203.935 142.745 204.465 ;
        RECT 143.005 203.725 143.335 204.250 ;
        RECT 143.505 203.855 143.675 204.465 ;
        RECT 143.845 203.810 144.175 204.245 ;
        RECT 143.845 203.725 144.225 203.810 ;
        RECT 143.135 203.555 143.335 203.725 ;
        RECT 144.000 203.685 144.225 203.725 ;
        RECT 142.090 203.225 142.965 203.555 ;
        RECT 143.135 203.225 143.885 203.555 ;
        RECT 140.900 202.085 141.150 202.415 ;
        RECT 142.090 202.385 142.260 203.225 ;
        RECT 143.135 203.020 143.325 203.225 ;
        RECT 144.055 203.105 144.225 203.685 ;
        RECT 144.010 203.055 144.225 203.105 ;
        RECT 142.430 202.645 143.325 203.020 ;
        RECT 143.835 202.975 144.225 203.055 ;
        RECT 144.395 203.790 144.655 204.295 ;
        RECT 144.835 204.085 145.165 204.465 ;
        RECT 145.345 203.915 145.515 204.295 ;
        RECT 144.395 202.990 144.565 203.790 ;
        RECT 144.850 203.745 145.515 203.915 ;
        RECT 145.775 203.790 146.035 204.295 ;
        RECT 146.215 204.085 146.545 204.465 ;
        RECT 146.725 203.915 146.895 204.295 ;
        RECT 144.850 203.490 145.020 203.745 ;
        RECT 144.735 203.160 145.020 203.490 ;
        RECT 145.255 203.195 145.585 203.565 ;
        RECT 144.850 203.015 145.020 203.160 ;
        RECT 141.375 202.215 142.260 202.385 ;
        RECT 142.440 201.915 142.755 202.415 ;
        RECT 142.985 202.085 143.325 202.645 ;
        RECT 143.495 201.915 143.665 202.925 ;
        RECT 143.835 202.130 144.165 202.975 ;
        RECT 144.395 202.085 144.665 202.990 ;
        RECT 144.850 202.845 145.515 203.015 ;
        RECT 144.835 201.915 145.165 202.675 ;
        RECT 145.345 202.085 145.515 202.845 ;
        RECT 145.775 202.990 145.945 203.790 ;
        RECT 146.230 203.745 146.895 203.915 ;
        RECT 146.230 203.490 146.400 203.745 ;
        RECT 148.075 203.740 148.365 204.465 ;
        RECT 148.540 203.725 148.795 204.295 ;
        RECT 148.965 204.065 149.295 204.465 ;
        RECT 149.720 203.930 150.250 204.295 ;
        RECT 149.720 203.895 149.895 203.930 ;
        RECT 148.965 203.725 149.895 203.895 ;
        RECT 146.115 203.160 146.400 203.490 ;
        RECT 146.635 203.195 146.965 203.565 ;
        RECT 146.230 203.015 146.400 203.160 ;
        RECT 145.775 202.085 146.045 202.990 ;
        RECT 146.230 202.845 146.895 203.015 ;
        RECT 146.215 201.915 146.545 202.675 ;
        RECT 146.725 202.085 146.895 202.845 ;
        RECT 148.075 201.915 148.365 203.080 ;
        RECT 148.540 203.055 148.710 203.725 ;
        RECT 148.965 203.555 149.135 203.725 ;
        RECT 148.880 203.225 149.135 203.555 ;
        RECT 149.360 203.225 149.555 203.555 ;
        RECT 148.540 202.085 148.875 203.055 ;
        RECT 149.045 201.915 149.215 203.055 ;
        RECT 149.385 202.255 149.555 203.225 ;
        RECT 149.725 202.595 149.895 203.725 ;
        RECT 150.065 202.935 150.235 203.735 ;
        RECT 150.440 203.445 150.715 204.295 ;
        RECT 150.435 203.275 150.715 203.445 ;
        RECT 150.440 203.135 150.715 203.275 ;
        RECT 150.885 202.935 151.075 204.295 ;
        RECT 151.255 203.930 151.765 204.465 ;
        RECT 151.985 203.655 152.230 204.260 ;
        RECT 152.675 203.790 152.935 204.295 ;
        RECT 153.115 204.085 153.445 204.465 ;
        RECT 153.625 203.915 153.795 204.295 ;
        RECT 151.275 203.485 152.505 203.655 ;
        RECT 150.065 202.765 151.075 202.935 ;
        RECT 151.245 202.920 151.995 203.110 ;
        RECT 149.725 202.425 150.850 202.595 ;
        RECT 151.245 202.255 151.415 202.920 ;
        RECT 152.165 202.675 152.505 203.485 ;
        RECT 149.385 202.085 151.415 202.255 ;
        RECT 151.585 201.915 151.755 202.675 ;
        RECT 151.990 202.265 152.505 202.675 ;
        RECT 152.675 202.990 152.855 203.790 ;
        RECT 153.130 203.745 153.795 203.915 ;
        RECT 153.130 203.490 153.300 203.745 ;
        RECT 154.975 203.715 156.185 204.465 ;
        RECT 153.025 203.160 153.300 203.490 ;
        RECT 153.525 203.195 153.865 203.565 ;
        RECT 153.130 203.015 153.300 203.160 ;
        RECT 152.675 202.085 152.945 202.990 ;
        RECT 153.130 202.845 153.805 203.015 ;
        RECT 153.115 201.915 153.445 202.675 ;
        RECT 153.625 202.085 153.805 202.845 ;
        RECT 154.975 203.005 155.495 203.545 ;
        RECT 155.665 203.175 156.185 203.715 ;
        RECT 154.975 201.915 156.185 203.005 ;
        RECT 70.710 201.745 156.270 201.915 ;
        RECT 70.795 200.655 72.005 201.745 ;
        RECT 72.175 200.655 73.845 201.745 ;
        RECT 74.105 201.075 74.275 201.575 ;
        RECT 74.445 201.245 74.775 201.745 ;
        RECT 74.105 200.905 74.770 201.075 ;
        RECT 70.795 199.945 71.315 200.485 ;
        RECT 71.485 200.115 72.005 200.655 ;
        RECT 72.175 199.965 72.925 200.485 ;
        RECT 73.095 200.135 73.845 200.655 ;
        RECT 74.020 200.085 74.370 200.735 ;
        RECT 70.795 199.195 72.005 199.945 ;
        RECT 72.175 199.195 73.845 199.965 ;
        RECT 74.540 199.915 74.770 200.905 ;
        RECT 74.105 199.745 74.770 199.915 ;
        RECT 74.105 199.455 74.275 199.745 ;
        RECT 74.445 199.195 74.775 199.575 ;
        RECT 74.945 199.455 75.130 201.575 ;
        RECT 75.370 201.285 75.635 201.745 ;
        RECT 75.805 201.150 76.055 201.575 ;
        RECT 76.265 201.300 77.370 201.470 ;
        RECT 75.750 201.020 76.055 201.150 ;
        RECT 75.300 199.825 75.580 200.775 ;
        RECT 75.750 199.915 75.920 201.020 ;
        RECT 76.090 200.235 76.330 200.830 ;
        RECT 76.500 200.765 77.030 201.130 ;
        RECT 76.500 200.065 76.670 200.765 ;
        RECT 77.200 200.685 77.370 201.300 ;
        RECT 77.540 200.945 77.710 201.745 ;
        RECT 77.880 201.245 78.130 201.575 ;
        RECT 78.355 201.275 79.240 201.445 ;
        RECT 77.200 200.595 77.710 200.685 ;
        RECT 75.750 199.785 75.975 199.915 ;
        RECT 76.145 199.845 76.670 200.065 ;
        RECT 76.840 200.425 77.710 200.595 ;
        RECT 75.385 199.195 75.635 199.655 ;
        RECT 75.805 199.645 75.975 199.785 ;
        RECT 76.840 199.645 77.010 200.425 ;
        RECT 77.540 200.355 77.710 200.425 ;
        RECT 77.220 200.175 77.420 200.205 ;
        RECT 77.880 200.175 78.050 201.245 ;
        RECT 78.220 200.355 78.410 201.075 ;
        RECT 77.220 199.875 78.050 200.175 ;
        RECT 78.580 200.145 78.900 201.105 ;
        RECT 75.805 199.475 76.140 199.645 ;
        RECT 76.335 199.475 77.010 199.645 ;
        RECT 77.330 199.195 77.700 199.695 ;
        RECT 77.880 199.645 78.050 199.875 ;
        RECT 78.435 199.815 78.900 200.145 ;
        RECT 79.070 200.435 79.240 201.275 ;
        RECT 79.420 201.245 79.735 201.745 ;
        RECT 79.965 201.015 80.305 201.575 ;
        RECT 79.410 200.640 80.305 201.015 ;
        RECT 80.475 200.735 80.645 201.745 ;
        RECT 80.115 200.435 80.305 200.640 ;
        RECT 80.815 200.685 81.145 201.530 ;
        RECT 82.385 200.815 82.555 201.575 ;
        RECT 82.735 200.985 83.065 201.745 ;
        RECT 80.815 200.605 81.205 200.685 ;
        RECT 82.385 200.645 83.050 200.815 ;
        RECT 83.235 200.670 83.505 201.575 ;
        RECT 80.990 200.555 81.205 200.605 ;
        RECT 79.070 200.105 79.945 200.435 ;
        RECT 80.115 200.105 80.865 200.435 ;
        RECT 79.070 199.645 79.240 200.105 ;
        RECT 80.115 199.935 80.315 200.105 ;
        RECT 81.035 199.975 81.205 200.555 ;
        RECT 82.880 200.500 83.050 200.645 ;
        RECT 82.315 200.095 82.645 200.465 ;
        RECT 82.880 200.170 83.165 200.500 ;
        RECT 80.980 199.935 81.205 199.975 ;
        RECT 77.880 199.475 78.285 199.645 ;
        RECT 78.455 199.475 79.240 199.645 ;
        RECT 79.515 199.195 79.725 199.725 ;
        RECT 79.985 199.410 80.315 199.935 ;
        RECT 80.825 199.850 81.205 199.935 ;
        RECT 82.880 199.915 83.050 200.170 ;
        RECT 80.485 199.195 80.655 199.805 ;
        RECT 80.825 199.415 81.155 199.850 ;
        RECT 82.385 199.745 83.050 199.915 ;
        RECT 83.335 199.870 83.505 200.670 ;
        RECT 83.675 200.580 83.965 201.745 ;
        RECT 84.195 200.685 84.525 201.530 ;
        RECT 84.695 200.735 84.865 201.745 ;
        RECT 85.035 201.015 85.375 201.575 ;
        RECT 85.605 201.245 85.920 201.745 ;
        RECT 86.100 201.275 86.985 201.445 ;
        RECT 84.135 200.605 84.525 200.685 ;
        RECT 85.035 200.640 85.930 201.015 ;
        RECT 84.135 200.555 84.350 200.605 ;
        RECT 84.135 199.975 84.305 200.555 ;
        RECT 85.035 200.435 85.225 200.640 ;
        RECT 86.100 200.435 86.270 201.275 ;
        RECT 87.210 201.245 87.460 201.575 ;
        RECT 84.475 200.105 85.225 200.435 ;
        RECT 85.395 200.105 86.270 200.435 ;
        RECT 84.135 199.935 84.360 199.975 ;
        RECT 85.025 199.935 85.225 200.105 ;
        RECT 82.385 199.365 82.555 199.745 ;
        RECT 82.735 199.195 83.065 199.575 ;
        RECT 83.245 199.365 83.505 199.870 ;
        RECT 83.675 199.195 83.965 199.920 ;
        RECT 84.135 199.850 84.515 199.935 ;
        RECT 84.185 199.415 84.515 199.850 ;
        RECT 84.685 199.195 84.855 199.805 ;
        RECT 85.025 199.410 85.355 199.935 ;
        RECT 85.615 199.195 85.825 199.725 ;
        RECT 86.100 199.645 86.270 200.105 ;
        RECT 86.440 200.145 86.760 201.105 ;
        RECT 86.930 200.355 87.120 201.075 ;
        RECT 87.290 200.175 87.460 201.245 ;
        RECT 87.630 200.945 87.800 201.745 ;
        RECT 87.970 201.300 89.075 201.470 ;
        RECT 87.970 200.685 88.140 201.300 ;
        RECT 89.285 201.150 89.535 201.575 ;
        RECT 89.705 201.285 89.970 201.745 ;
        RECT 88.310 200.765 88.840 201.130 ;
        RECT 89.285 201.020 89.590 201.150 ;
        RECT 87.630 200.595 88.140 200.685 ;
        RECT 87.630 200.425 88.500 200.595 ;
        RECT 87.630 200.355 87.800 200.425 ;
        RECT 87.920 200.175 88.120 200.205 ;
        RECT 86.440 199.815 86.905 200.145 ;
        RECT 87.290 199.875 88.120 200.175 ;
        RECT 87.290 199.645 87.460 199.875 ;
        RECT 86.100 199.475 86.885 199.645 ;
        RECT 87.055 199.475 87.460 199.645 ;
        RECT 87.640 199.195 88.010 199.695 ;
        RECT 88.330 199.645 88.500 200.425 ;
        RECT 88.670 200.065 88.840 200.765 ;
        RECT 89.010 200.235 89.250 200.830 ;
        RECT 88.670 199.845 89.195 200.065 ;
        RECT 89.420 199.915 89.590 201.020 ;
        RECT 89.365 199.785 89.590 199.915 ;
        RECT 89.760 199.825 90.040 200.775 ;
        RECT 89.365 199.645 89.535 199.785 ;
        RECT 88.330 199.475 89.005 199.645 ;
        RECT 89.200 199.475 89.535 199.645 ;
        RECT 89.705 199.195 89.955 199.655 ;
        RECT 90.210 199.455 90.395 201.575 ;
        RECT 90.565 201.245 90.895 201.745 ;
        RECT 91.065 201.075 91.235 201.575 ;
        RECT 90.570 200.905 91.235 201.075 ;
        RECT 92.045 201.075 92.215 201.575 ;
        RECT 92.385 201.245 92.715 201.745 ;
        RECT 92.045 200.905 92.710 201.075 ;
        RECT 90.570 199.915 90.800 200.905 ;
        RECT 90.970 200.085 91.320 200.735 ;
        RECT 91.960 200.085 92.310 200.735 ;
        RECT 92.480 199.915 92.710 200.905 ;
        RECT 90.570 199.745 91.235 199.915 ;
        RECT 90.565 199.195 90.895 199.575 ;
        RECT 91.065 199.455 91.235 199.745 ;
        RECT 92.045 199.745 92.710 199.915 ;
        RECT 92.045 199.455 92.215 199.745 ;
        RECT 92.385 199.195 92.715 199.575 ;
        RECT 92.885 199.455 93.070 201.575 ;
        RECT 93.310 201.285 93.575 201.745 ;
        RECT 93.745 201.150 93.995 201.575 ;
        RECT 94.205 201.300 95.310 201.470 ;
        RECT 93.690 201.020 93.995 201.150 ;
        RECT 93.240 199.825 93.520 200.775 ;
        RECT 93.690 199.915 93.860 201.020 ;
        RECT 94.030 200.235 94.270 200.830 ;
        RECT 94.440 200.765 94.970 201.130 ;
        RECT 94.440 200.065 94.610 200.765 ;
        RECT 95.140 200.685 95.310 201.300 ;
        RECT 95.480 200.945 95.650 201.745 ;
        RECT 95.820 201.245 96.070 201.575 ;
        RECT 96.295 201.275 97.180 201.445 ;
        RECT 95.140 200.595 95.650 200.685 ;
        RECT 93.690 199.785 93.915 199.915 ;
        RECT 94.085 199.845 94.610 200.065 ;
        RECT 94.780 200.425 95.650 200.595 ;
        RECT 93.325 199.195 93.575 199.655 ;
        RECT 93.745 199.645 93.915 199.785 ;
        RECT 94.780 199.645 94.950 200.425 ;
        RECT 95.480 200.355 95.650 200.425 ;
        RECT 95.160 200.175 95.360 200.205 ;
        RECT 95.820 200.175 95.990 201.245 ;
        RECT 96.160 200.355 96.350 201.075 ;
        RECT 95.160 199.875 95.990 200.175 ;
        RECT 96.520 200.145 96.840 201.105 ;
        RECT 93.745 199.475 94.080 199.645 ;
        RECT 94.275 199.475 94.950 199.645 ;
        RECT 95.270 199.195 95.640 199.695 ;
        RECT 95.820 199.645 95.990 199.875 ;
        RECT 96.375 199.815 96.840 200.145 ;
        RECT 97.010 200.435 97.180 201.275 ;
        RECT 97.360 201.245 97.675 201.745 ;
        RECT 97.905 201.015 98.245 201.575 ;
        RECT 97.350 200.640 98.245 201.015 ;
        RECT 98.415 200.735 98.585 201.745 ;
        RECT 98.055 200.435 98.245 200.640 ;
        RECT 98.755 200.685 99.085 201.530 ;
        RECT 99.315 200.985 99.830 201.395 ;
        RECT 100.065 200.985 100.235 201.745 ;
        RECT 100.405 201.405 102.435 201.575 ;
        RECT 98.755 200.605 99.145 200.685 ;
        RECT 98.930 200.555 99.145 200.605 ;
        RECT 97.010 200.105 97.885 200.435 ;
        RECT 98.055 200.105 98.805 200.435 ;
        RECT 97.010 199.645 97.180 200.105 ;
        RECT 98.055 199.935 98.255 200.105 ;
        RECT 98.975 199.975 99.145 200.555 ;
        RECT 99.315 200.175 99.655 200.985 ;
        RECT 100.405 200.740 100.575 201.405 ;
        RECT 100.970 201.065 102.095 201.235 ;
        RECT 99.825 200.550 100.575 200.740 ;
        RECT 100.745 200.725 101.755 200.895 ;
        RECT 99.315 200.005 100.545 200.175 ;
        RECT 98.920 199.935 99.145 199.975 ;
        RECT 95.820 199.475 96.225 199.645 ;
        RECT 96.395 199.475 97.180 199.645 ;
        RECT 97.455 199.195 97.665 199.725 ;
        RECT 97.925 199.410 98.255 199.935 ;
        RECT 98.765 199.850 99.145 199.935 ;
        RECT 98.425 199.195 98.595 199.805 ;
        RECT 98.765 199.415 99.095 199.850 ;
        RECT 99.590 199.400 99.835 200.005 ;
        RECT 100.055 199.195 100.565 199.730 ;
        RECT 100.745 199.365 100.935 200.725 ;
        RECT 101.105 200.045 101.380 200.525 ;
        RECT 101.105 199.875 101.385 200.045 ;
        RECT 101.585 199.925 101.755 200.725 ;
        RECT 101.925 199.935 102.095 201.065 ;
        RECT 102.265 200.435 102.435 201.405 ;
        RECT 102.605 200.605 102.775 201.745 ;
        RECT 102.945 200.605 103.280 201.575 ;
        RECT 102.265 200.105 102.460 200.435 ;
        RECT 102.685 200.105 102.940 200.435 ;
        RECT 102.685 199.935 102.855 200.105 ;
        RECT 103.110 199.935 103.280 200.605 ;
        RECT 101.105 199.365 101.380 199.875 ;
        RECT 101.925 199.765 102.855 199.935 ;
        RECT 101.925 199.730 102.100 199.765 ;
        RECT 101.570 199.365 102.100 199.730 ;
        RECT 102.525 199.195 102.855 199.595 ;
        RECT 103.025 199.365 103.280 199.935 ;
        RECT 104.375 201.025 104.835 201.575 ;
        RECT 105.025 201.025 105.355 201.745 ;
        RECT 104.375 199.655 104.625 201.025 ;
        RECT 105.555 200.855 105.855 201.405 ;
        RECT 106.025 201.075 106.305 201.745 ;
        RECT 104.915 200.685 105.855 200.855 ;
        RECT 104.915 200.435 105.085 200.685 ;
        RECT 106.225 200.435 106.490 200.795 ;
        RECT 106.685 200.605 107.015 201.745 ;
        RECT 107.545 200.775 107.875 201.560 ;
        RECT 107.195 200.605 107.875 200.775 ;
        RECT 108.095 200.605 108.325 201.745 ;
        RECT 104.795 200.105 105.085 200.435 ;
        RECT 105.255 200.185 105.595 200.435 ;
        RECT 105.815 200.185 106.490 200.435 ;
        RECT 106.675 200.185 107.025 200.435 ;
        RECT 104.915 200.015 105.085 200.105 ;
        RECT 104.915 199.825 106.305 200.015 ;
        RECT 107.195 200.005 107.365 200.605 ;
        RECT 108.495 200.595 108.825 201.575 ;
        RECT 108.995 200.605 109.205 201.745 ;
        RECT 107.535 200.185 107.885 200.435 ;
        RECT 108.075 200.185 108.405 200.435 ;
        RECT 104.375 199.365 104.935 199.655 ;
        RECT 105.105 199.195 105.355 199.655 ;
        RECT 105.975 199.465 106.305 199.825 ;
        RECT 106.685 199.195 106.955 200.005 ;
        RECT 107.125 199.365 107.455 200.005 ;
        RECT 107.625 199.195 107.865 200.005 ;
        RECT 108.095 199.195 108.325 200.015 ;
        RECT 108.575 199.995 108.825 200.595 ;
        RECT 109.435 200.580 109.725 201.745 ;
        RECT 110.815 200.140 111.095 201.575 ;
        RECT 111.265 200.970 111.975 201.745 ;
        RECT 112.145 200.800 112.475 201.575 ;
        RECT 111.325 200.585 112.475 200.800 ;
        RECT 108.495 199.365 108.825 199.995 ;
        RECT 108.995 199.195 109.205 200.015 ;
        RECT 109.435 199.195 109.725 199.920 ;
        RECT 110.815 199.365 111.155 200.140 ;
        RECT 111.325 200.015 111.610 200.585 ;
        RECT 111.795 200.185 112.265 200.415 ;
        RECT 112.670 200.385 112.885 201.500 ;
        RECT 113.065 201.025 113.395 201.745 ;
        RECT 114.585 201.075 114.755 201.575 ;
        RECT 114.925 201.245 115.255 201.745 ;
        RECT 114.585 200.905 115.250 201.075 ;
        RECT 113.175 200.385 113.405 200.725 ;
        RECT 112.435 200.205 112.885 200.385 ;
        RECT 112.435 200.185 112.765 200.205 ;
        RECT 113.075 200.185 113.405 200.385 ;
        RECT 114.500 200.085 114.850 200.735 ;
        RECT 111.325 199.825 112.035 200.015 ;
        RECT 111.735 199.685 112.035 199.825 ;
        RECT 112.225 199.825 113.405 200.015 ;
        RECT 115.020 199.915 115.250 200.905 ;
        RECT 112.225 199.745 112.555 199.825 ;
        RECT 111.735 199.675 112.050 199.685 ;
        RECT 111.735 199.665 112.060 199.675 ;
        RECT 111.735 199.660 112.070 199.665 ;
        RECT 111.325 199.195 111.495 199.655 ;
        RECT 111.735 199.650 112.075 199.660 ;
        RECT 111.735 199.645 112.080 199.650 ;
        RECT 111.735 199.635 112.085 199.645 ;
        RECT 111.735 199.630 112.090 199.635 ;
        RECT 111.735 199.365 112.095 199.630 ;
        RECT 112.725 199.195 112.895 199.655 ;
        RECT 113.065 199.365 113.405 199.825 ;
        RECT 114.585 199.745 115.250 199.915 ;
        RECT 114.585 199.455 114.755 199.745 ;
        RECT 114.925 199.195 115.255 199.575 ;
        RECT 115.425 199.455 115.610 201.575 ;
        RECT 115.850 201.285 116.115 201.745 ;
        RECT 116.285 201.150 116.535 201.575 ;
        RECT 116.745 201.300 117.850 201.470 ;
        RECT 116.230 201.020 116.535 201.150 ;
        RECT 115.780 199.825 116.060 200.775 ;
        RECT 116.230 199.915 116.400 201.020 ;
        RECT 116.570 200.235 116.810 200.830 ;
        RECT 116.980 200.765 117.510 201.130 ;
        RECT 116.980 200.065 117.150 200.765 ;
        RECT 117.680 200.685 117.850 201.300 ;
        RECT 118.020 200.945 118.190 201.745 ;
        RECT 118.360 201.245 118.610 201.575 ;
        RECT 118.835 201.275 119.720 201.445 ;
        RECT 117.680 200.595 118.190 200.685 ;
        RECT 116.230 199.785 116.455 199.915 ;
        RECT 116.625 199.845 117.150 200.065 ;
        RECT 117.320 200.425 118.190 200.595 ;
        RECT 115.865 199.195 116.115 199.655 ;
        RECT 116.285 199.645 116.455 199.785 ;
        RECT 117.320 199.645 117.490 200.425 ;
        RECT 118.020 200.355 118.190 200.425 ;
        RECT 117.700 200.175 117.900 200.205 ;
        RECT 118.360 200.175 118.530 201.245 ;
        RECT 118.700 200.355 118.890 201.075 ;
        RECT 117.700 199.875 118.530 200.175 ;
        RECT 119.060 200.145 119.380 201.105 ;
        RECT 116.285 199.475 116.620 199.645 ;
        RECT 116.815 199.475 117.490 199.645 ;
        RECT 117.810 199.195 118.180 199.695 ;
        RECT 118.360 199.645 118.530 199.875 ;
        RECT 118.915 199.815 119.380 200.145 ;
        RECT 119.550 200.435 119.720 201.275 ;
        RECT 119.900 201.245 120.215 201.745 ;
        RECT 120.445 201.015 120.785 201.575 ;
        RECT 119.890 200.640 120.785 201.015 ;
        RECT 120.955 200.735 121.125 201.745 ;
        RECT 120.595 200.435 120.785 200.640 ;
        RECT 121.295 200.685 121.625 201.530 ;
        RECT 121.295 200.605 121.685 200.685 ;
        RECT 121.470 200.555 121.685 200.605 ;
        RECT 119.550 200.105 120.425 200.435 ;
        RECT 120.595 200.105 121.345 200.435 ;
        RECT 119.550 199.645 119.720 200.105 ;
        RECT 120.595 199.935 120.795 200.105 ;
        RECT 121.515 199.975 121.685 200.555 ;
        RECT 121.460 199.935 121.685 199.975 ;
        RECT 118.360 199.475 118.765 199.645 ;
        RECT 118.935 199.475 119.720 199.645 ;
        RECT 119.995 199.195 120.205 199.725 ;
        RECT 120.465 199.410 120.795 199.935 ;
        RECT 121.305 199.850 121.685 199.935 ;
        RECT 121.855 200.140 122.135 201.575 ;
        RECT 122.305 200.970 123.015 201.745 ;
        RECT 123.185 200.800 123.515 201.575 ;
        RECT 122.365 200.585 123.515 200.800 ;
        RECT 120.965 199.195 121.135 199.805 ;
        RECT 121.305 199.415 121.635 199.850 ;
        RECT 121.855 199.365 122.195 200.140 ;
        RECT 122.365 200.015 122.650 200.585 ;
        RECT 122.835 200.185 123.305 200.415 ;
        RECT 123.710 200.385 123.925 201.500 ;
        RECT 124.105 201.025 124.435 201.745 ;
        RECT 125.075 200.985 125.590 201.395 ;
        RECT 125.825 200.985 125.995 201.745 ;
        RECT 126.165 201.405 128.195 201.575 ;
        RECT 124.215 200.385 124.445 200.725 ;
        RECT 123.475 200.205 123.925 200.385 ;
        RECT 123.475 200.185 123.805 200.205 ;
        RECT 124.115 200.185 124.445 200.385 ;
        RECT 125.075 200.175 125.415 200.985 ;
        RECT 126.165 200.740 126.335 201.405 ;
        RECT 126.730 201.065 127.855 201.235 ;
        RECT 125.585 200.550 126.335 200.740 ;
        RECT 126.505 200.725 127.515 200.895 ;
        RECT 122.365 199.825 123.075 200.015 ;
        RECT 122.775 199.685 123.075 199.825 ;
        RECT 123.265 199.825 124.445 200.015 ;
        RECT 125.075 200.005 126.305 200.175 ;
        RECT 123.265 199.745 123.595 199.825 ;
        RECT 122.775 199.675 123.090 199.685 ;
        RECT 122.775 199.665 123.100 199.675 ;
        RECT 122.775 199.660 123.110 199.665 ;
        RECT 122.365 199.195 122.535 199.655 ;
        RECT 122.775 199.650 123.115 199.660 ;
        RECT 122.775 199.645 123.120 199.650 ;
        RECT 122.775 199.635 123.125 199.645 ;
        RECT 122.775 199.630 123.130 199.635 ;
        RECT 122.775 199.365 123.135 199.630 ;
        RECT 123.765 199.195 123.935 199.655 ;
        RECT 124.105 199.365 124.445 199.825 ;
        RECT 125.350 199.400 125.595 200.005 ;
        RECT 125.815 199.195 126.325 199.730 ;
        RECT 126.505 199.365 126.695 200.725 ;
        RECT 126.865 200.045 127.140 200.525 ;
        RECT 126.865 199.875 127.145 200.045 ;
        RECT 127.345 199.925 127.515 200.725 ;
        RECT 127.685 199.935 127.855 201.065 ;
        RECT 128.025 200.435 128.195 201.405 ;
        RECT 128.365 200.605 128.535 201.745 ;
        RECT 128.705 200.605 129.040 201.575 ;
        RECT 128.025 200.105 128.220 200.435 ;
        RECT 128.445 200.105 128.700 200.435 ;
        RECT 128.445 199.935 128.615 200.105 ;
        RECT 128.870 199.935 129.040 200.605 ;
        RECT 126.865 199.365 127.140 199.875 ;
        RECT 127.685 199.765 128.615 199.935 ;
        RECT 127.685 199.730 127.860 199.765 ;
        RECT 127.330 199.365 127.860 199.730 ;
        RECT 128.285 199.195 128.615 199.595 ;
        RECT 128.785 199.365 129.040 199.935 ;
        RECT 129.215 200.140 129.495 201.575 ;
        RECT 129.665 200.970 130.375 201.745 ;
        RECT 130.545 200.800 130.875 201.575 ;
        RECT 129.725 200.585 130.875 200.800 ;
        RECT 129.215 199.365 129.555 200.140 ;
        RECT 129.725 200.015 130.010 200.585 ;
        RECT 130.195 200.185 130.665 200.415 ;
        RECT 131.070 200.385 131.285 201.500 ;
        RECT 131.465 201.025 131.795 201.745 ;
        RECT 131.575 200.385 131.805 200.725 ;
        RECT 130.835 200.205 131.285 200.385 ;
        RECT 130.835 200.185 131.165 200.205 ;
        RECT 131.475 200.185 131.805 200.385 ;
        RECT 132.435 200.140 132.715 201.575 ;
        RECT 132.885 200.970 133.595 201.745 ;
        RECT 133.765 200.800 134.095 201.575 ;
        RECT 132.945 200.585 134.095 200.800 ;
        RECT 129.725 199.825 130.435 200.015 ;
        RECT 130.135 199.685 130.435 199.825 ;
        RECT 130.625 199.825 131.805 200.015 ;
        RECT 130.625 199.745 130.955 199.825 ;
        RECT 130.135 199.675 130.450 199.685 ;
        RECT 130.135 199.665 130.460 199.675 ;
        RECT 130.135 199.660 130.470 199.665 ;
        RECT 129.725 199.195 129.895 199.655 ;
        RECT 130.135 199.650 130.475 199.660 ;
        RECT 130.135 199.645 130.480 199.650 ;
        RECT 130.135 199.635 130.485 199.645 ;
        RECT 130.135 199.630 130.490 199.635 ;
        RECT 130.135 199.365 130.495 199.630 ;
        RECT 131.125 199.195 131.295 199.655 ;
        RECT 131.465 199.365 131.805 199.825 ;
        RECT 132.435 199.365 132.775 200.140 ;
        RECT 132.945 200.015 133.230 200.585 ;
        RECT 133.415 200.185 133.885 200.415 ;
        RECT 134.290 200.385 134.505 201.500 ;
        RECT 134.685 201.025 135.015 201.745 ;
        RECT 134.795 200.385 135.025 200.725 ;
        RECT 135.195 200.580 135.485 201.745 ;
        RECT 135.660 200.605 135.995 201.575 ;
        RECT 136.165 200.605 136.335 201.745 ;
        RECT 136.505 201.405 138.535 201.575 ;
        RECT 134.055 200.205 134.505 200.385 ;
        RECT 134.055 200.185 134.385 200.205 ;
        RECT 134.695 200.185 135.025 200.385 ;
        RECT 132.945 199.825 133.655 200.015 ;
        RECT 133.355 199.685 133.655 199.825 ;
        RECT 133.845 199.825 135.025 200.015 ;
        RECT 135.660 199.935 135.830 200.605 ;
        RECT 136.505 200.435 136.675 201.405 ;
        RECT 136.000 200.105 136.255 200.435 ;
        RECT 136.480 200.105 136.675 200.435 ;
        RECT 136.845 201.065 137.970 201.235 ;
        RECT 136.085 199.935 136.255 200.105 ;
        RECT 136.845 199.935 137.015 201.065 ;
        RECT 133.845 199.745 134.175 199.825 ;
        RECT 133.355 199.675 133.670 199.685 ;
        RECT 133.355 199.665 133.680 199.675 ;
        RECT 133.355 199.660 133.690 199.665 ;
        RECT 132.945 199.195 133.115 199.655 ;
        RECT 133.355 199.650 133.695 199.660 ;
        RECT 133.355 199.645 133.700 199.650 ;
        RECT 133.355 199.635 133.705 199.645 ;
        RECT 133.355 199.630 133.710 199.635 ;
        RECT 133.355 199.365 133.715 199.630 ;
        RECT 134.345 199.195 134.515 199.655 ;
        RECT 134.685 199.365 135.025 199.825 ;
        RECT 135.195 199.195 135.485 199.920 ;
        RECT 135.660 199.365 135.915 199.935 ;
        RECT 136.085 199.765 137.015 199.935 ;
        RECT 137.185 200.725 138.195 200.895 ;
        RECT 137.185 199.925 137.355 200.725 ;
        RECT 137.560 200.385 137.835 200.525 ;
        RECT 137.555 200.215 137.835 200.385 ;
        RECT 136.840 199.730 137.015 199.765 ;
        RECT 136.085 199.195 136.415 199.595 ;
        RECT 136.840 199.365 137.370 199.730 ;
        RECT 137.560 199.365 137.835 200.215 ;
        RECT 138.005 199.365 138.195 200.725 ;
        RECT 138.365 200.740 138.535 201.405 ;
        RECT 138.705 200.985 138.875 201.745 ;
        RECT 139.110 200.985 139.625 201.395 ;
        RECT 139.800 201.320 140.135 201.745 ;
        RECT 140.305 201.140 140.490 201.545 ;
        RECT 138.365 200.550 139.115 200.740 ;
        RECT 139.285 200.175 139.625 200.985 ;
        RECT 138.395 200.005 139.625 200.175 ;
        RECT 139.825 200.965 140.490 201.140 ;
        RECT 140.695 200.965 141.025 201.745 ;
        RECT 138.375 199.195 138.885 199.730 ;
        RECT 139.105 199.400 139.350 200.005 ;
        RECT 139.825 199.935 140.165 200.965 ;
        RECT 141.195 200.775 141.465 201.545 ;
        RECT 140.335 200.605 141.465 200.775 ;
        RECT 140.335 200.105 140.585 200.605 ;
        RECT 139.825 199.765 140.510 199.935 ;
        RECT 140.765 199.855 141.125 200.435 ;
        RECT 139.800 199.195 140.135 199.595 ;
        RECT 140.305 199.365 140.510 199.765 ;
        RECT 141.295 199.695 141.465 200.605 ;
        RECT 142.095 200.985 142.610 201.395 ;
        RECT 142.845 200.985 143.015 201.745 ;
        RECT 143.185 201.405 145.215 201.575 ;
        RECT 142.095 200.175 142.435 200.985 ;
        RECT 143.185 200.740 143.355 201.405 ;
        RECT 143.750 201.065 144.875 201.235 ;
        RECT 142.605 200.550 143.355 200.740 ;
        RECT 143.525 200.725 144.535 200.895 ;
        RECT 142.095 200.005 143.325 200.175 ;
        RECT 140.720 199.195 140.995 199.675 ;
        RECT 141.205 199.365 141.465 199.695 ;
        RECT 142.370 199.400 142.615 200.005 ;
        RECT 142.835 199.195 143.345 199.730 ;
        RECT 143.525 199.365 143.715 200.725 ;
        RECT 143.885 200.045 144.160 200.525 ;
        RECT 143.885 199.875 144.165 200.045 ;
        RECT 144.365 199.925 144.535 200.725 ;
        RECT 144.705 199.935 144.875 201.065 ;
        RECT 145.045 200.435 145.215 201.405 ;
        RECT 145.385 200.605 145.555 201.745 ;
        RECT 145.725 200.605 146.060 201.575 ;
        RECT 146.325 201.075 146.495 201.575 ;
        RECT 146.665 201.245 146.995 201.745 ;
        RECT 146.325 200.905 146.990 201.075 ;
        RECT 145.045 200.105 145.240 200.435 ;
        RECT 145.465 200.105 145.720 200.435 ;
        RECT 145.465 199.935 145.635 200.105 ;
        RECT 145.890 199.935 146.060 200.605 ;
        RECT 146.240 200.085 146.590 200.735 ;
        RECT 143.885 199.365 144.160 199.875 ;
        RECT 144.705 199.765 145.635 199.935 ;
        RECT 144.705 199.730 144.880 199.765 ;
        RECT 144.350 199.365 144.880 199.730 ;
        RECT 145.305 199.195 145.635 199.595 ;
        RECT 145.805 199.365 146.060 199.935 ;
        RECT 146.760 199.915 146.990 200.905 ;
        RECT 146.325 199.745 146.990 199.915 ;
        RECT 146.325 199.455 146.495 199.745 ;
        RECT 146.665 199.195 146.995 199.575 ;
        RECT 147.165 199.455 147.350 201.575 ;
        RECT 147.590 201.285 147.855 201.745 ;
        RECT 148.025 201.150 148.275 201.575 ;
        RECT 148.485 201.300 149.590 201.470 ;
        RECT 147.970 201.020 148.275 201.150 ;
        RECT 147.520 199.825 147.800 200.775 ;
        RECT 147.970 199.915 148.140 201.020 ;
        RECT 148.310 200.235 148.550 200.830 ;
        RECT 148.720 200.765 149.250 201.130 ;
        RECT 148.720 200.065 148.890 200.765 ;
        RECT 149.420 200.685 149.590 201.300 ;
        RECT 149.760 200.945 149.930 201.745 ;
        RECT 150.100 201.245 150.350 201.575 ;
        RECT 150.575 201.275 151.460 201.445 ;
        RECT 149.420 200.595 149.930 200.685 ;
        RECT 147.970 199.785 148.195 199.915 ;
        RECT 148.365 199.845 148.890 200.065 ;
        RECT 149.060 200.425 149.930 200.595 ;
        RECT 147.605 199.195 147.855 199.655 ;
        RECT 148.025 199.645 148.195 199.785 ;
        RECT 149.060 199.645 149.230 200.425 ;
        RECT 149.760 200.355 149.930 200.425 ;
        RECT 149.440 200.175 149.640 200.205 ;
        RECT 150.100 200.175 150.270 201.245 ;
        RECT 150.440 200.355 150.630 201.075 ;
        RECT 149.440 199.875 150.270 200.175 ;
        RECT 150.800 200.145 151.120 201.105 ;
        RECT 148.025 199.475 148.360 199.645 ;
        RECT 148.555 199.475 149.230 199.645 ;
        RECT 149.550 199.195 149.920 199.695 ;
        RECT 150.100 199.645 150.270 199.875 ;
        RECT 150.655 199.815 151.120 200.145 ;
        RECT 151.290 200.435 151.460 201.275 ;
        RECT 151.640 201.245 151.955 201.745 ;
        RECT 152.185 201.015 152.525 201.575 ;
        RECT 151.630 200.640 152.525 201.015 ;
        RECT 152.695 200.735 152.865 201.745 ;
        RECT 152.335 200.435 152.525 200.640 ;
        RECT 153.035 200.685 153.365 201.530 ;
        RECT 153.035 200.605 153.425 200.685 ;
        RECT 153.595 200.655 154.805 201.745 ;
        RECT 153.210 200.555 153.425 200.605 ;
        RECT 151.290 200.105 152.165 200.435 ;
        RECT 152.335 200.105 153.085 200.435 ;
        RECT 151.290 199.645 151.460 200.105 ;
        RECT 152.335 199.935 152.535 200.105 ;
        RECT 153.255 199.975 153.425 200.555 ;
        RECT 153.200 199.935 153.425 199.975 ;
        RECT 150.100 199.475 150.505 199.645 ;
        RECT 150.675 199.475 151.460 199.645 ;
        RECT 151.735 199.195 151.945 199.725 ;
        RECT 152.205 199.410 152.535 199.935 ;
        RECT 153.045 199.850 153.425 199.935 ;
        RECT 153.595 199.945 154.115 200.485 ;
        RECT 154.285 200.115 154.805 200.655 ;
        RECT 154.975 200.655 156.185 201.745 ;
        RECT 154.975 200.115 155.495 200.655 ;
        RECT 155.665 199.945 156.185 200.485 ;
        RECT 152.705 199.195 152.875 199.805 ;
        RECT 153.045 199.415 153.375 199.850 ;
        RECT 153.595 199.195 154.805 199.945 ;
        RECT 154.975 199.195 156.185 199.945 ;
        RECT 70.710 199.025 156.270 199.195 ;
        RECT 70.795 198.275 72.005 199.025 ;
        RECT 70.795 197.735 71.315 198.275 ;
        RECT 72.175 198.255 74.765 199.025 ;
        RECT 71.485 197.565 72.005 198.105 ;
        RECT 72.175 197.735 73.385 198.255 ;
        RECT 73.555 197.565 74.765 198.085 ;
        RECT 70.795 196.475 72.005 197.565 ;
        RECT 72.175 196.475 74.765 197.565 ;
        RECT 74.935 198.080 75.275 198.855 ;
        RECT 75.445 198.565 75.615 199.025 ;
        RECT 75.855 198.590 76.215 198.855 ;
        RECT 75.855 198.585 76.210 198.590 ;
        RECT 75.855 198.575 76.205 198.585 ;
        RECT 75.855 198.570 76.200 198.575 ;
        RECT 75.855 198.560 76.195 198.570 ;
        RECT 76.845 198.565 77.015 199.025 ;
        RECT 75.855 198.555 76.190 198.560 ;
        RECT 75.855 198.545 76.180 198.555 ;
        RECT 75.855 198.535 76.170 198.545 ;
        RECT 75.855 198.395 76.155 198.535 ;
        RECT 75.445 198.205 76.155 198.395 ;
        RECT 76.345 198.395 76.675 198.475 ;
        RECT 77.185 198.395 77.525 198.855 ;
        RECT 76.345 198.205 77.525 198.395 ;
        RECT 77.715 198.295 78.045 199.025 ;
        RECT 74.935 196.645 75.215 198.080 ;
        RECT 75.445 197.635 75.730 198.205 ;
        RECT 78.215 198.115 78.425 198.735 ;
        RECT 78.605 198.315 79.035 198.845 ;
        RECT 75.915 197.805 76.385 198.035 ;
        RECT 76.555 198.015 76.885 198.035 ;
        RECT 76.555 197.835 77.005 198.015 ;
        RECT 77.195 197.835 77.525 198.035 ;
        RECT 75.445 197.420 76.595 197.635 ;
        RECT 75.385 196.475 76.095 197.250 ;
        RECT 76.265 196.645 76.595 197.420 ;
        RECT 76.790 196.720 77.005 197.835 ;
        RECT 77.295 197.495 77.525 197.835 ;
        RECT 77.730 197.765 78.020 198.115 ;
        RECT 78.215 197.765 78.610 198.115 ;
        RECT 78.790 198.065 79.035 198.315 ;
        RECT 79.215 198.245 79.445 199.025 ;
        RECT 79.625 198.395 80.005 198.845 ;
        RECT 78.790 197.765 79.325 198.065 ;
        RECT 79.625 197.945 79.855 198.395 ;
        RECT 80.455 198.205 80.715 199.025 ;
        RECT 80.885 198.205 81.215 198.625 ;
        RECT 81.395 198.540 82.185 198.805 ;
        RECT 77.785 197.385 78.825 197.585 ;
        RECT 77.185 196.475 77.515 197.195 ;
        RECT 77.785 196.655 77.955 197.385 ;
        RECT 78.135 196.475 78.465 197.205 ;
        RECT 78.635 196.655 78.825 197.385 ;
        RECT 78.995 196.655 79.325 197.765 ;
        RECT 79.515 197.265 79.855 197.945 ;
        RECT 80.035 197.445 80.265 198.135 ;
        RECT 80.965 198.115 81.215 198.205 ;
        RECT 79.515 197.065 80.275 197.265 ;
        RECT 80.455 197.155 80.795 198.035 ;
        RECT 80.965 197.865 81.760 198.115 ;
        RECT 79.515 196.475 79.845 196.885 ;
        RECT 80.015 196.675 80.275 197.065 ;
        RECT 80.455 196.475 80.715 196.985 ;
        RECT 80.965 196.645 81.135 197.865 ;
        RECT 81.930 197.685 82.185 198.540 ;
        RECT 82.355 198.385 82.555 198.805 ;
        RECT 82.745 198.565 83.075 199.025 ;
        RECT 82.355 197.865 82.765 198.385 ;
        RECT 83.245 198.375 83.505 198.855 ;
        RECT 82.935 197.685 83.165 198.115 ;
        RECT 81.375 197.515 83.165 197.685 ;
        RECT 81.375 197.150 81.625 197.515 ;
        RECT 81.795 197.155 82.125 197.345 ;
        RECT 82.345 197.220 83.060 197.515 ;
        RECT 83.335 197.345 83.505 198.375 ;
        RECT 83.765 198.475 83.935 198.855 ;
        RECT 84.115 198.645 84.445 199.025 ;
        RECT 83.765 198.305 84.430 198.475 ;
        RECT 84.625 198.350 84.885 198.855 ;
        RECT 83.695 197.755 84.035 198.125 ;
        RECT 84.260 198.050 84.430 198.305 ;
        RECT 84.260 197.720 84.535 198.050 ;
        RECT 84.260 197.575 84.430 197.720 ;
        RECT 81.795 196.980 81.990 197.155 ;
        RECT 81.375 196.475 81.990 196.980 ;
        RECT 82.160 196.645 82.635 196.985 ;
        RECT 82.805 196.475 83.020 197.020 ;
        RECT 83.230 196.645 83.505 197.345 ;
        RECT 83.755 197.405 84.430 197.575 ;
        RECT 84.705 197.550 84.885 198.350 ;
        RECT 83.755 196.645 83.935 197.405 ;
        RECT 84.115 196.475 84.445 197.235 ;
        RECT 84.615 196.645 84.885 197.550 ;
        RECT 85.975 198.350 86.235 198.855 ;
        RECT 86.415 198.645 86.745 199.025 ;
        RECT 86.925 198.475 87.095 198.855 ;
        RECT 85.975 197.550 86.155 198.350 ;
        RECT 86.430 198.305 87.095 198.475 ;
        RECT 87.355 198.350 87.615 198.855 ;
        RECT 87.795 198.645 88.125 199.025 ;
        RECT 88.305 198.475 88.475 198.855 ;
        RECT 86.430 198.050 86.600 198.305 ;
        RECT 86.325 197.720 86.600 198.050 ;
        RECT 86.825 197.755 87.165 198.125 ;
        RECT 86.430 197.575 86.600 197.720 ;
        RECT 85.975 196.645 86.245 197.550 ;
        RECT 86.430 197.405 87.105 197.575 ;
        RECT 86.415 196.475 86.745 197.235 ;
        RECT 86.925 196.645 87.105 197.405 ;
        RECT 87.355 197.550 87.535 198.350 ;
        RECT 87.810 198.305 88.475 198.475 ;
        RECT 88.735 198.350 88.995 198.855 ;
        RECT 89.175 198.645 89.505 199.025 ;
        RECT 89.685 198.475 89.855 198.855 ;
        RECT 90.120 198.625 90.455 199.025 ;
        RECT 87.810 198.050 87.980 198.305 ;
        RECT 87.705 197.720 87.980 198.050 ;
        RECT 88.205 197.755 88.545 198.125 ;
        RECT 87.810 197.575 87.980 197.720 ;
        RECT 87.355 196.645 87.625 197.550 ;
        RECT 87.810 197.405 88.485 197.575 ;
        RECT 87.795 196.475 88.125 197.235 ;
        RECT 88.305 196.645 88.485 197.405 ;
        RECT 88.735 197.550 88.915 198.350 ;
        RECT 89.190 198.305 89.855 198.475 ;
        RECT 90.625 198.455 90.830 198.855 ;
        RECT 91.040 198.545 91.315 199.025 ;
        RECT 91.525 198.525 91.785 198.855 ;
        RECT 89.190 198.050 89.360 198.305 ;
        RECT 90.145 198.285 90.830 198.455 ;
        RECT 89.085 197.720 89.360 198.050 ;
        RECT 89.585 197.755 89.925 198.125 ;
        RECT 89.190 197.575 89.360 197.720 ;
        RECT 88.735 196.645 89.005 197.550 ;
        RECT 89.190 197.405 89.865 197.575 ;
        RECT 89.175 196.475 89.505 197.235 ;
        RECT 89.685 196.645 89.865 197.405 ;
        RECT 90.145 197.255 90.485 198.285 ;
        RECT 90.655 197.615 90.905 198.115 ;
        RECT 91.085 197.785 91.445 198.365 ;
        RECT 91.615 197.615 91.785 198.525 ;
        RECT 90.655 197.445 91.785 197.615 ;
        RECT 90.145 197.080 90.810 197.255 ;
        RECT 90.120 196.475 90.455 196.900 ;
        RECT 90.625 196.675 90.810 197.080 ;
        RECT 91.015 196.475 91.345 197.255 ;
        RECT 91.515 196.675 91.785 197.445 ;
        RECT 91.965 198.300 92.295 198.810 ;
        RECT 92.465 198.625 92.795 199.025 ;
        RECT 93.845 198.455 94.175 198.795 ;
        RECT 94.345 198.625 94.675 199.025 ;
        RECT 95.265 198.475 95.435 198.855 ;
        RECT 95.615 198.645 95.945 199.025 ;
        RECT 91.965 197.535 92.155 198.300 ;
        RECT 92.465 198.285 94.830 198.455 ;
        RECT 95.265 198.305 95.930 198.475 ;
        RECT 96.125 198.350 96.385 198.855 ;
        RECT 92.465 198.115 92.635 198.285 ;
        RECT 92.325 197.785 92.635 198.115 ;
        RECT 92.805 197.785 93.110 198.115 ;
        RECT 91.965 196.685 92.295 197.535 ;
        RECT 92.465 196.475 92.715 197.615 ;
        RECT 92.895 197.455 93.110 197.785 ;
        RECT 93.285 197.455 93.570 198.115 ;
        RECT 93.765 197.455 94.030 198.115 ;
        RECT 94.245 197.455 94.490 198.115 ;
        RECT 94.660 197.285 94.830 198.285 ;
        RECT 95.195 197.755 95.535 198.125 ;
        RECT 95.760 198.050 95.930 198.305 ;
        RECT 95.760 197.720 96.035 198.050 ;
        RECT 95.760 197.575 95.930 197.720 ;
        RECT 92.905 197.115 94.195 197.285 ;
        RECT 92.905 196.695 93.155 197.115 ;
        RECT 93.385 196.475 93.715 196.945 ;
        RECT 93.945 196.695 94.195 197.115 ;
        RECT 94.375 197.115 94.830 197.285 ;
        RECT 95.255 197.405 95.930 197.575 ;
        RECT 96.205 197.550 96.385 198.350 ;
        RECT 96.555 198.300 96.845 199.025 ;
        RECT 97.105 198.475 97.275 198.855 ;
        RECT 97.455 198.645 97.785 199.025 ;
        RECT 97.105 198.305 97.770 198.475 ;
        RECT 97.965 198.350 98.225 198.855 ;
        RECT 97.035 197.755 97.375 198.125 ;
        RECT 97.600 198.050 97.770 198.305 ;
        RECT 97.600 197.720 97.875 198.050 ;
        RECT 94.375 196.685 94.705 197.115 ;
        RECT 95.255 196.645 95.435 197.405 ;
        RECT 95.615 196.475 95.945 197.235 ;
        RECT 96.115 196.645 96.385 197.550 ;
        RECT 96.555 196.475 96.845 197.640 ;
        RECT 97.600 197.575 97.770 197.720 ;
        RECT 97.095 197.405 97.770 197.575 ;
        RECT 98.045 197.550 98.225 198.350 ;
        RECT 98.395 198.225 98.705 199.025 ;
        RECT 98.910 198.225 99.605 198.855 ;
        RECT 99.775 198.255 101.445 199.025 ;
        RECT 102.075 198.395 102.415 198.855 ;
        RECT 102.585 198.565 102.755 199.025 ;
        RECT 103.385 198.590 103.745 198.855 ;
        RECT 103.390 198.585 103.745 198.590 ;
        RECT 103.395 198.575 103.745 198.585 ;
        RECT 103.400 198.570 103.745 198.575 ;
        RECT 103.405 198.560 103.745 198.570 ;
        RECT 103.985 198.565 104.155 199.025 ;
        RECT 103.410 198.555 103.745 198.560 ;
        RECT 103.420 198.545 103.745 198.555 ;
        RECT 103.430 198.535 103.745 198.545 ;
        RECT 102.925 198.395 103.255 198.475 ;
        RECT 98.405 197.785 98.740 198.055 ;
        RECT 98.910 197.625 99.080 198.225 ;
        RECT 99.250 197.785 99.585 198.035 ;
        RECT 99.775 197.735 100.525 198.255 ;
        RECT 102.075 198.205 103.255 198.395 ;
        RECT 103.445 198.395 103.745 198.535 ;
        RECT 103.445 198.205 104.155 198.395 ;
        RECT 97.095 196.645 97.275 197.405 ;
        RECT 97.455 196.475 97.785 197.235 ;
        RECT 97.955 196.645 98.225 197.550 ;
        RECT 98.395 196.475 98.675 197.615 ;
        RECT 98.845 196.645 99.175 197.625 ;
        RECT 99.345 196.475 99.605 197.615 ;
        RECT 100.695 197.565 101.445 198.085 ;
        RECT 99.775 196.475 101.445 197.565 ;
        RECT 102.075 197.835 102.405 198.035 ;
        RECT 102.715 198.015 103.045 198.035 ;
        RECT 102.595 197.835 103.045 198.015 ;
        RECT 102.075 197.495 102.305 197.835 ;
        RECT 102.085 196.475 102.415 197.195 ;
        RECT 102.595 196.720 102.810 197.835 ;
        RECT 103.215 197.805 103.685 198.035 ;
        RECT 103.870 197.635 104.155 198.205 ;
        RECT 104.325 198.080 104.665 198.855 ;
        RECT 105.040 198.245 105.540 198.855 ;
        RECT 103.005 197.420 104.155 197.635 ;
        RECT 103.005 196.645 103.335 197.420 ;
        RECT 103.505 196.475 104.215 197.250 ;
        RECT 104.385 196.645 104.665 198.080 ;
        RECT 104.835 197.785 105.185 198.035 ;
        RECT 105.370 197.615 105.540 198.245 ;
        RECT 106.170 198.375 106.500 198.855 ;
        RECT 106.670 198.565 106.895 199.025 ;
        RECT 107.065 198.375 107.395 198.855 ;
        RECT 106.170 198.205 107.395 198.375 ;
        RECT 107.585 198.225 107.835 199.025 ;
        RECT 108.005 198.225 108.345 198.855 ;
        RECT 105.710 197.835 106.040 198.035 ;
        RECT 106.210 197.835 106.540 198.035 ;
        RECT 106.710 197.835 107.130 198.035 ;
        RECT 107.305 197.865 108.000 198.035 ;
        RECT 107.305 197.615 107.475 197.865 ;
        RECT 108.170 197.615 108.345 198.225 ;
        RECT 108.515 198.255 112.025 199.025 ;
        RECT 113.115 198.350 113.375 198.855 ;
        RECT 113.555 198.645 113.885 199.025 ;
        RECT 114.065 198.475 114.235 198.855 ;
        RECT 108.515 197.735 110.165 198.255 ;
        RECT 105.040 197.445 107.475 197.615 ;
        RECT 105.040 196.645 105.370 197.445 ;
        RECT 105.540 196.475 105.870 197.275 ;
        RECT 106.170 196.645 106.500 197.445 ;
        RECT 107.145 196.475 107.395 197.275 ;
        RECT 107.665 196.475 107.835 197.615 ;
        RECT 108.005 196.645 108.345 197.615 ;
        RECT 110.335 197.565 112.025 198.085 ;
        RECT 108.515 196.475 112.025 197.565 ;
        RECT 113.115 197.550 113.295 198.350 ;
        RECT 113.570 198.305 114.235 198.475 ;
        RECT 115.045 198.475 115.215 198.855 ;
        RECT 115.395 198.645 115.725 199.025 ;
        RECT 115.045 198.305 115.710 198.475 ;
        RECT 115.905 198.350 116.165 198.855 ;
        RECT 113.570 198.050 113.740 198.305 ;
        RECT 113.465 197.720 113.740 198.050 ;
        RECT 113.965 197.755 114.305 198.125 ;
        RECT 114.975 197.755 115.315 198.125 ;
        RECT 115.540 198.050 115.710 198.305 ;
        RECT 113.570 197.575 113.740 197.720 ;
        RECT 115.540 197.720 115.815 198.050 ;
        RECT 115.540 197.575 115.710 197.720 ;
        RECT 113.115 196.645 113.385 197.550 ;
        RECT 113.570 197.405 114.245 197.575 ;
        RECT 113.555 196.475 113.885 197.235 ;
        RECT 114.065 196.645 114.245 197.405 ;
        RECT 115.035 197.405 115.710 197.575 ;
        RECT 115.985 197.550 116.165 198.350 ;
        RECT 115.035 196.645 115.215 197.405 ;
        RECT 115.395 196.475 115.725 197.235 ;
        RECT 115.895 196.645 116.165 197.550 ;
        RECT 116.335 198.080 116.675 198.855 ;
        RECT 116.845 198.565 117.015 199.025 ;
        RECT 117.255 198.590 117.615 198.855 ;
        RECT 117.255 198.585 117.610 198.590 ;
        RECT 117.255 198.575 117.605 198.585 ;
        RECT 117.255 198.570 117.600 198.575 ;
        RECT 117.255 198.560 117.595 198.570 ;
        RECT 118.245 198.565 118.415 199.025 ;
        RECT 117.255 198.555 117.590 198.560 ;
        RECT 117.255 198.545 117.580 198.555 ;
        RECT 117.255 198.535 117.570 198.545 ;
        RECT 117.255 198.395 117.555 198.535 ;
        RECT 116.845 198.205 117.555 198.395 ;
        RECT 117.745 198.395 118.075 198.475 ;
        RECT 118.585 198.395 118.925 198.855 ;
        RECT 117.745 198.205 118.925 198.395 ;
        RECT 119.095 198.255 121.685 199.025 ;
        RECT 122.315 198.300 122.605 199.025 ;
        RECT 116.335 196.645 116.615 198.080 ;
        RECT 116.845 197.635 117.130 198.205 ;
        RECT 117.315 197.805 117.785 198.035 ;
        RECT 117.955 198.015 118.285 198.035 ;
        RECT 117.955 197.835 118.405 198.015 ;
        RECT 118.595 197.835 118.925 198.035 ;
        RECT 116.845 197.420 117.995 197.635 ;
        RECT 116.785 196.475 117.495 197.250 ;
        RECT 117.665 196.645 117.995 197.420 ;
        RECT 118.190 196.720 118.405 197.835 ;
        RECT 118.695 197.495 118.925 197.835 ;
        RECT 119.095 197.735 120.305 198.255 ;
        RECT 120.475 197.565 121.685 198.085 ;
        RECT 122.775 198.080 123.115 198.855 ;
        RECT 123.285 198.565 123.455 199.025 ;
        RECT 123.695 198.590 124.055 198.855 ;
        RECT 123.695 198.585 124.050 198.590 ;
        RECT 123.695 198.575 124.045 198.585 ;
        RECT 123.695 198.570 124.040 198.575 ;
        RECT 123.695 198.560 124.035 198.570 ;
        RECT 124.685 198.565 124.855 199.025 ;
        RECT 123.695 198.555 124.030 198.560 ;
        RECT 123.695 198.545 124.020 198.555 ;
        RECT 123.695 198.535 124.010 198.545 ;
        RECT 123.695 198.395 123.995 198.535 ;
        RECT 123.285 198.205 123.995 198.395 ;
        RECT 124.185 198.395 124.515 198.475 ;
        RECT 125.025 198.395 125.365 198.855 ;
        RECT 124.185 198.205 125.365 198.395 ;
        RECT 126.465 198.215 126.735 199.025 ;
        RECT 126.905 198.215 127.235 198.855 ;
        RECT 127.405 198.215 127.645 199.025 ;
        RECT 127.835 198.285 128.095 198.855 ;
        RECT 128.265 198.625 128.650 199.025 ;
        RECT 128.820 198.455 129.075 198.855 ;
        RECT 128.265 198.285 129.075 198.455 ;
        RECT 129.265 198.285 129.510 198.855 ;
        RECT 129.680 198.625 130.065 199.025 ;
        RECT 130.235 198.455 130.490 198.855 ;
        RECT 129.680 198.285 130.490 198.455 ;
        RECT 130.680 198.285 131.105 198.855 ;
        RECT 131.275 198.625 131.660 199.025 ;
        RECT 131.830 198.455 132.265 198.855 ;
        RECT 131.275 198.285 132.265 198.455 ;
        RECT 132.450 198.455 132.705 198.805 ;
        RECT 132.875 198.625 133.205 199.025 ;
        RECT 133.375 198.455 133.545 198.805 ;
        RECT 133.715 198.625 134.095 199.025 ;
        RECT 132.450 198.285 134.115 198.455 ;
        RECT 134.285 198.350 134.560 198.695 ;
        RECT 118.585 196.475 118.915 197.195 ;
        RECT 119.095 196.475 121.685 197.565 ;
        RECT 122.315 196.475 122.605 197.640 ;
        RECT 122.775 196.645 123.055 198.080 ;
        RECT 123.285 197.635 123.570 198.205 ;
        RECT 123.755 197.805 124.225 198.035 ;
        RECT 124.395 198.015 124.725 198.035 ;
        RECT 124.395 197.835 124.845 198.015 ;
        RECT 125.035 197.835 125.365 198.035 ;
        RECT 123.285 197.420 124.435 197.635 ;
        RECT 123.225 196.475 123.935 197.250 ;
        RECT 124.105 196.645 124.435 197.420 ;
        RECT 124.630 196.720 124.845 197.835 ;
        RECT 125.135 197.495 125.365 197.835 ;
        RECT 126.455 197.785 126.805 198.035 ;
        RECT 126.975 197.615 127.145 198.215 ;
        RECT 127.315 197.785 127.665 198.035 ;
        RECT 127.835 197.615 128.020 198.285 ;
        RECT 128.265 198.115 128.615 198.285 ;
        RECT 129.265 198.115 129.435 198.285 ;
        RECT 129.680 198.115 130.030 198.285 ;
        RECT 130.680 198.115 131.030 198.285 ;
        RECT 131.275 198.115 131.610 198.285 ;
        RECT 133.945 198.115 134.115 198.285 ;
        RECT 128.190 197.785 128.615 198.115 ;
        RECT 125.025 196.475 125.355 197.195 ;
        RECT 126.465 196.475 126.795 197.615 ;
        RECT 126.975 197.445 127.655 197.615 ;
        RECT 127.325 196.660 127.655 197.445 ;
        RECT 127.835 196.645 128.095 197.615 ;
        RECT 128.265 197.265 128.615 197.785 ;
        RECT 128.785 197.615 129.435 198.115 ;
        RECT 129.605 197.785 130.030 198.115 ;
        RECT 128.785 197.435 129.510 197.615 ;
        RECT 128.265 197.070 129.075 197.265 ;
        RECT 128.265 196.475 128.650 196.900 ;
        RECT 128.820 196.645 129.075 197.070 ;
        RECT 129.265 196.645 129.510 197.435 ;
        RECT 129.680 197.265 130.030 197.785 ;
        RECT 130.200 197.615 131.030 198.115 ;
        RECT 131.200 197.785 131.610 198.115 ;
        RECT 130.200 197.435 131.105 197.615 ;
        RECT 129.680 197.070 130.510 197.265 ;
        RECT 129.680 196.475 130.065 196.900 ;
        RECT 130.235 196.645 130.510 197.070 ;
        RECT 130.680 196.645 131.105 197.435 ;
        RECT 131.275 197.240 131.610 197.785 ;
        RECT 131.780 197.410 132.265 198.115 ;
        RECT 132.435 197.785 132.780 198.115 ;
        RECT 132.950 197.785 133.775 198.115 ;
        RECT 133.945 197.785 134.220 198.115 ;
        RECT 132.455 197.325 132.780 197.615 ;
        RECT 132.950 197.495 133.145 197.785 ;
        RECT 133.945 197.615 134.115 197.785 ;
        RECT 134.390 197.615 134.560 198.350 ;
        RECT 133.455 197.445 134.115 197.615 ;
        RECT 133.455 197.325 133.625 197.445 ;
        RECT 131.275 197.070 132.265 197.240 ;
        RECT 132.455 197.155 133.625 197.325 ;
        RECT 131.275 196.475 131.660 196.900 ;
        RECT 131.830 196.645 132.265 197.070 ;
        RECT 132.435 196.695 133.625 196.985 ;
        RECT 133.795 196.475 134.075 197.275 ;
        RECT 134.285 196.645 134.560 197.615 ;
        RECT 134.735 198.350 134.995 198.855 ;
        RECT 135.175 198.645 135.505 199.025 ;
        RECT 135.685 198.475 135.855 198.855 ;
        RECT 134.735 197.550 134.905 198.350 ;
        RECT 135.190 198.305 135.855 198.475 ;
        RECT 135.190 198.050 135.360 198.305 ;
        RECT 135.075 197.720 135.360 198.050 ;
        RECT 135.595 197.755 135.925 198.125 ;
        RECT 136.575 198.080 136.915 198.855 ;
        RECT 137.085 198.565 137.255 199.025 ;
        RECT 137.495 198.590 137.855 198.855 ;
        RECT 137.495 198.585 137.850 198.590 ;
        RECT 137.495 198.575 137.845 198.585 ;
        RECT 137.495 198.570 137.840 198.575 ;
        RECT 137.495 198.560 137.835 198.570 ;
        RECT 138.485 198.565 138.655 199.025 ;
        RECT 137.495 198.555 137.830 198.560 ;
        RECT 137.495 198.545 137.820 198.555 ;
        RECT 137.495 198.535 137.810 198.545 ;
        RECT 137.495 198.395 137.795 198.535 ;
        RECT 137.085 198.205 137.795 198.395 ;
        RECT 137.985 198.395 138.315 198.475 ;
        RECT 138.825 198.395 139.165 198.855 ;
        RECT 137.985 198.205 139.165 198.395 ;
        RECT 135.190 197.575 135.360 197.720 ;
        RECT 134.735 196.645 135.005 197.550 ;
        RECT 135.190 197.405 135.855 197.575 ;
        RECT 135.175 196.475 135.505 197.235 ;
        RECT 135.685 196.645 135.855 197.405 ;
        RECT 136.575 196.645 136.855 198.080 ;
        RECT 137.085 197.635 137.370 198.205 ;
        RECT 139.335 198.080 139.675 198.855 ;
        RECT 139.845 198.565 140.015 199.025 ;
        RECT 140.255 198.590 140.615 198.855 ;
        RECT 140.255 198.585 140.610 198.590 ;
        RECT 140.255 198.575 140.605 198.585 ;
        RECT 140.255 198.570 140.600 198.575 ;
        RECT 140.255 198.560 140.595 198.570 ;
        RECT 141.245 198.565 141.415 199.025 ;
        RECT 140.255 198.555 140.590 198.560 ;
        RECT 140.255 198.545 140.580 198.555 ;
        RECT 140.255 198.535 140.570 198.545 ;
        RECT 140.255 198.395 140.555 198.535 ;
        RECT 139.845 198.205 140.555 198.395 ;
        RECT 140.745 198.395 141.075 198.475 ;
        RECT 141.585 198.395 141.925 198.855 ;
        RECT 140.745 198.205 141.925 198.395 ;
        RECT 142.185 198.475 142.355 198.855 ;
        RECT 142.535 198.645 142.865 199.025 ;
        RECT 142.185 198.305 142.850 198.475 ;
        RECT 143.045 198.350 143.305 198.855 ;
        RECT 137.555 197.805 138.025 198.035 ;
        RECT 138.195 198.015 138.525 198.035 ;
        RECT 138.195 197.835 138.645 198.015 ;
        RECT 138.835 197.835 139.165 198.035 ;
        RECT 137.085 197.420 138.235 197.635 ;
        RECT 137.025 196.475 137.735 197.250 ;
        RECT 137.905 196.645 138.235 197.420 ;
        RECT 138.430 196.720 138.645 197.835 ;
        RECT 138.935 197.495 139.165 197.835 ;
        RECT 138.825 196.475 139.155 197.195 ;
        RECT 139.335 196.645 139.615 198.080 ;
        RECT 139.845 197.635 140.130 198.205 ;
        RECT 140.315 197.805 140.785 198.035 ;
        RECT 140.955 198.015 141.285 198.035 ;
        RECT 140.955 197.835 141.405 198.015 ;
        RECT 141.595 197.835 141.925 198.035 ;
        RECT 139.845 197.420 140.995 197.635 ;
        RECT 139.785 196.475 140.495 197.250 ;
        RECT 140.665 196.645 140.995 197.420 ;
        RECT 141.190 196.720 141.405 197.835 ;
        RECT 141.695 197.495 141.925 197.835 ;
        RECT 142.115 197.755 142.455 198.125 ;
        RECT 142.680 198.050 142.850 198.305 ;
        RECT 142.680 197.720 142.955 198.050 ;
        RECT 142.680 197.575 142.850 197.720 ;
        RECT 142.175 197.405 142.850 197.575 ;
        RECT 143.125 197.550 143.305 198.350 ;
        RECT 143.475 198.255 145.145 199.025 ;
        RECT 145.405 198.475 145.575 198.855 ;
        RECT 145.755 198.645 146.085 199.025 ;
        RECT 145.405 198.305 146.070 198.475 ;
        RECT 146.265 198.350 146.525 198.855 ;
        RECT 143.475 197.735 144.225 198.255 ;
        RECT 144.395 197.565 145.145 198.085 ;
        RECT 145.335 197.755 145.665 198.125 ;
        RECT 145.900 198.050 146.070 198.305 ;
        RECT 145.900 197.720 146.185 198.050 ;
        RECT 145.900 197.575 146.070 197.720 ;
        RECT 141.585 196.475 141.915 197.195 ;
        RECT 142.175 196.645 142.355 197.405 ;
        RECT 142.535 196.475 142.865 197.235 ;
        RECT 143.035 196.645 143.305 197.550 ;
        RECT 143.475 196.475 145.145 197.565 ;
        RECT 145.405 197.405 146.070 197.575 ;
        RECT 146.355 197.550 146.525 198.350 ;
        RECT 145.405 196.645 145.575 197.405 ;
        RECT 145.755 196.475 146.085 197.235 ;
        RECT 146.255 196.645 146.525 197.550 ;
        RECT 146.695 198.350 146.955 198.855 ;
        RECT 147.135 198.645 147.465 199.025 ;
        RECT 147.645 198.475 147.815 198.855 ;
        RECT 146.695 197.550 146.865 198.350 ;
        RECT 147.150 198.305 147.815 198.475 ;
        RECT 147.150 198.050 147.320 198.305 ;
        RECT 148.075 198.300 148.365 199.025 ;
        RECT 148.535 198.255 151.125 199.025 ;
        RECT 147.035 197.720 147.320 198.050 ;
        RECT 147.555 197.755 147.885 198.125 ;
        RECT 148.535 197.735 149.745 198.255 ;
        RECT 151.815 198.205 152.025 199.025 ;
        RECT 152.195 198.225 152.525 198.855 ;
        RECT 147.150 197.575 147.320 197.720 ;
        RECT 146.695 196.645 146.965 197.550 ;
        RECT 147.150 197.405 147.815 197.575 ;
        RECT 147.135 196.475 147.465 197.235 ;
        RECT 147.645 196.645 147.815 197.405 ;
        RECT 148.075 196.475 148.365 197.640 ;
        RECT 149.915 197.565 151.125 198.085 ;
        RECT 152.195 197.625 152.445 198.225 ;
        RECT 152.695 198.205 152.925 199.025 ;
        RECT 153.135 198.350 153.395 198.855 ;
        RECT 153.575 198.645 153.905 199.025 ;
        RECT 154.085 198.475 154.255 198.855 ;
        RECT 152.615 197.785 152.945 198.035 ;
        RECT 148.535 196.475 151.125 197.565 ;
        RECT 151.815 196.475 152.025 197.615 ;
        RECT 152.195 196.645 152.525 197.625 ;
        RECT 152.695 196.475 152.925 197.615 ;
        RECT 153.135 197.550 153.315 198.350 ;
        RECT 153.590 198.305 154.255 198.475 ;
        RECT 153.590 198.050 153.760 198.305 ;
        RECT 154.975 198.275 156.185 199.025 ;
        RECT 153.485 197.720 153.760 198.050 ;
        RECT 153.985 197.755 154.325 198.125 ;
        RECT 153.590 197.575 153.760 197.720 ;
        RECT 153.135 196.645 153.405 197.550 ;
        RECT 153.590 197.405 154.265 197.575 ;
        RECT 153.575 196.475 153.905 197.235 ;
        RECT 154.085 196.645 154.265 197.405 ;
        RECT 154.975 197.565 155.495 198.105 ;
        RECT 155.665 197.735 156.185 198.275 ;
        RECT 154.975 196.475 156.185 197.565 ;
        RECT 70.710 196.305 156.270 196.475 ;
        RECT 70.795 195.215 72.005 196.305 ;
        RECT 72.265 195.635 72.435 196.135 ;
        RECT 72.605 195.805 72.935 196.305 ;
        RECT 72.265 195.465 72.930 195.635 ;
        RECT 70.795 194.505 71.315 195.045 ;
        RECT 71.485 194.675 72.005 195.215 ;
        RECT 72.180 194.645 72.530 195.295 ;
        RECT 70.795 193.755 72.005 194.505 ;
        RECT 72.700 194.475 72.930 195.465 ;
        RECT 72.265 194.305 72.930 194.475 ;
        RECT 72.265 194.015 72.435 194.305 ;
        RECT 72.605 193.755 72.935 194.135 ;
        RECT 73.105 194.015 73.290 196.135 ;
        RECT 73.530 195.845 73.795 196.305 ;
        RECT 73.965 195.710 74.215 196.135 ;
        RECT 74.425 195.860 75.530 196.030 ;
        RECT 73.910 195.580 74.215 195.710 ;
        RECT 73.460 194.385 73.740 195.335 ;
        RECT 73.910 194.475 74.080 195.580 ;
        RECT 74.250 194.795 74.490 195.390 ;
        RECT 74.660 195.325 75.190 195.690 ;
        RECT 74.660 194.625 74.830 195.325 ;
        RECT 75.360 195.245 75.530 195.860 ;
        RECT 75.700 195.505 75.870 196.305 ;
        RECT 76.040 195.805 76.290 196.135 ;
        RECT 76.515 195.835 77.400 196.005 ;
        RECT 75.360 195.155 75.870 195.245 ;
        RECT 73.910 194.345 74.135 194.475 ;
        RECT 74.305 194.405 74.830 194.625 ;
        RECT 75.000 194.985 75.870 195.155 ;
        RECT 73.545 193.755 73.795 194.215 ;
        RECT 73.965 194.205 74.135 194.345 ;
        RECT 75.000 194.205 75.170 194.985 ;
        RECT 75.700 194.915 75.870 194.985 ;
        RECT 75.380 194.735 75.580 194.765 ;
        RECT 76.040 194.735 76.210 195.805 ;
        RECT 76.380 194.915 76.570 195.635 ;
        RECT 75.380 194.435 76.210 194.735 ;
        RECT 76.740 194.705 77.060 195.665 ;
        RECT 73.965 194.035 74.300 194.205 ;
        RECT 74.495 194.035 75.170 194.205 ;
        RECT 75.490 193.755 75.860 194.255 ;
        RECT 76.040 194.205 76.210 194.435 ;
        RECT 76.595 194.375 77.060 194.705 ;
        RECT 77.230 194.995 77.400 195.835 ;
        RECT 77.580 195.805 77.895 196.305 ;
        RECT 78.125 195.575 78.465 196.135 ;
        RECT 77.570 195.200 78.465 195.575 ;
        RECT 78.635 195.295 78.805 196.305 ;
        RECT 78.275 194.995 78.465 195.200 ;
        RECT 78.975 195.245 79.305 196.090 ;
        RECT 78.975 195.165 79.365 195.245 ;
        RECT 79.535 195.215 81.205 196.305 ;
        RECT 79.150 195.115 79.365 195.165 ;
        RECT 77.230 194.665 78.105 194.995 ;
        RECT 78.275 194.665 79.025 194.995 ;
        RECT 77.230 194.205 77.400 194.665 ;
        RECT 78.275 194.495 78.475 194.665 ;
        RECT 79.195 194.535 79.365 195.115 ;
        RECT 79.140 194.495 79.365 194.535 ;
        RECT 76.040 194.035 76.445 194.205 ;
        RECT 76.615 194.035 77.400 194.205 ;
        RECT 77.675 193.755 77.885 194.285 ;
        RECT 78.145 193.970 78.475 194.495 ;
        RECT 78.985 194.410 79.365 194.495 ;
        RECT 79.535 194.525 80.285 195.045 ;
        RECT 80.455 194.695 81.205 195.215 ;
        RECT 81.375 195.435 81.650 196.135 ;
        RECT 81.820 195.760 82.075 196.305 ;
        RECT 82.245 195.795 82.725 196.135 ;
        RECT 82.900 195.750 83.505 196.305 ;
        RECT 82.890 195.650 83.505 195.750 ;
        RECT 82.890 195.625 83.075 195.650 ;
        RECT 78.645 193.755 78.815 194.365 ;
        RECT 78.985 193.975 79.315 194.410 ;
        RECT 79.535 193.755 81.205 194.525 ;
        RECT 81.375 194.405 81.545 195.435 ;
        RECT 81.820 195.305 82.575 195.555 ;
        RECT 82.745 195.380 83.075 195.625 ;
        RECT 81.820 195.270 82.590 195.305 ;
        RECT 81.820 195.260 82.605 195.270 ;
        RECT 81.715 195.245 82.610 195.260 ;
        RECT 81.715 195.230 82.630 195.245 ;
        RECT 81.715 195.220 82.650 195.230 ;
        RECT 81.715 195.210 82.675 195.220 ;
        RECT 81.715 195.180 82.745 195.210 ;
        RECT 81.715 195.150 82.765 195.180 ;
        RECT 81.715 195.120 82.785 195.150 ;
        RECT 81.715 195.095 82.815 195.120 ;
        RECT 81.715 195.060 82.850 195.095 ;
        RECT 81.715 195.055 82.880 195.060 ;
        RECT 81.715 194.660 81.945 195.055 ;
        RECT 82.490 195.050 82.880 195.055 ;
        RECT 82.515 195.040 82.880 195.050 ;
        RECT 82.530 195.035 82.880 195.040 ;
        RECT 82.545 195.030 82.880 195.035 ;
        RECT 83.245 195.030 83.505 195.480 ;
        RECT 83.675 195.140 83.965 196.305 ;
        RECT 84.145 195.245 84.475 196.095 ;
        RECT 82.545 195.025 83.505 195.030 ;
        RECT 82.555 195.015 83.505 195.025 ;
        RECT 82.565 195.010 83.505 195.015 ;
        RECT 82.575 195.000 83.505 195.010 ;
        RECT 82.580 194.990 83.505 195.000 ;
        RECT 82.585 194.985 83.505 194.990 ;
        RECT 82.595 194.970 83.505 194.985 ;
        RECT 82.600 194.955 83.505 194.970 ;
        RECT 82.610 194.930 83.505 194.955 ;
        RECT 82.115 194.460 82.445 194.885 ;
        RECT 81.375 193.925 81.635 194.405 ;
        RECT 81.805 193.755 82.055 194.295 ;
        RECT 82.225 193.975 82.445 194.460 ;
        RECT 82.615 194.860 83.505 194.930 ;
        RECT 82.615 194.135 82.785 194.860 ;
        RECT 82.955 194.305 83.505 194.690 ;
        RECT 84.145 194.480 84.335 195.245 ;
        RECT 84.645 195.165 84.895 196.305 ;
        RECT 85.085 195.665 85.335 196.085 ;
        RECT 85.565 195.835 85.895 196.305 ;
        RECT 86.125 195.665 86.375 196.085 ;
        RECT 85.085 195.495 86.375 195.665 ;
        RECT 86.555 195.665 86.885 196.095 ;
        RECT 86.555 195.495 87.010 195.665 ;
        RECT 85.075 194.995 85.290 195.325 ;
        RECT 84.505 194.665 84.815 194.995 ;
        RECT 84.985 194.665 85.290 194.995 ;
        RECT 85.465 194.665 85.750 195.325 ;
        RECT 85.945 194.665 86.210 195.325 ;
        RECT 86.425 194.665 86.670 195.325 ;
        RECT 84.645 194.495 84.815 194.665 ;
        RECT 86.840 194.495 87.010 195.495 ;
        RECT 82.615 193.965 83.505 194.135 ;
        RECT 83.675 193.755 83.965 194.480 ;
        RECT 84.145 193.970 84.475 194.480 ;
        RECT 84.645 194.325 87.010 194.495 ;
        RECT 87.355 195.505 87.795 196.135 ;
        RECT 87.355 194.495 87.665 195.505 ;
        RECT 87.970 195.455 88.285 196.305 ;
        RECT 88.455 195.965 89.885 196.135 ;
        RECT 88.455 195.285 88.625 195.965 ;
        RECT 87.835 195.115 88.625 195.285 ;
        RECT 87.835 194.665 88.005 195.115 ;
        RECT 88.795 194.995 88.995 195.795 ;
        RECT 88.175 194.665 88.565 194.945 ;
        RECT 88.750 194.665 88.995 194.995 ;
        RECT 89.195 194.665 89.445 195.795 ;
        RECT 89.635 195.335 89.885 195.965 ;
        RECT 90.065 195.505 90.395 196.305 ;
        RECT 91.120 195.685 91.295 196.135 ;
        RECT 91.465 195.865 91.795 196.305 ;
        RECT 92.100 195.715 92.270 196.135 ;
        RECT 92.505 195.895 93.175 196.305 ;
        RECT 93.390 195.715 93.560 196.135 ;
        RECT 93.760 195.895 94.090 196.305 ;
        RECT 91.120 195.515 91.750 195.685 ;
        RECT 89.635 195.165 90.405 195.335 ;
        RECT 89.660 194.665 90.065 194.995 ;
        RECT 90.235 194.495 90.405 195.165 ;
        RECT 91.035 194.665 91.400 195.345 ;
        RECT 91.580 194.995 91.750 195.515 ;
        RECT 92.100 195.545 94.115 195.715 ;
        RECT 91.580 194.665 91.930 194.995 ;
        RECT 91.580 194.495 91.750 194.665 ;
        RECT 84.645 193.755 84.975 194.155 ;
        RECT 86.025 193.985 86.355 194.325 ;
        RECT 86.525 193.755 86.855 194.155 ;
        RECT 87.355 193.935 87.795 194.495 ;
        RECT 87.965 193.755 88.415 194.495 ;
        RECT 88.585 194.325 89.745 194.495 ;
        RECT 88.585 193.925 88.755 194.325 ;
        RECT 88.925 193.755 89.345 194.155 ;
        RECT 89.515 193.925 89.745 194.325 ;
        RECT 89.915 193.925 90.405 194.495 ;
        RECT 91.120 194.325 91.750 194.495 ;
        RECT 91.120 193.925 91.295 194.325 ;
        RECT 92.100 194.255 92.270 195.545 ;
        RECT 91.465 193.755 91.795 194.135 ;
        RECT 92.040 193.925 92.270 194.255 ;
        RECT 92.470 194.090 92.750 195.365 ;
        RECT 92.975 194.265 93.245 195.365 ;
        RECT 93.435 194.335 93.775 195.365 ;
        RECT 93.945 194.995 94.115 195.545 ;
        RECT 94.285 195.165 94.545 196.135 ;
        RECT 93.945 194.665 94.205 194.995 ;
        RECT 94.375 194.475 94.545 195.165 ;
        RECT 92.935 194.095 93.245 194.265 ;
        RECT 92.975 194.090 93.245 194.095 ;
        RECT 93.705 193.755 94.035 194.135 ;
        RECT 94.205 194.010 94.545 194.475 ;
        RECT 94.715 195.165 94.975 196.135 ;
        RECT 95.170 195.895 95.500 196.305 ;
        RECT 95.700 195.715 95.870 196.135 ;
        RECT 96.085 195.895 96.755 196.305 ;
        RECT 96.990 195.715 97.160 196.135 ;
        RECT 97.465 195.865 97.795 196.305 ;
        RECT 95.145 195.545 97.160 195.715 ;
        RECT 97.965 195.685 98.140 196.135 ;
        RECT 94.715 194.475 94.885 195.165 ;
        RECT 95.145 194.995 95.315 195.545 ;
        RECT 95.055 194.665 95.315 194.995 ;
        RECT 94.715 194.010 95.055 194.475 ;
        RECT 95.485 194.335 95.825 195.365 ;
        RECT 96.015 195.285 96.285 195.365 ;
        RECT 96.015 195.115 96.325 195.285 ;
        RECT 94.205 193.965 94.540 194.010 ;
        RECT 94.720 193.965 95.055 194.010 ;
        RECT 95.225 193.755 95.555 194.135 ;
        RECT 96.015 194.090 96.285 195.115 ;
        RECT 96.510 194.090 96.790 195.365 ;
        RECT 96.990 194.255 97.160 195.545 ;
        RECT 97.510 195.515 98.140 195.685 ;
        RECT 98.970 195.675 99.255 196.135 ;
        RECT 99.425 195.845 99.695 196.305 ;
        RECT 97.510 194.995 97.680 195.515 ;
        RECT 98.970 195.455 99.925 195.675 ;
        RECT 97.330 194.665 97.680 194.995 ;
        RECT 97.860 194.665 98.225 195.345 ;
        RECT 98.855 194.725 99.545 195.285 ;
        RECT 97.510 194.495 97.680 194.665 ;
        RECT 99.715 194.555 99.925 195.455 ;
        RECT 97.510 194.325 98.140 194.495 ;
        RECT 96.990 193.925 97.220 194.255 ;
        RECT 97.465 193.755 97.795 194.135 ;
        RECT 97.965 193.925 98.140 194.325 ;
        RECT 98.970 194.385 99.925 194.555 ;
        RECT 100.095 195.285 100.495 196.135 ;
        RECT 100.685 195.675 100.965 196.135 ;
        RECT 101.485 195.845 101.810 196.305 ;
        RECT 100.685 195.455 101.810 195.675 ;
        RECT 100.095 194.725 101.190 195.285 ;
        RECT 101.360 194.995 101.810 195.455 ;
        RECT 101.980 195.165 102.365 196.135 ;
        RECT 103.000 195.925 103.335 196.305 ;
        RECT 98.970 193.925 99.255 194.385 ;
        RECT 99.425 193.755 99.695 194.215 ;
        RECT 100.095 193.925 100.495 194.725 ;
        RECT 101.360 194.665 101.915 194.995 ;
        RECT 101.360 194.555 101.810 194.665 ;
        RECT 100.685 194.385 101.810 194.555 ;
        RECT 102.085 194.495 102.365 195.165 ;
        RECT 100.685 193.925 100.965 194.385 ;
        RECT 101.485 193.755 101.810 194.215 ;
        RECT 101.980 193.925 102.365 194.495 ;
        RECT 102.995 194.435 103.235 195.745 ;
        RECT 103.505 195.335 103.755 196.135 ;
        RECT 103.975 195.585 104.305 196.305 ;
        RECT 104.490 195.335 104.740 196.135 ;
        RECT 105.205 195.505 105.535 196.305 ;
        RECT 105.705 195.875 106.045 196.135 ;
        RECT 103.405 195.165 105.595 195.335 ;
        RECT 103.405 194.255 103.575 195.165 ;
        RECT 105.280 194.995 105.595 195.165 ;
        RECT 103.080 193.925 103.575 194.255 ;
        RECT 103.795 194.030 104.145 194.995 ;
        RECT 104.325 194.025 104.625 194.995 ;
        RECT 104.805 194.025 105.085 194.995 ;
        RECT 105.280 194.745 105.610 194.995 ;
        RECT 105.265 193.755 105.535 194.555 ;
        RECT 105.785 194.475 106.045 195.875 ;
        RECT 106.215 195.165 106.475 196.305 ;
        RECT 106.715 195.795 108.330 196.125 ;
        RECT 106.725 194.995 106.895 195.555 ;
        RECT 107.155 195.455 108.330 195.625 ;
        RECT 108.500 195.505 108.780 196.305 ;
        RECT 107.155 195.165 107.485 195.455 ;
        RECT 108.160 195.335 108.330 195.455 ;
        RECT 107.655 194.995 107.900 195.285 ;
        RECT 108.160 195.165 108.820 195.335 ;
        RECT 108.990 195.165 109.265 196.135 ;
        RECT 108.650 194.995 108.820 195.165 ;
        RECT 106.220 194.745 106.555 194.995 ;
        RECT 106.725 194.665 107.440 194.995 ;
        RECT 107.655 194.665 108.480 194.995 ;
        RECT 108.650 194.665 108.925 194.995 ;
        RECT 106.725 194.575 106.975 194.665 ;
        RECT 105.705 193.965 106.045 194.475 ;
        RECT 106.215 193.755 106.475 194.575 ;
        RECT 106.645 194.155 106.975 194.575 ;
        RECT 108.650 194.495 108.820 194.665 ;
        RECT 107.155 194.325 108.820 194.495 ;
        RECT 109.095 194.430 109.265 195.165 ;
        RECT 109.435 195.140 109.725 196.305 ;
        RECT 109.895 195.795 111.085 196.085 ;
        RECT 109.915 195.455 111.085 195.625 ;
        RECT 111.255 195.505 111.535 196.305 ;
        RECT 109.915 195.165 110.240 195.455 ;
        RECT 110.915 195.335 111.085 195.455 ;
        RECT 110.410 194.995 110.605 195.285 ;
        RECT 110.915 195.165 111.575 195.335 ;
        RECT 111.745 195.165 112.020 196.135 ;
        RECT 112.195 195.870 117.540 196.305 ;
        RECT 117.715 195.870 123.060 196.305 ;
        RECT 123.700 195.880 124.035 196.305 ;
        RECT 111.405 194.995 111.575 195.165 ;
        RECT 109.895 194.665 110.240 194.995 ;
        RECT 110.410 194.665 111.235 194.995 ;
        RECT 111.405 194.665 111.680 194.995 ;
        RECT 111.405 194.495 111.575 194.665 ;
        RECT 107.155 193.925 107.415 194.325 ;
        RECT 107.585 193.755 107.915 194.155 ;
        RECT 108.085 193.975 108.255 194.325 ;
        RECT 108.425 193.755 108.800 194.155 ;
        RECT 108.990 194.085 109.265 194.430 ;
        RECT 109.435 193.755 109.725 194.480 ;
        RECT 109.910 194.325 111.575 194.495 ;
        RECT 111.850 194.430 112.020 195.165 ;
        RECT 109.910 193.975 110.165 194.325 ;
        RECT 110.335 193.755 110.665 194.155 ;
        RECT 110.835 193.975 111.005 194.325 ;
        RECT 111.175 193.755 111.555 194.155 ;
        RECT 111.745 194.085 112.020 194.430 ;
        RECT 113.780 194.300 114.120 195.130 ;
        RECT 115.600 194.620 115.950 195.870 ;
        RECT 119.300 194.300 119.640 195.130 ;
        RECT 121.120 194.620 121.470 195.870 ;
        RECT 124.205 195.700 124.390 196.105 ;
        RECT 123.725 195.525 124.390 195.700 ;
        RECT 124.595 195.525 124.925 196.305 ;
        RECT 123.725 194.495 124.065 195.525 ;
        RECT 125.095 195.335 125.365 196.105 ;
        RECT 124.235 195.165 125.365 195.335 ;
        RECT 125.595 195.245 125.925 196.090 ;
        RECT 126.095 195.295 126.265 196.305 ;
        RECT 126.435 195.575 126.775 196.135 ;
        RECT 127.005 195.805 127.320 196.305 ;
        RECT 127.500 195.835 128.385 196.005 ;
        RECT 124.235 194.665 124.485 195.165 ;
        RECT 123.725 194.325 124.410 194.495 ;
        RECT 124.665 194.415 125.025 194.995 ;
        RECT 112.195 193.755 117.540 194.300 ;
        RECT 117.715 193.755 123.060 194.300 ;
        RECT 123.700 193.755 124.035 194.155 ;
        RECT 124.205 193.925 124.410 194.325 ;
        RECT 125.195 194.255 125.365 195.165 ;
        RECT 125.535 195.165 125.925 195.245 ;
        RECT 126.435 195.200 127.330 195.575 ;
        RECT 125.535 195.115 125.750 195.165 ;
        RECT 125.535 194.535 125.705 195.115 ;
        RECT 126.435 194.995 126.625 195.200 ;
        RECT 127.500 194.995 127.670 195.835 ;
        RECT 128.610 195.805 128.860 196.135 ;
        RECT 125.875 194.665 126.625 194.995 ;
        RECT 126.795 194.665 127.670 194.995 ;
        RECT 125.535 194.495 125.760 194.535 ;
        RECT 126.425 194.495 126.625 194.665 ;
        RECT 125.535 194.410 125.915 194.495 ;
        RECT 124.620 193.755 124.895 194.235 ;
        RECT 125.105 193.925 125.365 194.255 ;
        RECT 125.585 193.975 125.915 194.410 ;
        RECT 126.085 193.755 126.255 194.365 ;
        RECT 126.425 193.970 126.755 194.495 ;
        RECT 127.015 193.755 127.225 194.285 ;
        RECT 127.500 194.205 127.670 194.665 ;
        RECT 127.840 194.705 128.160 195.665 ;
        RECT 128.330 194.915 128.520 195.635 ;
        RECT 128.690 194.735 128.860 195.805 ;
        RECT 129.030 195.505 129.200 196.305 ;
        RECT 129.370 195.860 130.475 196.030 ;
        RECT 129.370 195.245 129.540 195.860 ;
        RECT 130.685 195.710 130.935 196.135 ;
        RECT 131.105 195.845 131.370 196.305 ;
        RECT 129.710 195.325 130.240 195.690 ;
        RECT 130.685 195.580 130.990 195.710 ;
        RECT 129.030 195.155 129.540 195.245 ;
        RECT 129.030 194.985 129.900 195.155 ;
        RECT 129.030 194.915 129.200 194.985 ;
        RECT 129.320 194.735 129.520 194.765 ;
        RECT 127.840 194.375 128.305 194.705 ;
        RECT 128.690 194.435 129.520 194.735 ;
        RECT 128.690 194.205 128.860 194.435 ;
        RECT 127.500 194.035 128.285 194.205 ;
        RECT 128.455 194.035 128.860 194.205 ;
        RECT 129.040 193.755 129.410 194.255 ;
        RECT 129.730 194.205 129.900 194.985 ;
        RECT 130.070 194.625 130.240 195.325 ;
        RECT 130.410 194.795 130.650 195.390 ;
        RECT 130.070 194.405 130.595 194.625 ;
        RECT 130.820 194.475 130.990 195.580 ;
        RECT 130.765 194.345 130.990 194.475 ;
        RECT 131.160 194.385 131.440 195.335 ;
        RECT 130.765 194.205 130.935 194.345 ;
        RECT 129.730 194.035 130.405 194.205 ;
        RECT 130.600 194.035 130.935 194.205 ;
        RECT 131.105 193.755 131.355 194.215 ;
        RECT 131.610 194.015 131.795 196.135 ;
        RECT 131.965 195.805 132.295 196.305 ;
        RECT 132.465 195.635 132.635 196.135 ;
        RECT 131.970 195.465 132.635 195.635 ;
        RECT 131.970 194.475 132.200 195.465 ;
        RECT 132.370 194.645 132.720 195.295 ;
        RECT 132.895 195.230 133.165 196.135 ;
        RECT 133.335 195.545 133.665 196.305 ;
        RECT 133.845 195.375 134.025 196.135 ;
        RECT 131.970 194.305 132.635 194.475 ;
        RECT 131.965 193.755 132.295 194.135 ;
        RECT 132.465 194.015 132.635 194.305 ;
        RECT 132.895 194.430 133.075 195.230 ;
        RECT 133.350 195.205 134.025 195.375 ;
        RECT 133.350 195.060 133.520 195.205 ;
        RECT 135.195 195.140 135.485 196.305 ;
        RECT 135.735 195.375 135.915 196.135 ;
        RECT 136.095 195.545 136.425 196.305 ;
        RECT 135.735 195.205 136.410 195.375 ;
        RECT 136.595 195.230 136.865 196.135 ;
        RECT 133.245 194.730 133.520 195.060 ;
        RECT 136.240 195.060 136.410 195.205 ;
        RECT 133.350 194.475 133.520 194.730 ;
        RECT 133.745 194.655 134.085 195.025 ;
        RECT 135.675 194.655 136.015 195.025 ;
        RECT 136.240 194.730 136.515 195.060 ;
        RECT 132.895 193.925 133.155 194.430 ;
        RECT 133.350 194.305 134.015 194.475 ;
        RECT 133.335 193.755 133.665 194.135 ;
        RECT 133.845 193.925 134.015 194.305 ;
        RECT 135.195 193.755 135.485 194.480 ;
        RECT 136.240 194.475 136.410 194.730 ;
        RECT 135.745 194.305 136.410 194.475 ;
        RECT 136.685 194.430 136.865 195.230 ;
        RECT 137.115 195.375 137.295 196.135 ;
        RECT 137.475 195.545 137.805 196.305 ;
        RECT 137.115 195.205 137.790 195.375 ;
        RECT 137.975 195.230 138.245 196.135 ;
        RECT 139.335 195.795 139.595 196.305 ;
        RECT 137.620 195.060 137.790 195.205 ;
        RECT 137.055 194.655 137.395 195.025 ;
        RECT 137.620 194.730 137.895 195.060 ;
        RECT 137.620 194.475 137.790 194.730 ;
        RECT 135.745 193.925 135.915 194.305 ;
        RECT 136.095 193.755 136.425 194.135 ;
        RECT 136.605 193.925 136.865 194.430 ;
        RECT 137.125 194.305 137.790 194.475 ;
        RECT 138.065 194.430 138.245 195.230 ;
        RECT 139.335 194.745 139.675 195.625 ;
        RECT 139.845 194.915 140.015 196.135 ;
        RECT 140.255 195.800 140.870 196.305 ;
        RECT 140.255 195.265 140.505 195.630 ;
        RECT 140.675 195.625 140.870 195.800 ;
        RECT 141.040 195.795 141.515 196.135 ;
        RECT 141.685 195.760 141.900 196.305 ;
        RECT 140.675 195.435 141.005 195.625 ;
        RECT 141.225 195.265 141.940 195.560 ;
        RECT 142.110 195.435 142.385 196.135 ;
        RECT 140.255 195.095 142.045 195.265 ;
        RECT 139.845 194.665 140.640 194.915 ;
        RECT 139.845 194.575 140.095 194.665 ;
        RECT 137.125 193.925 137.295 194.305 ;
        RECT 137.475 193.755 137.805 194.135 ;
        RECT 137.985 193.925 138.245 194.430 ;
        RECT 139.335 193.755 139.595 194.575 ;
        RECT 139.765 194.155 140.095 194.575 ;
        RECT 140.810 194.240 141.065 195.095 ;
        RECT 140.275 193.975 141.065 194.240 ;
        RECT 141.235 194.395 141.645 194.915 ;
        RECT 141.815 194.665 142.045 195.095 ;
        RECT 142.215 194.405 142.385 195.435 ;
        RECT 142.555 195.215 145.145 196.305 ;
        RECT 141.235 193.975 141.435 194.395 ;
        RECT 141.625 193.755 141.955 194.215 ;
        RECT 142.125 193.925 142.385 194.405 ;
        RECT 142.555 194.525 143.765 195.045 ;
        RECT 143.935 194.695 145.145 195.215 ;
        RECT 145.405 195.375 145.575 196.135 ;
        RECT 145.755 195.545 146.085 196.305 ;
        RECT 145.405 195.205 146.070 195.375 ;
        RECT 146.255 195.230 146.525 196.135 ;
        RECT 147.245 195.635 147.415 196.135 ;
        RECT 147.585 195.805 147.915 196.305 ;
        RECT 147.245 195.465 147.910 195.635 ;
        RECT 145.900 195.060 146.070 195.205 ;
        RECT 145.335 194.655 145.665 195.025 ;
        RECT 145.900 194.730 146.185 195.060 ;
        RECT 142.555 193.755 145.145 194.525 ;
        RECT 145.900 194.475 146.070 194.730 ;
        RECT 145.405 194.305 146.070 194.475 ;
        RECT 146.355 194.430 146.525 195.230 ;
        RECT 147.160 194.645 147.510 195.295 ;
        RECT 147.680 194.475 147.910 195.465 ;
        RECT 145.405 193.925 145.575 194.305 ;
        RECT 145.755 193.755 146.085 194.135 ;
        RECT 146.265 193.925 146.525 194.430 ;
        RECT 147.245 194.305 147.910 194.475 ;
        RECT 147.245 194.015 147.415 194.305 ;
        RECT 147.585 193.755 147.915 194.135 ;
        RECT 148.085 194.015 148.270 196.135 ;
        RECT 148.510 195.845 148.775 196.305 ;
        RECT 148.945 195.710 149.195 196.135 ;
        RECT 149.405 195.860 150.510 196.030 ;
        RECT 148.890 195.580 149.195 195.710 ;
        RECT 148.440 194.385 148.720 195.335 ;
        RECT 148.890 194.475 149.060 195.580 ;
        RECT 149.230 194.795 149.470 195.390 ;
        RECT 149.640 195.325 150.170 195.690 ;
        RECT 149.640 194.625 149.810 195.325 ;
        RECT 150.340 195.245 150.510 195.860 ;
        RECT 150.680 195.505 150.850 196.305 ;
        RECT 151.020 195.805 151.270 196.135 ;
        RECT 151.495 195.835 152.380 196.005 ;
        RECT 150.340 195.155 150.850 195.245 ;
        RECT 148.890 194.345 149.115 194.475 ;
        RECT 149.285 194.405 149.810 194.625 ;
        RECT 149.980 194.985 150.850 195.155 ;
        RECT 148.525 193.755 148.775 194.215 ;
        RECT 148.945 194.205 149.115 194.345 ;
        RECT 149.980 194.205 150.150 194.985 ;
        RECT 150.680 194.915 150.850 194.985 ;
        RECT 150.360 194.735 150.560 194.765 ;
        RECT 151.020 194.735 151.190 195.805 ;
        RECT 151.360 194.915 151.550 195.635 ;
        RECT 150.360 194.435 151.190 194.735 ;
        RECT 151.720 194.705 152.040 195.665 ;
        RECT 148.945 194.035 149.280 194.205 ;
        RECT 149.475 194.035 150.150 194.205 ;
        RECT 150.470 193.755 150.840 194.255 ;
        RECT 151.020 194.205 151.190 194.435 ;
        RECT 151.575 194.375 152.040 194.705 ;
        RECT 152.210 194.995 152.380 195.835 ;
        RECT 152.560 195.805 152.875 196.305 ;
        RECT 153.105 195.575 153.445 196.135 ;
        RECT 152.550 195.200 153.445 195.575 ;
        RECT 153.615 195.295 153.785 196.305 ;
        RECT 153.255 194.995 153.445 195.200 ;
        RECT 153.955 195.245 154.285 196.090 ;
        RECT 153.955 195.165 154.345 195.245 ;
        RECT 154.130 195.115 154.345 195.165 ;
        RECT 152.210 194.665 153.085 194.995 ;
        RECT 153.255 194.665 154.005 194.995 ;
        RECT 152.210 194.205 152.380 194.665 ;
        RECT 153.255 194.495 153.455 194.665 ;
        RECT 154.175 194.535 154.345 195.115 ;
        RECT 154.975 195.215 156.185 196.305 ;
        RECT 154.975 194.675 155.495 195.215 ;
        RECT 154.120 194.495 154.345 194.535 ;
        RECT 155.665 194.505 156.185 195.045 ;
        RECT 151.020 194.035 151.425 194.205 ;
        RECT 151.595 194.035 152.380 194.205 ;
        RECT 152.655 193.755 152.865 194.285 ;
        RECT 153.125 193.970 153.455 194.495 ;
        RECT 153.965 194.410 154.345 194.495 ;
        RECT 153.625 193.755 153.795 194.365 ;
        RECT 153.965 193.975 154.295 194.410 ;
        RECT 154.975 193.755 156.185 194.505 ;
        RECT 70.710 193.585 156.270 193.755 ;
        RECT 70.795 192.835 72.005 193.585 ;
        RECT 70.795 192.295 71.315 192.835 ;
        RECT 72.175 192.815 74.765 193.585 ;
        RECT 74.940 193.055 75.230 193.405 ;
        RECT 75.425 193.225 75.755 193.585 ;
        RECT 75.925 193.055 76.155 193.360 ;
        RECT 74.940 192.885 76.155 193.055 ;
        RECT 76.345 192.905 76.515 193.280 ;
        RECT 76.800 193.195 77.130 193.585 ;
        RECT 77.300 193.025 77.525 193.405 ;
        RECT 71.485 192.125 72.005 192.665 ;
        RECT 72.175 192.295 73.385 192.815 ;
        RECT 76.345 192.735 76.545 192.905 ;
        RECT 76.345 192.715 76.515 192.735 ;
        RECT 73.555 192.125 74.765 192.645 ;
        RECT 75.000 192.565 75.260 192.675 ;
        RECT 74.995 192.395 75.260 192.565 ;
        RECT 75.000 192.345 75.260 192.395 ;
        RECT 75.440 192.345 75.825 192.675 ;
        RECT 75.995 192.545 76.515 192.715 ;
        RECT 70.795 191.035 72.005 192.125 ;
        RECT 72.175 191.035 74.765 192.125 ;
        RECT 74.940 191.035 75.260 192.175 ;
        RECT 75.440 191.295 75.635 192.345 ;
        RECT 75.995 192.165 76.165 192.545 ;
        RECT 75.815 191.885 76.165 192.165 ;
        RECT 76.355 192.015 76.600 192.375 ;
        RECT 76.785 192.345 77.025 192.995 ;
        RECT 77.195 192.845 77.525 193.025 ;
        RECT 77.195 192.175 77.370 192.845 ;
        RECT 77.725 192.675 77.955 193.295 ;
        RECT 78.135 192.855 78.435 193.585 ;
        RECT 78.615 192.835 79.825 193.585 ;
        RECT 80.005 192.860 80.335 193.370 ;
        RECT 80.505 193.185 80.835 193.585 ;
        RECT 81.885 193.015 82.215 193.355 ;
        RECT 82.385 193.185 82.715 193.585 ;
        RECT 77.540 192.345 77.955 192.675 ;
        RECT 78.135 192.345 78.430 192.675 ;
        RECT 78.615 192.295 79.135 192.835 ;
        RECT 76.785 191.985 77.370 192.175 ;
        RECT 75.815 191.205 76.145 191.885 ;
        RECT 76.345 191.035 76.600 191.835 ;
        RECT 76.785 191.215 77.060 191.985 ;
        RECT 77.540 191.815 78.435 192.145 ;
        RECT 79.305 192.125 79.825 192.665 ;
        RECT 77.230 191.645 78.435 191.815 ;
        RECT 77.230 191.215 77.560 191.645 ;
        RECT 77.730 191.035 77.925 191.475 ;
        RECT 78.105 191.215 78.435 191.645 ;
        RECT 78.615 191.035 79.825 192.125 ;
        RECT 80.005 192.095 80.195 192.860 ;
        RECT 80.505 192.845 82.870 193.015 ;
        RECT 80.505 192.675 80.675 192.845 ;
        RECT 80.365 192.345 80.675 192.675 ;
        RECT 80.845 192.345 81.150 192.675 ;
        RECT 80.005 191.245 80.335 192.095 ;
        RECT 80.505 191.035 80.755 192.175 ;
        RECT 80.935 192.015 81.150 192.345 ;
        RECT 81.325 192.015 81.610 192.675 ;
        RECT 81.805 192.015 82.070 192.675 ;
        RECT 82.285 192.015 82.530 192.675 ;
        RECT 82.700 191.845 82.870 192.845 ;
        RECT 80.945 191.675 82.235 191.845 ;
        RECT 80.945 191.255 81.195 191.675 ;
        RECT 81.425 191.035 81.755 191.505 ;
        RECT 81.985 191.255 82.235 191.675 ;
        RECT 82.415 191.675 82.870 191.845 ;
        RECT 83.215 192.845 83.475 193.415 ;
        RECT 83.645 193.185 84.030 193.585 ;
        RECT 84.200 193.015 84.455 193.415 ;
        RECT 83.645 192.845 84.455 193.015 ;
        RECT 84.645 192.845 84.890 193.415 ;
        RECT 85.060 193.185 85.445 193.585 ;
        RECT 85.615 193.015 85.870 193.415 ;
        RECT 85.060 192.845 85.870 193.015 ;
        RECT 86.060 192.845 86.485 193.415 ;
        RECT 86.655 193.185 87.040 193.585 ;
        RECT 87.210 193.015 87.645 193.415 ;
        RECT 86.655 192.845 87.645 193.015 ;
        RECT 88.360 193.035 88.535 193.325 ;
        RECT 88.705 193.205 89.035 193.585 ;
        RECT 88.360 192.865 88.855 193.035 ;
        RECT 89.210 192.905 89.425 193.275 ;
        RECT 89.660 193.135 90.260 193.305 ;
        RECT 83.215 192.175 83.400 192.845 ;
        RECT 83.645 192.675 83.995 192.845 ;
        RECT 84.645 192.675 84.815 192.845 ;
        RECT 85.060 192.675 85.410 192.845 ;
        RECT 86.060 192.675 86.410 192.845 ;
        RECT 86.655 192.675 86.990 192.845 ;
        RECT 83.570 192.345 83.995 192.675 ;
        RECT 82.415 191.245 82.745 191.675 ;
        RECT 83.215 191.205 83.475 192.175 ;
        RECT 83.645 191.825 83.995 192.345 ;
        RECT 84.165 192.175 84.815 192.675 ;
        RECT 84.985 192.345 85.410 192.675 ;
        RECT 84.165 191.995 84.890 192.175 ;
        RECT 83.645 191.630 84.455 191.825 ;
        RECT 83.645 191.035 84.030 191.460 ;
        RECT 84.200 191.205 84.455 191.630 ;
        RECT 84.645 191.205 84.890 191.995 ;
        RECT 85.060 191.825 85.410 192.345 ;
        RECT 85.580 192.175 86.410 192.675 ;
        RECT 86.580 192.345 86.990 192.675 ;
        RECT 85.580 191.995 86.485 192.175 ;
        RECT 85.060 191.630 85.890 191.825 ;
        RECT 85.060 191.035 85.445 191.460 ;
        RECT 85.615 191.205 85.890 191.630 ;
        RECT 86.060 191.205 86.485 191.995 ;
        RECT 86.655 191.800 86.990 192.345 ;
        RECT 87.160 191.970 87.645 192.675 ;
        RECT 88.335 191.925 88.515 192.695 ;
        RECT 88.685 191.885 88.855 192.865 ;
        RECT 89.025 192.575 89.425 192.905 ;
        RECT 89.595 192.635 89.920 192.965 ;
        RECT 89.410 192.225 89.580 192.385 ;
        RECT 89.195 192.055 89.580 192.225 ;
        RECT 89.750 192.095 89.920 192.635 ;
        RECT 90.090 192.435 90.260 193.135 ;
        RECT 90.640 193.125 90.970 193.585 ;
        RECT 91.175 193.205 91.605 193.375 ;
        RECT 90.430 192.655 90.805 192.955 ;
        RECT 90.090 192.265 90.430 192.435 ;
        RECT 90.600 192.350 90.805 192.655 ;
        RECT 90.975 192.350 91.265 192.955 ;
        RECT 91.435 192.610 91.605 193.205 ;
        RECT 91.775 192.995 92.010 193.325 ;
        RECT 89.750 191.885 90.090 192.095 ;
        RECT 86.655 191.630 87.645 191.800 ;
        RECT 88.685 191.755 90.090 191.885 ;
        RECT 86.655 191.035 87.040 191.460 ;
        RECT 87.210 191.205 87.645 191.630 ;
        RECT 88.365 191.715 90.090 191.755 ;
        RECT 88.365 191.585 88.855 191.715 ;
        RECT 88.365 191.295 88.535 191.585 ;
        RECT 90.260 191.545 90.430 192.265 ;
        RECT 91.435 192.280 91.670 192.610 ;
        RECT 91.435 192.180 91.605 192.280 ;
        RECT 91.335 192.010 91.605 192.180 ;
        RECT 91.335 191.885 91.505 192.010 ;
        RECT 91.160 191.715 91.505 191.885 ;
        RECT 91.840 191.860 92.010 192.995 ;
        RECT 88.705 191.035 89.035 191.415 ;
        RECT 89.600 191.375 90.430 191.545 ;
        RECT 90.785 191.035 91.015 191.615 ;
        RECT 91.755 191.545 92.010 191.860 ;
        RECT 91.495 191.375 92.010 191.545 ;
        RECT 92.180 191.545 92.370 193.325 ;
        RECT 92.585 193.085 92.790 193.415 ;
        RECT 92.985 193.125 93.315 193.585 ;
        RECT 93.515 193.205 94.410 193.375 ;
        RECT 92.585 192.105 92.755 193.085 ;
        RECT 92.935 192.275 93.305 192.955 ;
        RECT 93.515 192.105 93.685 193.205 ;
        RECT 92.585 191.935 93.685 192.105 ;
        RECT 92.585 191.775 92.775 191.935 ;
        RECT 92.180 191.375 92.705 191.545 ;
        RECT 92.945 191.035 93.290 191.665 ;
        RECT 93.515 191.515 93.685 191.935 ;
        RECT 93.855 192.635 94.475 192.965 ;
        RECT 94.725 192.675 95.035 193.295 ;
        RECT 95.205 192.855 95.455 193.585 ;
        RECT 95.625 192.945 95.955 193.405 ;
        RECT 93.855 191.685 94.145 192.635 ;
        RECT 94.725 192.595 95.135 192.675 ;
        RECT 94.315 192.025 94.655 192.425 ;
        RECT 94.825 192.345 95.135 192.595 ;
        RECT 95.305 192.345 95.615 192.675 ;
        RECT 95.305 192.175 95.475 192.345 ;
        RECT 95.785 192.175 95.955 192.945 ;
        RECT 96.125 192.785 96.380 193.585 ;
        RECT 96.555 192.860 96.845 193.585 ;
        RECT 94.865 192.005 95.475 192.175 ;
        RECT 94.865 191.545 95.035 192.005 ;
        RECT 95.645 191.835 95.955 192.175 ;
        RECT 93.515 191.345 94.465 191.515 ;
        RECT 94.715 191.375 95.035 191.545 ;
        RECT 95.205 191.035 95.375 191.835 ;
        RECT 95.545 191.215 95.955 191.835 ;
        RECT 96.125 191.035 96.375 192.175 ;
        RECT 96.555 191.035 96.845 192.200 ;
        RECT 97.015 191.205 97.275 193.415 ;
        RECT 97.445 193.205 97.775 193.585 ;
        RECT 97.985 192.675 98.180 193.250 ;
        RECT 98.450 192.675 98.635 193.255 ;
        RECT 97.445 191.755 97.615 192.675 ;
        RECT 97.925 192.345 98.180 192.675 ;
        RECT 98.405 192.345 98.635 192.675 ;
        RECT 98.885 193.245 100.365 193.415 ;
        RECT 98.885 192.345 99.055 193.245 ;
        RECT 99.225 192.745 99.775 193.075 ;
        RECT 99.965 192.915 100.365 193.245 ;
        RECT 100.545 193.205 100.875 193.585 ;
        RECT 101.185 193.085 101.445 193.415 ;
        RECT 97.985 192.035 98.180 192.345 ;
        RECT 98.450 192.035 98.635 192.345 ;
        RECT 99.225 191.755 99.395 192.745 ;
        RECT 99.965 192.435 100.135 192.915 ;
        RECT 100.715 192.725 100.925 192.905 ;
        RECT 100.305 192.555 100.925 192.725 ;
        RECT 97.445 191.585 99.395 191.755 ;
        RECT 99.565 192.265 100.135 192.435 ;
        RECT 101.275 192.385 101.445 193.085 ;
        RECT 99.565 191.755 99.735 192.265 ;
        RECT 100.315 192.215 101.445 192.385 ;
        RECT 100.315 192.095 100.485 192.215 ;
        RECT 99.905 191.925 100.485 192.095 ;
        RECT 99.565 191.585 100.305 191.755 ;
        RECT 100.755 191.715 101.105 192.045 ;
        RECT 97.445 191.035 97.775 191.415 ;
        RECT 98.200 191.205 98.370 191.585 ;
        RECT 98.630 191.035 98.960 191.415 ;
        RECT 99.155 191.205 99.325 191.585 ;
        RECT 99.535 191.035 99.865 191.415 ;
        RECT 100.115 191.205 100.305 191.585 ;
        RECT 101.275 191.535 101.445 192.215 ;
        RECT 100.545 191.035 100.875 191.415 ;
        RECT 101.185 191.205 101.445 191.535 ;
        RECT 102.075 192.845 102.390 193.220 ;
        RECT 102.645 192.845 102.815 193.585 ;
        RECT 103.065 193.015 103.235 193.220 ;
        RECT 103.460 193.185 103.835 193.585 ;
        RECT 104.005 193.015 104.175 193.365 ;
        RECT 104.360 193.185 104.690 193.585 ;
        RECT 104.860 193.015 105.030 193.365 ;
        RECT 105.200 193.185 105.580 193.585 ;
        RECT 103.065 192.845 103.565 193.015 ;
        RECT 104.005 192.845 105.600 193.015 ;
        RECT 105.770 192.910 106.045 193.255 ;
        RECT 102.075 191.805 102.245 192.845 ;
        RECT 102.415 191.975 102.765 192.675 ;
        RECT 102.935 192.345 103.225 192.675 ;
        RECT 103.395 192.595 103.565 192.845 ;
        RECT 105.430 192.675 105.600 192.845 ;
        RECT 103.395 192.425 103.820 192.595 ;
        RECT 103.395 192.145 103.565 192.425 ;
        RECT 104.215 192.255 104.385 192.675 ;
        RECT 104.605 192.345 105.260 192.675 ;
        RECT 105.430 192.345 105.705 192.675 ;
        RECT 102.980 191.975 103.565 192.145 ;
        RECT 103.735 192.085 104.385 192.255 ;
        RECT 105.430 192.175 105.600 192.345 ;
        RECT 105.875 192.175 106.045 192.910 ;
        RECT 106.300 193.035 106.475 193.325 ;
        RECT 106.645 193.205 106.975 193.585 ;
        RECT 106.300 192.865 106.795 193.035 ;
        RECT 107.150 192.905 107.365 193.275 ;
        RECT 107.600 193.135 108.200 193.305 ;
        RECT 103.735 191.805 103.905 192.085 ;
        RECT 104.940 192.005 105.600 192.175 ;
        RECT 104.940 191.885 105.110 192.005 ;
        RECT 102.075 191.635 103.905 191.805 ;
        RECT 104.075 191.715 105.110 191.885 ;
        RECT 102.075 191.215 102.335 191.635 ;
        RECT 104.075 191.465 104.245 191.715 ;
        RECT 102.505 191.035 102.835 191.465 ;
        RECT 103.500 191.295 104.245 191.465 ;
        RECT 104.470 191.215 105.110 191.545 ;
        RECT 105.280 191.035 105.560 191.835 ;
        RECT 105.770 191.205 106.045 192.175 ;
        RECT 106.275 191.925 106.455 192.695 ;
        RECT 106.625 191.885 106.795 192.865 ;
        RECT 106.965 192.575 107.365 192.905 ;
        RECT 107.535 192.635 107.860 192.965 ;
        RECT 107.350 192.225 107.520 192.385 ;
        RECT 107.135 192.055 107.520 192.225 ;
        RECT 107.690 192.095 107.860 192.635 ;
        RECT 108.030 192.435 108.200 193.135 ;
        RECT 108.580 193.125 108.910 193.585 ;
        RECT 109.115 193.205 109.545 193.375 ;
        RECT 108.370 192.655 108.745 192.955 ;
        RECT 108.030 192.265 108.370 192.435 ;
        RECT 108.540 192.350 108.745 192.655 ;
        RECT 108.915 192.350 109.205 192.955 ;
        RECT 109.375 192.610 109.545 193.205 ;
        RECT 109.715 192.995 109.950 193.325 ;
        RECT 107.690 191.885 108.030 192.095 ;
        RECT 106.625 191.755 108.030 191.885 ;
        RECT 106.305 191.715 108.030 191.755 ;
        RECT 106.305 191.585 106.795 191.715 ;
        RECT 106.305 191.295 106.475 191.585 ;
        RECT 108.200 191.545 108.370 192.265 ;
        RECT 109.375 192.280 109.610 192.610 ;
        RECT 109.375 192.180 109.545 192.280 ;
        RECT 109.275 192.010 109.545 192.180 ;
        RECT 109.275 191.885 109.445 192.010 ;
        RECT 109.100 191.715 109.445 191.885 ;
        RECT 109.780 191.860 109.950 192.995 ;
        RECT 106.645 191.035 106.975 191.415 ;
        RECT 107.540 191.375 108.370 191.545 ;
        RECT 108.725 191.035 108.955 191.615 ;
        RECT 109.695 191.545 109.950 191.860 ;
        RECT 109.435 191.375 109.950 191.545 ;
        RECT 110.120 191.545 110.310 193.325 ;
        RECT 110.525 193.085 110.730 193.415 ;
        RECT 110.925 193.125 111.255 193.585 ;
        RECT 111.455 193.205 112.350 193.375 ;
        RECT 110.525 192.105 110.695 193.085 ;
        RECT 110.875 192.275 111.245 192.955 ;
        RECT 111.455 192.105 111.625 193.205 ;
        RECT 110.525 191.935 111.625 192.105 ;
        RECT 110.525 191.775 110.715 191.935 ;
        RECT 110.120 191.375 110.645 191.545 ;
        RECT 110.885 191.035 111.230 191.665 ;
        RECT 111.455 191.515 111.625 191.935 ;
        RECT 111.795 192.635 112.415 192.965 ;
        RECT 112.665 192.675 112.975 193.295 ;
        RECT 113.145 192.855 113.395 193.585 ;
        RECT 113.565 192.945 113.895 193.405 ;
        RECT 111.795 191.685 112.085 192.635 ;
        RECT 112.665 192.595 113.075 192.675 ;
        RECT 112.255 192.025 112.595 192.425 ;
        RECT 112.765 192.345 113.075 192.595 ;
        RECT 113.245 192.345 113.555 192.675 ;
        RECT 113.245 192.175 113.415 192.345 ;
        RECT 113.725 192.175 113.895 192.945 ;
        RECT 114.065 192.785 114.320 193.585 ;
        RECT 114.955 193.085 115.215 193.415 ;
        RECT 115.425 193.105 115.700 193.585 ;
        RECT 114.955 192.175 115.125 193.085 ;
        RECT 115.910 193.015 116.115 193.415 ;
        RECT 116.285 193.185 116.620 193.585 ;
        RECT 115.295 192.345 115.655 192.925 ;
        RECT 115.910 192.845 116.595 193.015 ;
        RECT 115.835 192.175 116.085 192.675 ;
        RECT 112.805 192.005 113.415 192.175 ;
        RECT 112.805 191.545 112.975 192.005 ;
        RECT 113.585 191.835 113.895 192.175 ;
        RECT 111.455 191.345 112.405 191.515 ;
        RECT 112.655 191.375 112.975 191.545 ;
        RECT 113.145 191.035 113.315 191.835 ;
        RECT 113.485 191.215 113.895 191.835 ;
        RECT 114.065 191.035 114.315 192.175 ;
        RECT 114.955 192.005 116.085 192.175 ;
        RECT 114.955 191.235 115.225 192.005 ;
        RECT 116.255 191.815 116.595 192.845 ;
        RECT 116.795 192.815 118.465 193.585 ;
        RECT 118.635 192.910 118.905 193.255 ;
        RECT 119.095 193.185 119.475 193.585 ;
        RECT 119.645 193.015 119.815 193.365 ;
        RECT 119.985 193.185 120.315 193.585 ;
        RECT 120.515 193.015 120.685 193.365 ;
        RECT 120.885 193.085 121.215 193.585 ;
        RECT 116.795 192.295 117.545 192.815 ;
        RECT 117.715 192.125 118.465 192.645 ;
        RECT 115.395 191.035 115.725 191.815 ;
        RECT 115.930 191.640 116.595 191.815 ;
        RECT 115.930 191.235 116.115 191.640 ;
        RECT 116.285 191.035 116.620 191.460 ;
        RECT 116.795 191.035 118.465 192.125 ;
        RECT 118.635 192.175 118.805 192.910 ;
        RECT 119.075 192.845 120.685 193.015 ;
        RECT 119.075 192.675 119.245 192.845 ;
        RECT 118.975 192.345 119.245 192.675 ;
        RECT 119.415 192.345 119.820 192.675 ;
        RECT 119.075 192.175 119.245 192.345 ;
        RECT 119.990 192.225 120.700 192.675 ;
        RECT 120.870 192.345 121.220 192.915 ;
        RECT 122.315 192.860 122.605 193.585 ;
        RECT 122.865 193.035 123.035 193.415 ;
        RECT 123.215 193.205 123.545 193.585 ;
        RECT 122.865 192.865 123.530 193.035 ;
        RECT 123.725 192.910 123.985 193.415 ;
        RECT 122.795 192.315 123.135 192.685 ;
        RECT 123.360 192.610 123.530 192.865 ;
        RECT 123.360 192.280 123.635 192.610 ;
        RECT 118.635 191.205 118.905 192.175 ;
        RECT 119.075 192.005 119.800 192.175 ;
        RECT 119.990 192.055 120.705 192.225 ;
        RECT 119.630 191.885 119.800 192.005 ;
        RECT 120.900 191.885 121.220 192.175 ;
        RECT 119.115 191.035 119.395 191.835 ;
        RECT 119.630 191.715 121.220 191.885 ;
        RECT 119.565 191.255 121.220 191.545 ;
        RECT 122.315 191.035 122.605 192.200 ;
        RECT 123.360 192.135 123.530 192.280 ;
        RECT 122.855 191.965 123.530 192.135 ;
        RECT 123.805 192.110 123.985 192.910 ;
        RECT 124.155 192.815 125.825 193.585 ;
        RECT 126.455 193.125 127.015 193.415 ;
        RECT 127.185 193.125 127.435 193.585 ;
        RECT 124.155 192.295 124.905 192.815 ;
        RECT 125.075 192.125 125.825 192.645 ;
        RECT 122.855 191.205 123.035 191.965 ;
        RECT 123.215 191.035 123.545 191.795 ;
        RECT 123.715 191.205 123.985 192.110 ;
        RECT 124.155 191.035 125.825 192.125 ;
        RECT 126.455 191.755 126.705 193.125 ;
        RECT 128.055 192.955 128.385 193.315 ;
        RECT 126.995 192.765 128.385 192.955 ;
        RECT 128.755 192.765 129.015 193.585 ;
        RECT 129.185 192.765 129.515 193.185 ;
        RECT 129.695 193.100 130.485 193.365 ;
        RECT 126.995 192.675 127.165 192.765 ;
        RECT 126.875 192.345 127.165 192.675 ;
        RECT 129.265 192.675 129.515 192.765 ;
        RECT 127.335 192.345 127.675 192.595 ;
        RECT 127.895 192.345 128.570 192.595 ;
        RECT 126.995 192.095 127.165 192.345 ;
        RECT 126.995 191.925 127.935 192.095 ;
        RECT 128.305 191.985 128.570 192.345 ;
        RECT 126.455 191.205 126.915 191.755 ;
        RECT 127.105 191.035 127.435 191.755 ;
        RECT 127.635 191.375 127.935 191.925 ;
        RECT 128.755 191.715 129.095 192.595 ;
        RECT 129.265 192.425 130.060 192.675 ;
        RECT 128.105 191.035 128.385 191.705 ;
        RECT 128.755 191.035 129.015 191.545 ;
        RECT 129.265 191.205 129.435 192.425 ;
        RECT 130.230 192.245 130.485 193.100 ;
        RECT 130.655 192.945 130.855 193.365 ;
        RECT 131.045 193.125 131.375 193.585 ;
        RECT 130.655 192.425 131.065 192.945 ;
        RECT 131.545 192.935 131.805 193.415 ;
        RECT 131.235 192.245 131.465 192.675 ;
        RECT 129.675 192.075 131.465 192.245 ;
        RECT 129.675 191.710 129.925 192.075 ;
        RECT 130.095 191.715 130.425 191.905 ;
        RECT 130.645 191.780 131.360 192.075 ;
        RECT 131.635 191.905 131.805 192.935 ;
        RECT 132.065 193.035 132.235 193.415 ;
        RECT 132.415 193.205 132.745 193.585 ;
        RECT 132.065 192.865 132.730 193.035 ;
        RECT 132.925 192.910 133.185 193.415 ;
        RECT 131.995 192.315 132.335 192.685 ;
        RECT 132.560 192.610 132.730 192.865 ;
        RECT 132.560 192.280 132.835 192.610 ;
        RECT 132.560 192.135 132.730 192.280 ;
        RECT 130.095 191.540 130.290 191.715 ;
        RECT 129.675 191.035 130.290 191.540 ;
        RECT 130.460 191.205 130.935 191.545 ;
        RECT 131.105 191.035 131.320 191.580 ;
        RECT 131.530 191.205 131.805 191.905 ;
        RECT 132.055 191.965 132.730 192.135 ;
        RECT 133.005 192.110 133.185 192.910 ;
        RECT 133.355 192.815 135.945 193.585 ;
        RECT 136.600 193.195 136.930 193.585 ;
        RECT 137.100 193.025 137.325 193.405 ;
        RECT 133.355 192.295 134.565 192.815 ;
        RECT 134.735 192.125 135.945 192.645 ;
        RECT 136.585 192.345 136.825 192.995 ;
        RECT 136.995 192.845 137.325 193.025 ;
        RECT 136.995 192.175 137.170 192.845 ;
        RECT 137.525 192.675 137.755 193.295 ;
        RECT 137.935 192.855 138.235 193.585 ;
        RECT 139.425 193.035 139.595 193.325 ;
        RECT 139.765 193.205 140.095 193.585 ;
        RECT 139.425 192.865 140.090 193.035 ;
        RECT 137.340 192.345 137.755 192.675 ;
        RECT 137.935 192.345 138.230 192.675 ;
        RECT 132.055 191.205 132.235 191.965 ;
        RECT 132.415 191.035 132.745 191.795 ;
        RECT 132.915 191.205 133.185 192.110 ;
        RECT 133.355 191.035 135.945 192.125 ;
        RECT 136.585 191.985 137.170 192.175 ;
        RECT 136.585 191.215 136.860 191.985 ;
        RECT 137.340 191.815 138.235 192.145 ;
        RECT 139.340 192.045 139.690 192.695 ;
        RECT 139.860 191.875 140.090 192.865 ;
        RECT 137.030 191.645 138.235 191.815 ;
        RECT 137.030 191.215 137.360 191.645 ;
        RECT 137.530 191.035 137.725 191.475 ;
        RECT 137.905 191.215 138.235 191.645 ;
        RECT 139.425 191.705 140.090 191.875 ;
        RECT 139.425 191.205 139.595 191.705 ;
        RECT 139.765 191.035 140.095 191.535 ;
        RECT 140.265 191.205 140.450 193.325 ;
        RECT 140.705 193.125 140.955 193.585 ;
        RECT 141.125 193.135 141.460 193.305 ;
        RECT 141.655 193.135 142.330 193.305 ;
        RECT 141.125 192.995 141.295 193.135 ;
        RECT 140.620 192.005 140.900 192.955 ;
        RECT 141.070 192.865 141.295 192.995 ;
        RECT 141.070 191.760 141.240 192.865 ;
        RECT 141.465 192.715 141.990 192.935 ;
        RECT 141.410 191.950 141.650 192.545 ;
        RECT 141.820 192.015 141.990 192.715 ;
        RECT 142.160 192.355 142.330 193.135 ;
        RECT 142.650 193.085 143.020 193.585 ;
        RECT 143.200 193.135 143.605 193.305 ;
        RECT 143.775 193.135 144.560 193.305 ;
        RECT 143.200 192.905 143.370 193.135 ;
        RECT 142.540 192.605 143.370 192.905 ;
        RECT 143.755 192.635 144.220 192.965 ;
        RECT 142.540 192.575 142.740 192.605 ;
        RECT 142.860 192.355 143.030 192.425 ;
        RECT 142.160 192.185 143.030 192.355 ;
        RECT 142.520 192.095 143.030 192.185 ;
        RECT 141.070 191.630 141.375 191.760 ;
        RECT 141.820 191.650 142.350 192.015 ;
        RECT 140.690 191.035 140.955 191.495 ;
        RECT 141.125 191.205 141.375 191.630 ;
        RECT 142.520 191.480 142.690 192.095 ;
        RECT 141.585 191.310 142.690 191.480 ;
        RECT 142.860 191.035 143.030 191.835 ;
        RECT 143.200 191.535 143.370 192.605 ;
        RECT 143.540 191.705 143.730 192.425 ;
        RECT 143.900 191.675 144.220 192.635 ;
        RECT 144.390 192.675 144.560 193.135 ;
        RECT 144.835 193.055 145.045 193.585 ;
        RECT 145.305 192.845 145.635 193.370 ;
        RECT 145.805 192.975 145.975 193.585 ;
        RECT 146.145 192.930 146.475 193.365 ;
        RECT 146.145 192.845 146.525 192.930 ;
        RECT 145.435 192.675 145.635 192.845 ;
        RECT 146.300 192.805 146.525 192.845 ;
        RECT 144.390 192.345 145.265 192.675 ;
        RECT 145.435 192.345 146.185 192.675 ;
        RECT 143.200 191.205 143.450 191.535 ;
        RECT 144.390 191.505 144.560 192.345 ;
        RECT 145.435 192.140 145.625 192.345 ;
        RECT 146.355 192.225 146.525 192.805 ;
        RECT 146.310 192.175 146.525 192.225 ;
        RECT 144.730 191.765 145.625 192.140 ;
        RECT 146.135 192.095 146.525 192.175 ;
        RECT 146.695 192.910 146.955 193.415 ;
        RECT 147.135 193.205 147.465 193.585 ;
        RECT 147.645 193.035 147.815 193.415 ;
        RECT 146.695 192.110 146.875 192.910 ;
        RECT 147.150 192.865 147.815 193.035 ;
        RECT 147.150 192.610 147.320 192.865 ;
        RECT 148.075 192.860 148.365 193.585 ;
        RECT 148.535 193.040 153.880 193.585 ;
        RECT 147.045 192.280 147.320 192.610 ;
        RECT 147.545 192.315 147.885 192.685 ;
        RECT 147.150 192.135 147.320 192.280 ;
        RECT 150.120 192.210 150.460 193.040 ;
        RECT 154.975 192.835 156.185 193.585 ;
        RECT 143.675 191.335 144.560 191.505 ;
        RECT 144.740 191.035 145.055 191.535 ;
        RECT 145.285 191.205 145.625 191.765 ;
        RECT 145.795 191.035 145.965 192.045 ;
        RECT 146.135 191.250 146.465 192.095 ;
        RECT 146.695 191.205 146.965 192.110 ;
        RECT 147.150 191.965 147.825 192.135 ;
        RECT 147.135 191.035 147.465 191.795 ;
        RECT 147.645 191.205 147.825 191.965 ;
        RECT 148.075 191.035 148.365 192.200 ;
        RECT 151.940 191.470 152.290 192.720 ;
        RECT 154.975 192.125 155.495 192.665 ;
        RECT 155.665 192.295 156.185 192.835 ;
        RECT 148.535 191.035 153.880 191.470 ;
        RECT 154.975 191.035 156.185 192.125 ;
        RECT 70.710 190.865 156.270 191.035 ;
        RECT 70.795 189.775 72.005 190.865 ;
        RECT 72.175 190.430 77.520 190.865 ;
        RECT 70.795 189.065 71.315 189.605 ;
        RECT 71.485 189.235 72.005 189.775 ;
        RECT 70.795 188.315 72.005 189.065 ;
        RECT 73.760 188.860 74.100 189.690 ;
        RECT 75.580 189.180 75.930 190.430 ;
        RECT 77.695 189.775 80.285 190.865 ;
        RECT 77.695 189.085 78.905 189.605 ;
        RECT 79.075 189.255 80.285 189.775 ;
        RECT 80.915 190.145 81.375 190.695 ;
        RECT 81.565 190.145 81.895 190.865 ;
        RECT 72.175 188.315 77.520 188.860 ;
        RECT 77.695 188.315 80.285 189.085 ;
        RECT 80.915 188.775 81.165 190.145 ;
        RECT 82.095 189.975 82.395 190.525 ;
        RECT 82.565 190.195 82.845 190.865 ;
        RECT 81.455 189.805 82.395 189.975 ;
        RECT 81.455 189.555 81.625 189.805 ;
        RECT 82.765 189.555 83.030 189.915 ;
        RECT 83.675 189.700 83.965 190.865 ;
        RECT 84.215 189.935 84.395 190.695 ;
        RECT 84.575 190.105 84.905 190.865 ;
        RECT 84.215 189.765 84.890 189.935 ;
        RECT 85.075 189.790 85.345 190.695 ;
        RECT 84.720 189.620 84.890 189.765 ;
        RECT 81.335 189.225 81.625 189.555 ;
        RECT 81.795 189.305 82.135 189.555 ;
        RECT 82.355 189.305 83.030 189.555 ;
        RECT 81.455 189.135 81.625 189.225 ;
        RECT 84.155 189.215 84.495 189.585 ;
        RECT 84.720 189.290 84.995 189.620 ;
        RECT 81.455 188.945 82.845 189.135 ;
        RECT 80.915 188.485 81.475 188.775 ;
        RECT 81.645 188.315 81.895 188.775 ;
        RECT 82.515 188.585 82.845 188.945 ;
        RECT 83.675 188.315 83.965 189.040 ;
        RECT 84.720 189.035 84.890 189.290 ;
        RECT 84.225 188.865 84.890 189.035 ;
        RECT 85.165 188.990 85.345 189.790 ;
        RECT 85.525 189.725 85.855 190.865 ;
        RECT 86.385 189.895 86.715 190.680 ;
        RECT 86.035 189.725 86.715 189.895 ;
        RECT 86.905 189.805 87.235 190.655 ;
        RECT 85.515 189.305 85.865 189.555 ;
        RECT 86.035 189.125 86.205 189.725 ;
        RECT 86.375 189.305 86.725 189.555 ;
        RECT 84.225 188.485 84.395 188.865 ;
        RECT 84.575 188.315 84.905 188.695 ;
        RECT 85.085 188.485 85.345 188.990 ;
        RECT 85.525 188.315 85.795 189.125 ;
        RECT 85.965 188.485 86.295 189.125 ;
        RECT 86.465 188.315 86.705 189.125 ;
        RECT 86.905 189.040 87.095 189.805 ;
        RECT 87.405 189.725 87.655 190.865 ;
        RECT 87.845 190.225 88.095 190.645 ;
        RECT 88.325 190.395 88.655 190.865 ;
        RECT 88.885 190.225 89.135 190.645 ;
        RECT 87.845 190.055 89.135 190.225 ;
        RECT 89.315 190.225 89.645 190.655 ;
        RECT 89.315 190.055 89.770 190.225 ;
        RECT 87.835 189.555 88.050 189.885 ;
        RECT 87.265 189.225 87.575 189.555 ;
        RECT 87.745 189.225 88.050 189.555 ;
        RECT 88.225 189.225 88.510 189.885 ;
        RECT 88.705 189.225 88.970 189.885 ;
        RECT 89.185 189.225 89.430 189.885 ;
        RECT 87.405 189.055 87.575 189.225 ;
        RECT 89.600 189.055 89.770 190.055 ;
        RECT 90.195 189.935 90.375 190.695 ;
        RECT 90.555 190.105 90.885 190.865 ;
        RECT 90.195 189.765 90.870 189.935 ;
        RECT 91.055 189.790 91.325 190.695 ;
        RECT 90.700 189.620 90.870 189.765 ;
        RECT 90.135 189.215 90.475 189.585 ;
        RECT 90.700 189.290 90.975 189.620 ;
        RECT 86.905 188.530 87.235 189.040 ;
        RECT 87.405 188.885 89.770 189.055 ;
        RECT 90.700 189.035 90.870 189.290 ;
        RECT 87.405 188.315 87.735 188.715 ;
        RECT 88.785 188.545 89.115 188.885 ;
        RECT 90.205 188.865 90.870 189.035 ;
        RECT 91.145 188.990 91.325 189.790 ;
        RECT 91.585 189.755 91.835 190.865 ;
        RECT 92.015 189.895 92.275 190.695 ;
        RECT 92.445 190.065 92.775 190.865 ;
        RECT 92.945 189.895 93.135 190.695 ;
        RECT 93.305 190.070 93.635 190.865 ;
        RECT 93.805 189.895 93.985 190.695 ;
        RECT 94.165 190.065 94.495 190.865 ;
        RECT 94.720 190.505 95.910 190.695 ;
        RECT 94.720 190.065 94.980 190.505 ;
        RECT 95.225 189.895 95.415 190.335 ;
        RECT 92.015 189.725 95.415 189.895 ;
        RECT 95.650 189.915 95.910 190.505 ;
        RECT 96.080 190.085 96.340 190.865 ;
        RECT 96.510 189.915 96.770 190.695 ;
        RECT 95.650 189.745 96.770 189.915 ;
        RECT 97.015 189.775 98.225 190.865 ;
        RECT 91.495 189.305 91.835 189.585 ;
        RECT 92.015 189.135 92.275 189.725 ;
        RECT 92.455 189.305 93.200 189.555 ;
        RECT 93.610 189.305 94.595 189.555 ;
        RECT 94.775 189.305 95.865 189.555 ;
        RECT 96.045 189.305 96.845 189.555 ;
        RECT 89.285 188.315 89.615 188.715 ;
        RECT 90.205 188.485 90.375 188.865 ;
        RECT 90.555 188.315 90.885 188.695 ;
        RECT 91.065 188.485 91.325 188.990 ;
        RECT 91.585 188.675 91.845 189.095 ;
        RECT 92.015 188.845 92.345 189.135 ;
        RECT 92.525 188.965 93.685 189.135 ;
        RECT 92.525 188.675 92.710 188.965 ;
        RECT 93.335 188.850 93.685 188.965 ;
        RECT 93.860 188.885 96.845 189.070 ;
        RECT 91.585 188.490 92.710 188.675 ;
        RECT 92.880 188.760 93.170 188.795 ;
        RECT 92.880 188.675 93.185 188.760 ;
        RECT 94.290 188.675 94.620 188.715 ;
        RECT 92.880 188.485 94.620 188.675 ;
        RECT 94.790 188.595 94.980 188.885 ;
        RECT 95.650 188.880 96.845 188.885 ;
        RECT 95.150 188.315 95.480 188.715 ;
        RECT 95.650 188.595 95.840 188.880 ;
        RECT 96.010 188.315 96.340 188.710 ;
        RECT 96.510 188.595 96.845 188.880 ;
        RECT 97.015 189.065 97.535 189.605 ;
        RECT 97.705 189.235 98.225 189.775 ;
        RECT 98.395 190.265 98.655 190.685 ;
        RECT 98.825 190.435 99.155 190.865 ;
        RECT 99.820 190.435 100.565 190.605 ;
        RECT 98.395 190.095 100.225 190.265 ;
        RECT 97.015 188.315 98.225 189.065 ;
        RECT 98.395 189.055 98.565 190.095 ;
        RECT 98.735 189.225 99.085 189.925 ;
        RECT 99.300 189.755 99.885 189.925 ;
        RECT 99.255 189.225 99.545 189.555 ;
        RECT 99.715 189.475 99.885 189.755 ;
        RECT 100.055 189.815 100.225 190.095 ;
        RECT 100.395 190.185 100.565 190.435 ;
        RECT 100.790 190.355 101.430 190.685 ;
        RECT 100.395 190.015 101.430 190.185 ;
        RECT 101.600 190.065 101.880 190.865 ;
        RECT 101.260 189.895 101.430 190.015 ;
        RECT 100.055 189.645 100.705 189.815 ;
        RECT 101.260 189.725 101.920 189.895 ;
        RECT 102.090 189.725 102.365 190.695 ;
        RECT 102.615 189.935 102.795 190.695 ;
        RECT 102.975 190.105 103.305 190.865 ;
        RECT 102.615 189.765 103.290 189.935 ;
        RECT 103.475 189.790 103.745 190.695 ;
        RECT 99.715 189.305 100.140 189.475 ;
        RECT 99.715 189.055 99.885 189.305 ;
        RECT 100.535 189.225 100.705 189.645 ;
        RECT 101.750 189.555 101.920 189.725 ;
        RECT 100.925 189.225 101.580 189.555 ;
        RECT 101.750 189.225 102.025 189.555 ;
        RECT 101.750 189.055 101.920 189.225 ;
        RECT 98.395 188.680 98.710 189.055 ;
        RECT 98.965 188.315 99.135 189.055 ;
        RECT 99.385 188.885 99.885 189.055 ;
        RECT 100.325 188.885 101.920 189.055 ;
        RECT 102.195 188.990 102.365 189.725 ;
        RECT 103.120 189.620 103.290 189.765 ;
        RECT 102.555 189.215 102.895 189.585 ;
        RECT 103.120 189.290 103.395 189.620 ;
        RECT 103.120 189.035 103.290 189.290 ;
        RECT 99.385 188.680 99.555 188.885 ;
        RECT 99.780 188.315 100.155 188.715 ;
        RECT 100.325 188.535 100.495 188.885 ;
        RECT 100.680 188.315 101.010 188.715 ;
        RECT 101.180 188.535 101.350 188.885 ;
        RECT 101.520 188.315 101.900 188.715 ;
        RECT 102.090 188.645 102.365 188.990 ;
        RECT 102.625 188.865 103.290 189.035 ;
        RECT 103.565 188.990 103.745 189.790 ;
        RECT 102.625 188.485 102.795 188.865 ;
        RECT 102.975 188.315 103.305 188.695 ;
        RECT 103.485 188.485 103.745 188.990 ;
        RECT 103.915 189.725 104.190 190.695 ;
        RECT 104.400 190.065 104.680 190.865 ;
        RECT 104.850 190.355 105.490 190.685 ;
        RECT 105.715 190.435 106.460 190.605 ;
        RECT 107.125 190.435 107.455 190.865 ;
        RECT 105.715 190.185 105.885 190.435 ;
        RECT 107.625 190.265 107.885 190.685 ;
        RECT 104.850 190.015 105.885 190.185 ;
        RECT 106.055 190.095 107.885 190.265 ;
        RECT 104.850 189.895 105.020 190.015 ;
        RECT 104.360 189.725 105.020 189.895 ;
        RECT 106.055 189.815 106.225 190.095 ;
        RECT 103.915 188.990 104.085 189.725 ;
        RECT 104.360 189.555 104.530 189.725 ;
        RECT 105.575 189.645 106.225 189.815 ;
        RECT 106.395 189.755 106.980 189.925 ;
        RECT 104.255 189.225 104.530 189.555 ;
        RECT 104.700 189.225 105.355 189.555 ;
        RECT 105.575 189.225 105.745 189.645 ;
        RECT 106.395 189.475 106.565 189.755 ;
        RECT 106.140 189.305 106.565 189.475 ;
        RECT 104.360 189.055 104.530 189.225 ;
        RECT 106.395 189.055 106.565 189.305 ;
        RECT 106.735 189.225 107.025 189.555 ;
        RECT 107.195 189.225 107.545 189.925 ;
        RECT 107.715 189.055 107.885 190.095 ;
        RECT 108.055 189.775 109.265 190.865 ;
        RECT 103.915 188.645 104.190 188.990 ;
        RECT 104.360 188.885 105.955 189.055 ;
        RECT 106.395 188.885 106.895 189.055 ;
        RECT 104.380 188.315 104.760 188.715 ;
        RECT 104.930 188.535 105.100 188.885 ;
        RECT 105.270 188.315 105.600 188.715 ;
        RECT 105.785 188.535 105.955 188.885 ;
        RECT 106.125 188.315 106.500 188.715 ;
        RECT 106.725 188.680 106.895 188.885 ;
        RECT 107.145 188.315 107.315 189.055 ;
        RECT 107.570 188.680 107.885 189.055 ;
        RECT 108.055 189.065 108.575 189.605 ;
        RECT 108.745 189.235 109.265 189.775 ;
        RECT 109.435 189.700 109.725 190.865 ;
        RECT 109.895 189.790 110.165 190.695 ;
        RECT 110.335 190.105 110.665 190.865 ;
        RECT 110.845 189.935 111.025 190.695 ;
        RECT 108.055 188.315 109.265 189.065 ;
        RECT 109.435 188.315 109.725 189.040 ;
        RECT 109.895 188.990 110.075 189.790 ;
        RECT 110.350 189.765 111.025 189.935 ;
        RECT 112.275 189.935 112.455 190.695 ;
        RECT 112.635 190.105 112.965 190.865 ;
        RECT 112.275 189.765 112.950 189.935 ;
        RECT 113.135 189.790 113.405 190.695 ;
        RECT 114.125 190.315 114.295 190.605 ;
        RECT 114.465 190.485 114.795 190.865 ;
        RECT 115.360 190.355 116.190 190.525 ;
        RECT 114.125 190.185 114.615 190.315 ;
        RECT 114.125 190.145 115.850 190.185 ;
        RECT 114.445 190.015 115.850 190.145 ;
        RECT 110.350 189.620 110.520 189.765 ;
        RECT 110.245 189.290 110.520 189.620 ;
        RECT 112.780 189.620 112.950 189.765 ;
        RECT 110.350 189.035 110.520 189.290 ;
        RECT 110.745 189.215 111.085 189.585 ;
        RECT 112.215 189.215 112.555 189.585 ;
        RECT 112.780 189.290 113.055 189.620 ;
        RECT 112.780 189.035 112.950 189.290 ;
        RECT 109.895 188.485 110.155 188.990 ;
        RECT 110.350 188.865 111.015 189.035 ;
        RECT 110.335 188.315 110.665 188.695 ;
        RECT 110.845 188.485 111.015 188.865 ;
        RECT 112.285 188.865 112.950 189.035 ;
        RECT 113.225 188.990 113.405 189.790 ;
        RECT 114.095 189.205 114.275 189.975 ;
        RECT 114.445 189.035 114.615 190.015 ;
        RECT 114.955 189.675 115.340 189.845 ;
        RECT 115.170 189.515 115.340 189.675 ;
        RECT 115.510 189.805 115.850 190.015 ;
        RECT 112.285 188.485 112.455 188.865 ;
        RECT 112.635 188.315 112.965 188.695 ;
        RECT 113.145 188.485 113.405 188.990 ;
        RECT 114.120 188.865 114.615 189.035 ;
        RECT 114.785 188.995 115.185 189.325 ;
        RECT 115.510 189.265 115.680 189.805 ;
        RECT 116.020 189.635 116.190 190.355 ;
        RECT 116.545 190.285 116.775 190.865 ;
        RECT 117.255 190.355 117.770 190.525 ;
        RECT 116.920 190.015 117.265 190.185 ;
        RECT 117.515 190.040 117.770 190.355 ;
        RECT 117.095 189.890 117.265 190.015 ;
        RECT 117.095 189.720 117.365 189.890 ;
        RECT 114.120 188.575 114.295 188.865 ;
        RECT 114.465 188.315 114.795 188.695 ;
        RECT 114.970 188.625 115.185 188.995 ;
        RECT 115.355 188.935 115.680 189.265 ;
        RECT 115.850 189.465 116.190 189.635 ;
        RECT 117.195 189.620 117.365 189.720 ;
        RECT 115.850 188.765 116.020 189.465 ;
        RECT 116.360 189.245 116.565 189.550 ;
        RECT 116.190 188.945 116.565 189.245 ;
        RECT 116.735 188.945 117.025 189.550 ;
        RECT 117.195 189.290 117.430 189.620 ;
        RECT 115.420 188.595 116.020 188.765 ;
        RECT 116.400 188.315 116.730 188.775 ;
        RECT 117.195 188.695 117.365 189.290 ;
        RECT 117.600 188.905 117.770 190.040 ;
        RECT 116.935 188.525 117.365 188.695 ;
        RECT 117.535 188.575 117.770 188.905 ;
        RECT 117.940 190.355 118.465 190.525 ;
        RECT 117.940 188.575 118.130 190.355 ;
        RECT 118.705 190.235 119.050 190.865 ;
        RECT 119.275 190.385 120.225 190.555 ;
        RECT 118.345 189.965 118.535 190.125 ;
        RECT 119.275 189.965 119.445 190.385 ;
        RECT 120.475 190.355 120.795 190.525 ;
        RECT 118.345 189.795 119.445 189.965 ;
        RECT 118.345 188.815 118.515 189.795 ;
        RECT 118.695 188.945 119.065 189.625 ;
        RECT 118.345 188.485 118.550 188.815 ;
        RECT 118.745 188.315 119.075 188.775 ;
        RECT 119.275 188.695 119.445 189.795 ;
        RECT 119.615 189.265 119.905 190.215 ;
        RECT 120.625 189.895 120.795 190.355 ;
        RECT 120.965 190.065 121.135 190.865 ;
        RECT 121.305 190.065 121.715 190.685 ;
        RECT 120.075 189.475 120.415 189.875 ;
        RECT 120.625 189.725 121.235 189.895 ;
        RECT 121.405 189.725 121.715 190.065 ;
        RECT 121.885 189.725 122.135 190.865 ;
        RECT 122.315 189.995 122.590 190.695 ;
        RECT 122.760 190.320 123.015 190.865 ;
        RECT 123.185 190.355 123.665 190.695 ;
        RECT 123.840 190.310 124.445 190.865 ;
        RECT 123.830 190.210 124.445 190.310 ;
        RECT 123.830 190.185 124.015 190.210 ;
        RECT 121.065 189.555 121.235 189.725 ;
        RECT 120.585 189.305 120.895 189.555 ;
        RECT 119.615 188.935 120.235 189.265 ;
        RECT 120.485 189.225 120.895 189.305 ;
        RECT 121.065 189.225 121.375 189.555 ;
        RECT 119.275 188.525 120.170 188.695 ;
        RECT 120.485 188.605 120.795 189.225 ;
        RECT 120.965 188.315 121.215 189.045 ;
        RECT 121.545 188.955 121.715 189.725 ;
        RECT 121.385 188.495 121.715 188.955 ;
        RECT 121.885 188.315 122.140 189.115 ;
        RECT 122.315 188.965 122.485 189.995 ;
        RECT 122.760 189.865 123.515 190.115 ;
        RECT 123.685 189.940 124.015 190.185 ;
        RECT 122.760 189.830 123.530 189.865 ;
        RECT 122.760 189.820 123.545 189.830 ;
        RECT 122.655 189.805 123.550 189.820 ;
        RECT 122.655 189.790 123.570 189.805 ;
        RECT 122.655 189.780 123.590 189.790 ;
        RECT 122.655 189.770 123.615 189.780 ;
        RECT 122.655 189.740 123.685 189.770 ;
        RECT 122.655 189.710 123.705 189.740 ;
        RECT 122.655 189.680 123.725 189.710 ;
        RECT 122.655 189.655 123.755 189.680 ;
        RECT 122.655 189.620 123.790 189.655 ;
        RECT 122.655 189.615 123.820 189.620 ;
        RECT 122.655 189.220 122.885 189.615 ;
        RECT 123.430 189.610 123.820 189.615 ;
        RECT 123.455 189.600 123.820 189.610 ;
        RECT 123.470 189.595 123.820 189.600 ;
        RECT 123.485 189.590 123.820 189.595 ;
        RECT 124.185 189.590 124.445 190.040 ;
        RECT 123.485 189.585 124.445 189.590 ;
        RECT 123.495 189.575 124.445 189.585 ;
        RECT 123.505 189.570 124.445 189.575 ;
        RECT 123.515 189.560 124.445 189.570 ;
        RECT 123.520 189.550 124.445 189.560 ;
        RECT 123.525 189.545 124.445 189.550 ;
        RECT 123.535 189.530 124.445 189.545 ;
        RECT 123.540 189.515 124.445 189.530 ;
        RECT 123.550 189.490 124.445 189.515 ;
        RECT 123.055 189.020 123.385 189.445 ;
        RECT 122.315 188.485 122.575 188.965 ;
        RECT 122.745 188.315 122.995 188.855 ;
        RECT 123.165 188.535 123.385 189.020 ;
        RECT 123.555 189.420 124.445 189.490 ;
        RECT 124.615 189.895 124.885 190.665 ;
        RECT 125.055 190.085 125.385 190.865 ;
        RECT 125.590 190.260 125.775 190.665 ;
        RECT 125.945 190.440 126.280 190.865 ;
        RECT 125.590 190.085 126.255 190.260 ;
        RECT 124.615 189.725 125.745 189.895 ;
        RECT 123.555 188.695 123.725 189.420 ;
        RECT 123.895 188.865 124.445 189.250 ;
        RECT 124.615 188.815 124.785 189.725 ;
        RECT 124.955 188.975 125.315 189.555 ;
        RECT 125.495 189.225 125.745 189.725 ;
        RECT 125.915 189.055 126.255 190.085 ;
        RECT 125.570 188.885 126.255 189.055 ;
        RECT 126.455 189.790 126.725 190.695 ;
        RECT 126.895 190.105 127.225 190.865 ;
        RECT 127.405 189.935 127.585 190.695 ;
        RECT 126.455 188.990 126.635 189.790 ;
        RECT 126.910 189.765 127.585 189.935 ;
        RECT 127.835 189.790 128.105 190.695 ;
        RECT 128.275 190.105 128.605 190.865 ;
        RECT 128.785 189.935 128.965 190.695 ;
        RECT 126.910 189.620 127.080 189.765 ;
        RECT 126.805 189.290 127.080 189.620 ;
        RECT 126.910 189.035 127.080 189.290 ;
        RECT 127.305 189.215 127.645 189.585 ;
        RECT 123.555 188.525 124.445 188.695 ;
        RECT 124.615 188.485 124.875 188.815 ;
        RECT 125.085 188.315 125.360 188.795 ;
        RECT 125.570 188.485 125.775 188.885 ;
        RECT 125.945 188.315 126.280 188.715 ;
        RECT 126.455 188.485 126.715 188.990 ;
        RECT 126.910 188.865 127.575 189.035 ;
        RECT 126.895 188.315 127.225 188.695 ;
        RECT 127.405 188.485 127.575 188.865 ;
        RECT 127.835 188.990 128.015 189.790 ;
        RECT 128.290 189.765 128.965 189.935 ;
        RECT 129.295 189.935 129.475 190.695 ;
        RECT 129.655 190.105 129.985 190.865 ;
        RECT 129.295 189.765 129.970 189.935 ;
        RECT 130.155 189.790 130.425 190.695 ;
        RECT 128.290 189.620 128.460 189.765 ;
        RECT 128.185 189.290 128.460 189.620 ;
        RECT 129.800 189.620 129.970 189.765 ;
        RECT 128.290 189.035 128.460 189.290 ;
        RECT 128.685 189.215 129.025 189.585 ;
        RECT 129.235 189.215 129.575 189.585 ;
        RECT 129.800 189.290 130.075 189.620 ;
        RECT 129.800 189.035 129.970 189.290 ;
        RECT 127.835 188.485 128.095 188.990 ;
        RECT 128.290 188.865 128.955 189.035 ;
        RECT 128.275 188.315 128.605 188.695 ;
        RECT 128.785 188.485 128.955 188.865 ;
        RECT 129.305 188.865 129.970 189.035 ;
        RECT 130.245 188.990 130.425 189.790 ;
        RECT 129.305 188.485 129.475 188.865 ;
        RECT 129.655 188.315 129.985 188.695 ;
        RECT 130.165 188.485 130.425 188.990 ;
        RECT 130.595 190.145 131.055 190.695 ;
        RECT 131.245 190.145 131.575 190.865 ;
        RECT 130.595 188.775 130.845 190.145 ;
        RECT 131.775 189.975 132.075 190.525 ;
        RECT 132.245 190.195 132.525 190.865 ;
        RECT 131.135 189.805 132.075 189.975 ;
        RECT 131.135 189.555 131.305 189.805 ;
        RECT 132.445 189.555 132.710 189.915 ;
        RECT 131.015 189.225 131.305 189.555 ;
        RECT 131.475 189.305 131.815 189.555 ;
        RECT 132.035 189.305 132.710 189.555 ;
        RECT 132.895 189.790 133.165 190.695 ;
        RECT 133.335 190.105 133.665 190.865 ;
        RECT 133.845 189.935 134.025 190.695 ;
        RECT 131.135 189.135 131.305 189.225 ;
        RECT 131.135 188.945 132.525 189.135 ;
        RECT 130.595 188.485 131.155 188.775 ;
        RECT 131.325 188.315 131.575 188.775 ;
        RECT 132.195 188.585 132.525 188.945 ;
        RECT 132.895 188.990 133.075 189.790 ;
        RECT 133.350 189.765 134.025 189.935 ;
        RECT 133.350 189.620 133.520 189.765 ;
        RECT 135.195 189.700 135.485 190.865 ;
        RECT 135.660 190.065 135.915 190.865 ;
        RECT 136.115 190.015 136.445 190.695 ;
        RECT 133.245 189.290 133.520 189.620 ;
        RECT 133.350 189.035 133.520 189.290 ;
        RECT 133.745 189.215 134.085 189.585 ;
        RECT 135.660 189.525 135.905 189.885 ;
        RECT 136.095 189.735 136.445 190.015 ;
        RECT 136.095 189.355 136.265 189.735 ;
        RECT 136.625 189.555 136.820 190.605 ;
        RECT 137.000 189.725 137.320 190.865 ;
        RECT 137.530 190.075 138.065 190.695 ;
        RECT 135.745 189.185 136.265 189.355 ;
        RECT 136.435 189.225 136.820 189.555 ;
        RECT 137.000 189.505 137.260 189.555 ;
        RECT 137.000 189.335 137.265 189.505 ;
        RECT 137.000 189.225 137.260 189.335 ;
        RECT 132.895 188.485 133.155 188.990 ;
        RECT 133.350 188.865 134.015 189.035 ;
        RECT 133.335 188.315 133.665 188.695 ;
        RECT 133.845 188.485 134.015 188.865 ;
        RECT 135.195 188.315 135.485 189.040 ;
        RECT 135.745 188.620 135.915 189.185 ;
        RECT 137.530 189.055 137.845 190.075 ;
        RECT 138.235 190.065 138.565 190.865 ;
        RECT 139.885 190.195 140.055 190.695 ;
        RECT 140.225 190.365 140.555 190.865 ;
        RECT 139.050 189.895 139.440 190.070 ;
        RECT 139.885 190.025 140.550 190.195 ;
        RECT 138.015 189.725 139.440 189.895 ;
        RECT 138.015 189.225 138.185 189.725 ;
        RECT 136.105 188.845 137.320 189.015 ;
        RECT 136.105 188.540 136.335 188.845 ;
        RECT 136.505 188.315 136.835 188.675 ;
        RECT 137.030 188.495 137.320 188.845 ;
        RECT 137.530 188.485 138.145 189.055 ;
        RECT 138.435 188.995 138.700 189.555 ;
        RECT 138.870 188.825 139.040 189.725 ;
        RECT 139.210 188.995 139.565 189.555 ;
        RECT 139.800 189.205 140.150 189.855 ;
        RECT 140.320 189.035 140.550 190.025 ;
        RECT 139.885 188.865 140.550 189.035 ;
        RECT 138.315 188.315 138.530 188.825 ;
        RECT 138.760 188.495 139.040 188.825 ;
        RECT 139.220 188.315 139.460 188.825 ;
        RECT 139.885 188.575 140.055 188.865 ;
        RECT 140.225 188.315 140.555 188.695 ;
        RECT 140.725 188.575 140.910 190.695 ;
        RECT 141.150 190.405 141.415 190.865 ;
        RECT 141.585 190.270 141.835 190.695 ;
        RECT 142.045 190.420 143.150 190.590 ;
        RECT 141.530 190.140 141.835 190.270 ;
        RECT 141.080 188.945 141.360 189.895 ;
        RECT 141.530 189.035 141.700 190.140 ;
        RECT 141.870 189.355 142.110 189.950 ;
        RECT 142.280 189.885 142.810 190.250 ;
        RECT 142.280 189.185 142.450 189.885 ;
        RECT 142.980 189.805 143.150 190.420 ;
        RECT 143.320 190.065 143.490 190.865 ;
        RECT 143.660 190.365 143.910 190.695 ;
        RECT 144.135 190.395 145.020 190.565 ;
        RECT 142.980 189.715 143.490 189.805 ;
        RECT 141.530 188.905 141.755 189.035 ;
        RECT 141.925 188.965 142.450 189.185 ;
        RECT 142.620 189.545 143.490 189.715 ;
        RECT 141.165 188.315 141.415 188.775 ;
        RECT 141.585 188.765 141.755 188.905 ;
        RECT 142.620 188.765 142.790 189.545 ;
        RECT 143.320 189.475 143.490 189.545 ;
        RECT 143.000 189.295 143.200 189.325 ;
        RECT 143.660 189.295 143.830 190.365 ;
        RECT 144.000 189.475 144.190 190.195 ;
        RECT 143.000 188.995 143.830 189.295 ;
        RECT 144.360 189.265 144.680 190.225 ;
        RECT 141.585 188.595 141.920 188.765 ;
        RECT 142.115 188.595 142.790 188.765 ;
        RECT 143.110 188.315 143.480 188.815 ;
        RECT 143.660 188.765 143.830 188.995 ;
        RECT 144.215 188.935 144.680 189.265 ;
        RECT 144.850 189.555 145.020 190.395 ;
        RECT 145.200 190.365 145.515 190.865 ;
        RECT 145.745 190.135 146.085 190.695 ;
        RECT 145.190 189.760 146.085 190.135 ;
        RECT 146.255 189.855 146.425 190.865 ;
        RECT 145.895 189.555 146.085 189.760 ;
        RECT 146.595 189.805 146.925 190.650 ;
        RECT 147.155 190.015 147.535 190.695 ;
        RECT 148.125 190.015 148.295 190.865 ;
        RECT 148.465 190.185 148.795 190.695 ;
        RECT 148.965 190.355 149.135 190.865 ;
        RECT 149.305 190.185 149.705 190.695 ;
        RECT 148.465 190.015 149.705 190.185 ;
        RECT 146.595 189.725 146.985 189.805 ;
        RECT 146.770 189.675 146.985 189.725 ;
        RECT 144.850 189.225 145.725 189.555 ;
        RECT 145.895 189.225 146.645 189.555 ;
        RECT 144.850 188.765 145.020 189.225 ;
        RECT 145.895 189.055 146.095 189.225 ;
        RECT 146.815 189.095 146.985 189.675 ;
        RECT 146.760 189.055 146.985 189.095 ;
        RECT 143.660 188.595 144.065 188.765 ;
        RECT 144.235 188.595 145.020 188.765 ;
        RECT 145.295 188.315 145.505 188.845 ;
        RECT 145.765 188.530 146.095 189.055 ;
        RECT 146.605 188.970 146.985 189.055 ;
        RECT 147.155 189.055 147.325 190.015 ;
        RECT 147.495 189.675 148.800 189.845 ;
        RECT 149.885 189.765 150.205 190.695 ;
        RECT 147.495 189.225 147.740 189.675 ;
        RECT 147.910 189.305 148.460 189.505 ;
        RECT 148.630 189.475 148.800 189.675 ;
        RECT 149.575 189.595 150.205 189.765 ;
        RECT 151.295 189.790 151.565 190.695 ;
        RECT 151.735 190.105 152.065 190.865 ;
        RECT 152.245 189.935 152.425 190.695 ;
        RECT 148.630 189.305 149.005 189.475 ;
        RECT 149.175 189.055 149.405 189.555 ;
        RECT 146.265 188.315 146.435 188.925 ;
        RECT 146.605 188.535 146.935 188.970 ;
        RECT 147.155 188.885 149.405 189.055 ;
        RECT 147.205 188.315 147.535 188.705 ;
        RECT 147.705 188.565 147.875 188.885 ;
        RECT 149.575 188.715 149.745 189.595 ;
        RECT 148.045 188.315 148.375 188.705 ;
        RECT 148.790 188.545 149.745 188.715 ;
        RECT 149.915 188.315 150.205 189.150 ;
        RECT 151.295 188.990 151.475 189.790 ;
        RECT 151.750 189.765 152.425 189.935 ;
        RECT 152.675 189.790 152.945 190.695 ;
        RECT 153.115 190.105 153.445 190.865 ;
        RECT 153.625 189.935 153.805 190.695 ;
        RECT 151.750 189.620 151.920 189.765 ;
        RECT 151.645 189.290 151.920 189.620 ;
        RECT 151.750 189.035 151.920 189.290 ;
        RECT 152.145 189.215 152.485 189.585 ;
        RECT 151.295 188.485 151.555 188.990 ;
        RECT 151.750 188.865 152.415 189.035 ;
        RECT 151.735 188.315 152.065 188.695 ;
        RECT 152.245 188.485 152.415 188.865 ;
        RECT 152.675 188.990 152.855 189.790 ;
        RECT 153.130 189.765 153.805 189.935 ;
        RECT 154.975 189.775 156.185 190.865 ;
        RECT 153.130 189.620 153.300 189.765 ;
        RECT 153.025 189.290 153.300 189.620 ;
        RECT 153.130 189.035 153.300 189.290 ;
        RECT 153.525 189.215 153.865 189.585 ;
        RECT 154.975 189.235 155.495 189.775 ;
        RECT 155.665 189.065 156.185 189.605 ;
        RECT 152.675 188.485 152.935 188.990 ;
        RECT 153.130 188.865 153.795 189.035 ;
        RECT 153.115 188.315 153.445 188.695 ;
        RECT 153.625 188.485 153.795 188.865 ;
        RECT 154.975 188.315 156.185 189.065 ;
        RECT 70.710 188.145 156.270 188.315 ;
        RECT 70.795 187.395 72.005 188.145 ;
        RECT 72.725 187.595 72.895 187.885 ;
        RECT 73.065 187.765 73.395 188.145 ;
        RECT 72.725 187.425 73.390 187.595 ;
        RECT 70.795 186.855 71.315 187.395 ;
        RECT 71.485 186.685 72.005 187.225 ;
        RECT 70.795 185.595 72.005 186.685 ;
        RECT 72.640 186.605 72.990 187.255 ;
        RECT 73.160 186.435 73.390 187.425 ;
        RECT 72.725 186.265 73.390 186.435 ;
        RECT 72.725 185.765 72.895 186.265 ;
        RECT 73.065 185.595 73.395 186.095 ;
        RECT 73.565 185.765 73.750 187.885 ;
        RECT 74.005 187.685 74.255 188.145 ;
        RECT 74.425 187.695 74.760 187.865 ;
        RECT 74.955 187.695 75.630 187.865 ;
        RECT 74.425 187.555 74.595 187.695 ;
        RECT 73.920 186.565 74.200 187.515 ;
        RECT 74.370 187.425 74.595 187.555 ;
        RECT 74.370 186.320 74.540 187.425 ;
        RECT 74.765 187.275 75.290 187.495 ;
        RECT 74.710 186.510 74.950 187.105 ;
        RECT 75.120 186.575 75.290 187.275 ;
        RECT 75.460 186.915 75.630 187.695 ;
        RECT 75.950 187.645 76.320 188.145 ;
        RECT 76.500 187.695 76.905 187.865 ;
        RECT 77.075 187.695 77.860 187.865 ;
        RECT 76.500 187.465 76.670 187.695 ;
        RECT 75.840 187.165 76.670 187.465 ;
        RECT 77.055 187.195 77.520 187.525 ;
        RECT 75.840 187.135 76.040 187.165 ;
        RECT 76.160 186.915 76.330 186.985 ;
        RECT 75.460 186.745 76.330 186.915 ;
        RECT 75.820 186.655 76.330 186.745 ;
        RECT 74.370 186.190 74.675 186.320 ;
        RECT 75.120 186.210 75.650 186.575 ;
        RECT 73.990 185.595 74.255 186.055 ;
        RECT 74.425 185.765 74.675 186.190 ;
        RECT 75.820 186.040 75.990 186.655 ;
        RECT 74.885 185.870 75.990 186.040 ;
        RECT 76.160 185.595 76.330 186.395 ;
        RECT 76.500 186.095 76.670 187.165 ;
        RECT 76.840 186.265 77.030 186.985 ;
        RECT 77.200 186.235 77.520 187.195 ;
        RECT 77.690 187.235 77.860 187.695 ;
        RECT 78.135 187.615 78.345 188.145 ;
        RECT 78.605 187.405 78.935 187.930 ;
        RECT 79.105 187.535 79.275 188.145 ;
        RECT 79.445 187.490 79.775 187.925 ;
        RECT 79.445 187.405 79.825 187.490 ;
        RECT 78.735 187.235 78.935 187.405 ;
        RECT 79.600 187.365 79.825 187.405 ;
        RECT 77.690 186.905 78.565 187.235 ;
        RECT 78.735 186.905 79.485 187.235 ;
        RECT 76.500 185.765 76.750 186.095 ;
        RECT 77.690 186.065 77.860 186.905 ;
        RECT 78.735 186.700 78.925 186.905 ;
        RECT 79.655 186.785 79.825 187.365 ;
        RECT 79.610 186.735 79.825 186.785 ;
        RECT 78.030 186.325 78.925 186.700 ;
        RECT 79.435 186.655 79.825 186.735 ;
        RECT 79.995 187.470 80.255 187.975 ;
        RECT 80.435 187.765 80.765 188.145 ;
        RECT 80.945 187.595 81.115 187.975 ;
        RECT 79.995 186.670 80.175 187.470 ;
        RECT 80.450 187.425 81.115 187.595 ;
        RECT 81.375 187.495 81.635 187.975 ;
        RECT 81.805 187.605 82.055 188.145 ;
        RECT 80.450 187.170 80.620 187.425 ;
        RECT 80.345 186.840 80.620 187.170 ;
        RECT 80.845 186.875 81.185 187.245 ;
        RECT 80.450 186.695 80.620 186.840 ;
        RECT 76.975 185.895 77.860 186.065 ;
        RECT 78.040 185.595 78.355 186.095 ;
        RECT 78.585 185.765 78.925 186.325 ;
        RECT 79.095 185.595 79.265 186.605 ;
        RECT 79.435 185.810 79.765 186.655 ;
        RECT 79.995 185.765 80.265 186.670 ;
        RECT 80.450 186.525 81.125 186.695 ;
        RECT 80.435 185.595 80.765 186.355 ;
        RECT 80.945 185.765 81.125 186.525 ;
        RECT 81.375 186.465 81.545 187.495 ;
        RECT 82.225 187.440 82.445 187.925 ;
        RECT 81.715 186.845 81.945 187.240 ;
        RECT 82.115 187.015 82.445 187.440 ;
        RECT 82.615 187.765 83.505 187.935 ;
        RECT 82.615 187.040 82.785 187.765 ;
        RECT 83.765 187.595 83.935 187.975 ;
        RECT 84.115 187.765 84.445 188.145 ;
        RECT 82.955 187.210 83.505 187.595 ;
        RECT 83.765 187.425 84.430 187.595 ;
        RECT 84.625 187.470 84.885 187.975 ;
        RECT 82.615 186.970 83.505 187.040 ;
        RECT 82.610 186.945 83.505 186.970 ;
        RECT 82.600 186.930 83.505 186.945 ;
        RECT 82.595 186.915 83.505 186.930 ;
        RECT 82.585 186.910 83.505 186.915 ;
        RECT 82.580 186.900 83.505 186.910 ;
        RECT 82.575 186.890 83.505 186.900 ;
        RECT 82.565 186.885 83.505 186.890 ;
        RECT 82.555 186.875 83.505 186.885 ;
        RECT 83.695 186.875 84.035 187.245 ;
        RECT 84.260 187.170 84.430 187.425 ;
        RECT 82.545 186.870 83.505 186.875 ;
        RECT 82.545 186.865 82.880 186.870 ;
        RECT 82.530 186.860 82.880 186.865 ;
        RECT 82.515 186.850 82.880 186.860 ;
        RECT 82.490 186.845 82.880 186.850 ;
        RECT 81.715 186.840 82.880 186.845 ;
        RECT 81.715 186.805 82.850 186.840 ;
        RECT 81.715 186.780 82.815 186.805 ;
        RECT 81.715 186.750 82.785 186.780 ;
        RECT 81.715 186.720 82.765 186.750 ;
        RECT 81.715 186.690 82.745 186.720 ;
        RECT 81.715 186.680 82.675 186.690 ;
        RECT 81.715 186.670 82.650 186.680 ;
        RECT 81.715 186.655 82.630 186.670 ;
        RECT 81.715 186.640 82.610 186.655 ;
        RECT 81.820 186.630 82.605 186.640 ;
        RECT 81.820 186.595 82.590 186.630 ;
        RECT 81.375 185.765 81.650 186.465 ;
        RECT 81.820 186.345 82.575 186.595 ;
        RECT 82.745 186.275 83.075 186.520 ;
        RECT 83.245 186.420 83.505 186.870 ;
        RECT 84.260 186.840 84.535 187.170 ;
        RECT 84.260 186.695 84.430 186.840 ;
        RECT 83.755 186.525 84.430 186.695 ;
        RECT 84.705 186.670 84.885 187.470 ;
        RECT 85.145 187.595 85.315 187.975 ;
        RECT 85.495 187.765 85.825 188.145 ;
        RECT 85.145 187.425 85.810 187.595 ;
        RECT 86.005 187.470 86.265 187.975 ;
        RECT 85.075 186.875 85.415 187.245 ;
        RECT 85.640 187.170 85.810 187.425 ;
        RECT 85.640 186.840 85.915 187.170 ;
        RECT 85.640 186.695 85.810 186.840 ;
        RECT 82.890 186.250 83.075 186.275 ;
        RECT 82.890 186.150 83.505 186.250 ;
        RECT 81.820 185.595 82.075 186.140 ;
        RECT 82.245 185.765 82.725 186.105 ;
        RECT 82.900 185.595 83.505 186.150 ;
        RECT 83.755 185.765 83.935 186.525 ;
        RECT 84.115 185.595 84.445 186.355 ;
        RECT 84.615 185.765 84.885 186.670 ;
        RECT 85.135 186.525 85.810 186.695 ;
        RECT 86.085 186.670 86.265 187.470 ;
        RECT 85.135 185.765 85.315 186.525 ;
        RECT 85.495 185.595 85.825 186.355 ;
        RECT 85.995 185.765 86.265 186.670 ;
        RECT 87.390 187.405 88.005 187.975 ;
        RECT 88.175 187.635 88.390 188.145 ;
        RECT 88.620 187.635 88.900 187.965 ;
        RECT 89.080 187.635 89.320 188.145 ;
        RECT 87.390 186.385 87.705 187.405 ;
        RECT 87.875 186.735 88.045 187.235 ;
        RECT 88.295 186.905 88.560 187.465 ;
        RECT 88.730 186.735 88.900 187.635 ;
        RECT 90.665 187.595 90.835 187.975 ;
        RECT 91.015 187.765 91.345 188.145 ;
        RECT 89.070 186.905 89.425 187.465 ;
        RECT 90.665 187.425 91.330 187.595 ;
        RECT 91.525 187.470 91.785 187.975 ;
        RECT 90.595 186.875 90.935 187.245 ;
        RECT 91.160 187.170 91.330 187.425 ;
        RECT 91.160 186.840 91.435 187.170 ;
        RECT 87.875 186.565 89.300 186.735 ;
        RECT 91.160 186.695 91.330 186.840 ;
        RECT 87.390 185.765 87.925 186.385 ;
        RECT 88.095 185.595 88.425 186.395 ;
        RECT 88.910 186.390 89.300 186.565 ;
        RECT 90.655 186.525 91.330 186.695 ;
        RECT 91.605 186.670 91.785 187.470 ;
        RECT 90.655 185.765 90.835 186.525 ;
        RECT 91.015 185.595 91.345 186.355 ;
        RECT 91.515 185.765 91.785 186.670 ;
        RECT 91.955 187.405 92.215 187.975 ;
        RECT 92.385 187.745 92.770 188.145 ;
        RECT 92.940 187.575 93.195 187.975 ;
        RECT 92.385 187.405 93.195 187.575 ;
        RECT 93.385 187.405 93.630 187.975 ;
        RECT 93.800 187.745 94.185 188.145 ;
        RECT 94.355 187.575 94.610 187.975 ;
        RECT 93.800 187.405 94.610 187.575 ;
        RECT 94.800 187.405 95.225 187.975 ;
        RECT 95.395 187.745 95.780 188.145 ;
        RECT 95.950 187.575 96.385 187.975 ;
        RECT 95.395 187.405 96.385 187.575 ;
        RECT 96.555 187.420 96.845 188.145 ;
        RECT 97.015 187.470 97.275 187.975 ;
        RECT 97.455 187.765 97.785 188.145 ;
        RECT 97.965 187.595 98.135 187.975 ;
        RECT 91.955 186.735 92.140 187.405 ;
        RECT 92.385 187.235 92.735 187.405 ;
        RECT 93.385 187.235 93.555 187.405 ;
        RECT 93.800 187.235 94.150 187.405 ;
        RECT 94.800 187.235 95.150 187.405 ;
        RECT 95.395 187.235 95.730 187.405 ;
        RECT 92.310 186.905 92.735 187.235 ;
        RECT 91.955 185.765 92.215 186.735 ;
        RECT 92.385 186.385 92.735 186.905 ;
        RECT 92.905 186.735 93.555 187.235 ;
        RECT 93.725 186.905 94.150 187.235 ;
        RECT 92.905 186.555 93.630 186.735 ;
        RECT 92.385 186.190 93.195 186.385 ;
        RECT 92.385 185.595 92.770 186.020 ;
        RECT 92.940 185.765 93.195 186.190 ;
        RECT 93.385 185.765 93.630 186.555 ;
        RECT 93.800 186.385 94.150 186.905 ;
        RECT 94.320 186.735 95.150 187.235 ;
        RECT 95.320 186.905 95.730 187.235 ;
        RECT 94.320 186.555 95.225 186.735 ;
        RECT 93.800 186.190 94.630 186.385 ;
        RECT 93.800 185.595 94.185 186.020 ;
        RECT 94.355 185.765 94.630 186.190 ;
        RECT 94.800 185.765 95.225 186.555 ;
        RECT 95.395 186.360 95.730 186.905 ;
        RECT 95.900 186.530 96.385 187.235 ;
        RECT 95.395 186.190 96.385 186.360 ;
        RECT 95.395 185.595 95.780 186.020 ;
        RECT 95.950 185.765 96.385 186.190 ;
        RECT 96.555 185.595 96.845 186.760 ;
        RECT 97.015 186.670 97.195 187.470 ;
        RECT 97.470 187.425 98.135 187.595 ;
        RECT 97.470 187.170 97.640 187.425 ;
        RECT 98.395 187.395 99.605 188.145 ;
        RECT 99.860 187.595 100.035 187.885 ;
        RECT 100.205 187.765 100.535 188.145 ;
        RECT 99.860 187.425 100.355 187.595 ;
        RECT 100.710 187.465 100.925 187.835 ;
        RECT 101.160 187.695 101.760 187.865 ;
        RECT 97.365 186.840 97.640 187.170 ;
        RECT 97.865 186.875 98.205 187.245 ;
        RECT 98.395 186.855 98.915 187.395 ;
        RECT 97.470 186.695 97.640 186.840 ;
        RECT 97.015 185.765 97.285 186.670 ;
        RECT 97.470 186.525 98.145 186.695 ;
        RECT 99.085 186.685 99.605 187.225 ;
        RECT 97.455 185.595 97.785 186.355 ;
        RECT 97.965 185.765 98.145 186.525 ;
        RECT 98.395 185.595 99.605 186.685 ;
        RECT 99.835 186.485 100.015 187.255 ;
        RECT 100.185 186.445 100.355 187.425 ;
        RECT 100.525 187.135 100.925 187.465 ;
        RECT 101.095 187.195 101.420 187.525 ;
        RECT 100.910 186.785 101.080 186.945 ;
        RECT 100.695 186.615 101.080 186.785 ;
        RECT 101.250 186.655 101.420 187.195 ;
        RECT 101.590 186.995 101.760 187.695 ;
        RECT 102.140 187.685 102.470 188.145 ;
        RECT 102.675 187.765 103.105 187.935 ;
        RECT 101.930 187.215 102.305 187.515 ;
        RECT 101.590 186.825 101.930 186.995 ;
        RECT 102.100 186.910 102.305 187.215 ;
        RECT 102.475 186.910 102.765 187.515 ;
        RECT 102.935 187.170 103.105 187.765 ;
        RECT 103.275 187.555 103.510 187.885 ;
        RECT 101.250 186.445 101.590 186.655 ;
        RECT 100.185 186.315 101.590 186.445 ;
        RECT 99.865 186.275 101.590 186.315 ;
        RECT 99.865 186.145 100.355 186.275 ;
        RECT 99.865 185.855 100.035 186.145 ;
        RECT 101.760 186.105 101.930 186.825 ;
        RECT 102.935 186.840 103.170 187.170 ;
        RECT 102.935 186.740 103.105 186.840 ;
        RECT 102.835 186.570 103.105 186.740 ;
        RECT 102.835 186.445 103.005 186.570 ;
        RECT 102.660 186.275 103.005 186.445 ;
        RECT 103.340 186.420 103.510 187.555 ;
        RECT 100.205 185.595 100.535 185.975 ;
        RECT 101.100 185.935 101.930 186.105 ;
        RECT 102.285 185.595 102.515 186.175 ;
        RECT 103.255 186.105 103.510 186.420 ;
        RECT 102.995 185.935 103.510 186.105 ;
        RECT 103.680 186.105 103.870 187.885 ;
        RECT 104.085 187.645 104.290 187.975 ;
        RECT 104.485 187.685 104.815 188.145 ;
        RECT 105.015 187.765 105.910 187.935 ;
        RECT 104.085 186.665 104.255 187.645 ;
        RECT 104.435 186.835 104.805 187.515 ;
        RECT 105.015 186.665 105.185 187.765 ;
        RECT 104.085 186.495 105.185 186.665 ;
        RECT 104.085 186.335 104.275 186.495 ;
        RECT 103.680 185.935 104.205 186.105 ;
        RECT 104.445 185.595 104.790 186.225 ;
        RECT 105.015 186.075 105.185 186.495 ;
        RECT 105.355 187.195 105.975 187.525 ;
        RECT 106.225 187.235 106.535 187.855 ;
        RECT 106.705 187.415 106.955 188.145 ;
        RECT 107.125 187.505 107.455 187.965 ;
        RECT 105.355 186.245 105.645 187.195 ;
        RECT 106.225 187.155 106.635 187.235 ;
        RECT 105.815 186.585 106.155 186.985 ;
        RECT 106.325 186.905 106.635 187.155 ;
        RECT 106.805 186.905 107.115 187.235 ;
        RECT 106.805 186.735 106.975 186.905 ;
        RECT 107.285 186.735 107.455 187.505 ;
        RECT 107.625 187.345 107.880 188.145 ;
        RECT 108.140 187.595 108.315 187.885 ;
        RECT 108.485 187.765 108.815 188.145 ;
        RECT 108.140 187.425 108.635 187.595 ;
        RECT 108.990 187.465 109.205 187.835 ;
        RECT 109.440 187.695 110.040 187.865 ;
        RECT 106.365 186.565 106.975 186.735 ;
        RECT 106.365 186.105 106.535 186.565 ;
        RECT 107.145 186.395 107.455 186.735 ;
        RECT 105.015 185.905 105.965 186.075 ;
        RECT 106.215 185.935 106.535 186.105 ;
        RECT 106.705 185.595 106.875 186.395 ;
        RECT 107.045 185.775 107.455 186.395 ;
        RECT 107.625 185.595 107.875 186.735 ;
        RECT 108.115 186.485 108.295 187.255 ;
        RECT 108.465 186.445 108.635 187.425 ;
        RECT 108.805 187.135 109.205 187.465 ;
        RECT 109.375 187.195 109.700 187.525 ;
        RECT 109.190 186.785 109.360 186.945 ;
        RECT 108.975 186.615 109.360 186.785 ;
        RECT 109.530 186.655 109.700 187.195 ;
        RECT 109.870 186.995 110.040 187.695 ;
        RECT 110.420 187.685 110.750 188.145 ;
        RECT 110.955 187.765 111.385 187.935 ;
        RECT 110.210 187.215 110.585 187.515 ;
        RECT 109.870 186.825 110.210 186.995 ;
        RECT 110.380 186.910 110.585 187.215 ;
        RECT 110.755 186.910 111.045 187.515 ;
        RECT 111.215 187.170 111.385 187.765 ;
        RECT 111.555 187.555 111.790 187.885 ;
        RECT 109.530 186.445 109.870 186.655 ;
        RECT 108.465 186.315 109.870 186.445 ;
        RECT 108.145 186.275 109.870 186.315 ;
        RECT 108.145 186.145 108.635 186.275 ;
        RECT 108.145 185.855 108.315 186.145 ;
        RECT 110.040 186.105 110.210 186.825 ;
        RECT 111.215 186.840 111.450 187.170 ;
        RECT 111.215 186.740 111.385 186.840 ;
        RECT 111.115 186.570 111.385 186.740 ;
        RECT 111.115 186.445 111.285 186.570 ;
        RECT 110.940 186.275 111.285 186.445 ;
        RECT 111.620 186.420 111.790 187.555 ;
        RECT 108.485 185.595 108.815 185.975 ;
        RECT 109.380 185.935 110.210 186.105 ;
        RECT 110.565 185.595 110.795 186.175 ;
        RECT 111.535 186.105 111.790 186.420 ;
        RECT 111.275 185.935 111.790 186.105 ;
        RECT 111.960 186.105 112.150 187.885 ;
        RECT 112.365 187.645 112.570 187.975 ;
        RECT 112.765 187.685 113.095 188.145 ;
        RECT 113.295 187.765 114.190 187.935 ;
        RECT 112.365 186.665 112.535 187.645 ;
        RECT 112.715 186.835 113.085 187.515 ;
        RECT 113.295 186.665 113.465 187.765 ;
        RECT 112.365 186.495 113.465 186.665 ;
        RECT 112.365 186.335 112.555 186.495 ;
        RECT 111.960 185.935 112.485 186.105 ;
        RECT 112.725 185.595 113.070 186.225 ;
        RECT 113.295 186.075 113.465 186.495 ;
        RECT 113.635 187.195 114.255 187.525 ;
        RECT 114.505 187.235 114.815 187.855 ;
        RECT 114.985 187.415 115.235 188.145 ;
        RECT 115.405 187.505 115.735 187.965 ;
        RECT 113.635 186.245 113.925 187.195 ;
        RECT 114.505 187.155 114.915 187.235 ;
        RECT 114.095 186.585 114.435 186.985 ;
        RECT 114.605 186.905 114.915 187.155 ;
        RECT 115.085 186.905 115.395 187.235 ;
        RECT 115.085 186.735 115.255 186.905 ;
        RECT 115.565 186.735 115.735 187.505 ;
        RECT 115.905 187.345 116.160 188.145 ;
        RECT 116.335 187.470 116.595 187.975 ;
        RECT 116.775 187.765 117.105 188.145 ;
        RECT 117.285 187.595 117.455 187.975 ;
        RECT 114.645 186.565 115.255 186.735 ;
        RECT 114.645 186.105 114.815 186.565 ;
        RECT 115.425 186.395 115.735 186.735 ;
        RECT 113.295 185.905 114.245 186.075 ;
        RECT 114.495 185.935 114.815 186.105 ;
        RECT 114.985 185.595 115.155 186.395 ;
        RECT 115.325 185.775 115.735 186.395 ;
        RECT 115.905 185.595 116.155 186.735 ;
        RECT 116.335 186.670 116.515 187.470 ;
        RECT 116.790 187.425 117.455 187.595 ;
        RECT 116.790 187.170 116.960 187.425 ;
        RECT 117.715 187.405 118.030 187.780 ;
        RECT 118.285 187.405 118.455 188.145 ;
        RECT 118.705 187.575 118.875 187.780 ;
        RECT 119.100 187.745 119.475 188.145 ;
        RECT 119.645 187.575 119.815 187.925 ;
        RECT 120.000 187.745 120.330 188.145 ;
        RECT 120.500 187.575 120.670 187.925 ;
        RECT 120.840 187.745 121.220 188.145 ;
        RECT 118.705 187.405 119.205 187.575 ;
        RECT 119.645 187.405 121.240 187.575 ;
        RECT 121.410 187.470 121.685 187.815 ;
        RECT 116.685 186.840 116.960 187.170 ;
        RECT 117.185 186.875 117.525 187.245 ;
        RECT 116.790 186.695 116.960 186.840 ;
        RECT 116.335 185.765 116.605 186.670 ;
        RECT 116.790 186.525 117.465 186.695 ;
        RECT 116.775 185.595 117.105 186.355 ;
        RECT 117.285 185.765 117.465 186.525 ;
        RECT 117.715 186.365 117.885 187.405 ;
        RECT 118.055 186.535 118.405 187.235 ;
        RECT 118.575 186.905 118.865 187.235 ;
        RECT 119.035 187.155 119.205 187.405 ;
        RECT 121.070 187.235 121.240 187.405 ;
        RECT 119.035 186.985 119.460 187.155 ;
        RECT 119.035 186.705 119.205 186.985 ;
        RECT 119.855 186.815 120.025 187.235 ;
        RECT 120.245 186.905 120.900 187.235 ;
        RECT 121.070 186.905 121.345 187.235 ;
        RECT 118.620 186.535 119.205 186.705 ;
        RECT 119.375 186.645 120.025 186.815 ;
        RECT 121.070 186.735 121.240 186.905 ;
        RECT 121.515 186.735 121.685 187.470 ;
        RECT 122.315 187.420 122.605 188.145 ;
        RECT 122.775 187.470 123.035 187.975 ;
        RECT 123.215 187.765 123.545 188.145 ;
        RECT 123.725 187.595 123.895 187.975 ;
        RECT 124.615 187.635 124.920 188.145 ;
        RECT 119.375 186.365 119.545 186.645 ;
        RECT 120.580 186.565 121.240 186.735 ;
        RECT 120.580 186.445 120.750 186.565 ;
        RECT 117.715 186.195 119.545 186.365 ;
        RECT 119.715 186.275 120.750 186.445 ;
        RECT 117.715 185.775 117.975 186.195 ;
        RECT 119.715 186.025 119.885 186.275 ;
        RECT 118.145 185.595 118.475 186.025 ;
        RECT 119.140 185.855 119.885 186.025 ;
        RECT 120.075 185.935 120.750 186.105 ;
        RECT 120.110 185.775 120.750 185.935 ;
        RECT 120.920 185.595 121.200 186.395 ;
        RECT 121.410 185.765 121.685 186.735 ;
        RECT 122.315 185.595 122.605 186.760 ;
        RECT 122.775 186.670 122.955 187.470 ;
        RECT 123.230 187.425 123.895 187.595 ;
        RECT 123.230 187.170 123.400 187.425 ;
        RECT 123.125 186.840 123.400 187.170 ;
        RECT 123.625 186.875 123.965 187.245 ;
        RECT 124.615 186.905 124.930 187.465 ;
        RECT 125.100 187.155 125.350 187.965 ;
        RECT 125.520 187.620 125.780 188.145 ;
        RECT 125.960 187.155 126.210 187.965 ;
        RECT 126.380 187.585 126.640 188.145 ;
        RECT 126.810 187.495 127.070 187.950 ;
        RECT 127.240 187.665 127.500 188.145 ;
        RECT 127.670 187.495 127.930 187.950 ;
        RECT 128.100 187.665 128.360 188.145 ;
        RECT 128.530 187.495 128.790 187.950 ;
        RECT 128.960 187.665 129.205 188.145 ;
        RECT 129.375 187.495 129.650 187.950 ;
        RECT 129.820 187.665 130.065 188.145 ;
        RECT 130.235 187.495 130.495 187.950 ;
        RECT 130.675 187.665 130.925 188.145 ;
        RECT 131.095 187.495 131.355 187.950 ;
        RECT 131.535 187.665 131.785 188.145 ;
        RECT 131.955 187.495 132.215 187.950 ;
        RECT 132.395 187.665 132.655 188.145 ;
        RECT 132.825 187.495 133.085 187.950 ;
        RECT 133.255 187.665 133.555 188.145 ;
        RECT 133.900 187.595 134.075 187.885 ;
        RECT 134.245 187.765 134.575 188.145 ;
        RECT 126.810 187.325 133.555 187.495 ;
        RECT 133.900 187.425 134.395 187.595 ;
        RECT 134.750 187.465 134.965 187.835 ;
        RECT 135.200 187.695 135.800 187.865 ;
        RECT 125.100 186.905 132.220 187.155 ;
        RECT 123.230 186.695 123.400 186.840 ;
        RECT 122.775 185.765 123.045 186.670 ;
        RECT 123.230 186.525 123.905 186.695 ;
        RECT 123.215 185.595 123.545 186.355 ;
        RECT 123.725 185.765 123.905 186.525 ;
        RECT 124.625 185.595 124.920 186.405 ;
        RECT 125.100 185.765 125.345 186.905 ;
        RECT 125.520 185.595 125.780 186.405 ;
        RECT 125.960 185.770 126.210 186.905 ;
        RECT 132.390 186.735 133.555 187.325 ;
        RECT 126.810 186.510 133.555 186.735 ;
        RECT 126.810 186.495 132.215 186.510 ;
        RECT 126.380 185.600 126.640 186.395 ;
        RECT 126.810 185.770 127.070 186.495 ;
        RECT 127.240 185.600 127.500 186.325 ;
        RECT 127.670 185.770 127.930 186.495 ;
        RECT 128.100 185.600 128.360 186.325 ;
        RECT 128.530 185.770 128.790 186.495 ;
        RECT 128.960 185.600 129.220 186.325 ;
        RECT 129.390 185.770 129.650 186.495 ;
        RECT 129.820 185.600 130.065 186.325 ;
        RECT 130.235 185.770 130.495 186.495 ;
        RECT 130.680 185.600 130.925 186.325 ;
        RECT 131.095 185.770 131.355 186.495 ;
        RECT 131.540 185.600 131.785 186.325 ;
        RECT 131.955 185.770 132.215 186.495 ;
        RECT 132.400 185.600 132.655 186.325 ;
        RECT 132.825 185.770 133.115 186.510 ;
        RECT 133.875 186.485 134.055 187.255 ;
        RECT 134.225 186.445 134.395 187.425 ;
        RECT 134.565 187.135 134.965 187.465 ;
        RECT 135.135 187.195 135.460 187.525 ;
        RECT 134.950 186.785 135.120 186.945 ;
        RECT 134.735 186.615 135.120 186.785 ;
        RECT 135.290 186.655 135.460 187.195 ;
        RECT 135.630 186.995 135.800 187.695 ;
        RECT 136.180 187.685 136.510 188.145 ;
        RECT 136.715 187.765 137.145 187.935 ;
        RECT 135.970 187.215 136.345 187.515 ;
        RECT 135.630 186.825 135.970 186.995 ;
        RECT 136.140 186.910 136.345 187.215 ;
        RECT 136.515 186.910 136.805 187.515 ;
        RECT 136.975 187.170 137.145 187.765 ;
        RECT 137.315 187.555 137.550 187.885 ;
        RECT 135.290 186.445 135.630 186.655 ;
        RECT 126.380 185.595 132.655 185.600 ;
        RECT 133.285 185.595 133.555 186.340 ;
        RECT 134.225 186.315 135.630 186.445 ;
        RECT 133.905 186.275 135.630 186.315 ;
        RECT 133.905 186.145 134.395 186.275 ;
        RECT 133.905 185.855 134.075 186.145 ;
        RECT 135.800 186.105 135.970 186.825 ;
        RECT 136.975 186.840 137.210 187.170 ;
        RECT 136.975 186.740 137.145 186.840 ;
        RECT 136.875 186.570 137.145 186.740 ;
        RECT 136.875 186.445 137.045 186.570 ;
        RECT 136.700 186.275 137.045 186.445 ;
        RECT 137.380 186.420 137.550 187.555 ;
        RECT 134.245 185.595 134.575 185.975 ;
        RECT 135.140 185.935 135.970 186.105 ;
        RECT 136.325 185.595 136.555 186.175 ;
        RECT 137.295 186.105 137.550 186.420 ;
        RECT 137.035 185.935 137.550 186.105 ;
        RECT 137.720 186.105 137.910 187.885 ;
        RECT 138.125 187.645 138.330 187.975 ;
        RECT 138.525 187.685 138.855 188.145 ;
        RECT 139.055 187.765 139.950 187.935 ;
        RECT 138.125 186.665 138.295 187.645 ;
        RECT 138.475 186.835 138.845 187.515 ;
        RECT 139.055 186.665 139.225 187.765 ;
        RECT 138.125 186.495 139.225 186.665 ;
        RECT 138.125 186.335 138.315 186.495 ;
        RECT 137.720 185.935 138.245 186.105 ;
        RECT 138.485 185.595 138.830 186.225 ;
        RECT 139.055 186.075 139.225 186.495 ;
        RECT 139.395 187.195 140.015 187.525 ;
        RECT 140.265 187.235 140.575 187.855 ;
        RECT 140.745 187.415 140.995 188.145 ;
        RECT 141.165 187.505 141.495 187.965 ;
        RECT 139.395 186.245 139.685 187.195 ;
        RECT 140.265 187.155 140.675 187.235 ;
        RECT 139.855 186.585 140.195 186.985 ;
        RECT 140.365 186.905 140.675 187.155 ;
        RECT 140.845 186.905 141.155 187.235 ;
        RECT 140.845 186.735 141.015 186.905 ;
        RECT 141.325 186.735 141.495 187.505 ;
        RECT 141.665 187.345 141.920 188.145 ;
        RECT 142.095 187.575 142.530 187.975 ;
        RECT 142.700 187.745 143.085 188.145 ;
        RECT 142.095 187.405 143.085 187.575 ;
        RECT 143.255 187.405 143.680 187.975 ;
        RECT 143.870 187.575 144.125 187.975 ;
        RECT 144.295 187.745 144.680 188.145 ;
        RECT 143.870 187.405 144.680 187.575 ;
        RECT 144.850 187.405 145.095 187.975 ;
        RECT 145.285 187.575 145.540 187.975 ;
        RECT 145.710 187.745 146.095 188.145 ;
        RECT 145.285 187.405 146.095 187.575 ;
        RECT 146.265 187.405 146.525 187.975 ;
        RECT 142.750 187.235 143.085 187.405 ;
        RECT 143.330 187.235 143.680 187.405 ;
        RECT 144.330 187.235 144.680 187.405 ;
        RECT 144.925 187.235 145.095 187.405 ;
        RECT 145.745 187.235 146.095 187.405 ;
        RECT 140.405 186.565 141.015 186.735 ;
        RECT 140.405 186.105 140.575 186.565 ;
        RECT 141.185 186.395 141.495 186.735 ;
        RECT 139.055 185.905 140.005 186.075 ;
        RECT 140.255 185.935 140.575 186.105 ;
        RECT 140.745 185.595 140.915 186.395 ;
        RECT 141.085 185.775 141.495 186.395 ;
        RECT 141.665 185.595 141.915 186.735 ;
        RECT 142.095 186.530 142.580 187.235 ;
        RECT 142.750 186.905 143.160 187.235 ;
        RECT 142.750 186.360 143.085 186.905 ;
        RECT 143.330 186.735 144.160 187.235 ;
        RECT 142.095 186.190 143.085 186.360 ;
        RECT 143.255 186.555 144.160 186.735 ;
        RECT 144.330 186.905 144.755 187.235 ;
        RECT 142.095 185.765 142.530 186.190 ;
        RECT 142.700 185.595 143.085 186.020 ;
        RECT 143.255 185.765 143.680 186.555 ;
        RECT 144.330 186.385 144.680 186.905 ;
        RECT 144.925 186.735 145.575 187.235 ;
        RECT 143.850 186.190 144.680 186.385 ;
        RECT 144.850 186.555 145.575 186.735 ;
        RECT 145.745 186.905 146.170 187.235 ;
        RECT 143.850 185.765 144.125 186.190 ;
        RECT 144.295 185.595 144.680 186.020 ;
        RECT 144.850 185.765 145.095 186.555 ;
        RECT 145.745 186.385 146.095 186.905 ;
        RECT 146.340 186.735 146.525 187.405 ;
        RECT 145.285 186.190 146.095 186.385 ;
        RECT 145.285 185.765 145.540 186.190 ;
        RECT 145.710 185.595 146.095 186.020 ;
        RECT 146.265 185.765 146.525 186.735 ;
        RECT 146.695 187.470 146.955 187.975 ;
        RECT 147.135 187.765 147.465 188.145 ;
        RECT 147.645 187.595 147.815 187.975 ;
        RECT 146.695 186.670 146.865 187.470 ;
        RECT 147.150 187.425 147.815 187.595 ;
        RECT 147.150 187.170 147.320 187.425 ;
        RECT 148.075 187.420 148.365 188.145 ;
        RECT 148.535 187.685 149.095 187.975 ;
        RECT 149.265 187.685 149.515 188.145 ;
        RECT 147.035 186.840 147.320 187.170 ;
        RECT 147.555 186.875 147.885 187.245 ;
        RECT 147.150 186.695 147.320 186.840 ;
        RECT 146.695 185.765 146.965 186.670 ;
        RECT 147.150 186.525 147.815 186.695 ;
        RECT 147.135 185.595 147.465 186.355 ;
        RECT 147.645 185.765 147.815 186.525 ;
        RECT 148.075 185.595 148.365 186.760 ;
        RECT 148.535 186.315 148.785 187.685 ;
        RECT 150.135 187.515 150.465 187.875 ;
        RECT 149.075 187.325 150.465 187.515 ;
        RECT 150.835 187.470 151.095 187.975 ;
        RECT 151.275 187.765 151.605 188.145 ;
        RECT 151.785 187.595 151.955 187.975 ;
        RECT 149.075 187.235 149.245 187.325 ;
        RECT 148.955 186.905 149.245 187.235 ;
        RECT 149.415 186.905 149.755 187.155 ;
        RECT 149.975 186.905 150.650 187.155 ;
        RECT 149.075 186.655 149.245 186.905 ;
        RECT 149.075 186.485 150.015 186.655 ;
        RECT 150.385 186.545 150.650 186.905 ;
        RECT 150.835 186.670 151.015 187.470 ;
        RECT 151.290 187.425 151.955 187.595 ;
        RECT 152.215 187.470 152.475 187.975 ;
        RECT 152.655 187.765 152.985 188.145 ;
        RECT 153.165 187.595 153.335 187.975 ;
        RECT 151.290 187.170 151.460 187.425 ;
        RECT 151.185 186.840 151.460 187.170 ;
        RECT 151.685 186.875 152.025 187.245 ;
        RECT 151.290 186.695 151.460 186.840 ;
        RECT 148.535 185.765 148.995 186.315 ;
        RECT 149.185 185.595 149.515 186.315 ;
        RECT 149.715 185.935 150.015 186.485 ;
        RECT 150.185 185.595 150.465 186.265 ;
        RECT 150.835 185.765 151.105 186.670 ;
        RECT 151.290 186.525 151.965 186.695 ;
        RECT 151.275 185.595 151.605 186.355 ;
        RECT 151.785 185.765 151.965 186.525 ;
        RECT 152.215 186.670 152.395 187.470 ;
        RECT 152.670 187.425 153.335 187.595 ;
        RECT 153.595 187.470 153.855 187.975 ;
        RECT 154.035 187.765 154.365 188.145 ;
        RECT 154.545 187.595 154.715 187.975 ;
        RECT 152.670 187.170 152.840 187.425 ;
        RECT 152.565 186.840 152.840 187.170 ;
        RECT 153.065 186.875 153.405 187.245 ;
        RECT 152.670 186.695 152.840 186.840 ;
        RECT 152.215 185.765 152.485 186.670 ;
        RECT 152.670 186.525 153.345 186.695 ;
        RECT 152.655 185.595 152.985 186.355 ;
        RECT 153.165 185.765 153.345 186.525 ;
        RECT 153.595 186.670 153.765 187.470 ;
        RECT 154.050 187.425 154.715 187.595 ;
        RECT 154.050 187.170 154.220 187.425 ;
        RECT 154.975 187.395 156.185 188.145 ;
        RECT 153.935 186.840 154.220 187.170 ;
        RECT 154.455 186.875 154.785 187.245 ;
        RECT 154.050 186.695 154.220 186.840 ;
        RECT 153.595 185.765 153.865 186.670 ;
        RECT 154.050 186.525 154.715 186.695 ;
        RECT 154.035 185.595 154.365 186.355 ;
        RECT 154.545 185.765 154.715 186.525 ;
        RECT 154.975 186.685 155.495 187.225 ;
        RECT 155.665 186.855 156.185 187.395 ;
        RECT 154.975 185.595 156.185 186.685 ;
        RECT 70.710 185.425 156.270 185.595 ;
        RECT 70.795 184.335 72.005 185.425 ;
        RECT 72.175 184.335 73.845 185.425 ;
        RECT 70.795 183.625 71.315 184.165 ;
        RECT 71.485 183.795 72.005 184.335 ;
        RECT 72.175 183.645 72.925 184.165 ;
        RECT 73.095 183.815 73.845 184.335 ;
        RECT 74.485 184.455 74.815 185.240 ;
        RECT 74.485 184.285 75.165 184.455 ;
        RECT 75.345 184.285 75.675 185.425 ;
        RECT 75.860 184.625 76.115 185.425 ;
        RECT 76.315 184.575 76.645 185.255 ;
        RECT 74.475 183.865 74.825 184.115 ;
        RECT 74.995 183.685 75.165 184.285 ;
        RECT 75.335 183.865 75.685 184.115 ;
        RECT 75.860 184.085 76.105 184.445 ;
        RECT 76.295 184.295 76.645 184.575 ;
        RECT 76.295 183.915 76.465 184.295 ;
        RECT 76.825 184.115 77.020 185.165 ;
        RECT 77.200 184.285 77.520 185.425 ;
        RECT 77.695 184.335 80.285 185.425 ;
        RECT 80.455 184.915 80.715 185.425 ;
        RECT 75.945 183.745 76.465 183.915 ;
        RECT 76.635 183.785 77.020 184.115 ;
        RECT 77.200 184.065 77.460 184.115 ;
        RECT 77.200 183.895 77.465 184.065 ;
        RECT 77.200 183.785 77.460 183.895 ;
        RECT 75.945 183.725 76.115 183.745 ;
        RECT 70.795 182.875 72.005 183.625 ;
        RECT 72.175 182.875 73.845 183.645 ;
        RECT 74.495 182.875 74.735 183.685 ;
        RECT 74.905 183.045 75.235 183.685 ;
        RECT 75.405 182.875 75.675 183.685 ;
        RECT 75.915 183.555 76.115 183.725 ;
        RECT 77.695 183.645 78.905 184.165 ;
        RECT 79.075 183.815 80.285 184.335 ;
        RECT 80.455 183.865 80.795 184.745 ;
        RECT 80.965 184.035 81.135 185.255 ;
        RECT 81.375 184.920 81.990 185.425 ;
        RECT 81.375 184.385 81.625 184.750 ;
        RECT 81.795 184.745 81.990 184.920 ;
        RECT 82.160 184.915 82.635 185.255 ;
        RECT 82.805 184.880 83.020 185.425 ;
        RECT 81.795 184.555 82.125 184.745 ;
        RECT 82.345 184.385 83.060 184.680 ;
        RECT 83.230 184.555 83.505 185.255 ;
        RECT 81.375 184.215 83.165 184.385 ;
        RECT 80.965 183.785 81.760 184.035 ;
        RECT 80.965 183.695 81.215 183.785 ;
        RECT 75.945 183.180 76.115 183.555 ;
        RECT 76.305 183.405 77.520 183.575 ;
        RECT 76.305 183.100 76.535 183.405 ;
        RECT 76.705 182.875 77.035 183.235 ;
        RECT 77.230 183.055 77.520 183.405 ;
        RECT 77.695 182.875 80.285 183.645 ;
        RECT 80.455 182.875 80.715 183.695 ;
        RECT 80.885 183.275 81.215 183.695 ;
        RECT 81.930 183.360 82.185 184.215 ;
        RECT 81.395 183.095 82.185 183.360 ;
        RECT 82.355 183.515 82.765 184.035 ;
        RECT 82.935 183.785 83.165 184.215 ;
        RECT 83.335 183.525 83.505 184.555 ;
        RECT 83.675 184.260 83.965 185.425 ;
        RECT 84.225 184.755 84.395 185.255 ;
        RECT 84.565 184.925 84.895 185.425 ;
        RECT 84.225 184.585 84.890 184.755 ;
        RECT 84.140 183.765 84.490 184.415 ;
        RECT 82.355 183.095 82.555 183.515 ;
        RECT 82.745 182.875 83.075 183.335 ;
        RECT 83.245 183.045 83.505 183.525 ;
        RECT 83.675 182.875 83.965 183.600 ;
        RECT 84.660 183.595 84.890 184.585 ;
        RECT 84.225 183.425 84.890 183.595 ;
        RECT 84.225 183.135 84.395 183.425 ;
        RECT 84.565 182.875 84.895 183.255 ;
        RECT 85.065 183.135 85.250 185.255 ;
        RECT 85.490 184.965 85.755 185.425 ;
        RECT 85.925 184.830 86.175 185.255 ;
        RECT 86.385 184.980 87.490 185.150 ;
        RECT 85.870 184.700 86.175 184.830 ;
        RECT 85.420 183.505 85.700 184.455 ;
        RECT 85.870 183.595 86.040 184.700 ;
        RECT 86.210 183.915 86.450 184.510 ;
        RECT 86.620 184.445 87.150 184.810 ;
        RECT 86.620 183.745 86.790 184.445 ;
        RECT 87.320 184.365 87.490 184.980 ;
        RECT 87.660 184.625 87.830 185.425 ;
        RECT 88.000 184.925 88.250 185.255 ;
        RECT 88.475 184.955 89.360 185.125 ;
        RECT 87.320 184.275 87.830 184.365 ;
        RECT 85.870 183.465 86.095 183.595 ;
        RECT 86.265 183.525 86.790 183.745 ;
        RECT 86.960 184.105 87.830 184.275 ;
        RECT 85.505 182.875 85.755 183.335 ;
        RECT 85.925 183.325 86.095 183.465 ;
        RECT 86.960 183.325 87.130 184.105 ;
        RECT 87.660 184.035 87.830 184.105 ;
        RECT 87.340 183.855 87.540 183.885 ;
        RECT 88.000 183.855 88.170 184.925 ;
        RECT 88.340 184.035 88.530 184.755 ;
        RECT 87.340 183.555 88.170 183.855 ;
        RECT 88.700 183.825 89.020 184.785 ;
        RECT 85.925 183.155 86.260 183.325 ;
        RECT 86.455 183.155 87.130 183.325 ;
        RECT 87.450 182.875 87.820 183.375 ;
        RECT 88.000 183.325 88.170 183.555 ;
        RECT 88.555 183.495 89.020 183.825 ;
        RECT 89.190 184.115 89.360 184.955 ;
        RECT 89.540 184.925 89.855 185.425 ;
        RECT 90.085 184.695 90.425 185.255 ;
        RECT 89.530 184.320 90.425 184.695 ;
        RECT 90.595 184.415 90.765 185.425 ;
        RECT 90.235 184.115 90.425 184.320 ;
        RECT 90.935 184.365 91.265 185.210 ;
        RECT 90.935 184.285 91.325 184.365 ;
        RECT 91.110 184.235 91.325 184.285 ;
        RECT 89.190 183.785 90.065 184.115 ;
        RECT 90.235 183.785 90.985 184.115 ;
        RECT 89.190 183.325 89.360 183.785 ;
        RECT 90.235 183.615 90.435 183.785 ;
        RECT 91.155 183.655 91.325 184.235 ;
        RECT 91.100 183.615 91.325 183.655 ;
        RECT 88.000 183.155 88.405 183.325 ;
        RECT 88.575 183.155 89.360 183.325 ;
        RECT 89.635 182.875 89.845 183.405 ;
        RECT 90.105 183.090 90.435 183.615 ;
        RECT 90.945 183.530 91.325 183.615 ;
        RECT 92.415 184.350 92.685 185.255 ;
        RECT 92.855 184.665 93.185 185.425 ;
        RECT 93.365 184.495 93.545 185.255 ;
        RECT 93.795 184.830 94.230 185.255 ;
        RECT 94.400 185.000 94.785 185.425 ;
        RECT 93.795 184.660 94.785 184.830 ;
        RECT 92.415 183.550 92.595 184.350 ;
        RECT 92.870 184.325 93.545 184.495 ;
        RECT 92.870 184.180 93.040 184.325 ;
        RECT 92.765 183.850 93.040 184.180 ;
        RECT 92.870 183.595 93.040 183.850 ;
        RECT 93.265 183.775 93.605 184.145 ;
        RECT 93.795 183.785 94.280 184.490 ;
        RECT 94.450 184.115 94.785 184.660 ;
        RECT 94.955 184.465 95.380 185.255 ;
        RECT 95.550 184.830 95.825 185.255 ;
        RECT 95.995 185.000 96.380 185.425 ;
        RECT 95.550 184.635 96.380 184.830 ;
        RECT 94.955 184.285 95.860 184.465 ;
        RECT 94.450 183.785 94.860 184.115 ;
        RECT 95.030 183.785 95.860 184.285 ;
        RECT 96.030 184.115 96.380 184.635 ;
        RECT 96.550 184.465 96.795 185.255 ;
        RECT 96.985 184.830 97.240 185.255 ;
        RECT 97.410 185.000 97.795 185.425 ;
        RECT 96.985 184.635 97.795 184.830 ;
        RECT 96.550 184.285 97.275 184.465 ;
        RECT 96.030 183.785 96.455 184.115 ;
        RECT 96.625 183.785 97.275 184.285 ;
        RECT 97.445 184.115 97.795 184.635 ;
        RECT 97.965 184.285 98.225 185.255 ;
        RECT 97.445 183.785 97.870 184.115 ;
        RECT 94.450 183.615 94.785 183.785 ;
        RECT 95.030 183.615 95.380 183.785 ;
        RECT 96.030 183.615 96.380 183.785 ;
        RECT 96.625 183.615 96.795 183.785 ;
        RECT 97.445 183.615 97.795 183.785 ;
        RECT 98.040 183.615 98.225 184.285 ;
        RECT 90.605 182.875 90.775 183.485 ;
        RECT 90.945 183.095 91.275 183.530 ;
        RECT 92.415 183.045 92.675 183.550 ;
        RECT 92.870 183.425 93.535 183.595 ;
        RECT 92.855 182.875 93.185 183.255 ;
        RECT 93.365 183.045 93.535 183.425 ;
        RECT 93.795 183.445 94.785 183.615 ;
        RECT 93.795 183.045 94.230 183.445 ;
        RECT 94.400 182.875 94.785 183.275 ;
        RECT 94.955 183.045 95.380 183.615 ;
        RECT 95.570 183.445 96.380 183.615 ;
        RECT 95.570 183.045 95.825 183.445 ;
        RECT 95.995 182.875 96.380 183.275 ;
        RECT 96.550 183.045 96.795 183.615 ;
        RECT 96.985 183.445 97.795 183.615 ;
        RECT 96.985 183.045 97.240 183.445 ;
        RECT 97.410 182.875 97.795 183.275 ;
        RECT 97.965 183.045 98.225 183.615 ;
        RECT 98.400 184.285 98.735 185.255 ;
        RECT 98.905 184.285 99.075 185.425 ;
        RECT 99.245 185.085 101.275 185.255 ;
        RECT 98.400 183.615 98.570 184.285 ;
        RECT 99.245 184.115 99.415 185.085 ;
        RECT 98.740 183.785 98.995 184.115 ;
        RECT 99.220 183.785 99.415 184.115 ;
        RECT 99.585 184.745 100.710 184.915 ;
        RECT 98.825 183.615 98.995 183.785 ;
        RECT 99.585 183.615 99.755 184.745 ;
        RECT 98.400 183.045 98.655 183.615 ;
        RECT 98.825 183.445 99.755 183.615 ;
        RECT 99.925 184.405 100.935 184.575 ;
        RECT 99.925 183.605 100.095 184.405 ;
        RECT 100.300 184.065 100.575 184.205 ;
        RECT 100.295 183.895 100.575 184.065 ;
        RECT 99.580 183.410 99.755 183.445 ;
        RECT 98.825 182.875 99.155 183.275 ;
        RECT 99.580 183.045 100.110 183.410 ;
        RECT 100.300 183.045 100.575 183.895 ;
        RECT 100.745 183.045 100.935 184.405 ;
        RECT 101.105 184.420 101.275 185.085 ;
        RECT 101.445 184.665 101.615 185.425 ;
        RECT 101.850 184.665 102.365 185.075 ;
        RECT 101.105 184.230 101.855 184.420 ;
        RECT 102.025 183.855 102.365 184.665 ;
        RECT 102.615 184.495 102.795 185.255 ;
        RECT 102.975 184.665 103.305 185.425 ;
        RECT 102.615 184.325 103.290 184.495 ;
        RECT 103.475 184.350 103.745 185.255 ;
        RECT 103.915 184.990 109.260 185.425 ;
        RECT 103.120 184.180 103.290 184.325 ;
        RECT 101.135 183.685 102.365 183.855 ;
        RECT 102.555 183.775 102.895 184.145 ;
        RECT 103.120 183.850 103.395 184.180 ;
        RECT 101.115 182.875 101.625 183.410 ;
        RECT 101.845 183.080 102.090 183.685 ;
        RECT 103.120 183.595 103.290 183.850 ;
        RECT 102.625 183.425 103.290 183.595 ;
        RECT 103.565 183.550 103.745 184.350 ;
        RECT 102.625 183.045 102.795 183.425 ;
        RECT 102.975 182.875 103.305 183.255 ;
        RECT 103.485 183.045 103.745 183.550 ;
        RECT 105.500 183.420 105.840 184.250 ;
        RECT 107.320 183.740 107.670 184.990 ;
        RECT 109.435 184.260 109.725 185.425 ;
        RECT 109.900 185.000 110.235 185.425 ;
        RECT 110.405 184.820 110.590 185.225 ;
        RECT 109.925 184.645 110.590 184.820 ;
        RECT 110.795 184.645 111.125 185.425 ;
        RECT 109.925 183.615 110.265 184.645 ;
        RECT 111.295 184.455 111.565 185.225 ;
        RECT 110.435 184.285 111.565 184.455 ;
        RECT 111.735 184.335 115.245 185.425 ;
        RECT 110.435 183.785 110.685 184.285 ;
        RECT 103.915 182.875 109.260 183.420 ;
        RECT 109.435 182.875 109.725 183.600 ;
        RECT 109.925 183.445 110.610 183.615 ;
        RECT 110.865 183.535 111.225 184.115 ;
        RECT 109.900 182.875 110.235 183.275 ;
        RECT 110.405 183.045 110.610 183.445 ;
        RECT 111.395 183.375 111.565 184.285 ;
        RECT 110.820 182.875 111.095 183.355 ;
        RECT 111.305 183.045 111.565 183.375 ;
        RECT 111.735 183.645 113.385 184.165 ;
        RECT 113.555 183.815 115.245 184.335 ;
        RECT 115.415 184.350 115.685 185.255 ;
        RECT 115.855 184.665 116.185 185.425 ;
        RECT 116.365 184.495 116.545 185.255 ;
        RECT 116.885 184.875 117.055 185.165 ;
        RECT 117.225 185.045 117.555 185.425 ;
        RECT 118.120 184.915 118.950 185.085 ;
        RECT 116.885 184.745 117.375 184.875 ;
        RECT 116.885 184.705 118.610 184.745 ;
        RECT 117.205 184.575 118.610 184.705 ;
        RECT 111.735 182.875 115.245 183.645 ;
        RECT 115.415 183.550 115.595 184.350 ;
        RECT 115.870 184.325 116.545 184.495 ;
        RECT 115.870 184.180 116.040 184.325 ;
        RECT 115.765 183.850 116.040 184.180 ;
        RECT 115.870 183.595 116.040 183.850 ;
        RECT 116.265 183.775 116.605 184.145 ;
        RECT 116.855 183.765 117.035 184.535 ;
        RECT 117.205 183.595 117.375 184.575 ;
        RECT 117.715 184.235 118.100 184.405 ;
        RECT 117.930 184.075 118.100 184.235 ;
        RECT 118.270 184.365 118.610 184.575 ;
        RECT 115.415 183.045 115.675 183.550 ;
        RECT 115.870 183.425 116.535 183.595 ;
        RECT 115.855 182.875 116.185 183.255 ;
        RECT 116.365 183.045 116.535 183.425 ;
        RECT 116.880 183.425 117.375 183.595 ;
        RECT 117.545 183.555 117.945 183.885 ;
        RECT 118.270 183.825 118.440 184.365 ;
        RECT 118.780 184.195 118.950 184.915 ;
        RECT 119.305 184.845 119.535 185.425 ;
        RECT 120.015 184.915 120.530 185.085 ;
        RECT 119.680 184.575 120.025 184.745 ;
        RECT 120.275 184.600 120.530 184.915 ;
        RECT 119.855 184.450 120.025 184.575 ;
        RECT 119.855 184.280 120.125 184.450 ;
        RECT 116.880 183.135 117.055 183.425 ;
        RECT 117.225 182.875 117.555 183.255 ;
        RECT 117.730 183.185 117.945 183.555 ;
        RECT 118.115 183.495 118.440 183.825 ;
        RECT 118.610 184.025 118.950 184.195 ;
        RECT 119.955 184.180 120.125 184.280 ;
        RECT 118.610 183.325 118.780 184.025 ;
        RECT 119.120 183.805 119.325 184.110 ;
        RECT 118.950 183.505 119.325 183.805 ;
        RECT 119.495 183.505 119.785 184.110 ;
        RECT 119.955 183.850 120.190 184.180 ;
        RECT 118.180 183.155 118.780 183.325 ;
        RECT 119.160 182.875 119.490 183.335 ;
        RECT 119.955 183.255 120.125 183.850 ;
        RECT 120.360 183.465 120.530 184.600 ;
        RECT 119.695 183.085 120.125 183.255 ;
        RECT 120.295 183.135 120.530 183.465 ;
        RECT 120.700 184.915 121.225 185.085 ;
        RECT 120.700 183.135 120.890 184.915 ;
        RECT 121.465 184.795 121.810 185.425 ;
        RECT 122.035 184.945 122.985 185.115 ;
        RECT 121.105 184.525 121.295 184.685 ;
        RECT 122.035 184.525 122.205 184.945 ;
        RECT 123.235 184.915 123.555 185.085 ;
        RECT 121.105 184.355 122.205 184.525 ;
        RECT 121.105 183.375 121.275 184.355 ;
        RECT 121.455 183.505 121.825 184.185 ;
        RECT 121.105 183.045 121.310 183.375 ;
        RECT 121.505 182.875 121.835 183.335 ;
        RECT 122.035 183.255 122.205 184.355 ;
        RECT 122.375 183.825 122.665 184.775 ;
        RECT 123.385 184.455 123.555 184.915 ;
        RECT 123.725 184.625 123.895 185.425 ;
        RECT 124.065 184.625 124.475 185.245 ;
        RECT 122.835 184.035 123.175 184.435 ;
        RECT 123.385 184.285 123.995 184.455 ;
        RECT 124.165 184.285 124.475 184.625 ;
        RECT 124.645 184.285 124.895 185.425 ;
        RECT 125.075 184.335 126.285 185.425 ;
        RECT 123.825 184.115 123.995 184.285 ;
        RECT 123.345 183.865 123.655 184.115 ;
        RECT 122.375 183.495 122.995 183.825 ;
        RECT 123.245 183.785 123.655 183.865 ;
        RECT 123.825 183.785 124.135 184.115 ;
        RECT 122.035 183.085 122.930 183.255 ;
        RECT 123.245 183.165 123.555 183.785 ;
        RECT 123.725 182.875 123.975 183.605 ;
        RECT 124.305 183.515 124.475 184.285 ;
        RECT 124.145 183.055 124.475 183.515 ;
        RECT 124.645 182.875 124.900 183.675 ;
        RECT 125.075 183.625 125.595 184.165 ;
        RECT 125.765 183.795 126.285 184.335 ;
        RECT 126.535 184.495 126.715 185.255 ;
        RECT 126.895 184.665 127.225 185.425 ;
        RECT 126.535 184.325 127.210 184.495 ;
        RECT 127.395 184.350 127.665 185.255 ;
        RECT 127.040 184.180 127.210 184.325 ;
        RECT 126.475 183.775 126.815 184.145 ;
        RECT 127.040 183.850 127.315 184.180 ;
        RECT 125.075 182.875 126.285 183.625 ;
        RECT 127.040 183.595 127.210 183.850 ;
        RECT 126.545 183.425 127.210 183.595 ;
        RECT 127.485 183.550 127.665 184.350 ;
        RECT 126.545 183.045 126.715 183.425 ;
        RECT 126.895 182.875 127.225 183.255 ;
        RECT 127.405 183.045 127.665 183.550 ;
        RECT 127.835 184.350 128.105 185.255 ;
        RECT 128.275 184.665 128.605 185.425 ;
        RECT 128.785 184.495 128.965 185.255 ;
        RECT 127.835 183.550 128.015 184.350 ;
        RECT 128.290 184.325 128.965 184.495 ;
        RECT 130.145 184.365 130.475 185.215 ;
        RECT 128.290 184.180 128.460 184.325 ;
        RECT 128.185 183.850 128.460 184.180 ;
        RECT 130.145 184.235 130.365 184.365 ;
        RECT 130.645 184.285 130.895 185.425 ;
        RECT 131.085 184.785 131.335 185.205 ;
        RECT 131.565 184.955 131.895 185.425 ;
        RECT 132.125 184.785 132.375 185.205 ;
        RECT 131.085 184.615 132.375 184.785 ;
        RECT 132.555 184.785 132.885 185.215 ;
        RECT 132.555 184.615 133.010 184.785 ;
        RECT 128.290 183.595 128.460 183.850 ;
        RECT 128.685 183.775 129.025 184.145 ;
        RECT 130.145 183.600 130.335 184.235 ;
        RECT 131.075 184.115 131.290 184.445 ;
        RECT 130.505 183.785 130.815 184.115 ;
        RECT 130.985 183.785 131.290 184.115 ;
        RECT 131.465 183.785 131.750 184.445 ;
        RECT 131.945 183.785 132.210 184.445 ;
        RECT 132.425 183.785 132.670 184.445 ;
        RECT 130.645 183.615 130.815 183.785 ;
        RECT 132.840 183.615 133.010 184.615 ;
        RECT 133.355 184.335 135.025 185.425 ;
        RECT 127.835 183.045 128.095 183.550 ;
        RECT 128.290 183.425 128.955 183.595 ;
        RECT 128.275 182.875 128.605 183.255 ;
        RECT 128.785 183.045 128.955 183.425 ;
        RECT 130.145 183.090 130.475 183.600 ;
        RECT 130.645 183.445 133.010 183.615 ;
        RECT 133.355 183.645 134.105 184.165 ;
        RECT 134.275 183.815 135.025 184.335 ;
        RECT 135.195 184.260 135.485 185.425 ;
        RECT 135.655 184.350 135.925 185.255 ;
        RECT 136.095 184.665 136.425 185.425 ;
        RECT 136.605 184.495 136.785 185.255 ;
        RECT 137.035 184.830 137.470 185.255 ;
        RECT 137.640 185.000 138.025 185.425 ;
        RECT 137.035 184.660 138.025 184.830 ;
        RECT 130.645 182.875 130.975 183.275 ;
        RECT 132.025 183.105 132.355 183.445 ;
        RECT 132.525 182.875 132.855 183.275 ;
        RECT 133.355 182.875 135.025 183.645 ;
        RECT 135.195 182.875 135.485 183.600 ;
        RECT 135.655 183.550 135.835 184.350 ;
        RECT 136.110 184.325 136.785 184.495 ;
        RECT 136.110 184.180 136.280 184.325 ;
        RECT 136.005 183.850 136.280 184.180 ;
        RECT 136.110 183.595 136.280 183.850 ;
        RECT 136.505 183.775 136.845 184.145 ;
        RECT 137.035 183.785 137.520 184.490 ;
        RECT 137.690 184.115 138.025 184.660 ;
        RECT 138.195 184.465 138.620 185.255 ;
        RECT 138.790 184.830 139.065 185.255 ;
        RECT 139.235 185.000 139.620 185.425 ;
        RECT 138.790 184.635 139.620 184.830 ;
        RECT 138.195 184.285 139.100 184.465 ;
        RECT 137.690 183.785 138.100 184.115 ;
        RECT 138.270 183.785 139.100 184.285 ;
        RECT 139.270 184.115 139.620 184.635 ;
        RECT 139.790 184.465 140.035 185.255 ;
        RECT 140.225 184.830 140.480 185.255 ;
        RECT 140.650 185.000 141.035 185.425 ;
        RECT 140.225 184.635 141.035 184.830 ;
        RECT 139.790 184.285 140.515 184.465 ;
        RECT 139.270 183.785 139.695 184.115 ;
        RECT 139.865 183.785 140.515 184.285 ;
        RECT 140.685 184.115 141.035 184.635 ;
        RECT 141.205 184.285 141.465 185.255 ;
        RECT 142.095 184.830 142.530 185.255 ;
        RECT 142.700 185.000 143.085 185.425 ;
        RECT 142.095 184.660 143.085 184.830 ;
        RECT 140.685 183.785 141.110 184.115 ;
        RECT 137.690 183.615 138.025 183.785 ;
        RECT 138.270 183.615 138.620 183.785 ;
        RECT 139.270 183.615 139.620 183.785 ;
        RECT 139.865 183.615 140.035 183.785 ;
        RECT 140.685 183.615 141.035 183.785 ;
        RECT 141.280 183.615 141.465 184.285 ;
        RECT 142.095 183.785 142.580 184.490 ;
        RECT 142.750 184.115 143.085 184.660 ;
        RECT 143.255 184.465 143.680 185.255 ;
        RECT 143.850 184.830 144.125 185.255 ;
        RECT 144.295 185.000 144.680 185.425 ;
        RECT 143.850 184.635 144.680 184.830 ;
        RECT 143.255 184.285 144.160 184.465 ;
        RECT 142.750 183.785 143.160 184.115 ;
        RECT 143.330 183.785 144.160 184.285 ;
        RECT 144.330 184.115 144.680 184.635 ;
        RECT 144.850 184.465 145.095 185.255 ;
        RECT 145.285 184.830 145.540 185.255 ;
        RECT 145.710 185.000 146.095 185.425 ;
        RECT 145.285 184.635 146.095 184.830 ;
        RECT 144.850 184.285 145.575 184.465 ;
        RECT 144.330 183.785 144.755 184.115 ;
        RECT 144.925 183.785 145.575 184.285 ;
        RECT 145.745 184.115 146.095 184.635 ;
        RECT 146.265 184.285 146.525 185.255 ;
        RECT 147.245 184.755 147.415 185.255 ;
        RECT 147.585 184.925 147.915 185.425 ;
        RECT 147.245 184.585 147.910 184.755 ;
        RECT 145.745 183.785 146.170 184.115 ;
        RECT 142.750 183.615 143.085 183.785 ;
        RECT 143.330 183.615 143.680 183.785 ;
        RECT 144.330 183.615 144.680 183.785 ;
        RECT 144.925 183.615 145.095 183.785 ;
        RECT 145.745 183.615 146.095 183.785 ;
        RECT 146.340 183.615 146.525 184.285 ;
        RECT 147.160 183.765 147.510 184.415 ;
        RECT 135.655 183.045 135.915 183.550 ;
        RECT 136.110 183.425 136.775 183.595 ;
        RECT 136.095 182.875 136.425 183.255 ;
        RECT 136.605 183.045 136.775 183.425 ;
        RECT 137.035 183.445 138.025 183.615 ;
        RECT 137.035 183.045 137.470 183.445 ;
        RECT 137.640 182.875 138.025 183.275 ;
        RECT 138.195 183.045 138.620 183.615 ;
        RECT 138.810 183.445 139.620 183.615 ;
        RECT 138.810 183.045 139.065 183.445 ;
        RECT 139.235 182.875 139.620 183.275 ;
        RECT 139.790 183.045 140.035 183.615 ;
        RECT 140.225 183.445 141.035 183.615 ;
        RECT 140.225 183.045 140.480 183.445 ;
        RECT 140.650 182.875 141.035 183.275 ;
        RECT 141.205 183.045 141.465 183.615 ;
        RECT 142.095 183.445 143.085 183.615 ;
        RECT 142.095 183.045 142.530 183.445 ;
        RECT 142.700 182.875 143.085 183.275 ;
        RECT 143.255 183.045 143.680 183.615 ;
        RECT 143.870 183.445 144.680 183.615 ;
        RECT 143.870 183.045 144.125 183.445 ;
        RECT 144.295 182.875 144.680 183.275 ;
        RECT 144.850 183.045 145.095 183.615 ;
        RECT 145.285 183.445 146.095 183.615 ;
        RECT 145.285 183.045 145.540 183.445 ;
        RECT 145.710 182.875 146.095 183.275 ;
        RECT 146.265 183.045 146.525 183.615 ;
        RECT 147.680 183.595 147.910 184.585 ;
        RECT 147.245 183.425 147.910 183.595 ;
        RECT 147.245 183.135 147.415 183.425 ;
        RECT 147.585 182.875 147.915 183.255 ;
        RECT 148.085 183.135 148.270 185.255 ;
        RECT 148.510 184.965 148.775 185.425 ;
        RECT 148.945 184.830 149.195 185.255 ;
        RECT 149.405 184.980 150.510 185.150 ;
        RECT 148.890 184.700 149.195 184.830 ;
        RECT 148.440 183.505 148.720 184.455 ;
        RECT 148.890 183.595 149.060 184.700 ;
        RECT 149.230 183.915 149.470 184.510 ;
        RECT 149.640 184.445 150.170 184.810 ;
        RECT 149.640 183.745 149.810 184.445 ;
        RECT 150.340 184.365 150.510 184.980 ;
        RECT 150.680 184.625 150.850 185.425 ;
        RECT 151.020 184.925 151.270 185.255 ;
        RECT 151.495 184.955 152.380 185.125 ;
        RECT 150.340 184.275 150.850 184.365 ;
        RECT 148.890 183.465 149.115 183.595 ;
        RECT 149.285 183.525 149.810 183.745 ;
        RECT 149.980 184.105 150.850 184.275 ;
        RECT 148.525 182.875 148.775 183.335 ;
        RECT 148.945 183.325 149.115 183.465 ;
        RECT 149.980 183.325 150.150 184.105 ;
        RECT 150.680 184.035 150.850 184.105 ;
        RECT 150.360 183.855 150.560 183.885 ;
        RECT 151.020 183.855 151.190 184.925 ;
        RECT 151.360 184.035 151.550 184.755 ;
        RECT 150.360 183.555 151.190 183.855 ;
        RECT 151.720 183.825 152.040 184.785 ;
        RECT 148.945 183.155 149.280 183.325 ;
        RECT 149.475 183.155 150.150 183.325 ;
        RECT 150.470 182.875 150.840 183.375 ;
        RECT 151.020 183.325 151.190 183.555 ;
        RECT 151.575 183.495 152.040 183.825 ;
        RECT 152.210 184.115 152.380 184.955 ;
        RECT 152.560 184.925 152.875 185.425 ;
        RECT 153.105 184.695 153.445 185.255 ;
        RECT 152.550 184.320 153.445 184.695 ;
        RECT 153.615 184.415 153.785 185.425 ;
        RECT 153.255 184.115 153.445 184.320 ;
        RECT 153.955 184.365 154.285 185.210 ;
        RECT 153.955 184.285 154.345 184.365 ;
        RECT 154.130 184.235 154.345 184.285 ;
        RECT 152.210 183.785 153.085 184.115 ;
        RECT 153.255 183.785 154.005 184.115 ;
        RECT 152.210 183.325 152.380 183.785 ;
        RECT 153.255 183.615 153.455 183.785 ;
        RECT 154.175 183.655 154.345 184.235 ;
        RECT 154.975 184.335 156.185 185.425 ;
        RECT 154.975 183.795 155.495 184.335 ;
        RECT 154.120 183.615 154.345 183.655 ;
        RECT 155.665 183.625 156.185 184.165 ;
        RECT 151.020 183.155 151.425 183.325 ;
        RECT 151.595 183.155 152.380 183.325 ;
        RECT 152.655 182.875 152.865 183.405 ;
        RECT 153.125 183.090 153.455 183.615 ;
        RECT 153.965 183.530 154.345 183.615 ;
        RECT 153.625 182.875 153.795 183.485 ;
        RECT 153.965 183.095 154.295 183.530 ;
        RECT 154.975 182.875 156.185 183.625 ;
        RECT 70.710 182.705 156.270 182.875 ;
        RECT 70.795 181.955 72.005 182.705 ;
        RECT 72.265 182.155 72.435 182.445 ;
        RECT 72.605 182.325 72.935 182.705 ;
        RECT 72.265 181.985 72.930 182.155 ;
        RECT 70.795 181.415 71.315 181.955 ;
        RECT 71.485 181.245 72.005 181.785 ;
        RECT 70.795 180.155 72.005 181.245 ;
        RECT 72.180 181.165 72.530 181.815 ;
        RECT 72.700 180.995 72.930 181.985 ;
        RECT 72.265 180.825 72.930 180.995 ;
        RECT 72.265 180.325 72.435 180.825 ;
        RECT 72.605 180.155 72.935 180.655 ;
        RECT 73.105 180.325 73.290 182.445 ;
        RECT 73.545 182.245 73.795 182.705 ;
        RECT 73.965 182.255 74.300 182.425 ;
        RECT 74.495 182.255 75.170 182.425 ;
        RECT 73.965 182.115 74.135 182.255 ;
        RECT 73.460 181.125 73.740 182.075 ;
        RECT 73.910 181.985 74.135 182.115 ;
        RECT 73.910 180.880 74.080 181.985 ;
        RECT 74.305 181.835 74.830 182.055 ;
        RECT 74.250 181.070 74.490 181.665 ;
        RECT 74.660 181.135 74.830 181.835 ;
        RECT 75.000 181.475 75.170 182.255 ;
        RECT 75.490 182.205 75.860 182.705 ;
        RECT 76.040 182.255 76.445 182.425 ;
        RECT 76.615 182.255 77.400 182.425 ;
        RECT 76.040 182.025 76.210 182.255 ;
        RECT 75.380 181.725 76.210 182.025 ;
        RECT 76.595 181.755 77.060 182.085 ;
        RECT 75.380 181.695 75.580 181.725 ;
        RECT 75.700 181.475 75.870 181.545 ;
        RECT 75.000 181.305 75.870 181.475 ;
        RECT 75.360 181.215 75.870 181.305 ;
        RECT 73.910 180.750 74.215 180.880 ;
        RECT 74.660 180.770 75.190 181.135 ;
        RECT 73.530 180.155 73.795 180.615 ;
        RECT 73.965 180.325 74.215 180.750 ;
        RECT 75.360 180.600 75.530 181.215 ;
        RECT 74.425 180.430 75.530 180.600 ;
        RECT 75.700 180.155 75.870 180.955 ;
        RECT 76.040 180.655 76.210 181.725 ;
        RECT 76.380 180.825 76.570 181.545 ;
        RECT 76.740 180.795 77.060 181.755 ;
        RECT 77.230 181.795 77.400 182.255 ;
        RECT 77.675 182.175 77.885 182.705 ;
        RECT 78.145 181.965 78.475 182.490 ;
        RECT 78.645 182.095 78.815 182.705 ;
        RECT 78.985 182.050 79.315 182.485 ;
        RECT 78.985 181.965 79.365 182.050 ;
        RECT 78.275 181.795 78.475 181.965 ;
        RECT 79.140 181.925 79.365 181.965 ;
        RECT 77.230 181.465 78.105 181.795 ;
        RECT 78.275 181.465 79.025 181.795 ;
        RECT 76.040 180.325 76.290 180.655 ;
        RECT 77.230 180.625 77.400 181.465 ;
        RECT 78.275 181.260 78.465 181.465 ;
        RECT 79.195 181.345 79.365 181.925 ;
        RECT 79.535 181.935 82.125 182.705 ;
        RECT 82.845 182.155 83.015 182.535 ;
        RECT 83.195 182.325 83.525 182.705 ;
        RECT 82.845 181.985 83.510 182.155 ;
        RECT 83.705 182.030 83.965 182.535 ;
        RECT 79.535 181.415 80.745 181.935 ;
        RECT 79.150 181.295 79.365 181.345 ;
        RECT 77.570 180.885 78.465 181.260 ;
        RECT 78.975 181.215 79.365 181.295 ;
        RECT 80.915 181.245 82.125 181.765 ;
        RECT 82.775 181.435 83.105 181.805 ;
        RECT 83.340 181.730 83.510 181.985 ;
        RECT 83.340 181.400 83.625 181.730 ;
        RECT 83.340 181.255 83.510 181.400 ;
        RECT 76.515 180.455 77.400 180.625 ;
        RECT 77.580 180.155 77.895 180.655 ;
        RECT 78.125 180.325 78.465 180.885 ;
        RECT 78.635 180.155 78.805 181.165 ;
        RECT 78.975 180.370 79.305 181.215 ;
        RECT 79.535 180.155 82.125 181.245 ;
        RECT 82.845 181.085 83.510 181.255 ;
        RECT 83.795 181.230 83.965 182.030 ;
        RECT 84.655 181.885 84.865 182.705 ;
        RECT 85.035 181.905 85.365 182.535 ;
        RECT 85.035 181.305 85.285 181.905 ;
        RECT 85.535 181.885 85.765 182.705 ;
        RECT 85.975 182.030 86.235 182.535 ;
        RECT 86.415 182.325 86.745 182.705 ;
        RECT 86.925 182.155 87.095 182.535 ;
        RECT 85.455 181.465 85.785 181.715 ;
        RECT 82.845 180.325 83.015 181.085 ;
        RECT 83.195 180.155 83.525 180.915 ;
        RECT 83.695 180.325 83.965 181.230 ;
        RECT 84.655 180.155 84.865 181.295 ;
        RECT 85.035 180.325 85.365 181.305 ;
        RECT 85.535 180.155 85.765 181.295 ;
        RECT 85.975 181.230 86.155 182.030 ;
        RECT 86.430 181.985 87.095 182.155 ;
        RECT 86.430 181.730 86.600 181.985 ;
        RECT 87.355 181.965 87.615 182.535 ;
        RECT 87.785 182.305 88.170 182.705 ;
        RECT 88.340 182.135 88.595 182.535 ;
        RECT 87.785 181.965 88.595 182.135 ;
        RECT 88.785 181.965 89.030 182.535 ;
        RECT 89.200 182.305 89.585 182.705 ;
        RECT 89.755 182.135 90.010 182.535 ;
        RECT 89.200 181.965 90.010 182.135 ;
        RECT 90.200 181.965 90.625 182.535 ;
        RECT 90.795 182.305 91.180 182.705 ;
        RECT 91.350 182.135 91.785 182.535 ;
        RECT 90.795 181.965 91.785 182.135 ;
        RECT 91.955 182.135 92.390 182.535 ;
        RECT 92.560 182.305 92.945 182.705 ;
        RECT 91.955 181.965 92.945 182.135 ;
        RECT 93.115 181.965 93.540 182.535 ;
        RECT 93.730 182.135 93.985 182.535 ;
        RECT 94.155 182.305 94.540 182.705 ;
        RECT 93.730 181.965 94.540 182.135 ;
        RECT 94.710 181.965 94.955 182.535 ;
        RECT 95.145 182.135 95.400 182.535 ;
        RECT 95.570 182.305 95.955 182.705 ;
        RECT 95.145 181.965 95.955 182.135 ;
        RECT 96.125 181.965 96.385 182.535 ;
        RECT 96.555 181.980 96.845 182.705 ;
        RECT 97.015 182.245 97.575 182.535 ;
        RECT 97.745 182.245 97.995 182.705 ;
        RECT 86.325 181.400 86.600 181.730 ;
        RECT 86.825 181.435 87.165 181.805 ;
        RECT 86.430 181.255 86.600 181.400 ;
        RECT 87.355 181.295 87.540 181.965 ;
        RECT 87.785 181.795 88.135 181.965 ;
        RECT 88.785 181.795 88.955 181.965 ;
        RECT 89.200 181.795 89.550 181.965 ;
        RECT 90.200 181.795 90.550 181.965 ;
        RECT 90.795 181.795 91.130 181.965 ;
        RECT 92.610 181.795 92.945 181.965 ;
        RECT 93.190 181.795 93.540 181.965 ;
        RECT 94.190 181.795 94.540 181.965 ;
        RECT 94.785 181.795 94.955 181.965 ;
        RECT 95.605 181.795 95.955 181.965 ;
        RECT 87.710 181.465 88.135 181.795 ;
        RECT 85.975 180.325 86.245 181.230 ;
        RECT 86.430 181.085 87.105 181.255 ;
        RECT 86.415 180.155 86.745 180.915 ;
        RECT 86.925 180.325 87.105 181.085 ;
        RECT 87.355 180.325 87.615 181.295 ;
        RECT 87.785 180.945 88.135 181.465 ;
        RECT 88.305 181.295 88.955 181.795 ;
        RECT 89.125 181.465 89.550 181.795 ;
        RECT 88.305 181.115 89.030 181.295 ;
        RECT 87.785 180.750 88.595 180.945 ;
        RECT 87.785 180.155 88.170 180.580 ;
        RECT 88.340 180.325 88.595 180.750 ;
        RECT 88.785 180.325 89.030 181.115 ;
        RECT 89.200 180.945 89.550 181.465 ;
        RECT 89.720 181.295 90.550 181.795 ;
        RECT 90.720 181.465 91.130 181.795 ;
        RECT 89.720 181.115 90.625 181.295 ;
        RECT 89.200 180.750 90.030 180.945 ;
        RECT 89.200 180.155 89.585 180.580 ;
        RECT 89.755 180.325 90.030 180.750 ;
        RECT 90.200 180.325 90.625 181.115 ;
        RECT 90.795 180.920 91.130 181.465 ;
        RECT 91.300 181.090 91.785 181.795 ;
        RECT 91.955 181.090 92.440 181.795 ;
        RECT 92.610 181.465 93.020 181.795 ;
        RECT 92.610 180.920 92.945 181.465 ;
        RECT 93.190 181.295 94.020 181.795 ;
        RECT 90.795 180.750 91.785 180.920 ;
        RECT 90.795 180.155 91.180 180.580 ;
        RECT 91.350 180.325 91.785 180.750 ;
        RECT 91.955 180.750 92.945 180.920 ;
        RECT 93.115 181.115 94.020 181.295 ;
        RECT 94.190 181.465 94.615 181.795 ;
        RECT 91.955 180.325 92.390 180.750 ;
        RECT 92.560 180.155 92.945 180.580 ;
        RECT 93.115 180.325 93.540 181.115 ;
        RECT 94.190 180.945 94.540 181.465 ;
        RECT 94.785 181.295 95.435 181.795 ;
        RECT 93.710 180.750 94.540 180.945 ;
        RECT 94.710 181.115 95.435 181.295 ;
        RECT 95.605 181.465 96.030 181.795 ;
        RECT 93.710 180.325 93.985 180.750 ;
        RECT 94.155 180.155 94.540 180.580 ;
        RECT 94.710 180.325 94.955 181.115 ;
        RECT 95.605 180.945 95.955 181.465 ;
        RECT 96.200 181.295 96.385 181.965 ;
        RECT 95.145 180.750 95.955 180.945 ;
        RECT 95.145 180.325 95.400 180.750 ;
        RECT 95.570 180.155 95.955 180.580 ;
        RECT 96.125 180.325 96.385 181.295 ;
        RECT 96.555 180.155 96.845 181.320 ;
        RECT 97.015 180.875 97.265 182.245 ;
        RECT 98.615 182.075 98.945 182.435 ;
        RECT 97.555 181.885 98.945 182.075 ;
        RECT 99.315 182.135 99.750 182.535 ;
        RECT 99.920 182.305 100.305 182.705 ;
        RECT 99.315 181.965 100.305 182.135 ;
        RECT 100.475 181.965 100.900 182.535 ;
        RECT 101.090 182.135 101.345 182.535 ;
        RECT 101.515 182.305 101.900 182.705 ;
        RECT 101.090 181.965 101.900 182.135 ;
        RECT 102.070 181.965 102.315 182.535 ;
        RECT 102.505 182.135 102.760 182.535 ;
        RECT 102.930 182.305 103.315 182.705 ;
        RECT 102.505 181.965 103.315 182.135 ;
        RECT 103.485 181.965 103.745 182.535 ;
        RECT 97.555 181.795 97.725 181.885 ;
        RECT 99.970 181.795 100.305 181.965 ;
        RECT 100.550 181.795 100.900 181.965 ;
        RECT 101.550 181.795 101.900 181.965 ;
        RECT 102.145 181.795 102.315 181.965 ;
        RECT 102.965 181.795 103.315 181.965 ;
        RECT 97.435 181.465 97.725 181.795 ;
        RECT 97.895 181.465 98.235 181.715 ;
        RECT 98.455 181.465 99.130 181.715 ;
        RECT 97.555 181.215 97.725 181.465 ;
        RECT 97.555 181.045 98.495 181.215 ;
        RECT 98.865 181.105 99.130 181.465 ;
        RECT 99.315 181.090 99.800 181.795 ;
        RECT 99.970 181.465 100.380 181.795 ;
        RECT 97.015 180.325 97.475 180.875 ;
        RECT 97.665 180.155 97.995 180.875 ;
        RECT 98.195 180.495 98.495 181.045 ;
        RECT 99.970 180.920 100.305 181.465 ;
        RECT 100.550 181.295 101.380 181.795 ;
        RECT 98.665 180.155 98.945 180.825 ;
        RECT 99.315 180.750 100.305 180.920 ;
        RECT 100.475 181.115 101.380 181.295 ;
        RECT 101.550 181.465 101.975 181.795 ;
        RECT 99.315 180.325 99.750 180.750 ;
        RECT 99.920 180.155 100.305 180.580 ;
        RECT 100.475 180.325 100.900 181.115 ;
        RECT 101.550 180.945 101.900 181.465 ;
        RECT 102.145 181.295 102.795 181.795 ;
        RECT 101.070 180.750 101.900 180.945 ;
        RECT 102.070 181.115 102.795 181.295 ;
        RECT 102.965 181.465 103.390 181.795 ;
        RECT 101.070 180.325 101.345 180.750 ;
        RECT 101.515 180.155 101.900 180.580 ;
        RECT 102.070 180.325 102.315 181.115 ;
        RECT 102.965 180.945 103.315 181.465 ;
        RECT 103.560 181.295 103.745 181.965 ;
        RECT 102.505 180.750 103.315 180.945 ;
        RECT 102.505 180.325 102.760 180.750 ;
        RECT 102.930 180.155 103.315 180.580 ;
        RECT 103.485 180.325 103.745 181.295 ;
        RECT 103.920 182.230 104.255 182.490 ;
        RECT 104.425 182.305 104.755 182.705 ;
        RECT 104.925 182.305 106.540 182.475 ;
        RECT 103.920 180.875 104.175 182.230 ;
        RECT 104.925 182.135 105.095 182.305 ;
        RECT 104.535 181.965 105.095 182.135 ;
        RECT 104.535 181.795 104.705 181.965 ;
        RECT 104.400 181.465 104.705 181.795 ;
        RECT 104.900 181.685 105.150 181.795 ;
        RECT 105.360 181.685 105.630 182.125 ;
        RECT 105.820 182.025 106.110 182.125 ;
        RECT 105.815 181.855 106.110 182.025 ;
        RECT 104.895 181.515 105.150 181.685 ;
        RECT 105.355 181.515 105.630 181.685 ;
        RECT 104.900 181.465 105.150 181.515 ;
        RECT 105.360 181.465 105.630 181.515 ;
        RECT 105.820 181.465 106.110 181.855 ;
        RECT 106.280 181.465 106.700 182.130 ;
        RECT 107.085 181.985 107.415 182.705 ;
        RECT 107.595 182.245 108.155 182.535 ;
        RECT 108.325 182.245 108.575 182.705 ;
        RECT 107.010 181.465 107.360 181.795 ;
        RECT 104.535 181.295 104.705 181.465 ;
        RECT 107.155 181.345 107.360 181.465 ;
        RECT 104.535 181.125 106.905 181.295 ;
        RECT 107.155 181.175 107.365 181.345 ;
        RECT 103.920 180.365 104.255 180.875 ;
        RECT 104.505 180.155 104.835 180.955 ;
        RECT 105.080 180.745 106.505 180.915 ;
        RECT 105.080 180.325 105.365 180.745 ;
        RECT 105.620 180.155 105.950 180.575 ;
        RECT 106.175 180.495 106.505 180.745 ;
        RECT 106.735 180.665 106.905 181.125 ;
        RECT 107.165 180.495 107.335 180.995 ;
        RECT 106.175 180.325 107.335 180.495 ;
        RECT 107.595 180.875 107.845 182.245 ;
        RECT 109.195 182.075 109.525 182.435 ;
        RECT 108.135 181.885 109.525 182.075 ;
        RECT 109.895 182.030 110.155 182.535 ;
        RECT 110.335 182.325 110.665 182.705 ;
        RECT 110.845 182.155 111.015 182.535 ;
        RECT 111.275 182.160 116.620 182.705 ;
        RECT 116.795 182.160 122.140 182.705 ;
        RECT 108.135 181.795 108.305 181.885 ;
        RECT 108.015 181.465 108.305 181.795 ;
        RECT 108.475 181.465 108.815 181.715 ;
        RECT 109.035 181.465 109.710 181.715 ;
        RECT 108.135 181.215 108.305 181.465 ;
        RECT 108.135 181.045 109.075 181.215 ;
        RECT 109.445 181.105 109.710 181.465 ;
        RECT 109.895 181.230 110.075 182.030 ;
        RECT 110.350 181.985 111.015 182.155 ;
        RECT 110.350 181.730 110.520 181.985 ;
        RECT 110.245 181.400 110.520 181.730 ;
        RECT 110.745 181.435 111.085 181.805 ;
        RECT 110.350 181.255 110.520 181.400 ;
        RECT 112.860 181.330 113.200 182.160 ;
        RECT 107.595 180.325 108.055 180.875 ;
        RECT 108.245 180.155 108.575 180.875 ;
        RECT 108.775 180.495 109.075 181.045 ;
        RECT 109.245 180.155 109.525 180.825 ;
        RECT 109.895 180.325 110.165 181.230 ;
        RECT 110.350 181.085 111.025 181.255 ;
        RECT 110.335 180.155 110.665 180.915 ;
        RECT 110.845 180.325 111.025 181.085 ;
        RECT 114.680 180.590 115.030 181.840 ;
        RECT 118.380 181.330 118.720 182.160 ;
        RECT 122.315 181.980 122.605 182.705 ;
        RECT 122.775 181.935 124.445 182.705 ;
        RECT 125.165 182.155 125.335 182.445 ;
        RECT 125.505 182.325 125.835 182.705 ;
        RECT 125.165 181.985 125.830 182.155 ;
        RECT 120.200 180.590 120.550 181.840 ;
        RECT 122.775 181.415 123.525 181.935 ;
        RECT 111.275 180.155 116.620 180.590 ;
        RECT 116.795 180.155 122.140 180.590 ;
        RECT 122.315 180.155 122.605 181.320 ;
        RECT 123.695 181.245 124.445 181.765 ;
        RECT 122.775 180.155 124.445 181.245 ;
        RECT 125.080 181.165 125.430 181.815 ;
        RECT 125.600 180.995 125.830 181.985 ;
        RECT 125.165 180.825 125.830 180.995 ;
        RECT 125.165 180.325 125.335 180.825 ;
        RECT 125.505 180.155 125.835 180.655 ;
        RECT 126.005 180.325 126.190 182.445 ;
        RECT 126.445 182.245 126.695 182.705 ;
        RECT 126.865 182.255 127.200 182.425 ;
        RECT 127.395 182.255 128.070 182.425 ;
        RECT 126.865 182.115 127.035 182.255 ;
        RECT 126.360 181.125 126.640 182.075 ;
        RECT 126.810 181.985 127.035 182.115 ;
        RECT 126.810 180.880 126.980 181.985 ;
        RECT 127.205 181.835 127.730 182.055 ;
        RECT 127.150 181.070 127.390 181.665 ;
        RECT 127.560 181.135 127.730 181.835 ;
        RECT 127.900 181.475 128.070 182.255 ;
        RECT 128.390 182.205 128.760 182.705 ;
        RECT 128.940 182.255 129.345 182.425 ;
        RECT 129.515 182.255 130.300 182.425 ;
        RECT 128.940 182.025 129.110 182.255 ;
        RECT 128.280 181.725 129.110 182.025 ;
        RECT 129.495 181.755 129.960 182.085 ;
        RECT 128.280 181.695 128.480 181.725 ;
        RECT 128.600 181.475 128.770 181.545 ;
        RECT 127.900 181.305 128.770 181.475 ;
        RECT 128.260 181.215 128.770 181.305 ;
        RECT 126.810 180.750 127.115 180.880 ;
        RECT 127.560 180.770 128.090 181.135 ;
        RECT 126.430 180.155 126.695 180.615 ;
        RECT 126.865 180.325 127.115 180.750 ;
        RECT 128.260 180.600 128.430 181.215 ;
        RECT 127.325 180.430 128.430 180.600 ;
        RECT 128.600 180.155 128.770 180.955 ;
        RECT 128.940 180.655 129.110 181.725 ;
        RECT 129.280 180.825 129.470 181.545 ;
        RECT 129.640 180.795 129.960 181.755 ;
        RECT 130.130 181.795 130.300 182.255 ;
        RECT 130.575 182.175 130.785 182.705 ;
        RECT 131.045 181.965 131.375 182.490 ;
        RECT 131.545 182.095 131.715 182.705 ;
        RECT 131.885 182.050 132.215 182.485 ;
        RECT 131.885 181.965 132.265 182.050 ;
        RECT 131.175 181.795 131.375 181.965 ;
        RECT 132.040 181.925 132.265 181.965 ;
        RECT 130.130 181.465 131.005 181.795 ;
        RECT 131.175 181.465 131.925 181.795 ;
        RECT 128.940 180.325 129.190 180.655 ;
        RECT 130.130 180.625 130.300 181.465 ;
        RECT 131.175 181.260 131.365 181.465 ;
        RECT 132.095 181.345 132.265 181.925 ;
        RECT 132.435 181.935 135.945 182.705 ;
        RECT 132.435 181.415 134.085 181.935 ;
        RECT 136.585 181.895 136.855 182.705 ;
        RECT 137.025 181.895 137.355 182.535 ;
        RECT 137.525 181.895 137.765 182.705 ;
        RECT 137.960 182.200 138.295 182.705 ;
        RECT 138.465 182.135 138.705 182.510 ;
        RECT 138.985 182.375 139.155 182.520 ;
        RECT 138.985 182.180 139.360 182.375 ;
        RECT 139.720 182.210 140.115 182.705 ;
        RECT 132.050 181.295 132.265 181.345 ;
        RECT 130.470 180.885 131.365 181.260 ;
        RECT 131.875 181.215 132.265 181.295 ;
        RECT 134.255 181.245 135.945 181.765 ;
        RECT 136.575 181.465 136.925 181.715 ;
        RECT 137.095 181.295 137.265 181.895 ;
        RECT 137.435 181.465 137.785 181.715 ;
        RECT 129.415 180.455 130.300 180.625 ;
        RECT 130.480 180.155 130.795 180.655 ;
        RECT 131.025 180.325 131.365 180.885 ;
        RECT 131.535 180.155 131.705 181.165 ;
        RECT 131.875 180.370 132.205 181.215 ;
        RECT 132.435 180.155 135.945 181.245 ;
        RECT 136.585 180.155 136.915 181.295 ;
        RECT 137.095 181.125 137.775 181.295 ;
        RECT 138.015 181.175 138.315 182.025 ;
        RECT 138.485 181.985 138.705 182.135 ;
        RECT 138.485 181.655 139.020 181.985 ;
        RECT 139.190 181.845 139.360 182.180 ;
        RECT 140.285 182.015 140.525 182.535 ;
        RECT 137.445 180.340 137.775 181.125 ;
        RECT 138.485 181.005 138.720 181.655 ;
        RECT 139.190 181.485 140.175 181.845 ;
        RECT 138.045 180.775 138.720 181.005 ;
        RECT 138.890 181.465 140.175 181.485 ;
        RECT 138.890 181.315 139.750 181.465 ;
        RECT 140.350 181.345 140.525 182.015 ;
        RECT 140.805 182.155 140.975 182.445 ;
        RECT 141.145 182.325 141.475 182.705 ;
        RECT 140.805 181.985 141.470 182.155 ;
        RECT 138.045 180.345 138.215 180.775 ;
        RECT 138.385 180.155 138.715 180.605 ;
        RECT 138.890 180.370 139.175 181.315 ;
        RECT 140.315 181.210 140.525 181.345 ;
        RECT 139.350 180.835 140.045 181.145 ;
        RECT 139.355 180.155 140.040 180.625 ;
        RECT 140.220 180.425 140.525 181.210 ;
        RECT 140.720 181.165 141.070 181.815 ;
        RECT 141.240 180.995 141.470 181.985 ;
        RECT 140.805 180.825 141.470 180.995 ;
        RECT 140.805 180.325 140.975 180.825 ;
        RECT 141.145 180.155 141.475 180.655 ;
        RECT 141.645 180.325 141.830 182.445 ;
        RECT 142.085 182.245 142.335 182.705 ;
        RECT 142.505 182.255 142.840 182.425 ;
        RECT 143.035 182.255 143.710 182.425 ;
        RECT 142.505 182.115 142.675 182.255 ;
        RECT 142.000 181.125 142.280 182.075 ;
        RECT 142.450 181.985 142.675 182.115 ;
        RECT 142.450 180.880 142.620 181.985 ;
        RECT 142.845 181.835 143.370 182.055 ;
        RECT 142.790 181.070 143.030 181.665 ;
        RECT 143.200 181.135 143.370 181.835 ;
        RECT 143.540 181.475 143.710 182.255 ;
        RECT 144.030 182.205 144.400 182.705 ;
        RECT 144.580 182.255 144.985 182.425 ;
        RECT 145.155 182.255 145.940 182.425 ;
        RECT 144.580 182.025 144.750 182.255 ;
        RECT 143.920 181.725 144.750 182.025 ;
        RECT 145.135 181.755 145.600 182.085 ;
        RECT 143.920 181.695 144.120 181.725 ;
        RECT 144.240 181.475 144.410 181.545 ;
        RECT 143.540 181.305 144.410 181.475 ;
        RECT 143.900 181.215 144.410 181.305 ;
        RECT 142.450 180.750 142.755 180.880 ;
        RECT 143.200 180.770 143.730 181.135 ;
        RECT 142.070 180.155 142.335 180.615 ;
        RECT 142.505 180.325 142.755 180.750 ;
        RECT 143.900 180.600 144.070 181.215 ;
        RECT 142.965 180.430 144.070 180.600 ;
        RECT 144.240 180.155 144.410 180.955 ;
        RECT 144.580 180.655 144.750 181.725 ;
        RECT 144.920 180.825 145.110 181.545 ;
        RECT 145.280 180.795 145.600 181.755 ;
        RECT 145.770 181.795 145.940 182.255 ;
        RECT 146.215 182.175 146.425 182.705 ;
        RECT 146.685 181.965 147.015 182.490 ;
        RECT 147.185 182.095 147.355 182.705 ;
        RECT 147.525 182.050 147.855 182.485 ;
        RECT 147.525 181.965 147.905 182.050 ;
        RECT 148.075 181.980 148.365 182.705 ;
        RECT 146.815 181.795 147.015 181.965 ;
        RECT 147.680 181.925 147.905 181.965 ;
        RECT 145.770 181.465 146.645 181.795 ;
        RECT 146.815 181.465 147.565 181.795 ;
        RECT 144.580 180.325 144.830 180.655 ;
        RECT 145.770 180.625 145.940 181.465 ;
        RECT 146.815 181.260 147.005 181.465 ;
        RECT 147.735 181.345 147.905 181.925 ;
        RECT 149.455 181.870 149.745 182.705 ;
        RECT 149.915 182.305 150.870 182.475 ;
        RECT 151.285 182.315 151.615 182.705 ;
        RECT 149.915 181.425 150.085 182.305 ;
        RECT 151.785 182.135 151.955 182.455 ;
        RECT 152.125 182.315 152.455 182.705 ;
        RECT 152.675 182.245 153.235 182.535 ;
        RECT 153.405 182.245 153.655 182.705 ;
        RECT 150.255 181.965 152.505 182.135 ;
        RECT 150.255 181.465 150.485 181.965 ;
        RECT 150.655 181.545 151.030 181.715 ;
        RECT 147.690 181.295 147.905 181.345 ;
        RECT 146.110 180.885 147.005 181.260 ;
        RECT 147.515 181.215 147.905 181.295 ;
        RECT 145.055 180.455 145.940 180.625 ;
        RECT 146.120 180.155 146.435 180.655 ;
        RECT 146.665 180.325 147.005 180.885 ;
        RECT 147.175 180.155 147.345 181.165 ;
        RECT 147.515 180.370 147.845 181.215 ;
        RECT 148.075 180.155 148.365 181.320 ;
        RECT 149.455 181.255 150.085 181.425 ;
        RECT 150.860 181.345 151.030 181.545 ;
        RECT 151.200 181.515 151.750 181.715 ;
        RECT 151.920 181.345 152.165 181.795 ;
        RECT 149.455 180.325 149.775 181.255 ;
        RECT 150.860 181.175 152.165 181.345 ;
        RECT 152.335 181.005 152.505 181.965 ;
        RECT 149.955 180.835 151.195 181.005 ;
        RECT 149.955 180.325 150.355 180.835 ;
        RECT 150.525 180.155 150.695 180.665 ;
        RECT 150.865 180.325 151.195 180.835 ;
        RECT 151.365 180.155 151.535 181.005 ;
        RECT 152.125 180.325 152.505 181.005 ;
        RECT 152.675 180.875 152.925 182.245 ;
        RECT 154.275 182.075 154.605 182.435 ;
        RECT 153.215 181.885 154.605 182.075 ;
        RECT 154.975 181.955 156.185 182.705 ;
        RECT 153.215 181.795 153.385 181.885 ;
        RECT 153.095 181.465 153.385 181.795 ;
        RECT 153.555 181.465 153.895 181.715 ;
        RECT 154.115 181.465 154.790 181.715 ;
        RECT 153.215 181.215 153.385 181.465 ;
        RECT 153.215 181.045 154.155 181.215 ;
        RECT 154.525 181.105 154.790 181.465 ;
        RECT 154.975 181.245 155.495 181.785 ;
        RECT 155.665 181.415 156.185 181.955 ;
        RECT 152.675 180.325 153.135 180.875 ;
        RECT 153.325 180.155 153.655 180.875 ;
        RECT 153.855 180.495 154.155 181.045 ;
        RECT 154.325 180.155 154.605 180.825 ;
        RECT 154.975 180.155 156.185 181.245 ;
        RECT 70.710 179.985 156.270 180.155 ;
        RECT 70.795 178.895 72.005 179.985 ;
        RECT 72.175 178.895 74.765 179.985 ;
        RECT 70.795 178.185 71.315 178.725 ;
        RECT 71.485 178.355 72.005 178.895 ;
        RECT 72.175 178.205 73.385 178.725 ;
        RECT 73.555 178.375 74.765 178.895 ;
        RECT 74.945 179.015 75.275 179.800 ;
        RECT 74.945 178.845 75.625 179.015 ;
        RECT 75.805 178.845 76.135 179.985 ;
        RECT 76.775 179.115 77.050 179.815 ;
        RECT 77.220 179.440 77.475 179.985 ;
        RECT 77.645 179.475 78.125 179.815 ;
        RECT 78.300 179.430 78.905 179.985 ;
        RECT 78.290 179.330 78.905 179.430 ;
        RECT 78.290 179.305 78.475 179.330 ;
        RECT 74.935 178.425 75.285 178.675 ;
        RECT 75.455 178.245 75.625 178.845 ;
        RECT 75.795 178.425 76.145 178.675 ;
        RECT 70.795 177.435 72.005 178.185 ;
        RECT 72.175 177.435 74.765 178.205 ;
        RECT 74.955 177.435 75.195 178.245 ;
        RECT 75.365 177.605 75.695 178.245 ;
        RECT 75.865 177.435 76.135 178.245 ;
        RECT 76.775 178.085 76.945 179.115 ;
        RECT 77.220 178.985 77.975 179.235 ;
        RECT 78.145 179.060 78.475 179.305 ;
        RECT 79.080 179.185 79.335 179.985 ;
        RECT 77.220 178.950 77.990 178.985 ;
        RECT 77.220 178.940 78.005 178.950 ;
        RECT 77.115 178.925 78.010 178.940 ;
        RECT 77.115 178.910 78.030 178.925 ;
        RECT 77.115 178.900 78.050 178.910 ;
        RECT 77.115 178.890 78.075 178.900 ;
        RECT 77.115 178.860 78.145 178.890 ;
        RECT 77.115 178.830 78.165 178.860 ;
        RECT 77.115 178.800 78.185 178.830 ;
        RECT 77.115 178.775 78.215 178.800 ;
        RECT 77.115 178.740 78.250 178.775 ;
        RECT 77.115 178.735 78.280 178.740 ;
        RECT 77.115 178.340 77.345 178.735 ;
        RECT 77.890 178.730 78.280 178.735 ;
        RECT 77.915 178.720 78.280 178.730 ;
        RECT 77.930 178.715 78.280 178.720 ;
        RECT 77.945 178.710 78.280 178.715 ;
        RECT 78.645 178.710 78.905 179.160 ;
        RECT 79.535 179.135 79.865 179.815 ;
        RECT 77.945 178.705 78.905 178.710 ;
        RECT 77.955 178.695 78.905 178.705 ;
        RECT 77.965 178.690 78.905 178.695 ;
        RECT 77.975 178.680 78.905 178.690 ;
        RECT 77.980 178.670 78.905 178.680 ;
        RECT 77.985 178.665 78.905 178.670 ;
        RECT 77.995 178.650 78.905 178.665 ;
        RECT 78.000 178.635 78.905 178.650 ;
        RECT 79.080 178.645 79.325 179.005 ;
        RECT 79.515 178.855 79.865 179.135 ;
        RECT 78.010 178.610 78.905 178.635 ;
        RECT 77.515 178.140 77.845 178.565 ;
        RECT 76.775 177.605 77.035 178.085 ;
        RECT 77.205 177.435 77.455 177.975 ;
        RECT 77.625 177.655 77.845 178.140 ;
        RECT 78.015 178.540 78.905 178.610 ;
        RECT 78.015 177.815 78.185 178.540 ;
        RECT 79.515 178.475 79.685 178.855 ;
        RECT 80.045 178.675 80.240 179.725 ;
        RECT 80.420 178.845 80.740 179.985 ;
        RECT 80.915 178.895 83.505 179.985 ;
        RECT 78.355 177.985 78.905 178.370 ;
        RECT 79.165 178.305 79.685 178.475 ;
        RECT 79.855 178.345 80.240 178.675 ;
        RECT 80.420 178.625 80.680 178.675 ;
        RECT 80.420 178.455 80.685 178.625 ;
        RECT 80.420 178.345 80.680 178.455 ;
        RECT 79.165 177.945 79.335 178.305 ;
        RECT 80.915 178.205 82.125 178.725 ;
        RECT 82.295 178.375 83.505 178.895 ;
        RECT 83.675 178.820 83.965 179.985 ;
        RECT 84.135 178.895 85.805 179.985 ;
        RECT 84.135 178.205 84.885 178.725 ;
        RECT 85.055 178.375 85.805 178.895 ;
        RECT 86.435 178.910 86.705 179.815 ;
        RECT 86.875 179.225 87.205 179.985 ;
        RECT 87.385 179.055 87.565 179.815 ;
        RECT 78.015 177.645 78.905 177.815 ;
        RECT 79.135 177.775 79.335 177.945 ;
        RECT 79.165 177.740 79.335 177.775 ;
        RECT 79.525 177.965 80.740 178.135 ;
        RECT 79.525 177.660 79.755 177.965 ;
        RECT 79.925 177.435 80.255 177.795 ;
        RECT 80.450 177.615 80.740 177.965 ;
        RECT 80.915 177.435 83.505 178.205 ;
        RECT 83.675 177.435 83.965 178.160 ;
        RECT 84.135 177.435 85.805 178.205 ;
        RECT 86.435 178.110 86.615 178.910 ;
        RECT 86.890 178.885 87.565 179.055 ;
        RECT 87.815 179.135 88.075 179.815 ;
        RECT 88.245 179.205 88.495 179.985 ;
        RECT 88.745 179.435 88.995 179.815 ;
        RECT 89.165 179.605 89.520 179.985 ;
        RECT 90.525 179.595 90.860 179.815 ;
        RECT 90.125 179.435 90.355 179.475 ;
        RECT 88.745 179.235 90.355 179.435 ;
        RECT 88.745 179.225 89.580 179.235 ;
        RECT 90.170 179.145 90.355 179.235 ;
        RECT 86.890 178.740 87.060 178.885 ;
        RECT 86.785 178.410 87.060 178.740 ;
        RECT 86.890 178.155 87.060 178.410 ;
        RECT 87.285 178.335 87.625 178.705 ;
        RECT 86.435 177.605 86.695 178.110 ;
        RECT 86.890 177.985 87.555 178.155 ;
        RECT 86.875 177.435 87.205 177.815 ;
        RECT 87.385 177.605 87.555 177.985 ;
        RECT 87.815 177.935 87.985 179.135 ;
        RECT 89.685 179.035 90.015 179.065 ;
        RECT 88.215 178.975 90.015 179.035 ;
        RECT 90.605 178.975 90.860 179.595 ;
        RECT 91.125 179.240 91.395 179.985 ;
        RECT 92.025 179.980 98.300 179.985 ;
        RECT 91.565 179.070 91.855 179.810 ;
        RECT 92.025 179.255 92.280 179.980 ;
        RECT 92.465 179.085 92.725 179.810 ;
        RECT 92.895 179.255 93.140 179.980 ;
        RECT 93.325 179.085 93.585 179.810 ;
        RECT 93.755 179.255 94.000 179.980 ;
        RECT 94.185 179.085 94.445 179.810 ;
        RECT 94.615 179.255 94.860 179.980 ;
        RECT 95.030 179.085 95.290 179.810 ;
        RECT 95.460 179.255 95.720 179.980 ;
        RECT 95.890 179.085 96.150 179.810 ;
        RECT 96.320 179.255 96.580 179.980 ;
        RECT 96.750 179.085 97.010 179.810 ;
        RECT 97.180 179.255 97.440 179.980 ;
        RECT 97.610 179.085 97.870 179.810 ;
        RECT 98.040 179.185 98.300 179.980 ;
        RECT 92.465 179.070 97.870 179.085 ;
        RECT 88.155 178.865 90.860 178.975 ;
        RECT 91.125 178.965 97.870 179.070 ;
        RECT 88.155 178.830 88.355 178.865 ;
        RECT 88.155 178.255 88.325 178.830 ;
        RECT 89.685 178.805 90.860 178.865 ;
        RECT 91.095 178.845 97.870 178.965 ;
        RECT 91.095 178.795 92.290 178.845 ;
        RECT 88.555 178.390 88.965 178.695 ;
        RECT 89.135 178.425 89.465 178.635 ;
        RECT 88.155 178.135 88.425 178.255 ;
        RECT 88.155 178.090 89.000 178.135 ;
        RECT 88.245 177.965 89.000 178.090 ;
        RECT 89.255 178.025 89.465 178.425 ;
        RECT 89.710 178.425 90.185 178.635 ;
        RECT 90.375 178.425 90.865 178.625 ;
        RECT 89.710 178.025 89.930 178.425 ;
        RECT 91.125 178.255 92.290 178.795 ;
        RECT 98.470 178.675 98.720 179.810 ;
        RECT 98.900 179.175 99.160 179.985 ;
        RECT 99.335 178.675 99.580 179.815 ;
        RECT 99.760 179.175 100.055 179.985 ;
        RECT 100.235 178.895 103.745 179.985 ;
        RECT 92.460 178.425 99.580 178.675 ;
        RECT 87.815 177.605 88.075 177.935 ;
        RECT 88.830 177.815 89.000 177.965 ;
        RECT 88.245 177.435 88.575 177.795 ;
        RECT 88.830 177.605 90.130 177.815 ;
        RECT 90.405 177.435 90.860 178.200 ;
        RECT 91.125 178.085 97.870 178.255 ;
        RECT 91.125 177.435 91.425 177.915 ;
        RECT 91.595 177.630 91.855 178.085 ;
        RECT 92.025 177.435 92.285 177.915 ;
        RECT 92.465 177.630 92.725 178.085 ;
        RECT 92.895 177.435 93.145 177.915 ;
        RECT 93.325 177.630 93.585 178.085 ;
        RECT 93.755 177.435 94.005 177.915 ;
        RECT 94.185 177.630 94.445 178.085 ;
        RECT 94.615 177.435 94.860 177.915 ;
        RECT 95.030 177.630 95.305 178.085 ;
        RECT 95.475 177.435 95.720 177.915 ;
        RECT 95.890 177.630 96.150 178.085 ;
        RECT 96.320 177.435 96.580 177.915 ;
        RECT 96.750 177.630 97.010 178.085 ;
        RECT 97.180 177.435 97.440 177.915 ;
        RECT 97.610 177.630 97.870 178.085 ;
        RECT 98.040 177.435 98.300 177.995 ;
        RECT 98.470 177.615 98.720 178.425 ;
        RECT 98.900 177.435 99.160 177.960 ;
        RECT 99.330 177.615 99.580 178.425 ;
        RECT 99.750 178.115 100.065 178.675 ;
        RECT 100.235 178.205 101.885 178.725 ;
        RECT 102.055 178.375 103.745 178.895 ;
        RECT 104.835 179.015 105.125 179.815 ;
        RECT 105.295 179.185 105.530 179.985 ;
        RECT 105.715 179.645 107.250 179.815 ;
        RECT 105.715 179.015 106.045 179.645 ;
        RECT 104.835 178.845 106.045 179.015 ;
        RECT 104.835 178.345 105.080 178.675 ;
        RECT 99.760 177.435 100.065 177.945 ;
        RECT 100.235 177.435 103.745 178.205 ;
        RECT 105.250 178.175 105.420 178.845 ;
        RECT 106.215 178.675 106.450 179.420 ;
        RECT 105.590 178.345 105.990 178.675 ;
        RECT 106.160 178.345 106.450 178.675 ;
        RECT 106.640 178.675 106.910 179.420 ;
        RECT 107.080 179.015 107.250 179.645 ;
        RECT 107.420 179.185 107.825 179.985 ;
        RECT 107.080 178.845 107.825 179.015 ;
        RECT 106.640 178.345 106.980 178.675 ;
        RECT 107.150 178.345 107.485 178.675 ;
        RECT 107.655 178.345 107.825 178.845 ;
        RECT 107.995 178.420 108.345 179.815 ;
        RECT 109.435 178.820 109.725 179.985 ;
        RECT 110.815 178.845 111.085 179.815 ;
        RECT 111.295 179.185 111.575 179.985 ;
        RECT 111.745 179.475 113.400 179.765 ;
        RECT 111.810 179.135 113.400 179.305 ;
        RECT 111.810 179.015 111.980 179.135 ;
        RECT 111.255 178.845 111.980 179.015 ;
        RECT 104.835 177.605 105.420 178.175 ;
        RECT 105.670 178.005 107.065 178.175 ;
        RECT 105.670 177.660 106.000 178.005 ;
        RECT 106.215 177.435 106.590 177.835 ;
        RECT 106.770 177.660 107.065 178.005 ;
        RECT 107.235 177.435 107.905 178.175 ;
        RECT 108.075 177.605 108.345 178.420 ;
        RECT 109.435 177.435 109.725 178.160 ;
        RECT 110.815 178.110 110.985 178.845 ;
        RECT 111.255 178.675 111.425 178.845 ;
        RECT 112.170 178.795 112.885 178.965 ;
        RECT 113.080 178.845 113.400 179.135 ;
        RECT 113.575 178.845 113.845 179.815 ;
        RECT 114.055 179.185 114.335 179.985 ;
        RECT 114.505 179.475 116.160 179.765 ;
        RECT 114.570 179.135 116.160 179.305 ;
        RECT 114.570 179.015 114.740 179.135 ;
        RECT 114.015 178.845 114.740 179.015 ;
        RECT 111.155 178.345 111.425 178.675 ;
        RECT 111.595 178.345 112.000 178.675 ;
        RECT 112.170 178.345 112.880 178.795 ;
        RECT 111.255 178.175 111.425 178.345 ;
        RECT 110.815 177.765 111.085 178.110 ;
        RECT 111.255 178.005 112.865 178.175 ;
        RECT 113.050 178.105 113.400 178.675 ;
        RECT 113.575 178.110 113.745 178.845 ;
        RECT 114.015 178.675 114.185 178.845 ;
        RECT 113.915 178.345 114.185 178.675 ;
        RECT 114.355 178.345 114.760 178.675 ;
        RECT 114.930 178.345 115.640 178.965 ;
        RECT 115.840 178.845 116.160 179.135 ;
        RECT 114.015 178.175 114.185 178.345 ;
        RECT 111.275 177.435 111.655 177.835 ;
        RECT 111.825 177.655 111.995 178.005 ;
        RECT 112.165 177.435 112.495 177.835 ;
        RECT 112.695 177.655 112.865 178.005 ;
        RECT 113.065 177.435 113.395 177.935 ;
        RECT 113.575 177.765 113.845 178.110 ;
        RECT 114.015 178.005 115.625 178.175 ;
        RECT 115.810 178.105 116.160 178.675 ;
        RECT 114.035 177.435 114.415 177.835 ;
        RECT 114.585 177.655 114.755 178.005 ;
        RECT 114.925 177.435 115.255 177.835 ;
        RECT 115.455 177.655 115.625 178.005 ;
        RECT 115.825 177.435 116.155 177.935 ;
        RECT 116.345 177.615 116.605 179.805 ;
        RECT 116.775 179.255 117.115 179.985 ;
        RECT 117.295 179.075 117.565 179.805 ;
        RECT 116.795 178.855 117.565 179.075 ;
        RECT 117.745 179.095 117.975 179.805 ;
        RECT 118.145 179.275 118.475 179.985 ;
        RECT 118.645 179.095 118.905 179.805 ;
        RECT 119.295 179.645 120.905 179.815 ;
        RECT 119.295 179.145 119.545 179.645 ;
        RECT 117.745 178.855 118.905 179.095 ;
        RECT 119.715 178.975 119.965 179.475 ;
        RECT 120.135 179.305 120.905 179.645 ;
        RECT 121.075 179.485 121.380 179.985 ;
        RECT 121.550 179.305 121.800 179.815 ;
        RECT 121.970 179.485 122.220 179.985 ;
        RECT 122.390 179.475 122.705 179.815 ;
        RECT 122.910 179.645 124.000 179.815 ;
        RECT 122.910 179.485 123.160 179.645 ;
        RECT 123.750 179.485 124.000 179.645 ;
        RECT 124.170 179.485 124.420 179.985 ;
        RECT 124.590 179.485 124.870 179.815 ;
        RECT 123.755 179.475 123.925 179.485 ;
        RECT 124.675 179.475 124.845 179.485 ;
        RECT 122.390 179.305 122.600 179.475 ;
        RECT 123.330 179.305 123.580 179.475 ;
        RECT 120.135 179.135 122.600 179.305 ;
        RECT 122.770 179.135 124.870 179.305 ;
        RECT 116.795 178.185 117.085 178.855 ;
        RECT 119.095 178.765 119.965 178.975 ;
        RECT 122.770 178.965 122.940 179.135 ;
        RECT 120.205 178.795 122.940 178.965 ;
        RECT 123.110 178.795 124.285 178.965 ;
        RECT 117.265 178.365 117.730 178.675 ;
        RECT 117.910 178.365 118.435 178.675 ;
        RECT 116.795 177.985 118.025 178.185 ;
        RECT 116.865 177.435 117.535 177.805 ;
        RECT 117.715 177.615 118.025 177.985 ;
        RECT 118.205 177.725 118.435 178.365 ;
        RECT 118.615 178.345 118.915 178.675 ;
        RECT 119.095 178.255 119.505 178.765 ;
        RECT 120.205 178.595 120.375 178.795 ;
        RECT 123.110 178.625 123.280 178.795 ;
        RECT 124.115 178.625 124.285 178.795 ;
        RECT 119.715 178.425 120.375 178.595 ;
        RECT 120.900 178.425 121.570 178.625 ;
        RECT 121.760 178.425 123.280 178.625 ;
        RECT 123.450 178.425 123.945 178.625 ;
        RECT 124.115 178.425 124.445 178.625 ;
        RECT 120.535 178.255 120.705 178.285 ;
        RECT 124.700 178.255 124.870 179.135 ;
        RECT 118.615 177.435 118.905 178.165 ;
        RECT 119.095 178.075 121.365 178.255 ;
        RECT 119.675 177.995 120.005 178.075 ;
        RECT 121.035 177.995 121.365 178.075 ;
        RECT 121.590 178.075 122.680 178.255 ;
        RECT 119.335 177.435 119.505 177.905 ;
        RECT 120.175 177.435 120.345 177.905 ;
        RECT 121.590 177.825 121.840 178.075 ;
        RECT 120.610 177.605 121.840 177.825 ;
        RECT 122.010 177.435 122.180 177.905 ;
        RECT 122.350 177.605 122.680 178.075 ;
        RECT 123.290 178.075 124.870 178.255 ;
        RECT 125.075 178.910 125.345 179.815 ;
        RECT 125.515 179.225 125.845 179.985 ;
        RECT 126.025 179.055 126.205 179.815 ;
        RECT 125.075 178.110 125.255 178.910 ;
        RECT 125.530 178.885 126.205 179.055 ;
        RECT 125.530 178.740 125.700 178.885 ;
        RECT 126.465 178.845 126.795 179.985 ;
        RECT 127.325 179.015 127.655 179.800 ;
        RECT 127.840 179.185 128.095 179.985 ;
        RECT 128.295 179.135 128.625 179.815 ;
        RECT 126.975 178.845 127.655 179.015 ;
        RECT 125.425 178.410 125.700 178.740 ;
        RECT 125.530 178.155 125.700 178.410 ;
        RECT 125.925 178.335 126.265 178.705 ;
        RECT 126.455 178.425 126.805 178.675 ;
        RECT 126.975 178.245 127.145 178.845 ;
        RECT 127.315 178.425 127.665 178.675 ;
        RECT 127.840 178.645 128.085 179.005 ;
        RECT 128.275 178.855 128.625 179.135 ;
        RECT 128.275 178.475 128.445 178.855 ;
        RECT 128.805 178.675 129.000 179.725 ;
        RECT 129.180 178.845 129.500 179.985 ;
        RECT 130.595 178.910 130.865 179.815 ;
        RECT 131.035 179.225 131.365 179.985 ;
        RECT 131.545 179.055 131.725 179.815 ;
        RECT 127.925 178.305 128.445 178.475 ;
        RECT 128.615 178.345 129.000 178.675 ;
        RECT 129.180 178.625 129.440 178.675 ;
        RECT 129.180 178.455 129.445 178.625 ;
        RECT 129.180 178.345 129.440 178.455 ;
        RECT 127.925 178.285 128.095 178.305 ;
        RECT 122.950 177.435 123.120 177.905 ;
        RECT 123.290 177.605 123.620 178.075 ;
        RECT 123.790 177.435 123.960 177.905 ;
        RECT 124.130 177.605 124.460 178.075 ;
        RECT 124.630 177.435 124.800 177.905 ;
        RECT 125.075 177.605 125.335 178.110 ;
        RECT 125.530 177.985 126.195 178.155 ;
        RECT 125.515 177.435 125.845 177.815 ;
        RECT 126.025 177.605 126.195 177.985 ;
        RECT 126.465 177.435 126.735 178.245 ;
        RECT 126.905 177.605 127.235 178.245 ;
        RECT 127.405 177.435 127.645 178.245 ;
        RECT 127.895 178.115 128.095 178.285 ;
        RECT 127.925 177.740 128.095 178.115 ;
        RECT 128.285 177.965 129.500 178.135 ;
        RECT 128.285 177.660 128.515 177.965 ;
        RECT 128.685 177.435 129.015 177.795 ;
        RECT 129.210 177.615 129.500 177.965 ;
        RECT 130.595 178.110 130.775 178.910 ;
        RECT 131.050 178.885 131.725 179.055 ;
        RECT 131.975 179.115 132.250 179.815 ;
        RECT 132.420 179.440 132.675 179.985 ;
        RECT 132.845 179.475 133.325 179.815 ;
        RECT 133.500 179.430 134.105 179.985 ;
        RECT 133.490 179.330 134.105 179.430 ;
        RECT 133.490 179.305 133.675 179.330 ;
        RECT 131.050 178.740 131.220 178.885 ;
        RECT 130.945 178.410 131.220 178.740 ;
        RECT 131.050 178.155 131.220 178.410 ;
        RECT 131.445 178.335 131.785 178.705 ;
        RECT 130.595 177.605 130.855 178.110 ;
        RECT 131.050 177.985 131.715 178.155 ;
        RECT 131.035 177.435 131.365 177.815 ;
        RECT 131.545 177.605 131.715 177.985 ;
        RECT 131.975 178.085 132.145 179.115 ;
        RECT 132.420 178.985 133.175 179.235 ;
        RECT 133.345 179.060 133.675 179.305 ;
        RECT 132.420 178.950 133.190 178.985 ;
        RECT 132.420 178.940 133.205 178.950 ;
        RECT 132.315 178.925 133.210 178.940 ;
        RECT 132.315 178.910 133.230 178.925 ;
        RECT 132.315 178.900 133.250 178.910 ;
        RECT 132.315 178.890 133.275 178.900 ;
        RECT 132.315 178.860 133.345 178.890 ;
        RECT 132.315 178.830 133.365 178.860 ;
        RECT 132.315 178.800 133.385 178.830 ;
        RECT 132.315 178.775 133.415 178.800 ;
        RECT 132.315 178.740 133.450 178.775 ;
        RECT 132.315 178.735 133.480 178.740 ;
        RECT 132.315 178.340 132.545 178.735 ;
        RECT 133.090 178.730 133.480 178.735 ;
        RECT 133.115 178.720 133.480 178.730 ;
        RECT 133.130 178.715 133.480 178.720 ;
        RECT 133.145 178.710 133.480 178.715 ;
        RECT 133.845 178.710 134.105 179.160 ;
        RECT 135.195 178.820 135.485 179.985 ;
        RECT 135.655 179.475 135.915 179.985 ;
        RECT 133.145 178.705 134.105 178.710 ;
        RECT 133.155 178.695 134.105 178.705 ;
        RECT 133.165 178.690 134.105 178.695 ;
        RECT 133.175 178.680 134.105 178.690 ;
        RECT 133.180 178.670 134.105 178.680 ;
        RECT 133.185 178.665 134.105 178.670 ;
        RECT 133.195 178.650 134.105 178.665 ;
        RECT 133.200 178.635 134.105 178.650 ;
        RECT 133.210 178.610 134.105 178.635 ;
        RECT 132.715 178.140 133.045 178.565 ;
        RECT 131.975 177.605 132.235 178.085 ;
        RECT 132.405 177.435 132.655 177.975 ;
        RECT 132.825 177.655 133.045 178.140 ;
        RECT 133.215 178.540 134.105 178.610 ;
        RECT 133.215 177.815 133.385 178.540 ;
        RECT 135.655 178.425 135.995 179.305 ;
        RECT 136.165 178.595 136.335 179.815 ;
        RECT 136.575 179.480 137.190 179.985 ;
        RECT 136.575 178.945 136.825 179.310 ;
        RECT 136.995 179.305 137.190 179.480 ;
        RECT 137.360 179.475 137.835 179.815 ;
        RECT 138.005 179.440 138.220 179.985 ;
        RECT 136.995 179.115 137.325 179.305 ;
        RECT 137.545 178.945 138.260 179.240 ;
        RECT 138.430 179.115 138.705 179.815 ;
        RECT 136.575 178.775 138.365 178.945 ;
        RECT 133.555 177.985 134.105 178.370 ;
        RECT 136.165 178.345 136.960 178.595 ;
        RECT 136.165 178.255 136.415 178.345 ;
        RECT 133.215 177.645 134.105 177.815 ;
        RECT 135.195 177.435 135.485 178.160 ;
        RECT 135.655 177.435 135.915 178.255 ;
        RECT 136.085 177.835 136.415 178.255 ;
        RECT 137.130 177.920 137.385 178.775 ;
        RECT 136.595 177.655 137.385 177.920 ;
        RECT 137.555 178.075 137.965 178.595 ;
        RECT 138.135 178.345 138.365 178.775 ;
        RECT 138.535 178.085 138.705 179.115 ;
        RECT 137.555 177.655 137.755 178.075 ;
        RECT 137.945 177.435 138.275 177.895 ;
        RECT 138.445 177.605 138.705 178.085 ;
        RECT 138.875 179.115 139.150 179.815 ;
        RECT 139.320 179.440 139.575 179.985 ;
        RECT 139.745 179.475 140.225 179.815 ;
        RECT 140.400 179.430 141.005 179.985 ;
        RECT 140.390 179.330 141.005 179.430 ;
        RECT 140.390 179.305 140.575 179.330 ;
        RECT 138.875 178.085 139.045 179.115 ;
        RECT 139.320 178.985 140.075 179.235 ;
        RECT 140.245 179.060 140.575 179.305 ;
        RECT 139.320 178.950 140.090 178.985 ;
        RECT 139.320 178.940 140.105 178.950 ;
        RECT 139.215 178.925 140.110 178.940 ;
        RECT 139.215 178.910 140.130 178.925 ;
        RECT 139.215 178.900 140.150 178.910 ;
        RECT 139.215 178.890 140.175 178.900 ;
        RECT 139.215 178.860 140.245 178.890 ;
        RECT 139.215 178.830 140.265 178.860 ;
        RECT 139.215 178.800 140.285 178.830 ;
        RECT 139.215 178.775 140.315 178.800 ;
        RECT 139.215 178.740 140.350 178.775 ;
        RECT 139.215 178.735 140.380 178.740 ;
        RECT 139.215 178.340 139.445 178.735 ;
        RECT 139.990 178.730 140.380 178.735 ;
        RECT 140.015 178.720 140.380 178.730 ;
        RECT 140.030 178.715 140.380 178.720 ;
        RECT 140.045 178.710 140.380 178.715 ;
        RECT 140.745 178.710 141.005 179.160 ;
        RECT 141.360 179.015 141.750 179.190 ;
        RECT 142.235 179.185 142.565 179.985 ;
        RECT 142.735 179.195 143.270 179.815 ;
        RECT 141.360 178.845 142.785 179.015 ;
        RECT 140.045 178.705 141.005 178.710 ;
        RECT 140.055 178.695 141.005 178.705 ;
        RECT 140.065 178.690 141.005 178.695 ;
        RECT 140.075 178.680 141.005 178.690 ;
        RECT 140.080 178.670 141.005 178.680 ;
        RECT 140.085 178.665 141.005 178.670 ;
        RECT 140.095 178.650 141.005 178.665 ;
        RECT 140.100 178.635 141.005 178.650 ;
        RECT 140.110 178.610 141.005 178.635 ;
        RECT 139.615 178.140 139.945 178.565 ;
        RECT 138.875 177.605 139.135 178.085 ;
        RECT 139.305 177.435 139.555 177.975 ;
        RECT 139.725 177.655 139.945 178.140 ;
        RECT 140.115 178.540 141.005 178.610 ;
        RECT 140.115 177.815 140.285 178.540 ;
        RECT 140.455 177.985 141.005 178.370 ;
        RECT 141.235 178.115 141.590 178.675 ;
        RECT 141.760 177.945 141.930 178.845 ;
        RECT 142.100 178.115 142.365 178.675 ;
        RECT 142.615 178.345 142.785 178.845 ;
        RECT 142.955 178.175 143.270 179.195 ;
        RECT 144.485 179.315 144.655 179.815 ;
        RECT 144.825 179.485 145.155 179.985 ;
        RECT 144.485 179.145 145.150 179.315 ;
        RECT 144.400 178.325 144.750 178.975 ;
        RECT 140.115 177.645 141.005 177.815 ;
        RECT 141.340 177.435 141.580 177.945 ;
        RECT 141.760 177.615 142.040 177.945 ;
        RECT 142.270 177.435 142.485 177.945 ;
        RECT 142.655 177.605 143.270 178.175 ;
        RECT 144.920 178.155 145.150 179.145 ;
        RECT 144.485 177.985 145.150 178.155 ;
        RECT 144.485 177.695 144.655 177.985 ;
        RECT 144.825 177.435 145.155 177.815 ;
        RECT 145.325 177.695 145.510 179.815 ;
        RECT 145.750 179.525 146.015 179.985 ;
        RECT 146.185 179.390 146.435 179.815 ;
        RECT 146.645 179.540 147.750 179.710 ;
        RECT 146.130 179.260 146.435 179.390 ;
        RECT 145.680 178.065 145.960 179.015 ;
        RECT 146.130 178.155 146.300 179.260 ;
        RECT 146.470 178.475 146.710 179.070 ;
        RECT 146.880 179.005 147.410 179.370 ;
        RECT 146.880 178.305 147.050 179.005 ;
        RECT 147.580 178.925 147.750 179.540 ;
        RECT 147.920 179.185 148.090 179.985 ;
        RECT 148.260 179.485 148.510 179.815 ;
        RECT 148.735 179.515 149.620 179.685 ;
        RECT 147.580 178.835 148.090 178.925 ;
        RECT 146.130 178.025 146.355 178.155 ;
        RECT 146.525 178.085 147.050 178.305 ;
        RECT 147.220 178.665 148.090 178.835 ;
        RECT 145.765 177.435 146.015 177.895 ;
        RECT 146.185 177.885 146.355 178.025 ;
        RECT 147.220 177.885 147.390 178.665 ;
        RECT 147.920 178.595 148.090 178.665 ;
        RECT 147.600 178.415 147.800 178.445 ;
        RECT 148.260 178.415 148.430 179.485 ;
        RECT 148.600 178.595 148.790 179.315 ;
        RECT 147.600 178.115 148.430 178.415 ;
        RECT 148.960 178.385 149.280 179.345 ;
        RECT 146.185 177.715 146.520 177.885 ;
        RECT 146.715 177.715 147.390 177.885 ;
        RECT 147.710 177.435 148.080 177.935 ;
        RECT 148.260 177.885 148.430 178.115 ;
        RECT 148.815 178.055 149.280 178.385 ;
        RECT 149.450 178.675 149.620 179.515 ;
        RECT 149.800 179.485 150.115 179.985 ;
        RECT 150.345 179.255 150.685 179.815 ;
        RECT 149.790 178.880 150.685 179.255 ;
        RECT 150.855 178.975 151.025 179.985 ;
        RECT 150.495 178.675 150.685 178.880 ;
        RECT 151.195 178.925 151.525 179.770 ;
        RECT 151.195 178.845 151.585 178.925 ;
        RECT 151.755 178.895 154.345 179.985 ;
        RECT 151.370 178.795 151.585 178.845 ;
        RECT 149.450 178.345 150.325 178.675 ;
        RECT 150.495 178.345 151.245 178.675 ;
        RECT 149.450 177.885 149.620 178.345 ;
        RECT 150.495 178.175 150.695 178.345 ;
        RECT 151.415 178.215 151.585 178.795 ;
        RECT 151.360 178.175 151.585 178.215 ;
        RECT 148.260 177.715 148.665 177.885 ;
        RECT 148.835 177.715 149.620 177.885 ;
        RECT 149.895 177.435 150.105 177.965 ;
        RECT 150.365 177.650 150.695 178.175 ;
        RECT 151.205 178.090 151.585 178.175 ;
        RECT 151.755 178.205 152.965 178.725 ;
        RECT 153.135 178.375 154.345 178.895 ;
        RECT 154.975 178.895 156.185 179.985 ;
        RECT 154.975 178.355 155.495 178.895 ;
        RECT 150.865 177.435 151.035 178.045 ;
        RECT 151.205 177.655 151.535 178.090 ;
        RECT 151.755 177.435 154.345 178.205 ;
        RECT 155.665 178.185 156.185 178.725 ;
        RECT 154.975 177.435 156.185 178.185 ;
        RECT 70.710 177.265 156.270 177.435 ;
        RECT 70.795 176.515 72.005 177.265 ;
        RECT 70.795 175.975 71.315 176.515 ;
        RECT 72.175 176.495 75.685 177.265 ;
        RECT 76.315 176.805 76.875 177.095 ;
        RECT 77.045 176.805 77.295 177.265 ;
        RECT 71.485 175.805 72.005 176.345 ;
        RECT 72.175 175.975 73.825 176.495 ;
        RECT 73.995 175.805 75.685 176.325 ;
        RECT 70.795 174.715 72.005 175.805 ;
        RECT 72.175 174.715 75.685 175.805 ;
        RECT 76.315 175.435 76.565 176.805 ;
        RECT 77.915 176.635 78.245 176.995 ;
        RECT 76.855 176.445 78.245 176.635 ;
        RECT 78.620 176.735 78.910 177.085 ;
        RECT 79.105 176.905 79.435 177.265 ;
        RECT 79.605 176.735 79.835 177.040 ;
        RECT 78.620 176.565 79.835 176.735 ;
        RECT 76.855 176.355 77.025 176.445 ;
        RECT 80.025 176.395 80.195 176.960 ;
        RECT 81.005 176.715 81.175 177.005 ;
        RECT 81.345 176.885 81.675 177.265 ;
        RECT 81.005 176.545 81.670 176.715 ;
        RECT 76.735 176.025 77.025 176.355 ;
        RECT 77.195 176.025 77.535 176.275 ;
        RECT 77.755 176.025 78.430 176.275 ;
        RECT 78.680 176.245 78.940 176.355 ;
        RECT 78.675 176.075 78.940 176.245 ;
        RECT 78.680 176.025 78.940 176.075 ;
        RECT 79.120 176.025 79.505 176.355 ;
        RECT 79.675 176.225 80.195 176.395 ;
        RECT 76.855 175.775 77.025 176.025 ;
        RECT 76.855 175.605 77.795 175.775 ;
        RECT 78.165 175.665 78.430 176.025 ;
        RECT 76.315 174.885 76.775 175.435 ;
        RECT 76.965 174.715 77.295 175.435 ;
        RECT 77.495 175.055 77.795 175.605 ;
        RECT 77.965 174.715 78.245 175.385 ;
        RECT 78.620 174.715 78.940 175.855 ;
        RECT 79.120 174.975 79.315 176.025 ;
        RECT 79.675 175.845 79.845 176.225 ;
        RECT 79.495 175.565 79.845 175.845 ;
        RECT 80.035 175.695 80.280 176.055 ;
        RECT 80.920 175.725 81.270 176.375 ;
        RECT 79.495 174.885 79.825 175.565 ;
        RECT 81.440 175.555 81.670 176.545 ;
        RECT 80.025 174.715 80.280 175.515 ;
        RECT 81.005 175.385 81.670 175.555 ;
        RECT 81.005 174.885 81.175 175.385 ;
        RECT 81.345 174.715 81.675 175.215 ;
        RECT 81.845 174.885 82.030 177.005 ;
        RECT 82.285 176.805 82.535 177.265 ;
        RECT 82.705 176.815 83.040 176.985 ;
        RECT 83.235 176.815 83.910 176.985 ;
        RECT 82.705 176.675 82.875 176.815 ;
        RECT 82.200 175.685 82.480 176.635 ;
        RECT 82.650 176.545 82.875 176.675 ;
        RECT 82.650 175.440 82.820 176.545 ;
        RECT 83.045 176.395 83.570 176.615 ;
        RECT 82.990 175.630 83.230 176.225 ;
        RECT 83.400 175.695 83.570 176.395 ;
        RECT 83.740 176.035 83.910 176.815 ;
        RECT 84.230 176.765 84.600 177.265 ;
        RECT 84.780 176.815 85.185 176.985 ;
        RECT 85.355 176.815 86.140 176.985 ;
        RECT 84.780 176.585 84.950 176.815 ;
        RECT 84.120 176.285 84.950 176.585 ;
        RECT 85.335 176.315 85.800 176.645 ;
        RECT 84.120 176.255 84.320 176.285 ;
        RECT 84.440 176.035 84.610 176.105 ;
        RECT 83.740 175.865 84.610 176.035 ;
        RECT 84.100 175.775 84.610 175.865 ;
        RECT 82.650 175.310 82.955 175.440 ;
        RECT 83.400 175.330 83.930 175.695 ;
        RECT 82.270 174.715 82.535 175.175 ;
        RECT 82.705 174.885 82.955 175.310 ;
        RECT 84.100 175.160 84.270 175.775 ;
        RECT 83.165 174.990 84.270 175.160 ;
        RECT 84.440 174.715 84.610 175.515 ;
        RECT 84.780 175.215 84.950 176.285 ;
        RECT 85.120 175.385 85.310 176.105 ;
        RECT 85.480 175.355 85.800 176.315 ;
        RECT 85.970 176.355 86.140 176.815 ;
        RECT 86.415 176.735 86.625 177.265 ;
        RECT 86.885 176.525 87.215 177.050 ;
        RECT 87.385 176.655 87.555 177.265 ;
        RECT 87.725 176.610 88.055 177.045 ;
        RECT 88.360 176.765 88.855 177.095 ;
        RECT 87.725 176.525 88.105 176.610 ;
        RECT 87.015 176.355 87.215 176.525 ;
        RECT 87.880 176.485 88.105 176.525 ;
        RECT 85.970 176.025 86.845 176.355 ;
        RECT 87.015 176.025 87.765 176.355 ;
        RECT 84.780 174.885 85.030 175.215 ;
        RECT 85.970 175.185 86.140 176.025 ;
        RECT 87.015 175.820 87.205 176.025 ;
        RECT 87.935 175.905 88.105 176.485 ;
        RECT 87.890 175.855 88.105 175.905 ;
        RECT 86.310 175.445 87.205 175.820 ;
        RECT 87.715 175.775 88.105 175.855 ;
        RECT 85.255 175.015 86.140 175.185 ;
        RECT 86.320 174.715 86.635 175.215 ;
        RECT 86.865 174.885 87.205 175.445 ;
        RECT 87.375 174.715 87.545 175.725 ;
        RECT 87.715 174.930 88.045 175.775 ;
        RECT 88.275 175.275 88.515 176.585 ;
        RECT 88.685 175.855 88.855 176.765 ;
        RECT 89.075 176.025 89.425 176.990 ;
        RECT 89.605 176.025 89.905 176.995 ;
        RECT 90.085 176.025 90.365 176.995 ;
        RECT 90.545 176.465 90.815 177.265 ;
        RECT 90.985 176.545 91.325 177.055 ;
        RECT 90.560 176.025 90.890 176.275 ;
        RECT 90.560 175.855 90.875 176.025 ;
        RECT 88.685 175.685 90.875 175.855 ;
        RECT 88.280 174.715 88.615 175.095 ;
        RECT 88.785 174.885 89.035 175.685 ;
        RECT 89.255 174.715 89.585 175.435 ;
        RECT 89.770 174.885 90.020 175.685 ;
        RECT 90.485 174.715 90.815 175.515 ;
        RECT 91.065 175.145 91.325 176.545 ;
        RECT 91.495 176.525 91.770 177.265 ;
        RECT 91.990 176.695 92.180 176.855 ;
        RECT 92.525 176.705 92.695 177.095 ;
        RECT 92.900 176.865 93.230 177.095 ;
        RECT 91.990 176.525 92.300 176.695 ;
        RECT 92.525 176.525 92.765 176.705 ;
        RECT 92.130 176.355 92.300 176.525 ;
        RECT 90.985 174.885 91.325 175.145 ;
        RECT 91.495 176.005 91.945 176.355 ;
        RECT 91.495 174.905 91.765 176.005 ;
        RECT 92.130 175.815 92.425 176.355 ;
        RECT 91.935 175.645 92.425 175.815 ;
        RECT 92.595 175.895 92.765 176.525 ;
        RECT 92.980 176.615 93.150 176.865 ;
        RECT 93.405 176.795 93.575 177.265 ;
        RECT 93.745 176.615 94.075 177.080 ;
        RECT 92.980 176.445 94.075 176.615 ;
        RECT 94.345 176.715 94.515 177.095 ;
        RECT 94.695 176.885 95.025 177.265 ;
        RECT 94.345 176.545 95.010 176.715 ;
        RECT 95.205 176.590 95.465 177.095 ;
        RECT 92.935 176.065 93.435 176.275 ;
        RECT 93.605 176.065 94.085 176.275 ;
        RECT 94.275 175.995 94.615 176.365 ;
        RECT 94.840 176.290 95.010 176.545 ;
        RECT 94.840 175.960 95.115 176.290 ;
        RECT 92.595 175.725 93.205 175.895 ;
        RECT 94.840 175.815 95.010 175.960 ;
        RECT 91.935 175.140 92.210 175.645 ;
        RECT 92.380 174.715 92.710 175.475 ;
        RECT 92.880 174.885 93.205 175.725 ;
        RECT 93.680 174.715 94.055 175.815 ;
        RECT 94.335 175.645 95.010 175.815 ;
        RECT 95.285 175.790 95.465 176.590 ;
        RECT 96.555 176.540 96.845 177.265 ;
        RECT 97.105 176.715 97.275 177.095 ;
        RECT 97.455 176.885 97.785 177.265 ;
        RECT 97.105 176.545 97.770 176.715 ;
        RECT 97.965 176.590 98.225 177.095 ;
        RECT 97.035 175.995 97.375 176.365 ;
        RECT 97.600 176.290 97.770 176.545 ;
        RECT 97.600 175.960 97.875 176.290 ;
        RECT 94.335 174.885 94.515 175.645 ;
        RECT 94.695 174.715 95.025 175.475 ;
        RECT 95.195 174.885 95.465 175.790 ;
        RECT 96.555 174.715 96.845 175.880 ;
        RECT 97.600 175.815 97.770 175.960 ;
        RECT 97.095 175.645 97.770 175.815 ;
        RECT 98.045 175.790 98.225 176.590 ;
        RECT 98.395 176.495 100.985 177.265 ;
        RECT 98.395 175.975 99.605 176.495 ;
        RECT 101.655 176.445 101.885 177.265 ;
        RECT 102.055 176.465 102.385 177.095 ;
        RECT 99.775 175.805 100.985 176.325 ;
        RECT 101.635 176.025 101.965 176.275 ;
        RECT 102.135 175.865 102.385 176.465 ;
        RECT 102.555 176.445 102.765 177.265 ;
        RECT 103.095 176.615 103.425 177.095 ;
        RECT 103.595 176.805 103.925 177.265 ;
        RECT 104.140 176.615 104.470 177.095 ;
        RECT 104.670 176.805 105.000 177.265 ;
        RECT 105.225 176.615 105.395 176.935 ;
        RECT 103.095 176.445 105.395 176.615 ;
        RECT 105.565 176.635 105.895 177.080 ;
        RECT 106.165 176.805 106.335 177.265 ;
        RECT 105.565 176.445 106.315 176.635 ;
        RECT 106.625 176.465 106.965 177.095 ;
        RECT 107.135 176.465 107.445 177.265 ;
        RECT 107.650 176.465 108.345 177.095 ;
        RECT 108.515 176.495 111.105 177.265 ;
        RECT 111.275 176.590 111.545 176.935 ;
        RECT 111.735 176.865 112.115 177.265 ;
        RECT 112.285 176.695 112.455 177.045 ;
        RECT 112.625 176.865 112.955 177.265 ;
        RECT 113.155 176.695 113.325 177.045 ;
        RECT 113.525 176.765 113.855 177.265 ;
        RECT 105.945 176.275 106.315 176.445 ;
        RECT 103.055 176.025 103.565 176.275 ;
        RECT 97.095 174.885 97.275 175.645 ;
        RECT 97.455 174.715 97.785 175.475 ;
        RECT 97.955 174.885 98.225 175.790 ;
        RECT 98.395 174.715 100.985 175.805 ;
        RECT 101.655 174.715 101.885 175.855 ;
        RECT 102.055 174.885 102.385 175.865 ;
        RECT 102.555 174.715 102.765 175.855 ;
        RECT 103.115 174.715 103.445 175.835 ;
        RECT 103.775 174.960 104.145 176.275 ;
        RECT 104.315 174.960 104.645 176.275 ;
        RECT 104.855 174.960 105.185 176.275 ;
        RECT 105.355 176.065 105.775 176.275 ;
        RECT 105.945 176.065 106.525 176.275 ;
        RECT 105.945 175.895 106.205 176.065 ;
        RECT 106.695 175.895 106.965 176.465 ;
        RECT 107.145 176.025 107.480 176.295 ;
        RECT 105.455 175.605 106.205 175.895 ;
        RECT 105.455 174.885 105.705 175.605 ;
        RECT 105.875 174.715 106.205 175.435 ;
        RECT 106.440 174.885 106.965 175.895 ;
        RECT 107.650 175.865 107.820 176.465 ;
        RECT 107.990 176.025 108.325 176.275 ;
        RECT 108.515 175.975 109.725 176.495 ;
        RECT 107.135 174.715 107.415 175.855 ;
        RECT 107.585 174.885 107.915 175.865 ;
        RECT 108.085 174.715 108.345 175.855 ;
        RECT 109.895 175.805 111.105 176.325 ;
        RECT 108.515 174.715 111.105 175.805 ;
        RECT 111.275 175.855 111.445 176.590 ;
        RECT 111.715 176.525 113.325 176.695 ;
        RECT 111.715 176.355 111.885 176.525 ;
        RECT 111.615 176.025 111.885 176.355 ;
        RECT 112.055 176.025 112.460 176.355 ;
        RECT 111.715 175.855 111.885 176.025 ;
        RECT 112.630 175.905 113.340 176.355 ;
        RECT 113.510 176.025 113.860 176.595 ;
        RECT 114.040 176.590 114.315 176.935 ;
        RECT 114.505 176.865 114.885 177.265 ;
        RECT 115.055 176.695 115.225 177.045 ;
        RECT 115.395 176.865 115.725 177.265 ;
        RECT 115.895 176.695 116.150 177.045 ;
        RECT 111.275 174.885 111.545 175.855 ;
        RECT 111.715 175.685 112.440 175.855 ;
        RECT 112.630 175.735 113.345 175.905 ;
        RECT 114.040 175.855 114.210 176.590 ;
        RECT 114.485 176.525 116.150 176.695 ;
        RECT 114.485 176.355 114.655 176.525 ;
        RECT 116.335 176.495 119.845 177.265 ;
        RECT 120.015 176.805 120.575 177.095 ;
        RECT 120.745 176.805 120.995 177.265 ;
        RECT 114.380 176.025 114.655 176.355 ;
        RECT 114.825 176.025 115.650 176.355 ;
        RECT 115.820 176.025 116.165 176.355 ;
        RECT 114.485 175.855 114.655 176.025 ;
        RECT 112.270 175.565 112.440 175.685 ;
        RECT 113.540 175.565 113.860 175.855 ;
        RECT 111.755 174.715 112.035 175.515 ;
        RECT 112.270 175.395 113.860 175.565 ;
        RECT 112.205 174.935 113.860 175.225 ;
        RECT 114.040 174.885 114.315 175.855 ;
        RECT 114.485 175.685 115.145 175.855 ;
        RECT 115.455 175.735 115.650 176.025 ;
        RECT 116.335 175.975 117.985 176.495 ;
        RECT 114.975 175.565 115.145 175.685 ;
        RECT 115.820 175.565 116.145 175.855 ;
        RECT 118.155 175.805 119.845 176.325 ;
        RECT 114.525 174.715 114.805 175.515 ;
        RECT 114.975 175.395 116.145 175.565 ;
        RECT 114.975 174.935 116.165 175.225 ;
        RECT 116.335 174.715 119.845 175.805 ;
        RECT 120.015 175.435 120.265 176.805 ;
        RECT 121.615 176.635 121.945 176.995 ;
        RECT 120.555 176.445 121.945 176.635 ;
        RECT 122.315 176.540 122.605 177.265 ;
        RECT 122.775 176.515 123.985 177.265 ;
        RECT 124.175 176.875 125.350 177.095 ;
        RECT 120.555 176.355 120.725 176.445 ;
        RECT 120.435 176.025 120.725 176.355 ;
        RECT 120.895 176.025 121.235 176.275 ;
        RECT 121.455 176.025 122.130 176.275 ;
        RECT 120.555 175.775 120.725 176.025 ;
        RECT 120.555 175.605 121.495 175.775 ;
        RECT 121.865 175.665 122.130 176.025 ;
        RECT 122.775 175.975 123.295 176.515 ;
        RECT 124.155 176.455 124.930 176.705 ;
        RECT 125.100 176.625 125.350 176.875 ;
        RECT 125.520 176.795 125.690 177.265 ;
        RECT 125.860 176.625 126.190 177.095 ;
        RECT 120.015 174.885 120.475 175.435 ;
        RECT 120.665 174.715 120.995 175.435 ;
        RECT 121.195 175.055 121.495 175.605 ;
        RECT 121.665 174.715 121.945 175.385 ;
        RECT 122.315 174.715 122.605 175.880 ;
        RECT 123.465 175.805 123.985 176.345 ;
        RECT 122.775 174.715 123.985 175.805 ;
        RECT 124.155 175.565 124.385 176.455 ;
        RECT 125.100 176.445 126.190 176.625 ;
        RECT 126.500 176.445 126.670 177.265 ;
        RECT 126.840 176.625 127.170 177.095 ;
        RECT 127.340 176.795 127.510 177.265 ;
        RECT 127.680 176.625 128.045 177.095 ;
        RECT 128.215 176.795 128.385 177.265 ;
        RECT 128.655 176.875 129.965 177.045 ;
        RECT 129.075 176.625 129.405 176.705 ;
        RECT 126.840 176.445 129.405 176.625 ;
        RECT 124.555 176.065 125.030 176.275 ;
        RECT 125.325 176.075 126.775 176.275 ;
        RECT 124.860 175.905 125.030 176.065 ;
        RECT 127.000 176.065 128.025 176.275 ;
        RECT 128.705 176.105 129.365 176.275 ;
        RECT 127.000 175.905 127.170 176.065 ;
        RECT 124.860 175.735 127.170 175.905 ;
        RECT 128.705 175.895 128.875 176.105 ;
        RECT 129.575 175.935 129.965 176.875 ;
        RECT 130.135 176.755 130.440 177.265 ;
        RECT 130.135 176.025 130.450 176.585 ;
        RECT 130.620 176.275 130.870 177.085 ;
        RECT 131.040 176.740 131.300 177.265 ;
        RECT 131.480 176.275 131.730 177.085 ;
        RECT 131.900 176.705 132.160 177.265 ;
        RECT 132.330 176.615 132.590 177.070 ;
        RECT 132.760 176.785 133.020 177.265 ;
        RECT 133.190 176.615 133.450 177.070 ;
        RECT 133.620 176.785 133.880 177.265 ;
        RECT 134.050 176.615 134.310 177.070 ;
        RECT 134.480 176.785 134.725 177.265 ;
        RECT 134.895 176.615 135.170 177.070 ;
        RECT 135.340 176.785 135.585 177.265 ;
        RECT 135.755 176.615 136.015 177.070 ;
        RECT 136.195 176.785 136.445 177.265 ;
        RECT 136.615 176.615 136.875 177.070 ;
        RECT 137.055 176.785 137.305 177.265 ;
        RECT 137.475 176.615 137.735 177.070 ;
        RECT 137.915 176.785 138.175 177.265 ;
        RECT 138.345 176.615 138.605 177.070 ;
        RECT 138.775 176.785 139.075 177.265 ;
        RECT 132.330 176.445 139.075 176.615 ;
        RECT 130.620 176.025 137.740 176.275 ;
        RECT 137.910 176.245 139.075 176.445 ;
        RECT 139.335 176.495 141.005 177.265 ;
        RECT 141.635 176.525 141.895 177.095 ;
        RECT 142.065 176.865 142.450 177.265 ;
        RECT 142.620 176.695 142.875 177.095 ;
        RECT 142.065 176.525 142.875 176.695 ;
        RECT 143.065 176.525 143.310 177.095 ;
        RECT 143.480 176.865 143.865 177.265 ;
        RECT 144.035 176.695 144.290 177.095 ;
        RECT 143.480 176.525 144.290 176.695 ;
        RECT 144.480 176.525 144.905 177.095 ;
        RECT 145.075 176.865 145.460 177.265 ;
        RECT 145.630 176.695 146.065 177.095 ;
        RECT 146.325 176.925 146.495 176.960 ;
        RECT 146.295 176.755 146.495 176.925 ;
        RECT 145.075 176.525 146.065 176.695 ;
        RECT 137.910 176.075 139.105 176.245 ;
        RECT 127.380 175.725 128.875 175.895 ;
        RECT 129.115 175.725 129.965 175.935 ;
        RECT 127.380 175.565 127.550 175.725 ;
        RECT 124.155 175.395 127.550 175.565 ;
        RECT 129.115 175.555 129.365 175.725 ;
        RECT 124.155 175.385 126.150 175.395 ;
        RECT 124.155 174.885 124.470 175.385 ;
        RECT 124.640 174.715 124.890 175.215 ;
        RECT 125.060 174.885 125.310 175.385 ;
        RECT 125.480 174.715 125.730 175.215 ;
        RECT 125.900 174.885 126.150 175.385 ;
        RECT 127.795 175.385 129.365 175.555 ;
        RECT 127.795 175.225 128.005 175.385 ;
        RECT 129.115 175.225 129.365 175.385 ;
        RECT 126.460 174.885 126.710 175.225 ;
        RECT 126.880 174.715 127.130 175.215 ;
        RECT 127.300 175.055 127.625 175.225 ;
        RECT 128.175 175.055 128.425 175.215 ;
        RECT 127.300 174.885 128.425 175.055 ;
        RECT 128.695 174.715 128.945 175.215 ;
        RECT 129.535 174.715 129.965 175.555 ;
        RECT 130.145 174.715 130.440 175.525 ;
        RECT 130.620 174.885 130.865 176.025 ;
        RECT 131.040 174.715 131.300 175.525 ;
        RECT 131.480 174.890 131.730 176.025 ;
        RECT 137.910 175.855 139.075 176.075 ;
        RECT 139.335 175.975 140.085 176.495 ;
        RECT 132.330 175.630 139.075 175.855 ;
        RECT 140.255 175.805 141.005 176.325 ;
        RECT 132.330 175.615 137.735 175.630 ;
        RECT 131.900 174.720 132.160 175.515 ;
        RECT 132.330 174.890 132.590 175.615 ;
        RECT 132.760 174.720 133.020 175.445 ;
        RECT 133.190 174.890 133.450 175.615 ;
        RECT 133.620 174.720 133.880 175.445 ;
        RECT 134.050 174.890 134.310 175.615 ;
        RECT 134.480 174.720 134.740 175.445 ;
        RECT 134.910 174.890 135.170 175.615 ;
        RECT 135.340 174.720 135.585 175.445 ;
        RECT 135.755 174.890 136.015 175.615 ;
        RECT 136.200 174.720 136.445 175.445 ;
        RECT 136.615 174.890 136.875 175.615 ;
        RECT 137.060 174.720 137.305 175.445 ;
        RECT 137.475 174.890 137.735 175.615 ;
        RECT 137.920 174.720 138.175 175.445 ;
        RECT 138.345 174.890 138.635 175.630 ;
        RECT 131.900 174.715 138.175 174.720 ;
        RECT 138.805 174.715 139.075 175.460 ;
        RECT 139.335 174.715 141.005 175.805 ;
        RECT 141.635 175.855 141.820 176.525 ;
        RECT 142.065 176.355 142.415 176.525 ;
        RECT 143.065 176.355 143.235 176.525 ;
        RECT 143.480 176.355 143.830 176.525 ;
        RECT 144.480 176.355 144.830 176.525 ;
        RECT 145.075 176.355 145.410 176.525 ;
        RECT 146.325 176.395 146.495 176.755 ;
        RECT 146.685 176.735 146.915 177.040 ;
        RECT 147.085 176.905 147.415 177.265 ;
        RECT 147.610 176.735 147.900 177.085 ;
        RECT 146.685 176.565 147.900 176.735 ;
        RECT 148.075 176.540 148.365 177.265 ;
        RECT 148.535 176.590 148.795 177.095 ;
        RECT 148.975 176.885 149.305 177.265 ;
        RECT 149.485 176.715 149.655 177.095 ;
        RECT 141.990 176.025 142.415 176.355 ;
        RECT 141.635 174.885 141.895 175.855 ;
        RECT 142.065 175.505 142.415 176.025 ;
        RECT 142.585 175.855 143.235 176.355 ;
        RECT 143.405 176.025 143.830 176.355 ;
        RECT 142.585 175.675 143.310 175.855 ;
        RECT 142.065 175.310 142.875 175.505 ;
        RECT 142.065 174.715 142.450 175.140 ;
        RECT 142.620 174.885 142.875 175.310 ;
        RECT 143.065 174.885 143.310 175.675 ;
        RECT 143.480 175.505 143.830 176.025 ;
        RECT 144.000 175.855 144.830 176.355 ;
        RECT 145.000 176.025 145.410 176.355 ;
        RECT 144.000 175.675 144.905 175.855 ;
        RECT 143.480 175.310 144.310 175.505 ;
        RECT 143.480 174.715 143.865 175.140 ;
        RECT 144.035 174.885 144.310 175.310 ;
        RECT 144.480 174.885 144.905 175.675 ;
        RECT 145.075 175.480 145.410 176.025 ;
        RECT 145.580 175.650 146.065 176.355 ;
        RECT 146.325 176.225 146.845 176.395 ;
        RECT 146.240 175.695 146.485 176.055 ;
        RECT 146.675 175.845 146.845 176.225 ;
        RECT 147.015 176.025 147.400 176.355 ;
        RECT 147.580 176.245 147.840 176.355 ;
        RECT 147.580 176.075 147.845 176.245 ;
        RECT 147.580 176.025 147.840 176.075 ;
        RECT 146.675 175.565 147.025 175.845 ;
        RECT 145.075 175.310 146.065 175.480 ;
        RECT 145.075 174.715 145.460 175.140 ;
        RECT 145.630 174.885 146.065 175.310 ;
        RECT 146.240 174.715 146.495 175.515 ;
        RECT 146.695 174.885 147.025 175.565 ;
        RECT 147.205 174.975 147.400 176.025 ;
        RECT 147.580 174.715 147.900 175.855 ;
        RECT 148.075 174.715 148.365 175.880 ;
        RECT 148.535 175.790 148.705 176.590 ;
        RECT 148.990 176.545 149.655 176.715 ;
        RECT 148.990 176.290 149.160 176.545 ;
        RECT 150.395 176.535 150.685 177.265 ;
        RECT 148.875 175.960 149.160 176.290 ;
        RECT 149.395 175.995 149.725 176.365 ;
        RECT 150.385 176.025 150.685 176.355 ;
        RECT 150.865 176.335 151.095 176.975 ;
        RECT 151.275 176.715 151.585 177.085 ;
        RECT 151.765 176.895 152.435 177.265 ;
        RECT 151.275 176.515 152.505 176.715 ;
        RECT 150.865 176.025 151.390 176.335 ;
        RECT 151.570 176.025 152.035 176.335 ;
        RECT 148.990 175.815 149.160 175.960 ;
        RECT 152.215 175.845 152.505 176.515 ;
        RECT 148.535 174.885 148.805 175.790 ;
        RECT 148.990 175.645 149.655 175.815 ;
        RECT 148.975 174.715 149.305 175.475 ;
        RECT 149.485 174.885 149.655 175.645 ;
        RECT 150.395 175.605 151.555 175.845 ;
        RECT 150.395 174.895 150.655 175.605 ;
        RECT 150.825 174.715 151.155 175.425 ;
        RECT 151.325 174.895 151.555 175.605 ;
        RECT 151.735 175.625 152.505 175.845 ;
        RECT 151.735 174.895 152.005 175.625 ;
        RECT 152.185 174.715 152.525 175.445 ;
        RECT 152.695 174.895 152.955 177.085 ;
        RECT 153.135 176.495 154.805 177.265 ;
        RECT 154.975 176.515 156.185 177.265 ;
        RECT 153.135 175.975 153.885 176.495 ;
        RECT 154.055 175.805 154.805 176.325 ;
        RECT 153.135 174.715 154.805 175.805 ;
        RECT 154.975 175.805 155.495 176.345 ;
        RECT 155.665 175.975 156.185 176.515 ;
        RECT 154.975 174.715 156.185 175.805 ;
        RECT 70.710 174.545 156.270 174.715 ;
        RECT 70.795 173.455 72.005 174.545 ;
        RECT 72.175 173.455 74.765 174.545 ;
        RECT 70.795 172.745 71.315 173.285 ;
        RECT 71.485 172.915 72.005 173.455 ;
        RECT 72.175 172.765 73.385 173.285 ;
        RECT 73.555 172.935 74.765 173.455 ;
        RECT 75.405 173.575 75.735 174.360 ;
        RECT 75.405 173.405 76.085 173.575 ;
        RECT 76.265 173.405 76.595 174.545 ;
        RECT 76.775 174.110 82.120 174.545 ;
        RECT 75.395 172.985 75.745 173.235 ;
        RECT 75.915 172.805 76.085 173.405 ;
        RECT 76.255 172.985 76.605 173.235 ;
        RECT 70.795 171.995 72.005 172.745 ;
        RECT 72.175 171.995 74.765 172.765 ;
        RECT 75.415 171.995 75.655 172.805 ;
        RECT 75.825 172.165 76.155 172.805 ;
        RECT 76.325 171.995 76.595 172.805 ;
        RECT 78.360 172.540 78.700 173.370 ;
        RECT 80.180 172.860 80.530 174.110 ;
        RECT 82.295 173.455 83.505 174.545 ;
        RECT 82.295 172.745 82.815 173.285 ;
        RECT 82.985 172.915 83.505 173.455 ;
        RECT 83.675 173.380 83.965 174.545 ;
        RECT 84.135 173.455 85.345 174.545 ;
        RECT 84.135 172.745 84.655 173.285 ;
        RECT 84.825 172.915 85.345 173.455 ;
        RECT 85.515 173.405 85.775 174.375 ;
        RECT 85.945 174.120 86.330 174.545 ;
        RECT 86.500 173.950 86.755 174.375 ;
        RECT 85.945 173.755 86.755 173.950 ;
        RECT 76.775 171.995 82.120 172.540 ;
        RECT 82.295 171.995 83.505 172.745 ;
        RECT 83.675 171.995 83.965 172.720 ;
        RECT 84.135 171.995 85.345 172.745 ;
        RECT 85.515 172.735 85.700 173.405 ;
        RECT 85.945 173.235 86.295 173.755 ;
        RECT 86.945 173.585 87.190 174.375 ;
        RECT 87.360 174.120 87.745 174.545 ;
        RECT 87.915 173.950 88.190 174.375 ;
        RECT 85.870 172.905 86.295 173.235 ;
        RECT 86.465 173.405 87.190 173.585 ;
        RECT 87.360 173.755 88.190 173.950 ;
        RECT 86.465 172.905 87.115 173.405 ;
        RECT 87.360 173.235 87.710 173.755 ;
        RECT 88.360 173.585 88.785 174.375 ;
        RECT 88.955 174.120 89.340 174.545 ;
        RECT 89.510 173.950 89.945 174.375 ;
        RECT 87.285 172.905 87.710 173.235 ;
        RECT 87.880 173.405 88.785 173.585 ;
        RECT 88.955 173.780 89.945 173.950 ;
        RECT 87.880 172.905 88.710 173.405 ;
        RECT 88.955 173.235 89.290 173.780 ;
        RECT 88.880 172.905 89.290 173.235 ;
        RECT 89.460 172.905 89.945 173.610 ;
        RECT 90.575 173.405 90.850 174.375 ;
        RECT 91.060 173.745 91.340 174.545 ;
        RECT 91.510 174.205 93.560 174.325 ;
        RECT 91.510 174.035 93.565 174.205 ;
        RECT 91.510 173.695 93.140 173.865 ;
        RECT 91.510 173.575 91.680 173.695 ;
        RECT 91.020 173.405 91.680 173.575 ;
        RECT 85.945 172.735 86.295 172.905 ;
        RECT 86.945 172.735 87.115 172.905 ;
        RECT 87.360 172.735 87.710 172.905 ;
        RECT 88.360 172.735 88.710 172.905 ;
        RECT 88.955 172.735 89.290 172.905 ;
        RECT 85.515 172.165 85.775 172.735 ;
        RECT 85.945 172.565 86.755 172.735 ;
        RECT 85.945 171.995 86.330 172.395 ;
        RECT 86.500 172.165 86.755 172.565 ;
        RECT 86.945 172.165 87.190 172.735 ;
        RECT 87.360 172.565 88.170 172.735 ;
        RECT 87.360 171.995 87.745 172.395 ;
        RECT 87.915 172.165 88.170 172.565 ;
        RECT 88.360 172.165 88.785 172.735 ;
        RECT 88.955 172.565 89.945 172.735 ;
        RECT 88.955 171.995 89.340 172.395 ;
        RECT 89.510 172.165 89.945 172.565 ;
        RECT 90.575 172.670 90.745 173.405 ;
        RECT 91.020 173.235 91.190 173.405 ;
        RECT 90.915 172.905 91.190 173.235 ;
        RECT 91.360 172.905 91.740 173.235 ;
        RECT 91.910 172.905 92.650 173.525 ;
        RECT 92.820 173.405 93.140 173.695 ;
        RECT 93.335 173.235 93.575 173.830 ;
        RECT 93.745 173.470 94.085 174.545 ;
        RECT 95.180 174.165 95.515 174.545 ;
        RECT 92.920 172.905 93.575 173.235 ;
        RECT 91.020 172.735 91.190 172.905 ;
        RECT 90.575 172.325 90.850 172.670 ;
        RECT 91.020 172.565 92.605 172.735 ;
        RECT 91.040 171.995 91.420 172.395 ;
        RECT 91.590 172.215 91.760 172.565 ;
        RECT 91.930 171.995 92.260 172.395 ;
        RECT 92.435 172.215 92.605 172.565 ;
        RECT 92.805 171.995 93.135 172.495 ;
        RECT 93.330 172.215 93.575 172.905 ;
        RECT 93.745 172.665 94.085 173.235 ;
        RECT 95.175 172.675 95.415 173.985 ;
        RECT 95.685 173.575 95.935 174.375 ;
        RECT 96.155 173.825 96.485 174.545 ;
        RECT 96.670 173.575 96.920 174.375 ;
        RECT 97.385 173.745 97.715 174.545 ;
        RECT 97.885 174.115 98.225 174.375 ;
        RECT 95.585 173.405 97.775 173.575 ;
        RECT 95.585 172.495 95.755 173.405 ;
        RECT 97.460 173.235 97.775 173.405 ;
        RECT 93.745 171.995 94.085 172.495 ;
        RECT 95.260 172.165 95.755 172.495 ;
        RECT 95.975 172.270 96.325 173.235 ;
        RECT 96.505 172.265 96.805 173.235 ;
        RECT 96.985 172.265 97.265 173.235 ;
        RECT 97.460 172.985 97.790 173.235 ;
        RECT 97.445 171.995 97.715 172.795 ;
        RECT 97.965 172.715 98.225 174.115 ;
        RECT 97.885 172.205 98.225 172.715 ;
        RECT 98.400 173.825 98.735 174.335 ;
        RECT 98.400 172.470 98.655 173.825 ;
        RECT 98.985 173.745 99.315 174.545 ;
        RECT 99.560 173.955 99.845 174.375 ;
        RECT 100.100 174.125 100.430 174.545 ;
        RECT 100.655 174.205 101.815 174.375 ;
        RECT 100.655 173.955 100.985 174.205 ;
        RECT 99.560 173.785 100.985 173.955 ;
        RECT 101.215 173.575 101.385 174.035 ;
        RECT 101.645 173.705 101.815 174.205 ;
        RECT 99.015 173.405 101.385 173.575 ;
        RECT 102.995 173.695 103.255 174.375 ;
        RECT 103.425 173.765 103.675 174.545 ;
        RECT 103.925 173.995 104.175 174.375 ;
        RECT 104.345 174.165 104.700 174.545 ;
        RECT 105.705 174.155 106.040 174.375 ;
        RECT 105.305 173.995 105.535 174.035 ;
        RECT 103.925 173.795 105.535 173.995 ;
        RECT 103.925 173.785 104.760 173.795 ;
        RECT 105.350 173.705 105.535 173.795 ;
        RECT 99.015 173.235 99.185 173.405 ;
        RECT 101.635 173.355 101.845 173.525 ;
        RECT 101.635 173.235 101.840 173.355 ;
        RECT 98.880 172.905 99.185 173.235 ;
        RECT 99.380 173.185 99.630 173.235 ;
        RECT 99.375 173.015 99.630 173.185 ;
        RECT 99.380 172.905 99.630 173.015 ;
        RECT 99.015 172.735 99.185 172.905 ;
        RECT 99.840 172.845 100.110 173.235 ;
        RECT 100.300 172.845 100.590 173.235 ;
        RECT 99.015 172.565 99.575 172.735 ;
        RECT 99.835 172.675 100.110 172.845 ;
        RECT 100.295 172.675 100.590 172.845 ;
        RECT 99.840 172.575 100.110 172.675 ;
        RECT 100.300 172.575 100.590 172.675 ;
        RECT 100.760 172.570 101.180 173.235 ;
        RECT 101.490 172.905 101.840 173.235 ;
        RECT 98.400 172.210 98.735 172.470 ;
        RECT 99.405 172.395 99.575 172.565 ;
        RECT 98.905 171.995 99.235 172.395 ;
        RECT 99.405 172.225 101.020 172.395 ;
        RECT 101.565 171.995 101.895 172.715 ;
        RECT 102.995 172.495 103.165 173.695 ;
        RECT 104.865 173.595 105.195 173.625 ;
        RECT 103.395 173.535 105.195 173.595 ;
        RECT 105.785 173.535 106.040 174.155 ;
        RECT 103.335 173.425 106.040 173.535 ;
        RECT 106.295 173.615 106.475 174.375 ;
        RECT 106.655 173.785 106.985 174.545 ;
        RECT 106.295 173.445 106.970 173.615 ;
        RECT 107.155 173.470 107.425 174.375 ;
        RECT 103.335 173.390 103.535 173.425 ;
        RECT 103.335 172.815 103.505 173.390 ;
        RECT 104.865 173.365 106.040 173.425 ;
        RECT 106.800 173.300 106.970 173.445 ;
        RECT 103.735 172.950 104.145 173.255 ;
        RECT 104.315 172.985 104.645 173.195 ;
        RECT 103.335 172.695 103.605 172.815 ;
        RECT 103.335 172.650 104.180 172.695 ;
        RECT 103.425 172.525 104.180 172.650 ;
        RECT 104.435 172.585 104.645 172.985 ;
        RECT 104.890 172.985 105.365 173.195 ;
        RECT 105.555 172.985 106.045 173.185 ;
        RECT 104.890 172.585 105.110 172.985 ;
        RECT 106.235 172.895 106.575 173.265 ;
        RECT 106.800 172.970 107.075 173.300 ;
        RECT 102.995 172.165 103.255 172.495 ;
        RECT 104.010 172.375 104.180 172.525 ;
        RECT 103.425 171.995 103.755 172.355 ;
        RECT 104.010 172.165 105.310 172.375 ;
        RECT 105.585 171.995 106.040 172.760 ;
        RECT 106.800 172.715 106.970 172.970 ;
        RECT 106.305 172.545 106.970 172.715 ;
        RECT 107.245 172.670 107.425 173.470 ;
        RECT 107.595 173.455 109.265 174.545 ;
        RECT 106.305 172.165 106.475 172.545 ;
        RECT 106.655 171.995 106.985 172.375 ;
        RECT 107.165 172.165 107.425 172.670 ;
        RECT 107.595 172.765 108.345 173.285 ;
        RECT 108.515 172.935 109.265 173.455 ;
        RECT 109.435 173.380 109.725 174.545 ;
        RECT 110.445 173.800 110.715 174.545 ;
        RECT 111.345 174.540 117.620 174.545 ;
        RECT 110.885 173.630 111.175 174.370 ;
        RECT 111.345 173.815 111.600 174.540 ;
        RECT 111.785 173.645 112.045 174.370 ;
        RECT 112.215 173.815 112.460 174.540 ;
        RECT 112.645 173.645 112.905 174.370 ;
        RECT 113.075 173.815 113.320 174.540 ;
        RECT 113.505 173.645 113.765 174.370 ;
        RECT 113.935 173.815 114.180 174.540 ;
        RECT 114.350 173.645 114.610 174.370 ;
        RECT 114.780 173.815 115.040 174.540 ;
        RECT 115.210 173.645 115.470 174.370 ;
        RECT 115.640 173.815 115.900 174.540 ;
        RECT 116.070 173.645 116.330 174.370 ;
        RECT 116.500 173.815 116.760 174.540 ;
        RECT 116.930 173.645 117.190 174.370 ;
        RECT 117.360 173.745 117.620 174.540 ;
        RECT 111.785 173.630 117.190 173.645 ;
        RECT 110.445 173.405 117.190 173.630 ;
        RECT 110.445 172.815 111.610 173.405 ;
        RECT 117.790 173.235 118.040 174.370 ;
        RECT 118.220 173.735 118.480 174.545 ;
        RECT 118.655 173.235 118.900 174.375 ;
        RECT 119.080 173.735 119.375 174.545 ;
        RECT 119.555 174.110 124.900 174.545 ;
        RECT 125.075 174.110 130.420 174.545 ;
        RECT 111.780 172.985 118.900 173.235 ;
        RECT 107.595 171.995 109.265 172.765 ;
        RECT 109.435 171.995 109.725 172.720 ;
        RECT 110.445 172.645 117.190 172.815 ;
        RECT 110.445 171.995 110.745 172.475 ;
        RECT 110.915 172.190 111.175 172.645 ;
        RECT 111.345 171.995 111.605 172.475 ;
        RECT 111.785 172.190 112.045 172.645 ;
        RECT 112.215 171.995 112.465 172.475 ;
        RECT 112.645 172.190 112.905 172.645 ;
        RECT 113.075 171.995 113.325 172.475 ;
        RECT 113.505 172.190 113.765 172.645 ;
        RECT 113.935 171.995 114.180 172.475 ;
        RECT 114.350 172.190 114.625 172.645 ;
        RECT 114.795 171.995 115.040 172.475 ;
        RECT 115.210 172.190 115.470 172.645 ;
        RECT 115.640 171.995 115.900 172.475 ;
        RECT 116.070 172.190 116.330 172.645 ;
        RECT 116.500 171.995 116.760 172.475 ;
        RECT 116.930 172.190 117.190 172.645 ;
        RECT 117.360 171.995 117.620 172.555 ;
        RECT 117.790 172.175 118.040 172.985 ;
        RECT 118.220 171.995 118.480 172.520 ;
        RECT 118.650 172.175 118.900 172.985 ;
        RECT 119.070 172.675 119.385 173.235 ;
        RECT 121.140 172.540 121.480 173.370 ;
        RECT 122.960 172.860 123.310 174.110 ;
        RECT 126.660 172.540 127.000 173.370 ;
        RECT 128.480 172.860 128.830 174.110 ;
        RECT 131.055 173.825 131.515 174.375 ;
        RECT 131.705 173.825 132.035 174.545 ;
        RECT 119.080 171.995 119.385 172.505 ;
        RECT 119.555 171.995 124.900 172.540 ;
        RECT 125.075 171.995 130.420 172.540 ;
        RECT 131.055 172.455 131.305 173.825 ;
        RECT 132.235 173.655 132.535 174.205 ;
        RECT 132.705 173.875 132.985 174.545 ;
        RECT 131.595 173.485 132.535 173.655 ;
        RECT 131.595 173.235 131.765 173.485 ;
        RECT 132.905 173.235 133.170 173.595 ;
        RECT 133.365 173.575 133.695 174.360 ;
        RECT 133.365 173.405 134.045 173.575 ;
        RECT 134.225 173.405 134.555 174.545 ;
        RECT 131.475 172.905 131.765 173.235 ;
        RECT 131.935 172.985 132.275 173.235 ;
        RECT 132.495 172.985 133.170 173.235 ;
        RECT 133.355 172.985 133.705 173.235 ;
        RECT 131.595 172.815 131.765 172.905 ;
        RECT 131.595 172.625 132.985 172.815 ;
        RECT 133.875 172.805 134.045 173.405 ;
        RECT 135.195 173.380 135.485 174.545 ;
        RECT 135.655 173.825 136.115 174.375 ;
        RECT 136.305 173.825 136.635 174.545 ;
        RECT 134.215 172.985 134.565 173.235 ;
        RECT 131.055 172.165 131.615 172.455 ;
        RECT 131.785 171.995 132.035 172.455 ;
        RECT 132.655 172.265 132.985 172.625 ;
        RECT 133.375 171.995 133.615 172.805 ;
        RECT 133.785 172.165 134.115 172.805 ;
        RECT 134.285 171.995 134.555 172.805 ;
        RECT 135.195 171.995 135.485 172.720 ;
        RECT 135.655 172.455 135.905 173.825 ;
        RECT 136.835 173.655 137.135 174.205 ;
        RECT 137.305 173.875 137.585 174.545 ;
        RECT 136.195 173.485 137.135 173.655 ;
        RECT 136.195 173.235 136.365 173.485 ;
        RECT 137.505 173.235 137.770 173.595 ;
        RECT 137.955 173.455 139.625 174.545 ;
        RECT 139.795 174.035 140.055 174.545 ;
        RECT 136.075 172.905 136.365 173.235 ;
        RECT 136.535 172.985 136.875 173.235 ;
        RECT 137.095 172.985 137.770 173.235 ;
        RECT 136.195 172.815 136.365 172.905 ;
        RECT 136.195 172.625 137.585 172.815 ;
        RECT 135.655 172.165 136.215 172.455 ;
        RECT 136.385 171.995 136.635 172.455 ;
        RECT 137.255 172.265 137.585 172.625 ;
        RECT 137.955 172.765 138.705 173.285 ;
        RECT 138.875 172.935 139.625 173.455 ;
        RECT 139.795 172.985 140.135 173.865 ;
        RECT 140.305 173.155 140.475 174.375 ;
        RECT 140.715 174.040 141.330 174.545 ;
        RECT 140.715 173.505 140.965 173.870 ;
        RECT 141.135 173.865 141.330 174.040 ;
        RECT 141.500 174.035 141.975 174.375 ;
        RECT 142.145 174.000 142.360 174.545 ;
        RECT 141.135 173.675 141.465 173.865 ;
        RECT 141.685 173.505 142.400 173.800 ;
        RECT 142.570 173.675 142.845 174.375 ;
        RECT 140.715 173.335 142.505 173.505 ;
        RECT 140.305 172.905 141.100 173.155 ;
        RECT 140.305 172.815 140.555 172.905 ;
        RECT 137.955 171.995 139.625 172.765 ;
        RECT 139.795 171.995 140.055 172.815 ;
        RECT 140.225 172.395 140.555 172.815 ;
        RECT 141.270 172.480 141.525 173.335 ;
        RECT 140.735 172.215 141.525 172.480 ;
        RECT 141.695 172.635 142.105 173.155 ;
        RECT 142.275 172.905 142.505 173.335 ;
        RECT 142.675 172.645 142.845 173.675 ;
        RECT 143.200 173.575 143.590 173.750 ;
        RECT 144.075 173.745 144.405 174.545 ;
        RECT 144.575 173.755 145.110 174.375 ;
        RECT 143.200 173.405 144.625 173.575 ;
        RECT 143.075 172.675 143.430 173.235 ;
        RECT 141.695 172.215 141.895 172.635 ;
        RECT 142.085 171.995 142.415 172.455 ;
        RECT 142.585 172.165 142.845 172.645 ;
        RECT 143.600 172.505 143.770 173.405 ;
        RECT 143.940 172.675 144.205 173.235 ;
        RECT 144.455 172.905 144.625 173.405 ;
        RECT 144.795 172.735 145.110 173.755 ;
        RECT 143.180 171.995 143.420 172.505 ;
        RECT 143.600 172.175 143.880 172.505 ;
        RECT 144.110 171.995 144.325 172.505 ;
        RECT 144.495 172.165 145.110 172.735 ;
        RECT 145.315 173.470 145.585 174.375 ;
        RECT 145.755 173.785 146.085 174.545 ;
        RECT 146.265 173.615 146.445 174.375 ;
        RECT 145.315 172.670 145.495 173.470 ;
        RECT 145.770 173.445 146.445 173.615 ;
        RECT 146.695 173.455 149.285 174.545 ;
        RECT 149.455 174.035 149.755 174.545 ;
        RECT 149.925 173.865 150.255 174.375 ;
        RECT 150.425 174.035 151.055 174.545 ;
        RECT 151.635 174.035 152.015 174.205 ;
        RECT 152.185 174.035 152.485 174.545 ;
        RECT 151.845 173.865 152.015 174.035 ;
        RECT 145.770 173.300 145.940 173.445 ;
        RECT 145.665 172.970 145.940 173.300 ;
        RECT 145.770 172.715 145.940 172.970 ;
        RECT 146.165 172.895 146.505 173.265 ;
        RECT 146.695 172.765 147.905 173.285 ;
        RECT 148.075 172.935 149.285 173.455 ;
        RECT 149.455 173.695 151.675 173.865 ;
        RECT 145.315 172.165 145.575 172.670 ;
        RECT 145.770 172.545 146.435 172.715 ;
        RECT 145.755 171.995 146.085 172.375 ;
        RECT 146.265 172.165 146.435 172.545 ;
        RECT 146.695 171.995 149.285 172.765 ;
        RECT 149.455 172.735 149.625 173.695 ;
        RECT 149.795 173.355 151.335 173.525 ;
        RECT 149.795 172.905 150.040 173.355 ;
        RECT 150.300 172.985 150.995 173.185 ;
        RECT 151.165 173.155 151.335 173.355 ;
        RECT 151.505 173.495 151.675 173.695 ;
        RECT 151.845 173.665 152.505 173.865 ;
        RECT 151.505 173.325 152.165 173.495 ;
        RECT 151.165 172.985 151.765 173.155 ;
        RECT 151.995 172.905 152.165 173.325 ;
        RECT 149.455 172.190 149.920 172.735 ;
        RECT 150.425 171.995 150.595 172.815 ;
        RECT 150.765 172.735 151.675 172.815 ;
        RECT 152.335 172.735 152.505 173.665 ;
        RECT 152.675 173.455 154.345 174.545 ;
        RECT 150.765 172.645 152.015 172.735 ;
        RECT 150.765 172.165 151.095 172.645 ;
        RECT 151.505 172.565 152.015 172.645 ;
        RECT 151.265 171.995 151.615 172.385 ;
        RECT 151.785 172.165 152.015 172.565 ;
        RECT 152.185 172.255 152.505 172.735 ;
        RECT 152.675 172.765 153.425 173.285 ;
        RECT 153.595 172.935 154.345 173.455 ;
        RECT 154.975 173.455 156.185 174.545 ;
        RECT 154.975 172.915 155.495 173.455 ;
        RECT 152.675 171.995 154.345 172.765 ;
        RECT 155.665 172.745 156.185 173.285 ;
        RECT 154.975 171.995 156.185 172.745 ;
        RECT 70.710 171.825 156.270 171.995 ;
        RECT 70.795 171.075 72.005 171.825 ;
        RECT 72.265 171.275 72.435 171.565 ;
        RECT 72.605 171.445 72.935 171.825 ;
        RECT 72.265 171.105 72.930 171.275 ;
        RECT 70.795 170.535 71.315 171.075 ;
        RECT 71.485 170.365 72.005 170.905 ;
        RECT 70.795 169.275 72.005 170.365 ;
        RECT 72.180 170.285 72.530 170.935 ;
        RECT 72.700 170.115 72.930 171.105 ;
        RECT 72.265 169.945 72.930 170.115 ;
        RECT 72.265 169.445 72.435 169.945 ;
        RECT 72.605 169.275 72.935 169.775 ;
        RECT 73.105 169.445 73.290 171.565 ;
        RECT 73.545 171.365 73.795 171.825 ;
        RECT 73.965 171.375 74.300 171.545 ;
        RECT 74.495 171.375 75.170 171.545 ;
        RECT 73.965 171.235 74.135 171.375 ;
        RECT 73.460 170.245 73.740 171.195 ;
        RECT 73.910 171.105 74.135 171.235 ;
        RECT 73.910 170.000 74.080 171.105 ;
        RECT 74.305 170.955 74.830 171.175 ;
        RECT 74.250 170.190 74.490 170.785 ;
        RECT 74.660 170.255 74.830 170.955 ;
        RECT 75.000 170.595 75.170 171.375 ;
        RECT 75.490 171.325 75.860 171.825 ;
        RECT 76.040 171.375 76.445 171.545 ;
        RECT 76.615 171.375 77.400 171.545 ;
        RECT 76.040 171.145 76.210 171.375 ;
        RECT 75.380 170.845 76.210 171.145 ;
        RECT 76.595 170.875 77.060 171.205 ;
        RECT 75.380 170.815 75.580 170.845 ;
        RECT 75.700 170.595 75.870 170.665 ;
        RECT 75.000 170.425 75.870 170.595 ;
        RECT 75.360 170.335 75.870 170.425 ;
        RECT 73.910 169.870 74.215 170.000 ;
        RECT 74.660 169.890 75.190 170.255 ;
        RECT 73.530 169.275 73.795 169.735 ;
        RECT 73.965 169.445 74.215 169.870 ;
        RECT 75.360 169.720 75.530 170.335 ;
        RECT 74.425 169.550 75.530 169.720 ;
        RECT 75.700 169.275 75.870 170.075 ;
        RECT 76.040 169.775 76.210 170.845 ;
        RECT 76.380 169.945 76.570 170.665 ;
        RECT 76.740 169.915 77.060 170.875 ;
        RECT 77.230 170.915 77.400 171.375 ;
        RECT 77.675 171.295 77.885 171.825 ;
        RECT 78.145 171.085 78.475 171.610 ;
        RECT 78.645 171.215 78.815 171.825 ;
        RECT 78.985 171.170 79.315 171.605 ;
        RECT 79.625 171.275 79.795 171.565 ;
        RECT 79.965 171.445 80.295 171.825 ;
        RECT 78.985 171.085 79.365 171.170 ;
        RECT 79.625 171.105 80.290 171.275 ;
        RECT 78.275 170.915 78.475 171.085 ;
        RECT 79.140 171.045 79.365 171.085 ;
        RECT 77.230 170.585 78.105 170.915 ;
        RECT 78.275 170.585 79.025 170.915 ;
        RECT 76.040 169.445 76.290 169.775 ;
        RECT 77.230 169.745 77.400 170.585 ;
        RECT 78.275 170.380 78.465 170.585 ;
        RECT 79.195 170.465 79.365 171.045 ;
        RECT 79.150 170.415 79.365 170.465 ;
        RECT 77.570 170.005 78.465 170.380 ;
        RECT 78.975 170.335 79.365 170.415 ;
        RECT 76.515 169.575 77.400 169.745 ;
        RECT 77.580 169.275 77.895 169.775 ;
        RECT 78.125 169.445 78.465 170.005 ;
        RECT 78.635 169.275 78.805 170.285 ;
        RECT 78.975 169.490 79.305 170.335 ;
        RECT 79.540 170.285 79.890 170.935 ;
        RECT 80.060 170.115 80.290 171.105 ;
        RECT 79.625 169.945 80.290 170.115 ;
        RECT 79.625 169.445 79.795 169.945 ;
        RECT 79.965 169.275 80.295 169.775 ;
        RECT 80.465 169.445 80.650 171.565 ;
        RECT 80.905 171.365 81.155 171.825 ;
        RECT 81.325 171.375 81.660 171.545 ;
        RECT 81.855 171.375 82.530 171.545 ;
        RECT 81.325 171.235 81.495 171.375 ;
        RECT 80.820 170.245 81.100 171.195 ;
        RECT 81.270 171.105 81.495 171.235 ;
        RECT 81.270 170.000 81.440 171.105 ;
        RECT 81.665 170.955 82.190 171.175 ;
        RECT 81.610 170.190 81.850 170.785 ;
        RECT 82.020 170.255 82.190 170.955 ;
        RECT 82.360 170.595 82.530 171.375 ;
        RECT 82.850 171.325 83.220 171.825 ;
        RECT 83.400 171.375 83.805 171.545 ;
        RECT 83.975 171.375 84.760 171.545 ;
        RECT 83.400 171.145 83.570 171.375 ;
        RECT 82.740 170.845 83.570 171.145 ;
        RECT 83.955 170.875 84.420 171.205 ;
        RECT 82.740 170.815 82.940 170.845 ;
        RECT 83.060 170.595 83.230 170.665 ;
        RECT 82.360 170.425 83.230 170.595 ;
        RECT 82.720 170.335 83.230 170.425 ;
        RECT 81.270 169.870 81.575 170.000 ;
        RECT 82.020 169.890 82.550 170.255 ;
        RECT 80.890 169.275 81.155 169.735 ;
        RECT 81.325 169.445 81.575 169.870 ;
        RECT 82.720 169.720 82.890 170.335 ;
        RECT 81.785 169.550 82.890 169.720 ;
        RECT 83.060 169.275 83.230 170.075 ;
        RECT 83.400 169.775 83.570 170.845 ;
        RECT 83.740 169.945 83.930 170.665 ;
        RECT 84.100 169.915 84.420 170.875 ;
        RECT 84.590 170.915 84.760 171.375 ;
        RECT 85.035 171.295 85.245 171.825 ;
        RECT 85.505 171.085 85.835 171.610 ;
        RECT 86.005 171.215 86.175 171.825 ;
        RECT 86.345 171.170 86.675 171.605 ;
        RECT 86.895 171.350 87.235 171.610 ;
        RECT 86.345 171.085 86.725 171.170 ;
        RECT 85.635 170.915 85.835 171.085 ;
        RECT 86.500 171.045 86.725 171.085 ;
        RECT 84.590 170.585 85.465 170.915 ;
        RECT 85.635 170.585 86.385 170.915 ;
        RECT 83.400 169.445 83.650 169.775 ;
        RECT 84.590 169.745 84.760 170.585 ;
        RECT 85.635 170.380 85.825 170.585 ;
        RECT 86.555 170.465 86.725 171.045 ;
        RECT 86.510 170.415 86.725 170.465 ;
        RECT 84.930 170.005 85.825 170.380 ;
        RECT 86.335 170.335 86.725 170.415 ;
        RECT 83.875 169.575 84.760 169.745 ;
        RECT 84.940 169.275 85.255 169.775 ;
        RECT 85.485 169.445 85.825 170.005 ;
        RECT 85.995 169.275 86.165 170.285 ;
        RECT 86.335 169.490 86.665 170.335 ;
        RECT 86.895 169.745 87.155 171.350 ;
        RECT 87.405 171.345 87.735 171.825 ;
        RECT 87.925 171.175 88.340 171.610 ;
        RECT 88.510 171.310 89.460 171.495 ;
        RECT 87.325 171.100 88.340 171.175 ;
        RECT 87.325 171.005 88.145 171.100 ;
        RECT 87.325 170.085 87.495 171.005 ;
        RECT 87.815 170.275 88.145 170.835 ;
        RECT 88.345 170.805 88.725 170.915 ;
        RECT 88.335 170.635 88.725 170.805 ;
        RECT 88.345 170.585 88.725 170.635 ;
        RECT 89.035 170.585 89.255 171.310 ;
        RECT 89.690 170.915 89.895 171.515 ;
        RECT 90.065 171.100 90.405 171.825 ;
        RECT 90.590 171.255 90.845 171.605 ;
        RECT 91.015 171.425 91.345 171.825 ;
        RECT 91.515 171.255 91.685 171.605 ;
        RECT 91.855 171.425 92.235 171.825 ;
        RECT 90.590 171.085 92.255 171.255 ;
        RECT 92.425 171.150 92.700 171.495 ;
        RECT 93.420 171.325 93.915 171.655 ;
        RECT 92.085 170.915 92.255 171.085 ;
        RECT 88.345 170.290 88.645 170.585 ;
        RECT 89.515 170.285 89.895 170.915 ;
        RECT 90.125 170.285 90.380 170.915 ;
        RECT 90.575 170.585 90.920 170.915 ;
        RECT 91.090 170.585 91.915 170.915 ;
        RECT 92.085 170.585 92.360 170.915 ;
        RECT 90.595 170.125 90.920 170.415 ;
        RECT 91.090 170.295 91.285 170.585 ;
        RECT 92.085 170.415 92.255 170.585 ;
        RECT 92.530 170.415 92.700 171.150 ;
        RECT 91.595 170.245 92.255 170.415 ;
        RECT 91.595 170.125 91.765 170.245 ;
        RECT 87.325 169.915 88.175 170.085 ;
        RECT 86.895 169.485 87.235 169.745 ;
        RECT 87.405 169.275 87.655 169.735 ;
        RECT 87.845 169.485 88.175 169.915 ;
        RECT 88.345 169.945 90.315 170.115 ;
        RECT 90.595 169.955 91.765 170.125 ;
        RECT 88.345 169.445 88.515 169.945 ;
        RECT 88.725 169.275 88.975 169.735 ;
        RECT 89.185 169.445 89.355 169.945 ;
        RECT 89.655 169.275 89.905 169.735 ;
        RECT 90.145 169.445 90.315 169.945 ;
        RECT 90.575 169.495 91.765 169.785 ;
        RECT 91.935 169.275 92.215 170.075 ;
        RECT 92.425 169.445 92.700 170.415 ;
        RECT 93.335 169.835 93.575 171.145 ;
        RECT 93.745 170.415 93.915 171.325 ;
        RECT 94.135 170.585 94.485 171.550 ;
        RECT 94.665 170.585 94.965 171.555 ;
        RECT 95.145 170.585 95.425 171.555 ;
        RECT 95.605 171.025 95.875 171.825 ;
        RECT 96.045 171.105 96.385 171.615 ;
        RECT 95.620 170.585 95.950 170.835 ;
        RECT 95.620 170.415 95.935 170.585 ;
        RECT 93.745 170.245 95.935 170.415 ;
        RECT 93.340 169.275 93.675 169.655 ;
        RECT 93.845 169.445 94.095 170.245 ;
        RECT 94.315 169.275 94.645 169.995 ;
        RECT 94.830 169.445 95.080 170.245 ;
        RECT 95.545 169.275 95.875 170.075 ;
        RECT 96.125 169.705 96.385 171.105 ;
        RECT 96.555 171.100 96.845 171.825 ;
        RECT 97.015 171.445 97.905 171.615 ;
        RECT 97.015 170.890 97.565 171.275 ;
        RECT 97.735 170.720 97.905 171.445 ;
        RECT 97.015 170.650 97.905 170.720 ;
        RECT 98.075 171.120 98.295 171.605 ;
        RECT 98.465 171.285 98.715 171.825 ;
        RECT 98.885 171.175 99.145 171.655 ;
        RECT 98.075 170.695 98.405 171.120 ;
        RECT 97.015 170.625 97.910 170.650 ;
        RECT 97.015 170.610 97.920 170.625 ;
        RECT 97.015 170.595 97.925 170.610 ;
        RECT 97.015 170.590 97.935 170.595 ;
        RECT 97.015 170.580 97.940 170.590 ;
        RECT 97.015 170.570 97.945 170.580 ;
        RECT 97.015 170.565 97.955 170.570 ;
        RECT 97.015 170.555 97.965 170.565 ;
        RECT 97.015 170.550 97.975 170.555 ;
        RECT 96.045 169.445 96.385 169.705 ;
        RECT 96.555 169.275 96.845 170.440 ;
        RECT 97.015 170.100 97.275 170.550 ;
        RECT 97.640 170.545 97.975 170.550 ;
        RECT 97.640 170.540 97.990 170.545 ;
        RECT 97.640 170.530 98.005 170.540 ;
        RECT 97.640 170.525 98.030 170.530 ;
        RECT 98.575 170.525 98.805 170.920 ;
        RECT 97.640 170.520 98.805 170.525 ;
        RECT 97.670 170.485 98.805 170.520 ;
        RECT 97.705 170.460 98.805 170.485 ;
        RECT 97.735 170.430 98.805 170.460 ;
        RECT 97.755 170.400 98.805 170.430 ;
        RECT 97.775 170.370 98.805 170.400 ;
        RECT 97.845 170.360 98.805 170.370 ;
        RECT 97.870 170.350 98.805 170.360 ;
        RECT 97.890 170.335 98.805 170.350 ;
        RECT 97.910 170.320 98.805 170.335 ;
        RECT 97.915 170.310 98.700 170.320 ;
        RECT 97.930 170.275 98.700 170.310 ;
        RECT 97.445 169.955 97.775 170.200 ;
        RECT 97.945 170.025 98.700 170.275 ;
        RECT 98.975 170.145 99.145 171.175 ;
        RECT 97.445 169.930 97.630 169.955 ;
        RECT 97.015 169.830 97.630 169.930 ;
        RECT 97.015 169.275 97.620 169.830 ;
        RECT 97.795 169.445 98.275 169.785 ;
        RECT 98.445 169.275 98.700 169.820 ;
        RECT 98.870 169.445 99.145 170.145 ;
        RECT 99.315 171.085 99.780 171.630 ;
        RECT 99.315 170.125 99.485 171.085 ;
        RECT 100.285 171.005 100.455 171.825 ;
        RECT 100.625 171.175 100.955 171.655 ;
        RECT 101.125 171.435 101.475 171.825 ;
        RECT 101.645 171.255 101.875 171.655 ;
        RECT 101.365 171.175 101.875 171.255 ;
        RECT 100.625 171.085 101.875 171.175 ;
        RECT 102.045 171.085 102.365 171.565 ;
        RECT 100.625 171.005 101.535 171.085 ;
        RECT 99.655 170.465 99.900 170.915 ;
        RECT 100.160 170.635 100.855 170.835 ;
        RECT 101.025 170.665 101.625 170.835 ;
        RECT 101.025 170.465 101.195 170.665 ;
        RECT 101.855 170.495 102.025 170.915 ;
        RECT 99.655 170.295 101.195 170.465 ;
        RECT 101.365 170.325 102.025 170.495 ;
        RECT 101.365 170.125 101.535 170.325 ;
        RECT 102.195 170.155 102.365 171.085 ;
        RECT 99.315 169.955 101.535 170.125 ;
        RECT 101.705 169.955 102.365 170.155 ;
        RECT 102.570 171.085 103.185 171.655 ;
        RECT 103.355 171.315 103.570 171.825 ;
        RECT 103.800 171.315 104.080 171.645 ;
        RECT 104.260 171.315 104.500 171.825 ;
        RECT 102.570 170.065 102.885 171.085 ;
        RECT 103.055 170.415 103.225 170.915 ;
        RECT 103.475 170.585 103.740 171.145 ;
        RECT 103.910 170.415 104.080 171.315 ;
        RECT 104.250 170.585 104.605 171.145 ;
        RECT 104.835 171.025 105.145 171.825 ;
        RECT 105.350 171.025 106.045 171.655 ;
        RECT 106.215 171.075 107.425 171.825 ;
        RECT 107.595 171.350 107.935 171.610 ;
        RECT 104.845 170.585 105.180 170.855 ;
        RECT 105.350 170.465 105.520 171.025 ;
        RECT 105.690 170.585 106.025 170.835 ;
        RECT 106.215 170.535 106.735 171.075 ;
        RECT 105.350 170.425 105.525 170.465 ;
        RECT 103.055 170.245 104.480 170.415 ;
        RECT 99.315 169.275 99.615 169.785 ;
        RECT 99.785 169.445 100.115 169.955 ;
        RECT 101.705 169.785 101.875 169.955 ;
        RECT 100.285 169.275 100.915 169.785 ;
        RECT 101.495 169.615 101.875 169.785 ;
        RECT 102.045 169.275 102.345 169.785 ;
        RECT 102.570 169.445 103.105 170.065 ;
        RECT 103.275 169.275 103.605 170.075 ;
        RECT 104.090 170.070 104.480 170.245 ;
        RECT 104.835 169.275 105.115 170.415 ;
        RECT 105.285 169.445 105.615 170.425 ;
        RECT 105.785 169.275 106.045 170.415 ;
        RECT 106.905 170.365 107.425 170.905 ;
        RECT 106.215 169.275 107.425 170.365 ;
        RECT 107.595 169.745 107.855 171.350 ;
        RECT 108.105 171.345 108.435 171.825 ;
        RECT 108.625 171.175 109.040 171.610 ;
        RECT 109.210 171.310 110.160 171.495 ;
        RECT 108.025 171.100 109.040 171.175 ;
        RECT 108.025 171.005 108.845 171.100 ;
        RECT 108.025 170.085 108.195 171.005 ;
        RECT 108.515 170.275 108.845 170.835 ;
        RECT 109.045 170.805 109.425 170.915 ;
        RECT 109.735 170.805 109.955 171.310 ;
        RECT 110.390 170.915 110.595 171.515 ;
        RECT 110.765 171.100 111.105 171.825 ;
        RECT 111.735 171.150 112.005 171.495 ;
        RECT 112.195 171.425 112.575 171.825 ;
        RECT 112.745 171.255 112.915 171.605 ;
        RECT 113.085 171.425 113.415 171.825 ;
        RECT 113.615 171.255 113.785 171.605 ;
        RECT 113.985 171.325 114.315 171.825 ;
        RECT 109.035 170.635 109.425 170.805 ;
        RECT 109.725 170.635 109.955 170.805 ;
        RECT 109.045 170.585 109.425 170.635 ;
        RECT 109.735 170.585 109.955 170.635 ;
        RECT 109.045 170.290 109.345 170.585 ;
        RECT 110.215 170.285 110.595 170.915 ;
        RECT 110.825 170.285 111.080 170.915 ;
        RECT 111.735 170.415 111.905 171.150 ;
        RECT 112.175 171.085 113.785 171.255 ;
        RECT 112.175 170.915 112.345 171.085 ;
        RECT 112.075 170.585 112.345 170.915 ;
        RECT 112.515 170.585 112.920 170.915 ;
        RECT 112.175 170.415 112.345 170.585 ;
        RECT 113.090 170.465 113.800 170.915 ;
        RECT 113.970 170.585 114.320 171.155 ;
        RECT 114.495 171.150 114.755 171.655 ;
        RECT 114.935 171.445 115.265 171.825 ;
        RECT 115.445 171.275 115.615 171.655 ;
        RECT 108.025 169.915 108.875 170.085 ;
        RECT 107.595 169.485 107.935 169.745 ;
        RECT 108.105 169.275 108.355 169.735 ;
        RECT 108.545 169.485 108.875 169.915 ;
        RECT 109.045 169.945 111.015 170.115 ;
        RECT 109.045 169.445 109.215 169.945 ;
        RECT 109.425 169.275 109.675 169.735 ;
        RECT 109.885 169.445 110.055 169.945 ;
        RECT 110.355 169.275 110.605 169.735 ;
        RECT 110.845 169.445 111.015 169.945 ;
        RECT 111.735 169.445 112.005 170.415 ;
        RECT 112.175 170.245 112.900 170.415 ;
        RECT 113.090 170.295 113.805 170.465 ;
        RECT 112.730 170.125 112.900 170.245 ;
        RECT 114.000 170.125 114.320 170.415 ;
        RECT 112.215 169.275 112.495 170.075 ;
        RECT 112.730 169.955 114.320 170.125 ;
        RECT 114.495 170.350 114.675 171.150 ;
        RECT 114.950 171.105 115.615 171.275 ;
        RECT 114.950 170.850 115.120 171.105 ;
        RECT 115.935 171.005 116.145 171.825 ;
        RECT 116.315 171.025 116.645 171.655 ;
        RECT 114.845 170.520 115.120 170.850 ;
        RECT 115.345 170.555 115.685 170.925 ;
        RECT 114.950 170.375 115.120 170.520 ;
        RECT 116.315 170.425 116.565 171.025 ;
        RECT 116.815 171.005 117.045 171.825 ;
        RECT 118.200 171.435 118.530 171.825 ;
        RECT 118.700 171.265 118.925 171.645 ;
        RECT 116.735 170.585 117.065 170.835 ;
        RECT 118.185 170.585 118.425 171.235 ;
        RECT 118.595 171.085 118.925 171.265 ;
        RECT 112.665 169.495 114.320 169.785 ;
        RECT 114.495 169.445 114.765 170.350 ;
        RECT 114.950 170.205 115.625 170.375 ;
        RECT 114.935 169.275 115.265 170.035 ;
        RECT 115.445 169.445 115.625 170.205 ;
        RECT 115.935 169.275 116.145 170.415 ;
        RECT 116.315 169.445 116.645 170.425 ;
        RECT 118.595 170.415 118.770 171.085 ;
        RECT 119.125 170.915 119.355 171.535 ;
        RECT 119.535 171.095 119.835 171.825 ;
        RECT 120.475 171.025 120.785 171.825 ;
        RECT 120.990 171.025 121.685 171.655 ;
        RECT 122.315 171.100 122.605 171.825 ;
        RECT 122.865 171.275 123.035 171.565 ;
        RECT 123.205 171.445 123.535 171.825 ;
        RECT 122.865 171.105 123.530 171.275 ;
        RECT 120.990 170.975 121.165 171.025 ;
        RECT 118.940 170.585 119.355 170.915 ;
        RECT 119.535 170.585 119.830 170.915 ;
        RECT 120.485 170.585 120.820 170.855 ;
        RECT 120.990 170.425 121.160 170.975 ;
        RECT 121.330 170.585 121.665 170.835 ;
        RECT 116.815 169.275 117.045 170.415 ;
        RECT 118.185 170.225 118.770 170.415 ;
        RECT 118.185 169.455 118.460 170.225 ;
        RECT 118.940 170.055 119.835 170.385 ;
        RECT 118.630 169.885 119.835 170.055 ;
        RECT 118.630 169.455 118.960 169.885 ;
        RECT 119.130 169.275 119.325 169.715 ;
        RECT 119.505 169.455 119.835 169.885 ;
        RECT 120.475 169.275 120.755 170.415 ;
        RECT 120.925 169.445 121.255 170.425 ;
        RECT 121.425 169.275 121.685 170.415 ;
        RECT 122.315 169.275 122.605 170.440 ;
        RECT 122.780 170.285 123.130 170.935 ;
        RECT 123.300 170.115 123.530 171.105 ;
        RECT 122.865 169.945 123.530 170.115 ;
        RECT 122.865 169.445 123.035 169.945 ;
        RECT 123.205 169.275 123.535 169.775 ;
        RECT 123.705 169.445 123.890 171.565 ;
        RECT 124.145 171.365 124.395 171.825 ;
        RECT 124.565 171.375 124.900 171.545 ;
        RECT 125.095 171.375 125.770 171.545 ;
        RECT 124.565 171.235 124.735 171.375 ;
        RECT 124.060 170.245 124.340 171.195 ;
        RECT 124.510 171.105 124.735 171.235 ;
        RECT 124.510 170.000 124.680 171.105 ;
        RECT 124.905 170.955 125.430 171.175 ;
        RECT 124.850 170.190 125.090 170.785 ;
        RECT 125.260 170.255 125.430 170.955 ;
        RECT 125.600 170.595 125.770 171.375 ;
        RECT 126.090 171.325 126.460 171.825 ;
        RECT 126.640 171.375 127.045 171.545 ;
        RECT 127.215 171.375 128.000 171.545 ;
        RECT 126.640 171.145 126.810 171.375 ;
        RECT 125.980 170.845 126.810 171.145 ;
        RECT 127.195 170.875 127.660 171.205 ;
        RECT 125.980 170.815 126.180 170.845 ;
        RECT 126.300 170.595 126.470 170.665 ;
        RECT 125.600 170.425 126.470 170.595 ;
        RECT 125.960 170.335 126.470 170.425 ;
        RECT 124.510 169.870 124.815 170.000 ;
        RECT 125.260 169.890 125.790 170.255 ;
        RECT 124.130 169.275 124.395 169.735 ;
        RECT 124.565 169.445 124.815 169.870 ;
        RECT 125.960 169.720 126.130 170.335 ;
        RECT 125.025 169.550 126.130 169.720 ;
        RECT 126.300 169.275 126.470 170.075 ;
        RECT 126.640 169.775 126.810 170.845 ;
        RECT 126.980 169.945 127.170 170.665 ;
        RECT 127.340 169.915 127.660 170.875 ;
        RECT 127.830 170.915 128.000 171.375 ;
        RECT 128.275 171.295 128.485 171.825 ;
        RECT 128.745 171.085 129.075 171.610 ;
        RECT 129.245 171.215 129.415 171.825 ;
        RECT 129.585 171.170 129.915 171.605 ;
        RECT 129.585 171.085 129.965 171.170 ;
        RECT 128.875 170.915 129.075 171.085 ;
        RECT 129.740 171.045 129.965 171.085 ;
        RECT 127.830 170.585 128.705 170.915 ;
        RECT 128.875 170.585 129.625 170.915 ;
        RECT 126.640 169.445 126.890 169.775 ;
        RECT 127.830 169.745 128.000 170.585 ;
        RECT 128.875 170.380 129.065 170.585 ;
        RECT 129.795 170.465 129.965 171.045 ;
        RECT 129.750 170.415 129.965 170.465 ;
        RECT 128.170 170.005 129.065 170.380 ;
        RECT 129.575 170.335 129.965 170.415 ;
        RECT 130.135 171.150 130.395 171.655 ;
        RECT 130.575 171.445 130.905 171.825 ;
        RECT 131.085 171.275 131.255 171.655 ;
        RECT 130.135 170.350 130.315 171.150 ;
        RECT 130.590 171.105 131.255 171.275 ;
        RECT 131.515 171.150 131.775 171.655 ;
        RECT 131.955 171.445 132.285 171.825 ;
        RECT 132.465 171.275 132.635 171.655 ;
        RECT 130.590 170.850 130.760 171.105 ;
        RECT 130.485 170.520 130.760 170.850 ;
        RECT 130.985 170.555 131.325 170.925 ;
        RECT 130.590 170.375 130.760 170.520 ;
        RECT 127.115 169.575 128.000 169.745 ;
        RECT 128.180 169.275 128.495 169.775 ;
        RECT 128.725 169.445 129.065 170.005 ;
        RECT 129.235 169.275 129.405 170.285 ;
        RECT 129.575 169.490 129.905 170.335 ;
        RECT 130.135 169.445 130.405 170.350 ;
        RECT 130.590 170.205 131.265 170.375 ;
        RECT 130.575 169.275 130.905 170.035 ;
        RECT 131.085 169.445 131.265 170.205 ;
        RECT 131.515 170.350 131.695 171.150 ;
        RECT 131.970 171.105 132.635 171.275 ;
        RECT 131.970 170.850 132.140 171.105 ;
        RECT 132.895 171.055 134.565 171.825 ;
        RECT 135.285 171.275 135.455 171.655 ;
        RECT 135.635 171.445 135.965 171.825 ;
        RECT 135.285 171.105 135.950 171.275 ;
        RECT 136.145 171.150 136.405 171.655 ;
        RECT 131.865 170.520 132.140 170.850 ;
        RECT 132.365 170.555 132.705 170.925 ;
        RECT 132.895 170.535 133.645 171.055 ;
        RECT 131.970 170.375 132.140 170.520 ;
        RECT 131.515 169.445 131.785 170.350 ;
        RECT 131.970 170.205 132.645 170.375 ;
        RECT 133.815 170.365 134.565 170.885 ;
        RECT 135.215 170.555 135.555 170.925 ;
        RECT 135.780 170.850 135.950 171.105 ;
        RECT 135.780 170.520 136.055 170.850 ;
        RECT 135.780 170.375 135.950 170.520 ;
        RECT 131.955 169.275 132.285 170.035 ;
        RECT 132.465 169.445 132.645 170.205 ;
        RECT 132.895 169.275 134.565 170.365 ;
        RECT 135.275 170.205 135.950 170.375 ;
        RECT 136.225 170.350 136.405 171.150 ;
        RECT 136.575 171.075 137.785 171.825 ;
        RECT 138.155 171.195 138.485 171.555 ;
        RECT 139.105 171.365 139.355 171.825 ;
        RECT 139.525 171.365 140.085 171.655 ;
        RECT 136.575 170.535 137.095 171.075 ;
        RECT 138.155 171.005 139.545 171.195 ;
        RECT 139.375 170.915 139.545 171.005 ;
        RECT 137.265 170.365 137.785 170.905 ;
        RECT 135.275 169.445 135.455 170.205 ;
        RECT 135.635 169.275 135.965 170.035 ;
        RECT 136.135 169.445 136.405 170.350 ;
        RECT 136.575 169.275 137.785 170.365 ;
        RECT 137.970 170.585 138.645 170.835 ;
        RECT 138.865 170.585 139.205 170.835 ;
        RECT 139.375 170.585 139.665 170.915 ;
        RECT 137.970 170.225 138.235 170.585 ;
        RECT 139.375 170.335 139.545 170.585 ;
        RECT 138.605 170.165 139.545 170.335 ;
        RECT 138.155 169.275 138.435 169.945 ;
        RECT 138.605 169.615 138.905 170.165 ;
        RECT 139.835 169.995 140.085 171.365 ;
        RECT 140.255 171.055 143.765 171.825 ;
        RECT 140.255 170.535 141.905 171.055 ;
        RECT 143.995 171.005 144.205 171.825 ;
        RECT 144.375 171.025 144.705 171.655 ;
        RECT 142.075 170.365 143.765 170.885 ;
        RECT 144.375 170.425 144.625 171.025 ;
        RECT 144.875 171.005 145.105 171.825 ;
        RECT 144.795 170.585 145.125 170.835 ;
        RECT 139.105 169.275 139.435 169.995 ;
        RECT 139.625 169.445 140.085 169.995 ;
        RECT 140.255 169.275 143.765 170.365 ;
        RECT 143.995 169.275 144.205 170.415 ;
        RECT 144.375 169.445 144.705 170.425 ;
        RECT 144.875 169.275 145.105 170.415 ;
        RECT 145.325 169.455 145.585 171.645 ;
        RECT 145.845 171.455 146.515 171.825 ;
        RECT 146.695 171.275 147.005 171.645 ;
        RECT 145.775 171.075 147.005 171.275 ;
        RECT 145.775 170.405 146.065 171.075 ;
        RECT 147.185 170.895 147.415 171.535 ;
        RECT 147.595 171.095 147.885 171.825 ;
        RECT 148.075 171.100 148.365 171.825 ;
        RECT 148.535 171.085 149.000 171.630 ;
        RECT 146.245 170.585 146.710 170.895 ;
        RECT 146.890 170.585 147.415 170.895 ;
        RECT 147.595 170.585 147.895 170.915 ;
        RECT 145.775 170.185 146.545 170.405 ;
        RECT 145.755 169.275 146.095 170.005 ;
        RECT 146.275 169.455 146.545 170.185 ;
        RECT 146.725 170.165 147.885 170.405 ;
        RECT 146.725 169.455 146.955 170.165 ;
        RECT 147.125 169.275 147.455 169.985 ;
        RECT 147.625 169.455 147.885 170.165 ;
        RECT 148.075 169.275 148.365 170.440 ;
        RECT 148.535 170.125 148.705 171.085 ;
        RECT 149.505 171.005 149.675 171.825 ;
        RECT 149.845 171.175 150.175 171.655 ;
        RECT 150.345 171.435 150.695 171.825 ;
        RECT 150.865 171.255 151.095 171.655 ;
        RECT 150.585 171.175 151.095 171.255 ;
        RECT 149.845 171.085 151.095 171.175 ;
        RECT 151.265 171.085 151.585 171.565 ;
        RECT 149.845 171.005 150.755 171.085 ;
        RECT 148.875 170.465 149.120 170.915 ;
        RECT 149.380 170.635 150.075 170.835 ;
        RECT 150.245 170.665 150.845 170.835 ;
        RECT 150.245 170.465 150.415 170.665 ;
        RECT 151.075 170.495 151.245 170.915 ;
        RECT 148.875 170.295 150.415 170.465 ;
        RECT 150.585 170.325 151.245 170.495 ;
        RECT 150.585 170.125 150.755 170.325 ;
        RECT 151.415 170.155 151.585 171.085 ;
        RECT 151.765 171.015 152.035 171.825 ;
        RECT 152.205 171.015 152.535 171.655 ;
        RECT 152.705 171.015 152.945 171.825 ;
        RECT 151.755 170.585 152.105 170.835 ;
        RECT 152.275 170.415 152.445 171.015 ;
        RECT 153.175 171.005 153.405 171.825 ;
        RECT 153.575 171.025 153.905 171.655 ;
        RECT 152.615 170.585 152.965 170.835 ;
        RECT 153.155 170.585 153.485 170.835 ;
        RECT 153.655 170.425 153.905 171.025 ;
        RECT 154.075 171.005 154.285 171.825 ;
        RECT 154.975 171.075 156.185 171.825 ;
        RECT 148.535 169.955 150.755 170.125 ;
        RECT 150.925 169.955 151.585 170.155 ;
        RECT 148.535 169.275 148.835 169.785 ;
        RECT 149.005 169.445 149.335 169.955 ;
        RECT 150.925 169.785 151.095 169.955 ;
        RECT 149.505 169.275 150.135 169.785 ;
        RECT 150.715 169.615 151.095 169.785 ;
        RECT 151.265 169.275 151.565 169.785 ;
        RECT 151.765 169.275 152.095 170.415 ;
        RECT 152.275 170.245 152.955 170.415 ;
        RECT 152.625 169.460 152.955 170.245 ;
        RECT 153.175 169.275 153.405 170.415 ;
        RECT 153.575 169.445 153.905 170.425 ;
        RECT 154.075 169.275 154.285 170.415 ;
        RECT 154.975 170.365 155.495 170.905 ;
        RECT 155.665 170.535 156.185 171.075 ;
        RECT 154.975 169.275 156.185 170.365 ;
        RECT 70.710 169.105 156.270 169.275 ;
        RECT 70.795 168.015 72.005 169.105 ;
        RECT 72.265 168.435 72.435 168.935 ;
        RECT 72.605 168.605 72.935 169.105 ;
        RECT 72.265 168.265 72.930 168.435 ;
        RECT 70.795 167.305 71.315 167.845 ;
        RECT 71.485 167.475 72.005 168.015 ;
        RECT 72.180 167.445 72.530 168.095 ;
        RECT 70.795 166.555 72.005 167.305 ;
        RECT 72.700 167.275 72.930 168.265 ;
        RECT 72.265 167.105 72.930 167.275 ;
        RECT 72.265 166.815 72.435 167.105 ;
        RECT 72.605 166.555 72.935 166.935 ;
        RECT 73.105 166.815 73.290 168.935 ;
        RECT 73.530 168.645 73.795 169.105 ;
        RECT 73.965 168.510 74.215 168.935 ;
        RECT 74.425 168.660 75.530 168.830 ;
        RECT 73.910 168.380 74.215 168.510 ;
        RECT 73.460 167.185 73.740 168.135 ;
        RECT 73.910 167.275 74.080 168.380 ;
        RECT 74.250 167.595 74.490 168.190 ;
        RECT 74.660 168.125 75.190 168.490 ;
        RECT 74.660 167.425 74.830 168.125 ;
        RECT 75.360 168.045 75.530 168.660 ;
        RECT 75.700 168.305 75.870 169.105 ;
        RECT 76.040 168.605 76.290 168.935 ;
        RECT 76.515 168.635 77.400 168.805 ;
        RECT 75.360 167.955 75.870 168.045 ;
        RECT 73.910 167.145 74.135 167.275 ;
        RECT 74.305 167.205 74.830 167.425 ;
        RECT 75.000 167.785 75.870 167.955 ;
        RECT 73.545 166.555 73.795 167.015 ;
        RECT 73.965 167.005 74.135 167.145 ;
        RECT 75.000 167.005 75.170 167.785 ;
        RECT 75.700 167.715 75.870 167.785 ;
        RECT 75.380 167.535 75.580 167.565 ;
        RECT 76.040 167.535 76.210 168.605 ;
        RECT 76.380 167.715 76.570 168.435 ;
        RECT 75.380 167.235 76.210 167.535 ;
        RECT 76.740 167.505 77.060 168.465 ;
        RECT 73.965 166.835 74.300 167.005 ;
        RECT 74.495 166.835 75.170 167.005 ;
        RECT 75.490 166.555 75.860 167.055 ;
        RECT 76.040 167.005 76.210 167.235 ;
        RECT 76.595 167.175 77.060 167.505 ;
        RECT 77.230 167.795 77.400 168.635 ;
        RECT 77.580 168.605 77.895 169.105 ;
        RECT 78.125 168.375 78.465 168.935 ;
        RECT 77.570 168.000 78.465 168.375 ;
        RECT 78.635 168.095 78.805 169.105 ;
        RECT 78.275 167.795 78.465 168.000 ;
        RECT 78.975 168.045 79.305 168.890 ;
        RECT 79.615 168.175 79.795 168.935 ;
        RECT 79.975 168.345 80.305 169.105 ;
        RECT 78.975 167.965 79.365 168.045 ;
        RECT 79.615 168.005 80.290 168.175 ;
        RECT 80.475 168.030 80.745 168.935 ;
        RECT 79.150 167.915 79.365 167.965 ;
        RECT 77.230 167.465 78.105 167.795 ;
        RECT 78.275 167.465 79.025 167.795 ;
        RECT 77.230 167.005 77.400 167.465 ;
        RECT 78.275 167.295 78.475 167.465 ;
        RECT 79.195 167.335 79.365 167.915 ;
        RECT 80.120 167.860 80.290 168.005 ;
        RECT 79.555 167.455 79.895 167.825 ;
        RECT 80.120 167.530 80.395 167.860 ;
        RECT 79.140 167.295 79.365 167.335 ;
        RECT 76.040 166.835 76.445 167.005 ;
        RECT 76.615 166.835 77.400 167.005 ;
        RECT 77.675 166.555 77.885 167.085 ;
        RECT 78.145 166.770 78.475 167.295 ;
        RECT 78.985 167.210 79.365 167.295 ;
        RECT 80.120 167.275 80.290 167.530 ;
        RECT 78.645 166.555 78.815 167.165 ;
        RECT 78.985 166.775 79.315 167.210 ;
        RECT 79.625 167.105 80.290 167.275 ;
        RECT 80.565 167.230 80.745 168.030 ;
        RECT 80.955 167.965 81.185 169.105 ;
        RECT 81.355 167.955 81.685 168.935 ;
        RECT 81.855 167.965 82.065 169.105 ;
        RECT 82.295 168.015 83.505 169.105 ;
        RECT 80.935 167.545 81.265 167.795 ;
        RECT 79.625 166.725 79.795 167.105 ;
        RECT 79.975 166.555 80.305 166.935 ;
        RECT 80.485 166.725 80.745 167.230 ;
        RECT 80.955 166.555 81.185 167.375 ;
        RECT 81.435 167.355 81.685 167.955 ;
        RECT 81.355 166.725 81.685 167.355 ;
        RECT 81.855 166.555 82.065 167.375 ;
        RECT 82.295 167.305 82.815 167.845 ;
        RECT 82.985 167.475 83.505 168.015 ;
        RECT 83.675 167.940 83.965 169.105 ;
        RECT 84.135 168.015 86.725 169.105 ;
        RECT 84.135 167.325 85.345 167.845 ;
        RECT 85.515 167.495 86.725 168.015 ;
        RECT 86.975 168.175 87.155 168.935 ;
        RECT 87.335 168.345 87.665 169.105 ;
        RECT 86.975 168.005 87.650 168.175 ;
        RECT 87.835 168.030 88.105 168.935 ;
        RECT 87.480 167.860 87.650 168.005 ;
        RECT 86.915 167.455 87.255 167.825 ;
        RECT 87.480 167.530 87.755 167.860 ;
        RECT 82.295 166.555 83.505 167.305 ;
        RECT 83.675 166.555 83.965 167.280 ;
        RECT 84.135 166.555 86.725 167.325 ;
        RECT 87.480 167.275 87.650 167.530 ;
        RECT 86.985 167.105 87.650 167.275 ;
        RECT 87.925 167.230 88.105 168.030 ;
        RECT 88.285 167.965 88.615 169.105 ;
        RECT 89.145 168.135 89.475 168.920 ;
        RECT 90.205 168.360 90.475 169.105 ;
        RECT 91.105 169.100 97.380 169.105 ;
        RECT 90.645 168.190 90.935 168.930 ;
        RECT 91.105 168.375 91.360 169.100 ;
        RECT 91.545 168.205 91.805 168.930 ;
        RECT 91.975 168.375 92.220 169.100 ;
        RECT 92.405 168.205 92.665 168.930 ;
        RECT 92.835 168.375 93.080 169.100 ;
        RECT 93.265 168.205 93.525 168.930 ;
        RECT 93.695 168.375 93.940 169.100 ;
        RECT 94.110 168.205 94.370 168.930 ;
        RECT 94.540 168.375 94.800 169.100 ;
        RECT 94.970 168.205 95.230 168.930 ;
        RECT 95.400 168.375 95.660 169.100 ;
        RECT 95.830 168.205 96.090 168.930 ;
        RECT 96.260 168.375 96.520 169.100 ;
        RECT 96.690 168.205 96.950 168.930 ;
        RECT 97.120 168.305 97.380 169.100 ;
        RECT 91.545 168.190 96.950 168.205 ;
        RECT 88.795 167.965 89.475 168.135 ;
        RECT 90.205 167.965 96.950 168.190 ;
        RECT 88.275 167.545 88.625 167.795 ;
        RECT 88.795 167.365 88.965 167.965 ;
        RECT 89.135 167.545 89.485 167.795 ;
        RECT 90.205 167.375 91.370 167.965 ;
        RECT 97.550 167.795 97.800 168.930 ;
        RECT 97.980 168.295 98.240 169.105 ;
        RECT 98.415 167.795 98.660 168.935 ;
        RECT 98.840 168.295 99.135 169.105 ;
        RECT 99.320 168.385 99.655 168.895 ;
        RECT 91.540 167.545 98.660 167.795 ;
        RECT 86.985 166.725 87.155 167.105 ;
        RECT 87.335 166.555 87.665 166.935 ;
        RECT 87.845 166.725 88.105 167.230 ;
        RECT 88.285 166.555 88.555 167.365 ;
        RECT 88.725 166.725 89.055 167.365 ;
        RECT 89.225 166.555 89.465 167.365 ;
        RECT 90.205 167.205 96.950 167.375 ;
        RECT 90.205 166.555 90.505 167.035 ;
        RECT 90.675 166.750 90.935 167.205 ;
        RECT 91.105 166.555 91.365 167.035 ;
        RECT 91.545 166.750 91.805 167.205 ;
        RECT 91.975 166.555 92.225 167.035 ;
        RECT 92.405 166.750 92.665 167.205 ;
        RECT 92.835 166.555 93.085 167.035 ;
        RECT 93.265 166.750 93.525 167.205 ;
        RECT 93.695 166.555 93.940 167.035 ;
        RECT 94.110 166.750 94.385 167.205 ;
        RECT 94.555 166.555 94.800 167.035 ;
        RECT 94.970 166.750 95.230 167.205 ;
        RECT 95.400 166.555 95.660 167.035 ;
        RECT 95.830 166.750 96.090 167.205 ;
        RECT 96.260 166.555 96.520 167.035 ;
        RECT 96.690 166.750 96.950 167.205 ;
        RECT 97.120 166.555 97.380 167.115 ;
        RECT 97.550 166.735 97.800 167.545 ;
        RECT 97.980 166.555 98.240 167.080 ;
        RECT 98.410 166.735 98.660 167.545 ;
        RECT 98.830 167.235 99.145 167.795 ;
        RECT 98.840 166.555 99.145 167.065 ;
        RECT 99.320 167.030 99.575 168.385 ;
        RECT 99.905 168.305 100.235 169.105 ;
        RECT 100.480 168.515 100.765 168.935 ;
        RECT 101.020 168.685 101.350 169.105 ;
        RECT 101.575 168.765 102.735 168.935 ;
        RECT 101.575 168.515 101.905 168.765 ;
        RECT 100.480 168.345 101.905 168.515 ;
        RECT 102.135 168.135 102.305 168.595 ;
        RECT 102.565 168.265 102.735 168.765 ;
        RECT 102.995 168.670 108.340 169.105 ;
        RECT 99.935 167.965 102.305 168.135 ;
        RECT 99.935 167.795 100.105 167.965 ;
        RECT 102.555 167.915 102.765 168.085 ;
        RECT 102.555 167.795 102.760 167.915 ;
        RECT 99.800 167.465 100.105 167.795 ;
        RECT 100.300 167.745 100.550 167.795 ;
        RECT 100.295 167.575 100.550 167.745 ;
        RECT 100.300 167.465 100.550 167.575 ;
        RECT 99.935 167.295 100.105 167.465 ;
        RECT 100.760 167.405 101.030 167.795 ;
        RECT 101.220 167.745 101.510 167.795 ;
        RECT 101.215 167.575 101.510 167.745 ;
        RECT 99.935 167.125 100.495 167.295 ;
        RECT 100.755 167.235 101.030 167.405 ;
        RECT 100.760 167.135 101.030 167.235 ;
        RECT 101.220 167.135 101.510 167.575 ;
        RECT 101.680 167.130 102.100 167.795 ;
        RECT 102.410 167.465 102.760 167.795 ;
        RECT 99.320 166.770 99.655 167.030 ;
        RECT 100.325 166.955 100.495 167.125 ;
        RECT 99.825 166.555 100.155 166.955 ;
        RECT 100.325 166.785 101.940 166.955 ;
        RECT 102.485 166.555 102.815 167.275 ;
        RECT 104.580 167.100 104.920 167.930 ;
        RECT 106.400 167.420 106.750 168.670 ;
        RECT 109.435 167.940 109.725 169.105 ;
        RECT 109.895 168.015 113.405 169.105 ;
        RECT 109.895 167.325 111.545 167.845 ;
        RECT 111.715 167.495 113.405 168.015 ;
        RECT 113.655 168.175 113.835 168.935 ;
        RECT 114.015 168.345 114.345 169.105 ;
        RECT 113.655 168.005 114.330 168.175 ;
        RECT 114.515 168.030 114.785 168.935 ;
        RECT 114.160 167.860 114.330 168.005 ;
        RECT 113.595 167.455 113.935 167.825 ;
        RECT 114.160 167.530 114.435 167.860 ;
        RECT 102.995 166.555 108.340 167.100 ;
        RECT 109.435 166.555 109.725 167.280 ;
        RECT 109.895 166.555 113.405 167.325 ;
        RECT 114.160 167.275 114.330 167.530 ;
        RECT 113.665 167.105 114.330 167.275 ;
        RECT 114.605 167.230 114.785 168.030 ;
        RECT 114.955 168.015 116.625 169.105 ;
        RECT 116.885 168.765 118.045 168.935 ;
        RECT 116.885 168.265 117.055 168.765 ;
        RECT 117.315 168.135 117.485 168.595 ;
        RECT 117.715 168.515 118.045 168.765 ;
        RECT 118.270 168.685 118.600 169.105 ;
        RECT 118.855 168.515 119.140 168.935 ;
        RECT 117.715 168.345 119.140 168.515 ;
        RECT 119.385 168.305 119.715 169.105 ;
        RECT 119.965 168.385 120.300 168.895 ;
        RECT 113.665 166.725 113.835 167.105 ;
        RECT 114.015 166.555 114.345 166.935 ;
        RECT 114.525 166.725 114.785 167.230 ;
        RECT 114.955 167.325 115.705 167.845 ;
        RECT 115.875 167.495 116.625 168.015 ;
        RECT 116.860 167.795 117.065 168.085 ;
        RECT 117.315 167.965 119.685 168.135 ;
        RECT 119.515 167.795 119.685 167.965 ;
        RECT 116.860 167.745 117.210 167.795 ;
        RECT 116.855 167.575 117.210 167.745 ;
        RECT 116.860 167.465 117.210 167.575 ;
        RECT 114.955 166.555 116.625 167.325 ;
        RECT 116.805 166.555 117.135 167.275 ;
        RECT 117.520 167.130 117.940 167.795 ;
        RECT 118.110 167.745 118.400 167.795 ;
        RECT 118.590 167.745 118.860 167.795 ;
        RECT 119.070 167.745 119.320 167.795 ;
        RECT 118.110 167.575 118.405 167.745 ;
        RECT 118.590 167.575 118.865 167.745 ;
        RECT 119.070 167.575 119.325 167.745 ;
        RECT 118.110 167.135 118.400 167.575 ;
        RECT 118.590 167.135 118.860 167.575 ;
        RECT 119.070 167.465 119.320 167.575 ;
        RECT 119.515 167.465 119.820 167.795 ;
        RECT 119.515 167.295 119.685 167.465 ;
        RECT 119.125 167.125 119.685 167.295 ;
        RECT 119.125 166.955 119.295 167.125 ;
        RECT 120.045 167.030 120.300 168.385 ;
        RECT 120.565 168.435 120.735 168.935 ;
        RECT 120.905 168.605 121.235 169.105 ;
        RECT 120.565 168.265 121.230 168.435 ;
        RECT 120.480 167.445 120.830 168.095 ;
        RECT 121.000 167.275 121.230 168.265 ;
        RECT 117.680 166.785 119.295 166.955 ;
        RECT 119.465 166.555 119.795 166.955 ;
        RECT 119.965 166.770 120.300 167.030 ;
        RECT 120.565 167.105 121.230 167.275 ;
        RECT 120.565 166.815 120.735 167.105 ;
        RECT 120.905 166.555 121.235 166.935 ;
        RECT 121.405 166.815 121.590 168.935 ;
        RECT 121.830 168.645 122.095 169.105 ;
        RECT 122.265 168.510 122.515 168.935 ;
        RECT 122.725 168.660 123.830 168.830 ;
        RECT 122.210 168.380 122.515 168.510 ;
        RECT 121.760 167.185 122.040 168.135 ;
        RECT 122.210 167.275 122.380 168.380 ;
        RECT 122.550 167.595 122.790 168.190 ;
        RECT 122.960 168.125 123.490 168.490 ;
        RECT 122.960 167.425 123.130 168.125 ;
        RECT 123.660 168.045 123.830 168.660 ;
        RECT 124.000 168.305 124.170 169.105 ;
        RECT 124.340 168.605 124.590 168.935 ;
        RECT 124.815 168.635 125.700 168.805 ;
        RECT 123.660 167.955 124.170 168.045 ;
        RECT 122.210 167.145 122.435 167.275 ;
        RECT 122.605 167.205 123.130 167.425 ;
        RECT 123.300 167.785 124.170 167.955 ;
        RECT 121.845 166.555 122.095 167.015 ;
        RECT 122.265 167.005 122.435 167.145 ;
        RECT 123.300 167.005 123.470 167.785 ;
        RECT 124.000 167.715 124.170 167.785 ;
        RECT 123.680 167.535 123.880 167.565 ;
        RECT 124.340 167.535 124.510 168.605 ;
        RECT 124.680 167.715 124.870 168.435 ;
        RECT 123.680 167.235 124.510 167.535 ;
        RECT 125.040 167.505 125.360 168.465 ;
        RECT 122.265 166.835 122.600 167.005 ;
        RECT 122.795 166.835 123.470 167.005 ;
        RECT 123.790 166.555 124.160 167.055 ;
        RECT 124.340 167.005 124.510 167.235 ;
        RECT 124.895 167.175 125.360 167.505 ;
        RECT 125.530 167.795 125.700 168.635 ;
        RECT 125.880 168.605 126.195 169.105 ;
        RECT 126.425 168.375 126.765 168.935 ;
        RECT 125.870 168.000 126.765 168.375 ;
        RECT 126.935 168.095 127.105 169.105 ;
        RECT 126.575 167.795 126.765 168.000 ;
        RECT 127.275 168.045 127.605 168.890 ;
        RECT 127.775 168.190 127.945 169.105 ;
        RECT 127.275 167.965 127.665 168.045 ;
        RECT 127.450 167.915 127.665 167.965 ;
        RECT 125.530 167.465 126.405 167.795 ;
        RECT 126.575 167.465 127.325 167.795 ;
        RECT 125.530 167.005 125.700 167.465 ;
        RECT 126.575 167.295 126.775 167.465 ;
        RECT 127.495 167.335 127.665 167.915 ;
        RECT 127.440 167.295 127.665 167.335 ;
        RECT 124.340 166.835 124.745 167.005 ;
        RECT 124.915 166.835 125.700 167.005 ;
        RECT 125.975 166.555 126.185 167.085 ;
        RECT 126.445 166.770 126.775 167.295 ;
        RECT 127.285 167.210 127.665 167.295 ;
        RECT 128.295 167.965 128.565 168.935 ;
        RECT 128.775 168.305 129.055 169.105 ;
        RECT 129.225 168.595 130.880 168.885 ;
        RECT 129.290 168.255 130.880 168.425 ;
        RECT 129.290 168.135 129.460 168.255 ;
        RECT 128.735 167.965 129.460 168.135 ;
        RECT 128.295 167.230 128.465 167.965 ;
        RECT 128.735 167.795 128.905 167.965 ;
        RECT 128.635 167.465 128.905 167.795 ;
        RECT 129.075 167.465 129.480 167.795 ;
        RECT 129.650 167.465 130.360 168.085 ;
        RECT 130.560 167.965 130.880 168.255 ;
        RECT 131.135 168.175 131.315 168.935 ;
        RECT 131.495 168.345 131.825 169.105 ;
        RECT 131.135 168.005 131.810 168.175 ;
        RECT 131.995 168.030 132.265 168.935 ;
        RECT 131.640 167.860 131.810 168.005 ;
        RECT 128.735 167.295 128.905 167.465 ;
        RECT 126.945 166.555 127.115 167.165 ;
        RECT 127.285 166.775 127.615 167.210 ;
        RECT 127.785 166.555 127.955 167.070 ;
        RECT 128.295 166.885 128.565 167.230 ;
        RECT 128.735 167.125 130.345 167.295 ;
        RECT 130.530 167.225 130.880 167.795 ;
        RECT 131.075 167.455 131.415 167.825 ;
        RECT 131.640 167.530 131.915 167.860 ;
        RECT 131.640 167.275 131.810 167.530 ;
        RECT 128.755 166.555 129.135 166.955 ;
        RECT 129.305 166.775 129.475 167.125 ;
        RECT 129.645 166.555 129.975 166.955 ;
        RECT 130.175 166.775 130.345 167.125 ;
        RECT 131.145 167.105 131.810 167.275 ;
        RECT 132.085 167.230 132.265 168.030 ;
        RECT 132.435 168.015 133.645 169.105 ;
        RECT 130.545 166.555 130.875 167.055 ;
        RECT 131.145 166.725 131.315 167.105 ;
        RECT 131.495 166.555 131.825 166.935 ;
        RECT 132.005 166.725 132.265 167.230 ;
        RECT 132.435 167.305 132.955 167.845 ;
        RECT 133.125 167.475 133.645 168.015 ;
        RECT 133.815 168.030 134.085 168.935 ;
        RECT 134.255 168.345 134.585 169.105 ;
        RECT 134.765 168.175 134.945 168.935 ;
        RECT 132.435 166.555 133.645 167.305 ;
        RECT 133.815 167.230 133.995 168.030 ;
        RECT 134.270 168.005 134.945 168.175 ;
        RECT 134.270 167.860 134.440 168.005 ;
        RECT 135.195 167.940 135.485 169.105 ;
        RECT 135.840 168.135 136.230 168.310 ;
        RECT 136.715 168.305 137.045 169.105 ;
        RECT 137.215 168.315 137.750 168.935 ;
        RECT 135.840 167.965 137.265 168.135 ;
        RECT 134.165 167.530 134.440 167.860 ;
        RECT 134.270 167.275 134.440 167.530 ;
        RECT 134.665 167.455 135.005 167.825 ;
        RECT 133.815 166.725 134.075 167.230 ;
        RECT 134.270 167.105 134.935 167.275 ;
        RECT 134.255 166.555 134.585 166.935 ;
        RECT 134.765 166.725 134.935 167.105 ;
        RECT 135.195 166.555 135.485 167.280 ;
        RECT 135.715 167.235 136.070 167.795 ;
        RECT 136.240 167.065 136.410 167.965 ;
        RECT 136.580 167.235 136.845 167.795 ;
        RECT 137.095 167.465 137.265 167.965 ;
        RECT 137.435 167.295 137.750 168.315 ;
        RECT 138.620 168.135 138.950 168.935 ;
        RECT 139.120 168.305 139.450 169.105 ;
        RECT 139.750 168.135 140.080 168.935 ;
        RECT 140.725 168.305 140.975 169.105 ;
        RECT 138.620 167.965 141.055 168.135 ;
        RECT 141.245 167.965 141.415 169.105 ;
        RECT 141.585 167.965 141.925 168.935 ;
        RECT 142.185 168.435 142.355 168.935 ;
        RECT 142.525 168.605 142.855 169.105 ;
        RECT 142.185 168.265 142.850 168.435 ;
        RECT 138.415 167.545 138.765 167.795 ;
        RECT 138.950 167.335 139.120 167.965 ;
        RECT 139.290 167.545 139.620 167.745 ;
        RECT 139.790 167.545 140.120 167.745 ;
        RECT 140.290 167.545 140.710 167.745 ;
        RECT 140.885 167.715 141.055 167.965 ;
        RECT 140.885 167.545 141.580 167.715 ;
        RECT 141.750 167.405 141.925 167.965 ;
        RECT 142.100 167.445 142.450 168.095 ;
        RECT 135.820 166.555 136.060 167.065 ;
        RECT 136.240 166.735 136.520 167.065 ;
        RECT 136.750 166.555 136.965 167.065 ;
        RECT 137.135 166.725 137.750 167.295 ;
        RECT 138.620 166.725 139.120 167.335 ;
        RECT 139.750 167.205 140.975 167.375 ;
        RECT 141.695 167.355 141.925 167.405 ;
        RECT 139.750 166.725 140.080 167.205 ;
        RECT 140.250 166.555 140.475 167.015 ;
        RECT 140.645 166.725 140.975 167.205 ;
        RECT 141.165 166.555 141.415 167.355 ;
        RECT 141.585 166.725 141.925 167.355 ;
        RECT 142.620 167.275 142.850 168.265 ;
        RECT 142.185 167.105 142.850 167.275 ;
        RECT 142.185 166.815 142.355 167.105 ;
        RECT 142.525 166.555 142.855 166.935 ;
        RECT 143.025 166.815 143.210 168.935 ;
        RECT 143.450 168.645 143.715 169.105 ;
        RECT 143.885 168.510 144.135 168.935 ;
        RECT 144.345 168.660 145.450 168.830 ;
        RECT 143.830 168.380 144.135 168.510 ;
        RECT 143.380 167.185 143.660 168.135 ;
        RECT 143.830 167.275 144.000 168.380 ;
        RECT 144.170 167.595 144.410 168.190 ;
        RECT 144.580 168.125 145.110 168.490 ;
        RECT 144.580 167.425 144.750 168.125 ;
        RECT 145.280 168.045 145.450 168.660 ;
        RECT 145.620 168.305 145.790 169.105 ;
        RECT 145.960 168.605 146.210 168.935 ;
        RECT 146.435 168.635 147.320 168.805 ;
        RECT 145.280 167.955 145.790 168.045 ;
        RECT 143.830 167.145 144.055 167.275 ;
        RECT 144.225 167.205 144.750 167.425 ;
        RECT 144.920 167.785 145.790 167.955 ;
        RECT 143.465 166.555 143.715 167.015 ;
        RECT 143.885 167.005 144.055 167.145 ;
        RECT 144.920 167.005 145.090 167.785 ;
        RECT 145.620 167.715 145.790 167.785 ;
        RECT 145.300 167.535 145.500 167.565 ;
        RECT 145.960 167.535 146.130 168.605 ;
        RECT 146.300 167.715 146.490 168.435 ;
        RECT 145.300 167.235 146.130 167.535 ;
        RECT 146.660 167.505 146.980 168.465 ;
        RECT 143.885 166.835 144.220 167.005 ;
        RECT 144.415 166.835 145.090 167.005 ;
        RECT 145.410 166.555 145.780 167.055 ;
        RECT 145.960 167.005 146.130 167.235 ;
        RECT 146.515 167.175 146.980 167.505 ;
        RECT 147.150 167.795 147.320 168.635 ;
        RECT 147.500 168.605 147.815 169.105 ;
        RECT 148.045 168.375 148.385 168.935 ;
        RECT 147.490 168.000 148.385 168.375 ;
        RECT 148.555 168.095 148.725 169.105 ;
        RECT 148.195 167.795 148.385 168.000 ;
        RECT 148.895 168.045 149.225 168.890 ;
        RECT 150.375 168.510 150.810 168.935 ;
        RECT 150.980 168.680 151.365 169.105 ;
        RECT 150.375 168.340 151.365 168.510 ;
        RECT 148.895 167.965 149.285 168.045 ;
        RECT 149.070 167.915 149.285 167.965 ;
        RECT 147.150 167.465 148.025 167.795 ;
        RECT 148.195 167.465 148.945 167.795 ;
        RECT 147.150 167.005 147.320 167.465 ;
        RECT 148.195 167.295 148.395 167.465 ;
        RECT 149.115 167.335 149.285 167.915 ;
        RECT 150.375 167.465 150.860 168.170 ;
        RECT 151.030 167.795 151.365 168.340 ;
        RECT 151.535 168.145 151.960 168.935 ;
        RECT 152.130 168.510 152.405 168.935 ;
        RECT 152.575 168.680 152.960 169.105 ;
        RECT 152.130 168.315 152.960 168.510 ;
        RECT 151.535 167.965 152.440 168.145 ;
        RECT 151.030 167.465 151.440 167.795 ;
        RECT 151.610 167.465 152.440 167.965 ;
        RECT 152.610 167.795 152.960 168.315 ;
        RECT 153.130 168.145 153.375 168.935 ;
        RECT 153.565 168.510 153.820 168.935 ;
        RECT 153.990 168.680 154.375 169.105 ;
        RECT 153.565 168.315 154.375 168.510 ;
        RECT 153.130 167.965 153.855 168.145 ;
        RECT 152.610 167.465 153.035 167.795 ;
        RECT 153.205 167.465 153.855 167.965 ;
        RECT 154.025 167.795 154.375 168.315 ;
        RECT 154.545 167.965 154.805 168.935 ;
        RECT 154.025 167.465 154.450 167.795 ;
        RECT 149.060 167.295 149.285 167.335 ;
        RECT 151.030 167.295 151.365 167.465 ;
        RECT 151.610 167.295 151.960 167.465 ;
        RECT 152.610 167.295 152.960 167.465 ;
        RECT 153.205 167.295 153.375 167.465 ;
        RECT 154.025 167.295 154.375 167.465 ;
        RECT 154.620 167.295 154.805 167.965 ;
        RECT 154.975 168.015 156.185 169.105 ;
        RECT 154.975 167.475 155.495 168.015 ;
        RECT 155.665 167.305 156.185 167.845 ;
        RECT 145.960 166.835 146.365 167.005 ;
        RECT 146.535 166.835 147.320 167.005 ;
        RECT 147.595 166.555 147.805 167.085 ;
        RECT 148.065 166.770 148.395 167.295 ;
        RECT 148.905 167.210 149.285 167.295 ;
        RECT 148.565 166.555 148.735 167.165 ;
        RECT 148.905 166.775 149.235 167.210 ;
        RECT 150.375 167.125 151.365 167.295 ;
        RECT 150.375 166.725 150.810 167.125 ;
        RECT 150.980 166.555 151.365 166.955 ;
        RECT 151.535 166.725 151.960 167.295 ;
        RECT 152.150 167.125 152.960 167.295 ;
        RECT 152.150 166.725 152.405 167.125 ;
        RECT 152.575 166.555 152.960 166.955 ;
        RECT 153.130 166.725 153.375 167.295 ;
        RECT 153.565 167.125 154.375 167.295 ;
        RECT 153.565 166.725 153.820 167.125 ;
        RECT 153.990 166.555 154.375 166.955 ;
        RECT 154.545 166.725 154.805 167.295 ;
        RECT 154.975 166.555 156.185 167.305 ;
        RECT 70.710 166.385 156.270 166.555 ;
        RECT 70.795 165.635 72.005 166.385 ;
        RECT 70.795 165.095 71.315 165.635 ;
        RECT 72.175 165.615 75.685 166.385 ;
        RECT 76.865 165.835 77.035 166.125 ;
        RECT 77.205 166.005 77.535 166.385 ;
        RECT 76.865 165.665 77.530 165.835 ;
        RECT 71.485 164.925 72.005 165.465 ;
        RECT 72.175 165.095 73.825 165.615 ;
        RECT 73.995 164.925 75.685 165.445 ;
        RECT 70.795 163.835 72.005 164.925 ;
        RECT 72.175 163.835 75.685 164.925 ;
        RECT 76.780 164.845 77.130 165.495 ;
        RECT 77.300 164.675 77.530 165.665 ;
        RECT 76.865 164.505 77.530 164.675 ;
        RECT 76.865 164.005 77.035 164.505 ;
        RECT 77.205 163.835 77.535 164.335 ;
        RECT 77.705 164.005 77.890 166.125 ;
        RECT 78.145 165.925 78.395 166.385 ;
        RECT 78.565 165.935 78.900 166.105 ;
        RECT 79.095 165.935 79.770 166.105 ;
        RECT 78.565 165.795 78.735 165.935 ;
        RECT 78.060 164.805 78.340 165.755 ;
        RECT 78.510 165.665 78.735 165.795 ;
        RECT 78.510 164.560 78.680 165.665 ;
        RECT 78.905 165.515 79.430 165.735 ;
        RECT 78.850 164.750 79.090 165.345 ;
        RECT 79.260 164.815 79.430 165.515 ;
        RECT 79.600 165.155 79.770 165.935 ;
        RECT 80.090 165.885 80.460 166.385 ;
        RECT 80.640 165.935 81.045 166.105 ;
        RECT 81.215 165.935 82.000 166.105 ;
        RECT 80.640 165.705 80.810 165.935 ;
        RECT 79.980 165.405 80.810 165.705 ;
        RECT 81.195 165.435 81.660 165.765 ;
        RECT 79.980 165.375 80.180 165.405 ;
        RECT 80.300 165.155 80.470 165.225 ;
        RECT 79.600 164.985 80.470 165.155 ;
        RECT 79.960 164.895 80.470 164.985 ;
        RECT 78.510 164.430 78.815 164.560 ;
        RECT 79.260 164.450 79.790 164.815 ;
        RECT 78.130 163.835 78.395 164.295 ;
        RECT 78.565 164.005 78.815 164.430 ;
        RECT 79.960 164.280 80.130 164.895 ;
        RECT 79.025 164.110 80.130 164.280 ;
        RECT 80.300 163.835 80.470 164.635 ;
        RECT 80.640 164.335 80.810 165.405 ;
        RECT 80.980 164.505 81.170 165.225 ;
        RECT 81.340 164.475 81.660 165.435 ;
        RECT 81.830 165.475 82.000 165.935 ;
        RECT 82.275 165.855 82.485 166.385 ;
        RECT 82.745 165.645 83.075 166.170 ;
        RECT 83.245 165.775 83.415 166.385 ;
        RECT 83.585 165.730 83.915 166.165 ;
        RECT 84.185 165.730 84.515 166.165 ;
        RECT 84.685 165.775 84.855 166.385 ;
        RECT 83.585 165.645 83.965 165.730 ;
        RECT 82.875 165.475 83.075 165.645 ;
        RECT 83.740 165.605 83.965 165.645 ;
        RECT 81.830 165.145 82.705 165.475 ;
        RECT 82.875 165.145 83.625 165.475 ;
        RECT 80.640 164.005 80.890 164.335 ;
        RECT 81.830 164.305 82.000 165.145 ;
        RECT 82.875 164.940 83.065 165.145 ;
        RECT 83.795 165.025 83.965 165.605 ;
        RECT 83.750 164.975 83.965 165.025 ;
        RECT 82.170 164.565 83.065 164.940 ;
        RECT 83.575 164.895 83.965 164.975 ;
        RECT 84.135 165.645 84.515 165.730 ;
        RECT 85.025 165.645 85.355 166.170 ;
        RECT 85.615 165.855 85.825 166.385 ;
        RECT 86.100 165.935 86.885 166.105 ;
        RECT 87.055 165.935 87.460 166.105 ;
        RECT 84.135 165.605 84.360 165.645 ;
        RECT 84.135 165.025 84.305 165.605 ;
        RECT 85.025 165.475 85.225 165.645 ;
        RECT 86.100 165.475 86.270 165.935 ;
        RECT 84.475 165.145 85.225 165.475 ;
        RECT 85.395 165.145 86.270 165.475 ;
        RECT 84.135 164.975 84.350 165.025 ;
        RECT 84.135 164.895 84.525 164.975 ;
        RECT 81.115 164.135 82.000 164.305 ;
        RECT 82.180 163.835 82.495 164.335 ;
        RECT 82.725 164.005 83.065 164.565 ;
        RECT 83.235 163.835 83.405 164.845 ;
        RECT 83.575 164.050 83.905 164.895 ;
        RECT 84.195 164.050 84.525 164.895 ;
        RECT 85.035 164.940 85.225 165.145 ;
        RECT 84.695 163.835 84.865 164.845 ;
        RECT 85.035 164.565 85.930 164.940 ;
        RECT 85.035 164.005 85.375 164.565 ;
        RECT 85.605 163.835 85.920 164.335 ;
        RECT 86.100 164.305 86.270 165.145 ;
        RECT 86.440 165.435 86.905 165.765 ;
        RECT 87.290 165.705 87.460 165.935 ;
        RECT 87.640 165.885 88.010 166.385 ;
        RECT 88.330 165.935 89.005 166.105 ;
        RECT 89.200 165.935 89.535 166.105 ;
        RECT 86.440 164.475 86.760 165.435 ;
        RECT 87.290 165.405 88.120 165.705 ;
        RECT 86.930 164.505 87.120 165.225 ;
        RECT 87.290 164.335 87.460 165.405 ;
        RECT 87.920 165.375 88.120 165.405 ;
        RECT 87.630 165.155 87.800 165.225 ;
        RECT 88.330 165.155 88.500 165.935 ;
        RECT 89.365 165.795 89.535 165.935 ;
        RECT 89.705 165.925 89.955 166.385 ;
        RECT 87.630 164.985 88.500 165.155 ;
        RECT 88.670 165.515 89.195 165.735 ;
        RECT 89.365 165.665 89.590 165.795 ;
        RECT 87.630 164.895 88.140 164.985 ;
        RECT 86.100 164.135 86.985 164.305 ;
        RECT 87.210 164.005 87.460 164.335 ;
        RECT 87.630 163.835 87.800 164.635 ;
        RECT 87.970 164.280 88.140 164.895 ;
        RECT 88.670 164.815 88.840 165.515 ;
        RECT 88.310 164.450 88.840 164.815 ;
        RECT 89.010 164.750 89.250 165.345 ;
        RECT 89.420 164.560 89.590 165.665 ;
        RECT 89.760 164.805 90.040 165.755 ;
        RECT 89.285 164.430 89.590 164.560 ;
        RECT 87.970 164.110 89.075 164.280 ;
        RECT 89.285 164.005 89.535 164.430 ;
        RECT 89.705 163.835 89.970 164.295 ;
        RECT 90.210 164.005 90.395 166.125 ;
        RECT 90.565 166.005 90.895 166.385 ;
        RECT 91.065 165.835 91.235 166.125 ;
        RECT 90.570 165.665 91.235 165.835 ;
        RECT 91.495 165.815 91.930 166.215 ;
        RECT 92.100 165.985 92.485 166.385 ;
        RECT 90.570 164.675 90.800 165.665 ;
        RECT 91.495 165.645 92.485 165.815 ;
        RECT 92.655 165.645 93.080 166.215 ;
        RECT 93.270 165.815 93.525 166.215 ;
        RECT 93.695 165.985 94.080 166.385 ;
        RECT 93.270 165.645 94.080 165.815 ;
        RECT 94.250 165.645 94.495 166.215 ;
        RECT 94.685 165.815 94.940 166.215 ;
        RECT 95.110 165.985 95.495 166.385 ;
        RECT 94.685 165.645 95.495 165.815 ;
        RECT 95.665 165.645 95.925 166.215 ;
        RECT 96.555 165.660 96.845 166.385 ;
        RECT 90.970 164.845 91.320 165.495 ;
        RECT 92.150 165.475 92.485 165.645 ;
        RECT 92.730 165.475 93.080 165.645 ;
        RECT 93.730 165.475 94.080 165.645 ;
        RECT 94.325 165.475 94.495 165.645 ;
        RECT 95.145 165.475 95.495 165.645 ;
        RECT 91.495 164.770 91.980 165.475 ;
        RECT 92.150 165.145 92.560 165.475 ;
        RECT 90.570 164.505 91.235 164.675 ;
        RECT 92.150 164.600 92.485 165.145 ;
        RECT 92.730 164.975 93.560 165.475 ;
        RECT 90.565 163.835 90.895 164.335 ;
        RECT 91.065 164.005 91.235 164.505 ;
        RECT 91.495 164.430 92.485 164.600 ;
        RECT 92.655 164.795 93.560 164.975 ;
        RECT 93.730 165.145 94.155 165.475 ;
        RECT 91.495 164.005 91.930 164.430 ;
        RECT 92.100 163.835 92.485 164.260 ;
        RECT 92.655 164.005 93.080 164.795 ;
        RECT 93.730 164.625 94.080 165.145 ;
        RECT 94.325 164.975 94.975 165.475 ;
        RECT 93.250 164.430 94.080 164.625 ;
        RECT 94.250 164.795 94.975 164.975 ;
        RECT 95.145 165.145 95.570 165.475 ;
        RECT 93.250 164.005 93.525 164.430 ;
        RECT 93.695 163.835 94.080 164.260 ;
        RECT 94.250 164.005 94.495 164.795 ;
        RECT 95.145 164.625 95.495 165.145 ;
        RECT 95.740 164.975 95.925 165.645 ;
        RECT 97.485 165.575 97.755 166.385 ;
        RECT 97.925 165.575 98.255 166.215 ;
        RECT 98.425 165.575 98.665 166.385 ;
        RECT 98.890 165.645 99.505 166.215 ;
        RECT 99.675 165.875 99.890 166.385 ;
        RECT 100.120 165.875 100.400 166.205 ;
        RECT 100.580 165.875 100.820 166.385 ;
        RECT 101.160 165.910 101.495 166.170 ;
        RECT 101.665 165.985 101.995 166.385 ;
        RECT 102.165 165.985 103.780 166.155 ;
        RECT 97.475 165.145 97.825 165.395 ;
        RECT 94.685 164.430 95.495 164.625 ;
        RECT 94.685 164.005 94.940 164.430 ;
        RECT 95.110 163.835 95.495 164.260 ;
        RECT 95.665 164.005 95.925 164.975 ;
        RECT 96.555 163.835 96.845 165.000 ;
        RECT 97.995 164.975 98.165 165.575 ;
        RECT 98.335 165.145 98.685 165.395 ;
        RECT 97.485 163.835 97.815 164.975 ;
        RECT 97.995 164.805 98.675 164.975 ;
        RECT 98.345 164.020 98.675 164.805 ;
        RECT 98.890 164.625 99.205 165.645 ;
        RECT 99.375 164.975 99.545 165.475 ;
        RECT 99.795 165.145 100.060 165.705 ;
        RECT 100.230 164.975 100.400 165.875 ;
        RECT 100.570 165.145 100.925 165.705 ;
        RECT 99.375 164.805 100.800 164.975 ;
        RECT 98.890 164.005 99.425 164.625 ;
        RECT 99.595 163.835 99.925 164.635 ;
        RECT 100.410 164.630 100.800 164.805 ;
        RECT 101.160 164.555 101.415 165.910 ;
        RECT 102.165 165.815 102.335 165.985 ;
        RECT 101.775 165.645 102.335 165.815 ;
        RECT 101.775 165.475 101.945 165.645 ;
        RECT 101.640 165.145 101.945 165.475 ;
        RECT 102.140 165.365 102.390 165.475 ;
        RECT 102.600 165.365 102.870 165.805 ;
        RECT 103.060 165.705 103.350 165.805 ;
        RECT 103.055 165.535 103.350 165.705 ;
        RECT 102.135 165.195 102.390 165.365 ;
        RECT 102.595 165.195 102.870 165.365 ;
        RECT 102.140 165.145 102.390 165.195 ;
        RECT 102.600 165.145 102.870 165.195 ;
        RECT 103.060 165.145 103.350 165.535 ;
        RECT 103.520 165.145 103.940 165.810 ;
        RECT 104.325 165.665 104.655 166.385 ;
        RECT 104.875 165.565 105.105 166.385 ;
        RECT 105.275 165.585 105.605 166.215 ;
        RECT 104.250 165.145 104.600 165.475 ;
        RECT 104.855 165.145 105.185 165.395 ;
        RECT 101.775 164.975 101.945 165.145 ;
        RECT 104.395 165.025 104.600 165.145 ;
        RECT 101.775 164.805 104.145 164.975 ;
        RECT 104.395 164.855 104.605 165.025 ;
        RECT 105.355 164.985 105.605 165.585 ;
        RECT 105.775 165.565 105.985 166.385 ;
        RECT 106.215 165.615 107.885 166.385 ;
        RECT 108.055 165.815 108.490 166.215 ;
        RECT 108.660 165.985 109.045 166.385 ;
        RECT 108.055 165.645 109.045 165.815 ;
        RECT 109.215 165.645 109.640 166.215 ;
        RECT 109.830 165.815 110.085 166.215 ;
        RECT 110.255 165.985 110.640 166.385 ;
        RECT 109.830 165.645 110.640 165.815 ;
        RECT 110.810 165.645 111.055 166.215 ;
        RECT 111.245 165.815 111.500 166.215 ;
        RECT 111.670 165.985 112.055 166.385 ;
        RECT 111.245 165.645 112.055 165.815 ;
        RECT 112.225 165.645 112.485 166.215 ;
        RECT 106.215 165.095 106.965 165.615 ;
        RECT 108.710 165.475 109.045 165.645 ;
        RECT 109.290 165.475 109.640 165.645 ;
        RECT 110.290 165.475 110.640 165.645 ;
        RECT 110.885 165.475 111.055 165.645 ;
        RECT 111.705 165.475 112.055 165.645 ;
        RECT 101.160 164.045 101.495 164.555 ;
        RECT 101.745 163.835 102.075 164.635 ;
        RECT 102.320 164.425 103.745 164.595 ;
        RECT 102.320 164.005 102.605 164.425 ;
        RECT 102.860 163.835 103.190 164.255 ;
        RECT 103.415 164.175 103.745 164.425 ;
        RECT 103.975 164.345 104.145 164.805 ;
        RECT 104.405 164.175 104.575 164.675 ;
        RECT 103.415 164.005 104.575 164.175 ;
        RECT 104.875 163.835 105.105 164.975 ;
        RECT 105.275 164.005 105.605 164.985 ;
        RECT 105.775 163.835 105.985 164.975 ;
        RECT 107.135 164.925 107.885 165.445 ;
        RECT 106.215 163.835 107.885 164.925 ;
        RECT 108.055 164.770 108.540 165.475 ;
        RECT 108.710 165.145 109.120 165.475 ;
        RECT 108.710 164.600 109.045 165.145 ;
        RECT 109.290 164.975 110.120 165.475 ;
        RECT 108.055 164.430 109.045 164.600 ;
        RECT 109.215 164.795 110.120 164.975 ;
        RECT 110.290 165.145 110.715 165.475 ;
        RECT 108.055 164.005 108.490 164.430 ;
        RECT 108.660 163.835 109.045 164.260 ;
        RECT 109.215 164.005 109.640 164.795 ;
        RECT 110.290 164.625 110.640 165.145 ;
        RECT 110.885 164.975 111.535 165.475 ;
        RECT 109.810 164.430 110.640 164.625 ;
        RECT 110.810 164.795 111.535 164.975 ;
        RECT 111.705 165.145 112.130 165.475 ;
        RECT 109.810 164.005 110.085 164.430 ;
        RECT 110.255 163.835 110.640 164.260 ;
        RECT 110.810 164.005 111.055 164.795 ;
        RECT 111.705 164.625 112.055 165.145 ;
        RECT 112.300 164.975 112.485 165.645 ;
        RECT 111.245 164.430 112.055 164.625 ;
        RECT 111.245 164.005 111.500 164.430 ;
        RECT 111.670 163.835 112.055 164.260 ;
        RECT 112.225 164.005 112.485 164.975 ;
        RECT 112.655 165.585 112.995 166.215 ;
        RECT 113.165 165.585 113.415 166.385 ;
        RECT 113.605 165.735 113.935 166.215 ;
        RECT 114.105 165.925 114.330 166.385 ;
        RECT 114.500 165.735 114.830 166.215 ;
        RECT 112.655 165.535 112.885 165.585 ;
        RECT 113.605 165.565 114.830 165.735 ;
        RECT 115.460 165.605 115.960 166.215 ;
        RECT 116.335 165.615 118.005 166.385 ;
        RECT 118.640 165.620 119.095 166.385 ;
        RECT 119.370 166.005 120.670 166.215 ;
        RECT 120.925 166.025 121.255 166.385 ;
        RECT 120.500 165.855 120.670 166.005 ;
        RECT 121.425 165.885 121.685 166.215 ;
        RECT 121.455 165.875 121.685 165.885 ;
        RECT 112.655 164.975 112.830 165.535 ;
        RECT 113.000 165.225 113.695 165.395 ;
        RECT 113.525 164.975 113.695 165.225 ;
        RECT 113.870 165.195 114.290 165.395 ;
        RECT 114.460 165.195 114.790 165.395 ;
        RECT 114.960 165.195 115.290 165.395 ;
        RECT 115.460 164.975 115.630 165.605 ;
        RECT 115.815 165.145 116.165 165.395 ;
        RECT 116.335 165.095 117.085 165.615 ;
        RECT 112.655 164.005 112.995 164.975 ;
        RECT 113.165 163.835 113.335 164.975 ;
        RECT 113.525 164.805 115.960 164.975 ;
        RECT 117.255 164.925 118.005 165.445 ;
        RECT 119.570 165.395 119.790 165.795 ;
        RECT 118.635 165.195 119.125 165.395 ;
        RECT 119.315 165.185 119.790 165.395 ;
        RECT 120.035 165.395 120.245 165.795 ;
        RECT 120.500 165.730 121.255 165.855 ;
        RECT 120.500 165.685 121.345 165.730 ;
        RECT 121.075 165.565 121.345 165.685 ;
        RECT 120.035 165.185 120.365 165.395 ;
        RECT 120.535 165.125 120.945 165.430 ;
        RECT 113.605 163.835 113.855 164.635 ;
        RECT 114.500 164.005 114.830 164.805 ;
        RECT 115.130 163.835 115.460 164.635 ;
        RECT 115.630 164.005 115.960 164.805 ;
        RECT 116.335 163.835 118.005 164.925 ;
        RECT 118.640 164.955 119.815 165.015 ;
        RECT 121.175 164.990 121.345 165.565 ;
        RECT 121.145 164.955 121.345 164.990 ;
        RECT 118.640 164.845 121.345 164.955 ;
        RECT 118.640 164.225 118.895 164.845 ;
        RECT 119.485 164.785 121.285 164.845 ;
        RECT 119.485 164.755 119.815 164.785 ;
        RECT 121.515 164.685 121.685 165.875 ;
        RECT 122.315 165.660 122.605 166.385 ;
        RECT 122.810 165.645 123.425 166.215 ;
        RECT 123.595 165.875 123.810 166.385 ;
        RECT 124.040 165.875 124.320 166.205 ;
        RECT 124.500 165.875 124.740 166.385 ;
        RECT 119.145 164.585 119.330 164.675 ;
        RECT 119.920 164.585 120.755 164.595 ;
        RECT 119.145 164.385 120.755 164.585 ;
        RECT 119.145 164.345 119.375 164.385 ;
        RECT 118.640 164.005 118.975 164.225 ;
        RECT 119.980 163.835 120.335 164.215 ;
        RECT 120.505 164.005 120.755 164.385 ;
        RECT 121.005 163.835 121.255 164.615 ;
        RECT 121.425 164.005 121.685 164.685 ;
        RECT 122.315 163.835 122.605 165.000 ;
        RECT 122.810 164.625 123.125 165.645 ;
        RECT 123.295 164.975 123.465 165.475 ;
        RECT 123.715 165.145 123.980 165.705 ;
        RECT 124.150 164.975 124.320 165.875 ;
        RECT 125.075 165.735 125.335 166.215 ;
        RECT 125.505 165.845 125.755 166.385 ;
        RECT 124.490 165.145 124.845 165.705 ;
        RECT 123.295 164.805 124.720 164.975 ;
        RECT 122.810 164.005 123.345 164.625 ;
        RECT 123.515 163.835 123.845 164.635 ;
        RECT 124.330 164.630 124.720 164.805 ;
        RECT 125.075 164.705 125.245 165.735 ;
        RECT 125.925 165.705 126.145 166.165 ;
        RECT 125.895 165.680 126.145 165.705 ;
        RECT 125.415 165.085 125.645 165.480 ;
        RECT 125.815 165.255 126.145 165.680 ;
        RECT 126.315 166.005 127.205 166.175 ;
        RECT 126.315 165.280 126.485 166.005 ;
        RECT 126.655 165.450 127.205 165.835 ;
        RECT 127.375 165.615 129.045 166.385 ;
        RECT 126.315 165.210 127.205 165.280 ;
        RECT 126.310 165.185 127.205 165.210 ;
        RECT 126.300 165.170 127.205 165.185 ;
        RECT 126.295 165.155 127.205 165.170 ;
        RECT 126.285 165.150 127.205 165.155 ;
        RECT 126.280 165.140 127.205 165.150 ;
        RECT 126.275 165.130 127.205 165.140 ;
        RECT 126.265 165.125 127.205 165.130 ;
        RECT 126.255 165.115 127.205 165.125 ;
        RECT 126.245 165.110 127.205 165.115 ;
        RECT 126.245 165.105 126.580 165.110 ;
        RECT 126.230 165.100 126.580 165.105 ;
        RECT 126.215 165.090 126.580 165.100 ;
        RECT 126.190 165.085 126.580 165.090 ;
        RECT 125.415 165.080 126.580 165.085 ;
        RECT 125.415 165.045 126.550 165.080 ;
        RECT 125.415 165.020 126.515 165.045 ;
        RECT 125.415 164.990 126.485 165.020 ;
        RECT 125.415 164.960 126.465 164.990 ;
        RECT 125.415 164.930 126.445 164.960 ;
        RECT 125.415 164.920 126.375 164.930 ;
        RECT 125.415 164.910 126.350 164.920 ;
        RECT 125.415 164.895 126.330 164.910 ;
        RECT 125.415 164.880 126.310 164.895 ;
        RECT 125.520 164.870 126.305 164.880 ;
        RECT 125.520 164.835 126.290 164.870 ;
        RECT 125.075 164.005 125.350 164.705 ;
        RECT 125.520 164.585 126.275 164.835 ;
        RECT 126.445 164.515 126.775 164.760 ;
        RECT 126.945 164.660 127.205 165.110 ;
        RECT 127.375 165.095 128.125 165.615 ;
        RECT 129.685 165.575 129.955 166.385 ;
        RECT 130.125 165.575 130.455 166.215 ;
        RECT 130.625 165.575 130.865 166.385 ;
        RECT 131.055 165.635 132.265 166.385 ;
        RECT 132.435 165.815 132.870 166.215 ;
        RECT 133.040 165.985 133.425 166.385 ;
        RECT 132.435 165.645 133.425 165.815 ;
        RECT 133.595 165.645 134.020 166.215 ;
        RECT 134.210 165.815 134.465 166.215 ;
        RECT 134.635 165.985 135.020 166.385 ;
        RECT 134.210 165.645 135.020 165.815 ;
        RECT 135.190 165.645 135.435 166.215 ;
        RECT 135.625 165.815 135.880 166.215 ;
        RECT 136.050 165.985 136.435 166.385 ;
        RECT 135.625 165.645 136.435 165.815 ;
        RECT 136.605 165.645 136.865 166.215 ;
        RECT 137.035 165.815 137.470 166.215 ;
        RECT 137.640 165.985 138.025 166.385 ;
        RECT 137.035 165.645 138.025 165.815 ;
        RECT 138.195 165.645 138.620 166.215 ;
        RECT 138.810 165.815 139.065 166.215 ;
        RECT 139.235 165.985 139.620 166.385 ;
        RECT 138.810 165.645 139.620 165.815 ;
        RECT 139.790 165.645 140.035 166.215 ;
        RECT 140.225 165.815 140.480 166.215 ;
        RECT 140.650 165.985 141.035 166.385 ;
        RECT 140.225 165.645 141.035 165.815 ;
        RECT 141.205 165.645 141.465 166.215 ;
        RECT 141.725 165.835 141.895 166.215 ;
        RECT 142.075 166.005 142.405 166.385 ;
        RECT 141.725 165.665 142.390 165.835 ;
        RECT 142.585 165.710 142.845 166.215 ;
        RECT 128.295 164.925 129.045 165.445 ;
        RECT 129.675 165.145 130.025 165.395 ;
        RECT 130.195 164.975 130.365 165.575 ;
        RECT 130.535 165.145 130.885 165.395 ;
        RECT 131.055 165.095 131.575 165.635 ;
        RECT 133.090 165.475 133.425 165.645 ;
        RECT 133.670 165.475 134.020 165.645 ;
        RECT 134.670 165.475 135.020 165.645 ;
        RECT 135.265 165.475 135.435 165.645 ;
        RECT 136.085 165.475 136.435 165.645 ;
        RECT 126.590 164.490 126.775 164.515 ;
        RECT 126.590 164.390 127.205 164.490 ;
        RECT 125.520 163.835 125.775 164.380 ;
        RECT 125.945 164.005 126.425 164.345 ;
        RECT 126.600 163.835 127.205 164.390 ;
        RECT 127.375 163.835 129.045 164.925 ;
        RECT 129.685 163.835 130.015 164.975 ;
        RECT 130.195 164.805 130.875 164.975 ;
        RECT 131.745 164.925 132.265 165.465 ;
        RECT 130.545 164.020 130.875 164.805 ;
        RECT 131.055 163.835 132.265 164.925 ;
        RECT 132.435 164.770 132.920 165.475 ;
        RECT 133.090 165.145 133.500 165.475 ;
        RECT 133.090 164.600 133.425 165.145 ;
        RECT 133.670 164.975 134.500 165.475 ;
        RECT 132.435 164.430 133.425 164.600 ;
        RECT 133.595 164.795 134.500 164.975 ;
        RECT 134.670 165.145 135.095 165.475 ;
        RECT 132.435 164.005 132.870 164.430 ;
        RECT 133.040 163.835 133.425 164.260 ;
        RECT 133.595 164.005 134.020 164.795 ;
        RECT 134.670 164.625 135.020 165.145 ;
        RECT 135.265 164.975 135.915 165.475 ;
        RECT 134.190 164.430 135.020 164.625 ;
        RECT 135.190 164.795 135.915 164.975 ;
        RECT 136.085 165.145 136.510 165.475 ;
        RECT 134.190 164.005 134.465 164.430 ;
        RECT 134.635 163.835 135.020 164.260 ;
        RECT 135.190 164.005 135.435 164.795 ;
        RECT 136.085 164.625 136.435 165.145 ;
        RECT 136.680 164.975 136.865 165.645 ;
        RECT 137.690 165.475 138.025 165.645 ;
        RECT 138.270 165.475 138.620 165.645 ;
        RECT 139.270 165.475 139.620 165.645 ;
        RECT 139.865 165.475 140.035 165.645 ;
        RECT 140.685 165.475 141.035 165.645 ;
        RECT 135.625 164.430 136.435 164.625 ;
        RECT 135.625 164.005 135.880 164.430 ;
        RECT 136.050 163.835 136.435 164.260 ;
        RECT 136.605 164.005 136.865 164.975 ;
        RECT 137.035 164.770 137.520 165.475 ;
        RECT 137.690 165.145 138.100 165.475 ;
        RECT 137.690 164.600 138.025 165.145 ;
        RECT 138.270 164.975 139.100 165.475 ;
        RECT 137.035 164.430 138.025 164.600 ;
        RECT 138.195 164.795 139.100 164.975 ;
        RECT 139.270 165.145 139.695 165.475 ;
        RECT 137.035 164.005 137.470 164.430 ;
        RECT 137.640 163.835 138.025 164.260 ;
        RECT 138.195 164.005 138.620 164.795 ;
        RECT 139.270 164.625 139.620 165.145 ;
        RECT 139.865 164.975 140.515 165.475 ;
        RECT 138.790 164.430 139.620 164.625 ;
        RECT 139.790 164.795 140.515 164.975 ;
        RECT 140.685 165.145 141.110 165.475 ;
        RECT 138.790 164.005 139.065 164.430 ;
        RECT 139.235 163.835 139.620 164.260 ;
        RECT 139.790 164.005 140.035 164.795 ;
        RECT 140.685 164.625 141.035 165.145 ;
        RECT 141.280 164.975 141.465 165.645 ;
        RECT 141.655 165.115 141.995 165.485 ;
        RECT 142.220 165.410 142.390 165.665 ;
        RECT 140.225 164.430 141.035 164.625 ;
        RECT 140.225 164.005 140.480 164.430 ;
        RECT 140.650 163.835 141.035 164.260 ;
        RECT 141.205 164.005 141.465 164.975 ;
        RECT 142.220 165.080 142.495 165.410 ;
        RECT 142.220 164.935 142.390 165.080 ;
        RECT 141.715 164.765 142.390 164.935 ;
        RECT 142.665 164.910 142.845 165.710 ;
        RECT 143.075 165.565 143.285 166.385 ;
        RECT 143.455 165.585 143.785 166.215 ;
        RECT 143.455 164.985 143.705 165.585 ;
        RECT 143.955 165.565 144.185 166.385 ;
        RECT 144.395 165.615 146.065 166.385 ;
        RECT 143.875 165.145 144.205 165.395 ;
        RECT 144.395 165.095 145.145 165.615 ;
        RECT 146.755 165.565 146.965 166.385 ;
        RECT 147.135 165.585 147.465 166.215 ;
        RECT 141.715 164.005 141.895 164.765 ;
        RECT 142.075 163.835 142.405 164.595 ;
        RECT 142.575 164.005 142.845 164.910 ;
        RECT 143.075 163.835 143.285 164.975 ;
        RECT 143.455 164.005 143.785 164.985 ;
        RECT 143.955 163.835 144.185 164.975 ;
        RECT 145.315 164.925 146.065 165.445 ;
        RECT 147.135 164.985 147.385 165.585 ;
        RECT 147.635 165.565 147.865 166.385 ;
        RECT 148.075 165.660 148.365 166.385 ;
        RECT 148.535 165.645 148.795 166.215 ;
        RECT 148.965 165.985 149.350 166.385 ;
        RECT 149.520 165.815 149.775 166.215 ;
        RECT 148.965 165.645 149.775 165.815 ;
        RECT 149.965 165.645 150.210 166.215 ;
        RECT 150.380 165.985 150.765 166.385 ;
        RECT 150.935 165.815 151.190 166.215 ;
        RECT 150.380 165.645 151.190 165.815 ;
        RECT 151.380 165.645 151.805 166.215 ;
        RECT 151.975 165.985 152.360 166.385 ;
        RECT 152.530 165.815 152.965 166.215 ;
        RECT 151.975 165.645 152.965 165.815 ;
        RECT 153.225 165.835 153.395 166.215 ;
        RECT 153.575 166.005 153.905 166.385 ;
        RECT 153.225 165.665 153.890 165.835 ;
        RECT 154.085 165.710 154.345 166.215 ;
        RECT 147.555 165.145 147.885 165.395 ;
        RECT 144.395 163.835 146.065 164.925 ;
        RECT 146.755 163.835 146.965 164.975 ;
        RECT 147.135 164.005 147.465 164.985 ;
        RECT 147.635 163.835 147.865 164.975 ;
        RECT 148.075 163.835 148.365 165.000 ;
        RECT 148.535 164.975 148.720 165.645 ;
        RECT 148.965 165.475 149.315 165.645 ;
        RECT 149.965 165.475 150.135 165.645 ;
        RECT 150.380 165.475 150.730 165.645 ;
        RECT 151.380 165.475 151.730 165.645 ;
        RECT 151.975 165.475 152.310 165.645 ;
        RECT 148.890 165.145 149.315 165.475 ;
        RECT 148.535 164.005 148.795 164.975 ;
        RECT 148.965 164.625 149.315 165.145 ;
        RECT 149.485 164.975 150.135 165.475 ;
        RECT 150.305 165.145 150.730 165.475 ;
        RECT 149.485 164.795 150.210 164.975 ;
        RECT 148.965 164.430 149.775 164.625 ;
        RECT 148.965 163.835 149.350 164.260 ;
        RECT 149.520 164.005 149.775 164.430 ;
        RECT 149.965 164.005 150.210 164.795 ;
        RECT 150.380 164.625 150.730 165.145 ;
        RECT 150.900 164.975 151.730 165.475 ;
        RECT 151.900 165.145 152.310 165.475 ;
        RECT 150.900 164.795 151.805 164.975 ;
        RECT 150.380 164.430 151.210 164.625 ;
        RECT 150.380 163.835 150.765 164.260 ;
        RECT 150.935 164.005 151.210 164.430 ;
        RECT 151.380 164.005 151.805 164.795 ;
        RECT 151.975 164.600 152.310 165.145 ;
        RECT 152.480 164.770 152.965 165.475 ;
        RECT 153.155 165.115 153.495 165.485 ;
        RECT 153.720 165.410 153.890 165.665 ;
        RECT 153.720 165.080 153.995 165.410 ;
        RECT 153.720 164.935 153.890 165.080 ;
        RECT 153.215 164.765 153.890 164.935 ;
        RECT 154.165 164.910 154.345 165.710 ;
        RECT 154.975 165.635 156.185 166.385 ;
        RECT 151.975 164.430 152.965 164.600 ;
        RECT 151.975 163.835 152.360 164.260 ;
        RECT 152.530 164.005 152.965 164.430 ;
        RECT 153.215 164.005 153.395 164.765 ;
        RECT 153.575 163.835 153.905 164.595 ;
        RECT 154.075 164.005 154.345 164.910 ;
        RECT 154.975 164.925 155.495 165.465 ;
        RECT 155.665 165.095 156.185 165.635 ;
        RECT 154.975 163.835 156.185 164.925 ;
        RECT 70.710 163.665 156.270 163.835 ;
        RECT 70.795 162.575 72.005 163.665 ;
        RECT 72.235 162.605 72.565 163.450 ;
        RECT 72.735 162.655 72.905 163.665 ;
        RECT 73.075 162.935 73.415 163.495 ;
        RECT 73.645 163.165 73.960 163.665 ;
        RECT 74.140 163.195 75.025 163.365 ;
        RECT 70.795 161.865 71.315 162.405 ;
        RECT 71.485 162.035 72.005 162.575 ;
        RECT 72.175 162.525 72.565 162.605 ;
        RECT 73.075 162.560 73.970 162.935 ;
        RECT 72.175 162.475 72.390 162.525 ;
        RECT 72.175 161.895 72.345 162.475 ;
        RECT 73.075 162.355 73.265 162.560 ;
        RECT 74.140 162.355 74.310 163.195 ;
        RECT 75.250 163.165 75.500 163.495 ;
        RECT 72.515 162.025 73.265 162.355 ;
        RECT 73.435 162.025 74.310 162.355 ;
        RECT 70.795 161.115 72.005 161.865 ;
        RECT 72.175 161.855 72.400 161.895 ;
        RECT 73.065 161.855 73.265 162.025 ;
        RECT 72.175 161.770 72.555 161.855 ;
        RECT 72.225 161.335 72.555 161.770 ;
        RECT 72.725 161.115 72.895 161.725 ;
        RECT 73.065 161.330 73.395 161.855 ;
        RECT 73.655 161.115 73.865 161.645 ;
        RECT 74.140 161.565 74.310 162.025 ;
        RECT 74.480 162.065 74.800 163.025 ;
        RECT 74.970 162.275 75.160 162.995 ;
        RECT 75.330 162.095 75.500 163.165 ;
        RECT 75.670 162.865 75.840 163.665 ;
        RECT 76.010 163.220 77.115 163.390 ;
        RECT 76.010 162.605 76.180 163.220 ;
        RECT 77.325 163.070 77.575 163.495 ;
        RECT 77.745 163.205 78.010 163.665 ;
        RECT 76.350 162.685 76.880 163.050 ;
        RECT 77.325 162.940 77.630 163.070 ;
        RECT 75.670 162.515 76.180 162.605 ;
        RECT 75.670 162.345 76.540 162.515 ;
        RECT 75.670 162.275 75.840 162.345 ;
        RECT 75.960 162.095 76.160 162.125 ;
        RECT 74.480 161.735 74.945 162.065 ;
        RECT 75.330 161.795 76.160 162.095 ;
        RECT 75.330 161.565 75.500 161.795 ;
        RECT 74.140 161.395 74.925 161.565 ;
        RECT 75.095 161.395 75.500 161.565 ;
        RECT 75.680 161.115 76.050 161.615 ;
        RECT 76.370 161.565 76.540 162.345 ;
        RECT 76.710 161.985 76.880 162.685 ;
        RECT 77.050 162.155 77.290 162.750 ;
        RECT 76.710 161.765 77.235 161.985 ;
        RECT 77.460 161.835 77.630 162.940 ;
        RECT 77.405 161.705 77.630 161.835 ;
        RECT 77.800 161.745 78.080 162.695 ;
        RECT 77.405 161.565 77.575 161.705 ;
        RECT 76.370 161.395 77.045 161.565 ;
        RECT 77.240 161.395 77.575 161.565 ;
        RECT 77.745 161.115 77.995 161.575 ;
        RECT 78.250 161.375 78.435 163.495 ;
        RECT 78.605 163.165 78.935 163.665 ;
        RECT 79.105 162.995 79.275 163.495 ;
        RECT 78.610 162.825 79.275 162.995 ;
        RECT 78.610 161.835 78.840 162.825 ;
        RECT 79.010 162.005 79.360 162.655 ;
        RECT 79.535 162.575 83.045 163.665 ;
        RECT 79.535 161.885 81.185 162.405 ;
        RECT 81.355 162.055 83.045 162.575 ;
        RECT 83.675 162.500 83.965 163.665 ;
        RECT 84.135 162.575 86.725 163.665 ;
        RECT 87.095 163.325 88.705 163.495 ;
        RECT 87.095 162.825 87.345 163.325 ;
        RECT 87.515 162.655 87.765 163.155 ;
        RECT 87.935 162.985 88.705 163.325 ;
        RECT 88.875 163.165 89.180 163.665 ;
        RECT 89.350 162.985 89.600 163.495 ;
        RECT 89.770 163.165 90.020 163.665 ;
        RECT 90.190 163.155 90.505 163.495 ;
        RECT 90.710 163.325 91.800 163.495 ;
        RECT 90.710 163.165 90.960 163.325 ;
        RECT 91.550 163.165 91.800 163.325 ;
        RECT 91.970 163.165 92.220 163.665 ;
        RECT 92.390 163.165 92.670 163.495 ;
        RECT 91.555 163.155 91.725 163.165 ;
        RECT 92.475 163.155 92.645 163.165 ;
        RECT 90.190 162.985 90.400 163.155 ;
        RECT 91.130 162.985 91.380 163.155 ;
        RECT 92.875 163.065 93.135 163.485 ;
        RECT 93.305 163.235 93.635 163.665 ;
        RECT 94.300 163.235 95.045 163.405 ;
        RECT 87.935 162.815 90.400 162.985 ;
        RECT 90.570 162.815 92.670 162.985 ;
        RECT 84.135 161.885 85.345 162.405 ;
        RECT 85.515 162.055 86.725 162.575 ;
        RECT 86.895 162.445 87.765 162.655 ;
        RECT 90.570 162.645 90.740 162.815 ;
        RECT 88.005 162.475 90.740 162.645 ;
        RECT 90.910 162.475 92.085 162.645 ;
        RECT 86.895 161.935 87.305 162.445 ;
        RECT 88.005 162.275 88.175 162.475 ;
        RECT 90.910 162.305 91.080 162.475 ;
        RECT 91.915 162.305 92.085 162.475 ;
        RECT 87.515 162.105 88.175 162.275 ;
        RECT 88.700 162.105 89.370 162.305 ;
        RECT 89.560 162.105 91.080 162.305 ;
        RECT 91.250 162.105 91.745 162.305 ;
        RECT 91.915 162.105 92.245 162.305 ;
        RECT 92.500 161.935 92.670 162.815 ;
        RECT 78.610 161.665 79.275 161.835 ;
        RECT 78.605 161.115 78.935 161.495 ;
        RECT 79.105 161.375 79.275 161.665 ;
        RECT 79.535 161.115 83.045 161.885 ;
        RECT 83.675 161.115 83.965 161.840 ;
        RECT 84.135 161.115 86.725 161.885 ;
        RECT 86.895 161.755 89.165 161.935 ;
        RECT 87.475 161.675 87.805 161.755 ;
        RECT 88.835 161.675 89.165 161.755 ;
        RECT 89.390 161.755 90.480 161.935 ;
        RECT 87.135 161.115 87.305 161.585 ;
        RECT 87.975 161.115 88.145 161.585 ;
        RECT 89.390 161.505 89.640 161.755 ;
        RECT 88.410 161.285 89.640 161.505 ;
        RECT 89.810 161.115 89.980 161.585 ;
        RECT 90.150 161.285 90.480 161.755 ;
        RECT 91.090 161.755 92.670 161.935 ;
        RECT 92.875 162.895 94.705 163.065 ;
        RECT 92.875 161.855 93.045 162.895 ;
        RECT 93.215 162.025 93.565 162.725 ;
        RECT 93.780 162.555 94.365 162.725 ;
        RECT 93.735 162.025 94.025 162.355 ;
        RECT 94.195 162.275 94.365 162.555 ;
        RECT 94.535 162.615 94.705 162.895 ;
        RECT 94.875 162.985 95.045 163.235 ;
        RECT 95.270 163.155 95.910 163.485 ;
        RECT 94.875 162.815 95.910 162.985 ;
        RECT 96.080 162.865 96.360 163.665 ;
        RECT 95.740 162.695 95.910 162.815 ;
        RECT 94.535 162.445 95.185 162.615 ;
        RECT 95.740 162.525 96.400 162.695 ;
        RECT 96.570 162.525 96.845 163.495 ;
        RECT 94.195 162.105 94.620 162.275 ;
        RECT 94.195 161.855 94.365 162.105 ;
        RECT 95.015 162.025 95.185 162.445 ;
        RECT 96.230 162.355 96.400 162.525 ;
        RECT 95.405 162.025 96.060 162.355 ;
        RECT 96.230 162.025 96.505 162.355 ;
        RECT 96.230 161.855 96.400 162.025 ;
        RECT 90.750 161.115 90.920 161.585 ;
        RECT 91.090 161.285 91.420 161.755 ;
        RECT 91.590 161.115 91.760 161.585 ;
        RECT 91.930 161.285 92.260 161.755 ;
        RECT 92.430 161.115 92.600 161.585 ;
        RECT 92.875 161.480 93.190 161.855 ;
        RECT 93.445 161.115 93.615 161.855 ;
        RECT 93.865 161.685 94.365 161.855 ;
        RECT 94.805 161.685 96.400 161.855 ;
        RECT 96.675 161.790 96.845 162.525 ;
        RECT 93.865 161.480 94.035 161.685 ;
        RECT 94.260 161.115 94.635 161.515 ;
        RECT 94.805 161.335 94.975 161.685 ;
        RECT 95.160 161.115 95.490 161.515 ;
        RECT 95.660 161.335 95.830 161.685 ;
        RECT 96.000 161.115 96.380 161.515 ;
        RECT 96.570 161.445 96.845 161.790 ;
        RECT 97.015 161.395 97.295 163.495 ;
        RECT 97.485 162.905 98.270 163.665 ;
        RECT 98.665 162.835 99.050 163.495 ;
        RECT 98.665 162.735 99.075 162.835 ;
        RECT 97.465 162.525 99.075 162.735 ;
        RECT 99.375 162.645 99.575 163.435 ;
        RECT 97.465 161.925 97.740 162.525 ;
        RECT 99.245 162.475 99.575 162.645 ;
        RECT 99.745 162.485 100.065 163.665 ;
        RECT 100.255 162.610 100.560 163.395 ;
        RECT 100.740 163.195 101.425 163.665 ;
        RECT 100.735 162.675 101.430 162.985 ;
        RECT 100.255 162.475 100.465 162.610 ;
        RECT 101.605 162.505 101.890 163.450 ;
        RECT 102.065 163.215 102.395 163.665 ;
        RECT 102.565 163.045 102.735 163.475 ;
        RECT 99.245 162.355 99.425 162.475 ;
        RECT 97.910 162.105 98.265 162.355 ;
        RECT 98.460 162.305 98.925 162.355 ;
        RECT 98.455 162.135 98.925 162.305 ;
        RECT 98.460 162.105 98.925 162.135 ;
        RECT 99.095 162.105 99.425 162.355 ;
        RECT 99.600 162.105 100.065 162.305 ;
        RECT 97.465 161.745 98.715 161.925 ;
        RECT 98.350 161.675 98.715 161.745 ;
        RECT 98.885 161.725 100.065 161.895 ;
        RECT 97.525 161.115 97.695 161.575 ;
        RECT 98.885 161.505 99.215 161.725 ;
        RECT 97.965 161.325 99.215 161.505 ;
        RECT 99.385 161.115 99.555 161.555 ;
        RECT 99.725 161.310 100.065 161.725 ;
        RECT 100.255 161.805 100.430 162.475 ;
        RECT 101.030 162.355 101.890 162.505 ;
        RECT 100.605 162.335 101.890 162.355 ;
        RECT 102.060 162.815 102.735 163.045 ;
        RECT 100.605 161.975 101.590 162.335 ;
        RECT 102.060 162.165 102.295 162.815 ;
        RECT 100.255 161.285 100.495 161.805 ;
        RECT 101.420 161.640 101.590 161.975 ;
        RECT 101.760 161.835 102.295 162.165 ;
        RECT 102.075 161.685 102.295 161.835 ;
        RECT 102.465 161.795 102.765 162.645 ;
        RECT 103.035 162.525 103.265 163.665 ;
        RECT 103.435 162.515 103.765 163.495 ;
        RECT 103.935 162.525 104.145 163.665 ;
        RECT 104.385 162.695 104.715 163.480 ;
        RECT 104.385 162.525 105.065 162.695 ;
        RECT 105.245 162.525 105.575 163.665 ;
        RECT 103.015 162.105 103.345 162.355 ;
        RECT 100.665 161.115 101.060 161.610 ;
        RECT 101.420 161.445 101.795 161.640 ;
        RECT 101.625 161.300 101.795 161.445 ;
        RECT 102.075 161.310 102.315 161.685 ;
        RECT 102.485 161.115 102.820 161.620 ;
        RECT 103.035 161.115 103.265 161.935 ;
        RECT 103.515 161.915 103.765 162.515 ;
        RECT 104.375 162.105 104.725 162.355 ;
        RECT 103.435 161.285 103.765 161.915 ;
        RECT 103.935 161.115 104.145 161.935 ;
        RECT 104.895 161.925 105.065 162.525 ;
        RECT 105.235 162.105 105.585 162.355 ;
        RECT 104.395 161.115 104.635 161.925 ;
        RECT 104.805 161.285 105.135 161.925 ;
        RECT 105.305 161.115 105.575 161.925 ;
        RECT 106.225 161.295 106.485 163.485 ;
        RECT 106.655 162.935 106.995 163.665 ;
        RECT 107.175 162.755 107.445 163.485 ;
        RECT 106.675 162.535 107.445 162.755 ;
        RECT 107.625 162.775 107.855 163.485 ;
        RECT 108.025 162.955 108.355 163.665 ;
        RECT 108.525 162.775 108.785 163.485 ;
        RECT 107.625 162.535 108.785 162.775 ;
        RECT 106.675 161.865 106.965 162.535 ;
        RECT 109.435 162.500 109.725 163.665 ;
        RECT 110.355 163.070 110.790 163.495 ;
        RECT 110.960 163.240 111.345 163.665 ;
        RECT 110.355 162.900 111.345 163.070 ;
        RECT 107.145 162.045 107.610 162.355 ;
        RECT 107.790 162.045 108.315 162.355 ;
        RECT 106.675 161.665 107.905 161.865 ;
        RECT 106.745 161.115 107.415 161.485 ;
        RECT 107.595 161.295 107.905 161.665 ;
        RECT 108.085 161.405 108.315 162.045 ;
        RECT 108.495 162.025 108.795 162.355 ;
        RECT 110.355 162.025 110.840 162.730 ;
        RECT 111.010 162.355 111.345 162.900 ;
        RECT 111.515 162.705 111.940 163.495 ;
        RECT 112.110 163.070 112.385 163.495 ;
        RECT 112.555 163.240 112.940 163.665 ;
        RECT 112.110 162.875 112.940 163.070 ;
        RECT 111.515 162.525 112.420 162.705 ;
        RECT 111.010 162.025 111.420 162.355 ;
        RECT 111.590 162.025 112.420 162.525 ;
        RECT 112.590 162.355 112.940 162.875 ;
        RECT 113.110 162.705 113.355 163.495 ;
        RECT 113.545 163.070 113.800 163.495 ;
        RECT 113.970 163.240 114.355 163.665 ;
        RECT 113.545 162.875 114.355 163.070 ;
        RECT 113.110 162.525 113.835 162.705 ;
        RECT 112.590 162.025 113.015 162.355 ;
        RECT 113.185 162.025 113.835 162.525 ;
        RECT 114.005 162.355 114.355 162.875 ;
        RECT 114.525 162.525 114.785 163.495 ;
        RECT 114.955 162.525 115.215 163.665 ;
        RECT 114.005 162.025 114.430 162.355 ;
        RECT 111.010 161.855 111.345 162.025 ;
        RECT 111.590 161.855 111.940 162.025 ;
        RECT 112.590 161.855 112.940 162.025 ;
        RECT 113.185 161.855 113.355 162.025 ;
        RECT 114.005 161.855 114.355 162.025 ;
        RECT 114.600 161.855 114.785 162.525 ;
        RECT 115.385 162.515 115.715 163.495 ;
        RECT 115.885 162.525 116.165 163.665 ;
        RECT 116.795 163.195 117.135 163.455 ;
        RECT 117.305 163.205 117.555 163.665 ;
        RECT 114.975 162.105 115.310 162.355 ;
        RECT 115.480 161.915 115.650 162.515 ;
        RECT 115.820 162.085 116.155 162.355 ;
        RECT 108.495 161.115 108.785 161.845 ;
        RECT 109.435 161.115 109.725 161.840 ;
        RECT 110.355 161.685 111.345 161.855 ;
        RECT 110.355 161.285 110.790 161.685 ;
        RECT 110.960 161.115 111.345 161.515 ;
        RECT 111.515 161.285 111.940 161.855 ;
        RECT 112.130 161.685 112.940 161.855 ;
        RECT 112.130 161.285 112.385 161.685 ;
        RECT 112.555 161.115 112.940 161.515 ;
        RECT 113.110 161.285 113.355 161.855 ;
        RECT 113.545 161.685 114.355 161.855 ;
        RECT 113.545 161.285 113.800 161.685 ;
        RECT 113.970 161.115 114.355 161.515 ;
        RECT 114.525 161.285 114.785 161.855 ;
        RECT 114.955 161.285 115.650 161.915 ;
        RECT 115.855 161.115 116.165 161.915 ;
        RECT 116.795 161.590 117.055 163.195 ;
        RECT 117.745 163.025 118.075 163.455 ;
        RECT 117.225 162.855 118.075 163.025 ;
        RECT 118.245 162.995 118.415 163.495 ;
        RECT 118.625 163.205 118.875 163.665 ;
        RECT 119.085 162.995 119.255 163.495 ;
        RECT 119.555 163.205 119.805 163.665 ;
        RECT 120.045 162.995 120.215 163.495 ;
        RECT 117.225 161.935 117.395 162.855 ;
        RECT 118.245 162.825 120.215 162.995 ;
        RECT 117.715 162.105 118.045 162.665 ;
        RECT 118.245 162.355 118.545 162.650 ;
        RECT 118.245 162.305 118.625 162.355 ;
        RECT 118.235 162.135 118.625 162.305 ;
        RECT 118.245 162.025 118.625 162.135 ;
        RECT 117.225 161.840 118.045 161.935 ;
        RECT 117.225 161.765 118.240 161.840 ;
        RECT 116.795 161.330 117.135 161.590 ;
        RECT 117.305 161.115 117.635 161.595 ;
        RECT 117.825 161.330 118.240 161.765 ;
        RECT 118.935 161.630 119.155 162.355 ;
        RECT 119.415 162.025 119.795 162.655 ;
        RECT 120.025 162.025 120.280 162.655 ;
        RECT 120.475 162.575 123.065 163.665 ;
        RECT 118.410 161.445 119.360 161.630 ;
        RECT 119.590 161.425 119.795 162.025 ;
        RECT 120.475 161.885 121.685 162.405 ;
        RECT 121.855 162.055 123.065 162.575 ;
        RECT 123.270 162.875 123.805 163.495 ;
        RECT 119.965 161.115 120.305 161.840 ;
        RECT 120.475 161.115 123.065 161.885 ;
        RECT 123.270 161.855 123.585 162.875 ;
        RECT 123.975 162.865 124.305 163.665 ;
        RECT 124.790 162.695 125.180 162.870 ;
        RECT 123.755 162.525 125.180 162.695 ;
        RECT 125.535 162.590 125.805 163.495 ;
        RECT 125.975 162.905 126.305 163.665 ;
        RECT 126.485 162.735 126.665 163.495 ;
        RECT 126.915 163.230 132.260 163.665 ;
        RECT 123.755 162.025 123.925 162.525 ;
        RECT 123.270 161.285 123.885 161.855 ;
        RECT 124.175 161.795 124.440 162.355 ;
        RECT 124.610 161.625 124.780 162.525 ;
        RECT 124.950 161.795 125.305 162.355 ;
        RECT 125.535 161.790 125.715 162.590 ;
        RECT 125.990 162.565 126.665 162.735 ;
        RECT 125.990 162.420 126.160 162.565 ;
        RECT 125.885 162.090 126.160 162.420 ;
        RECT 125.990 161.835 126.160 162.090 ;
        RECT 126.385 162.015 126.725 162.385 ;
        RECT 124.055 161.115 124.270 161.625 ;
        RECT 124.500 161.295 124.780 161.625 ;
        RECT 124.960 161.115 125.200 161.625 ;
        RECT 125.535 161.285 125.795 161.790 ;
        RECT 125.990 161.665 126.655 161.835 ;
        RECT 125.975 161.115 126.305 161.495 ;
        RECT 126.485 161.285 126.655 161.665 ;
        RECT 128.500 161.660 128.840 162.490 ;
        RECT 130.320 161.980 130.670 163.230 ;
        RECT 132.435 162.575 135.025 163.665 ;
        RECT 132.435 161.885 133.645 162.405 ;
        RECT 133.815 162.055 135.025 162.575 ;
        RECT 135.195 162.500 135.485 163.665 ;
        RECT 135.810 162.655 136.110 163.495 ;
        RECT 136.305 162.825 136.555 163.665 ;
        RECT 137.145 163.075 137.950 163.495 ;
        RECT 136.725 162.905 138.290 163.075 ;
        RECT 136.725 162.655 136.895 162.905 ;
        RECT 135.810 162.485 136.895 162.655 ;
        RECT 135.655 162.025 135.985 162.315 ;
        RECT 126.915 161.115 132.260 161.660 ;
        RECT 132.435 161.115 135.025 161.885 ;
        RECT 136.155 161.855 136.325 162.485 ;
        RECT 137.065 162.355 137.385 162.735 ;
        RECT 136.495 162.105 136.825 162.315 ;
        RECT 137.005 162.105 137.385 162.355 ;
        RECT 137.575 162.315 137.950 162.735 ;
        RECT 138.120 162.655 138.290 162.905 ;
        RECT 138.460 162.825 138.790 163.665 ;
        RECT 138.960 162.905 139.625 163.495 ;
        RECT 139.795 163.230 145.140 163.665 ;
        RECT 138.120 162.485 139.040 162.655 ;
        RECT 138.870 162.315 139.040 162.485 ;
        RECT 137.575 162.305 138.060 162.315 ;
        RECT 137.555 162.135 138.060 162.305 ;
        RECT 137.575 162.105 138.060 162.135 ;
        RECT 138.250 162.105 138.700 162.315 ;
        RECT 138.870 162.105 139.205 162.315 ;
        RECT 139.375 161.935 139.625 162.905 ;
        RECT 135.195 161.115 135.485 161.840 ;
        RECT 135.815 161.675 136.325 161.855 ;
        RECT 136.730 161.765 138.430 161.935 ;
        RECT 136.730 161.675 137.115 161.765 ;
        RECT 135.815 161.285 136.145 161.675 ;
        RECT 136.315 161.335 137.500 161.505 ;
        RECT 137.760 161.115 137.930 161.585 ;
        RECT 138.100 161.300 138.430 161.765 ;
        RECT 138.600 161.115 138.770 161.935 ;
        RECT 138.940 161.295 139.625 161.935 ;
        RECT 141.380 161.660 141.720 162.490 ;
        RECT 143.200 161.980 143.550 163.230 ;
        RECT 145.315 162.575 146.985 163.665 ;
        RECT 147.705 162.995 147.875 163.495 ;
        RECT 148.045 163.165 148.375 163.665 ;
        RECT 147.705 162.825 148.370 162.995 ;
        RECT 145.315 161.885 146.065 162.405 ;
        RECT 146.235 162.055 146.985 162.575 ;
        RECT 147.620 162.005 147.970 162.655 ;
        RECT 139.795 161.115 145.140 161.660 ;
        RECT 145.315 161.115 146.985 161.885 ;
        RECT 148.140 161.835 148.370 162.825 ;
        RECT 147.705 161.665 148.370 161.835 ;
        RECT 147.705 161.375 147.875 161.665 ;
        RECT 148.045 161.115 148.375 161.495 ;
        RECT 148.545 161.375 148.730 163.495 ;
        RECT 148.970 163.205 149.235 163.665 ;
        RECT 149.405 163.070 149.655 163.495 ;
        RECT 149.865 163.220 150.970 163.390 ;
        RECT 149.350 162.940 149.655 163.070 ;
        RECT 148.900 161.745 149.180 162.695 ;
        RECT 149.350 161.835 149.520 162.940 ;
        RECT 149.690 162.155 149.930 162.750 ;
        RECT 150.100 162.685 150.630 163.050 ;
        RECT 150.100 161.985 150.270 162.685 ;
        RECT 150.800 162.605 150.970 163.220 ;
        RECT 151.140 162.865 151.310 163.665 ;
        RECT 151.480 163.165 151.730 163.495 ;
        RECT 151.955 163.195 152.840 163.365 ;
        RECT 150.800 162.515 151.310 162.605 ;
        RECT 149.350 161.705 149.575 161.835 ;
        RECT 149.745 161.765 150.270 161.985 ;
        RECT 150.440 162.345 151.310 162.515 ;
        RECT 148.985 161.115 149.235 161.575 ;
        RECT 149.405 161.565 149.575 161.705 ;
        RECT 150.440 161.565 150.610 162.345 ;
        RECT 151.140 162.275 151.310 162.345 ;
        RECT 150.820 162.095 151.020 162.125 ;
        RECT 151.480 162.095 151.650 163.165 ;
        RECT 151.820 162.275 152.010 162.995 ;
        RECT 150.820 161.795 151.650 162.095 ;
        RECT 152.180 162.065 152.500 163.025 ;
        RECT 149.405 161.395 149.740 161.565 ;
        RECT 149.935 161.395 150.610 161.565 ;
        RECT 150.930 161.115 151.300 161.615 ;
        RECT 151.480 161.565 151.650 161.795 ;
        RECT 152.035 161.735 152.500 162.065 ;
        RECT 152.670 162.355 152.840 163.195 ;
        RECT 153.020 163.165 153.335 163.665 ;
        RECT 153.565 162.935 153.905 163.495 ;
        RECT 153.010 162.560 153.905 162.935 ;
        RECT 154.075 162.655 154.245 163.665 ;
        RECT 153.715 162.355 153.905 162.560 ;
        RECT 154.415 162.605 154.745 163.450 ;
        RECT 154.415 162.525 154.805 162.605 ;
        RECT 154.590 162.475 154.805 162.525 ;
        RECT 152.670 162.025 153.545 162.355 ;
        RECT 153.715 162.025 154.465 162.355 ;
        RECT 152.670 161.565 152.840 162.025 ;
        RECT 153.715 161.855 153.915 162.025 ;
        RECT 154.635 161.895 154.805 162.475 ;
        RECT 154.975 162.575 156.185 163.665 ;
        RECT 154.975 162.035 155.495 162.575 ;
        RECT 154.580 161.855 154.805 161.895 ;
        RECT 155.665 161.865 156.185 162.405 ;
        RECT 151.480 161.395 151.885 161.565 ;
        RECT 152.055 161.395 152.840 161.565 ;
        RECT 153.115 161.115 153.325 161.645 ;
        RECT 153.585 161.330 153.915 161.855 ;
        RECT 154.425 161.770 154.805 161.855 ;
        RECT 154.085 161.115 154.255 161.725 ;
        RECT 154.425 161.335 154.755 161.770 ;
        RECT 154.975 161.115 156.185 161.865 ;
        RECT 70.710 160.945 156.270 161.115 ;
        RECT 70.795 160.195 72.005 160.945 ;
        RECT 70.795 159.655 71.315 160.195 ;
        RECT 72.175 160.175 75.685 160.945 ;
        RECT 75.860 160.415 76.150 160.765 ;
        RECT 76.345 160.585 76.675 160.945 ;
        RECT 76.845 160.415 77.075 160.720 ;
        RECT 75.860 160.245 77.075 160.415 ;
        RECT 71.485 159.485 72.005 160.025 ;
        RECT 72.175 159.655 73.825 160.175 ;
        RECT 77.265 160.075 77.435 160.640 ;
        RECT 73.995 159.485 75.685 160.005 ;
        RECT 75.920 159.925 76.180 160.035 ;
        RECT 75.915 159.755 76.180 159.925 ;
        RECT 75.920 159.705 76.180 159.755 ;
        RECT 76.360 159.705 76.745 160.035 ;
        RECT 76.915 159.905 77.435 160.075 ;
        RECT 77.695 160.205 78.160 160.750 ;
        RECT 70.795 158.395 72.005 159.485 ;
        RECT 72.175 158.395 75.685 159.485 ;
        RECT 75.860 158.395 76.180 159.535 ;
        RECT 76.360 158.655 76.555 159.705 ;
        RECT 76.915 159.525 77.085 159.905 ;
        RECT 76.735 159.245 77.085 159.525 ;
        RECT 77.275 159.375 77.520 159.735 ;
        RECT 77.695 159.245 77.865 160.205 ;
        RECT 78.665 160.125 78.835 160.945 ;
        RECT 79.005 160.295 79.335 160.775 ;
        RECT 79.505 160.555 79.855 160.945 ;
        RECT 80.025 160.375 80.255 160.775 ;
        RECT 79.745 160.295 80.255 160.375 ;
        RECT 79.005 160.205 80.255 160.295 ;
        RECT 80.425 160.205 80.745 160.685 ;
        RECT 79.005 160.125 79.915 160.205 ;
        RECT 78.035 159.585 78.280 160.035 ;
        RECT 78.540 159.755 79.235 159.955 ;
        RECT 79.405 159.785 80.005 159.955 ;
        RECT 79.405 159.585 79.575 159.785 ;
        RECT 80.235 159.615 80.405 160.035 ;
        RECT 78.035 159.415 79.575 159.585 ;
        RECT 79.745 159.445 80.405 159.615 ;
        RECT 79.745 159.245 79.915 159.445 ;
        RECT 80.575 159.275 80.745 160.205 ;
        RECT 76.735 158.565 77.065 159.245 ;
        RECT 77.265 158.395 77.520 159.195 ;
        RECT 77.695 159.075 79.915 159.245 ;
        RECT 80.085 159.075 80.745 159.275 ;
        RECT 80.950 160.205 81.565 160.775 ;
        RECT 81.735 160.435 81.950 160.945 ;
        RECT 82.180 160.435 82.460 160.765 ;
        RECT 82.640 160.435 82.880 160.945 ;
        RECT 80.950 159.185 81.265 160.205 ;
        RECT 81.435 159.535 81.605 160.035 ;
        RECT 81.855 159.705 82.120 160.265 ;
        RECT 82.290 159.535 82.460 160.435 ;
        RECT 83.305 160.395 83.475 160.775 ;
        RECT 83.655 160.565 83.985 160.945 ;
        RECT 82.630 159.705 82.985 160.265 ;
        RECT 83.305 160.225 83.970 160.395 ;
        RECT 84.165 160.270 84.425 160.775 ;
        RECT 83.235 159.675 83.575 160.045 ;
        RECT 83.800 159.970 83.970 160.225 ;
        RECT 83.800 159.640 84.075 159.970 ;
        RECT 81.435 159.365 82.860 159.535 ;
        RECT 83.800 159.495 83.970 159.640 ;
        RECT 77.695 158.395 77.995 158.905 ;
        RECT 78.165 158.565 78.495 159.075 ;
        RECT 80.085 158.905 80.255 159.075 ;
        RECT 78.665 158.395 79.295 158.905 ;
        RECT 79.875 158.735 80.255 158.905 ;
        RECT 80.425 158.395 80.725 158.905 ;
        RECT 80.950 158.565 81.485 159.185 ;
        RECT 81.655 158.395 81.985 159.195 ;
        RECT 82.470 159.190 82.860 159.365 ;
        RECT 83.295 159.325 83.970 159.495 ;
        RECT 84.245 159.470 84.425 160.270 ;
        RECT 84.595 160.175 88.105 160.945 ;
        RECT 88.365 160.395 88.535 160.775 ;
        RECT 88.715 160.565 89.045 160.945 ;
        RECT 88.365 160.225 89.030 160.395 ;
        RECT 89.225 160.270 89.485 160.775 ;
        RECT 84.595 159.655 86.245 160.175 ;
        RECT 86.415 159.485 88.105 160.005 ;
        RECT 88.295 159.675 88.635 160.045 ;
        RECT 88.860 159.970 89.030 160.225 ;
        RECT 88.860 159.640 89.135 159.970 ;
        RECT 88.860 159.495 89.030 159.640 ;
        RECT 83.295 158.565 83.475 159.325 ;
        RECT 83.655 158.395 83.985 159.155 ;
        RECT 84.155 158.565 84.425 159.470 ;
        RECT 84.595 158.395 88.105 159.485 ;
        RECT 88.355 159.325 89.030 159.495 ;
        RECT 89.305 159.470 89.485 160.270 ;
        RECT 89.745 160.395 89.915 160.775 ;
        RECT 90.095 160.565 90.425 160.945 ;
        RECT 89.745 160.225 90.410 160.395 ;
        RECT 90.605 160.270 90.865 160.775 ;
        RECT 91.035 160.445 91.375 160.945 ;
        RECT 89.675 159.675 90.015 160.045 ;
        RECT 90.240 159.970 90.410 160.225 ;
        RECT 90.240 159.640 90.515 159.970 ;
        RECT 90.240 159.495 90.410 159.640 ;
        RECT 88.355 158.565 88.535 159.325 ;
        RECT 88.715 158.395 89.045 159.155 ;
        RECT 89.215 158.565 89.485 159.470 ;
        RECT 89.735 159.325 90.410 159.495 ;
        RECT 90.685 159.470 90.865 160.270 ;
        RECT 91.035 159.705 91.375 160.275 ;
        RECT 91.545 160.035 91.790 160.725 ;
        RECT 91.985 160.445 92.315 160.945 ;
        RECT 92.515 160.375 92.685 160.725 ;
        RECT 92.860 160.545 93.190 160.945 ;
        RECT 93.360 160.375 93.530 160.725 ;
        RECT 93.700 160.545 94.080 160.945 ;
        RECT 92.515 160.205 94.100 160.375 ;
        RECT 94.270 160.270 94.545 160.615 ;
        RECT 93.930 160.035 94.100 160.205 ;
        RECT 91.545 159.705 92.200 160.035 ;
        RECT 89.735 158.565 89.915 159.325 ;
        RECT 90.095 158.395 90.425 159.155 ;
        RECT 90.595 158.565 90.865 159.470 ;
        RECT 91.035 158.395 91.375 159.470 ;
        RECT 91.545 159.110 91.785 159.705 ;
        RECT 91.980 159.245 92.300 159.535 ;
        RECT 92.470 159.415 93.210 160.035 ;
        RECT 93.380 159.705 93.760 160.035 ;
        RECT 93.930 159.705 94.205 160.035 ;
        RECT 93.930 159.535 94.100 159.705 ;
        RECT 94.375 159.535 94.545 160.270 ;
        RECT 94.805 160.395 94.975 160.775 ;
        RECT 95.155 160.565 95.485 160.945 ;
        RECT 94.805 160.225 95.470 160.395 ;
        RECT 95.665 160.270 95.925 160.775 ;
        RECT 94.735 159.675 95.075 160.045 ;
        RECT 95.300 159.970 95.470 160.225 ;
        RECT 93.440 159.365 94.100 159.535 ;
        RECT 93.440 159.245 93.610 159.365 ;
        RECT 91.980 159.075 93.610 159.245 ;
        RECT 91.560 158.615 93.610 158.905 ;
        RECT 93.780 158.395 94.060 159.195 ;
        RECT 94.270 158.565 94.545 159.535 ;
        RECT 95.300 159.640 95.575 159.970 ;
        RECT 95.300 159.495 95.470 159.640 ;
        RECT 94.795 159.325 95.470 159.495 ;
        RECT 95.745 159.470 95.925 160.270 ;
        RECT 96.555 160.220 96.845 160.945 ;
        RECT 97.475 160.565 98.365 160.735 ;
        RECT 97.475 160.010 98.025 160.395 ;
        RECT 98.195 159.840 98.365 160.565 ;
        RECT 97.475 159.770 98.365 159.840 ;
        RECT 98.535 160.240 98.755 160.725 ;
        RECT 98.925 160.405 99.175 160.945 ;
        RECT 99.345 160.295 99.605 160.775 ;
        RECT 99.775 160.565 100.665 160.735 ;
        RECT 98.535 159.815 98.865 160.240 ;
        RECT 97.475 159.745 98.370 159.770 ;
        RECT 97.475 159.730 98.380 159.745 ;
        RECT 97.475 159.715 98.385 159.730 ;
        RECT 97.475 159.710 98.395 159.715 ;
        RECT 97.475 159.700 98.400 159.710 ;
        RECT 97.475 159.690 98.405 159.700 ;
        RECT 97.475 159.685 98.415 159.690 ;
        RECT 97.475 159.675 98.425 159.685 ;
        RECT 97.475 159.670 98.435 159.675 ;
        RECT 94.795 158.565 94.975 159.325 ;
        RECT 95.155 158.395 95.485 159.155 ;
        RECT 95.655 158.565 95.925 159.470 ;
        RECT 96.555 158.395 96.845 159.560 ;
        RECT 97.475 159.220 97.735 159.670 ;
        RECT 98.100 159.665 98.435 159.670 ;
        RECT 98.100 159.660 98.450 159.665 ;
        RECT 98.100 159.650 98.465 159.660 ;
        RECT 98.100 159.645 98.490 159.650 ;
        RECT 99.035 159.645 99.265 160.040 ;
        RECT 98.100 159.640 99.265 159.645 ;
        RECT 98.130 159.605 99.265 159.640 ;
        RECT 98.165 159.580 99.265 159.605 ;
        RECT 98.195 159.550 99.265 159.580 ;
        RECT 98.215 159.520 99.265 159.550 ;
        RECT 98.235 159.490 99.265 159.520 ;
        RECT 98.305 159.480 99.265 159.490 ;
        RECT 98.330 159.470 99.265 159.480 ;
        RECT 98.350 159.455 99.265 159.470 ;
        RECT 98.370 159.440 99.265 159.455 ;
        RECT 98.375 159.430 99.160 159.440 ;
        RECT 98.390 159.395 99.160 159.430 ;
        RECT 97.905 159.075 98.235 159.320 ;
        RECT 98.405 159.145 99.160 159.395 ;
        RECT 99.435 159.265 99.605 160.295 ;
        RECT 99.775 160.010 100.325 160.395 ;
        RECT 100.495 159.840 100.665 160.565 ;
        RECT 97.905 159.050 98.090 159.075 ;
        RECT 97.475 158.950 98.090 159.050 ;
        RECT 97.475 158.395 98.080 158.950 ;
        RECT 98.255 158.565 98.735 158.905 ;
        RECT 98.905 158.395 99.160 158.940 ;
        RECT 99.330 158.565 99.605 159.265 ;
        RECT 99.775 159.770 100.665 159.840 ;
        RECT 100.835 160.265 101.055 160.725 ;
        RECT 101.225 160.405 101.475 160.945 ;
        RECT 101.645 160.295 101.905 160.775 ;
        RECT 100.835 160.240 101.085 160.265 ;
        RECT 100.835 159.815 101.165 160.240 ;
        RECT 99.775 159.745 100.670 159.770 ;
        RECT 99.775 159.730 100.680 159.745 ;
        RECT 99.775 159.715 100.685 159.730 ;
        RECT 99.775 159.710 100.695 159.715 ;
        RECT 99.775 159.700 100.700 159.710 ;
        RECT 99.775 159.690 100.705 159.700 ;
        RECT 99.775 159.685 100.715 159.690 ;
        RECT 99.775 159.675 100.725 159.685 ;
        RECT 99.775 159.670 100.735 159.675 ;
        RECT 99.775 159.220 100.035 159.670 ;
        RECT 100.400 159.665 100.735 159.670 ;
        RECT 100.400 159.660 100.750 159.665 ;
        RECT 100.400 159.650 100.765 159.660 ;
        RECT 100.400 159.645 100.790 159.650 ;
        RECT 101.335 159.645 101.565 160.040 ;
        RECT 100.400 159.640 101.565 159.645 ;
        RECT 100.430 159.605 101.565 159.640 ;
        RECT 100.465 159.580 101.565 159.605 ;
        RECT 100.495 159.550 101.565 159.580 ;
        RECT 100.515 159.520 101.565 159.550 ;
        RECT 100.535 159.490 101.565 159.520 ;
        RECT 100.605 159.480 101.565 159.490 ;
        RECT 100.630 159.470 101.565 159.480 ;
        RECT 100.650 159.455 101.565 159.470 ;
        RECT 100.670 159.440 101.565 159.455 ;
        RECT 100.675 159.430 101.460 159.440 ;
        RECT 100.690 159.395 101.460 159.430 ;
        RECT 100.205 159.075 100.535 159.320 ;
        RECT 100.705 159.145 101.460 159.395 ;
        RECT 101.735 159.265 101.905 160.295 ;
        RECT 102.075 160.175 105.585 160.945 ;
        RECT 105.755 160.205 106.015 160.775 ;
        RECT 106.185 160.545 106.570 160.945 ;
        RECT 106.740 160.375 106.995 160.775 ;
        RECT 106.185 160.205 106.995 160.375 ;
        RECT 107.185 160.205 107.430 160.775 ;
        RECT 107.600 160.545 107.985 160.945 ;
        RECT 108.155 160.375 108.410 160.775 ;
        RECT 107.600 160.205 108.410 160.375 ;
        RECT 108.600 160.205 109.025 160.775 ;
        RECT 109.195 160.545 109.580 160.945 ;
        RECT 109.750 160.375 110.185 160.775 ;
        RECT 110.355 160.400 115.700 160.945 ;
        RECT 109.195 160.205 110.185 160.375 ;
        RECT 102.075 159.655 103.725 160.175 ;
        RECT 103.895 159.485 105.585 160.005 ;
        RECT 100.205 159.050 100.390 159.075 ;
        RECT 99.775 158.950 100.390 159.050 ;
        RECT 99.775 158.395 100.380 158.950 ;
        RECT 100.555 158.565 101.035 158.905 ;
        RECT 101.205 158.395 101.460 158.940 ;
        RECT 101.630 158.565 101.905 159.265 ;
        RECT 102.075 158.395 105.585 159.485 ;
        RECT 105.755 159.535 105.940 160.205 ;
        RECT 106.185 160.035 106.535 160.205 ;
        RECT 107.185 160.035 107.355 160.205 ;
        RECT 107.600 160.035 107.950 160.205 ;
        RECT 108.600 160.035 108.950 160.205 ;
        RECT 109.195 160.035 109.530 160.205 ;
        RECT 106.110 159.705 106.535 160.035 ;
        RECT 105.755 158.565 106.015 159.535 ;
        RECT 106.185 159.185 106.535 159.705 ;
        RECT 106.705 159.535 107.355 160.035 ;
        RECT 107.525 159.705 107.950 160.035 ;
        RECT 106.705 159.355 107.430 159.535 ;
        RECT 106.185 158.990 106.995 159.185 ;
        RECT 106.185 158.395 106.570 158.820 ;
        RECT 106.740 158.565 106.995 158.990 ;
        RECT 107.185 158.565 107.430 159.355 ;
        RECT 107.600 159.185 107.950 159.705 ;
        RECT 108.120 159.535 108.950 160.035 ;
        RECT 109.120 159.705 109.530 160.035 ;
        RECT 108.120 159.355 109.025 159.535 ;
        RECT 107.600 158.990 108.430 159.185 ;
        RECT 107.600 158.395 107.985 158.820 ;
        RECT 108.155 158.565 108.430 158.990 ;
        RECT 108.600 158.565 109.025 159.355 ;
        RECT 109.195 159.160 109.530 159.705 ;
        RECT 109.700 159.330 110.185 160.035 ;
        RECT 111.940 159.570 112.280 160.400 ;
        RECT 115.875 160.175 119.385 160.945 ;
        RECT 109.195 158.990 110.185 159.160 ;
        RECT 109.195 158.395 109.580 158.820 ;
        RECT 109.750 158.565 110.185 158.990 ;
        RECT 113.760 158.830 114.110 160.080 ;
        RECT 115.875 159.655 117.525 160.175 ;
        RECT 119.555 160.145 119.865 160.945 ;
        RECT 120.070 160.145 120.765 160.775 ;
        RECT 120.935 160.270 121.195 160.775 ;
        RECT 121.375 160.565 121.705 160.945 ;
        RECT 121.885 160.395 122.055 160.775 ;
        RECT 117.695 159.485 119.385 160.005 ;
        RECT 119.565 159.705 119.900 159.975 ;
        RECT 120.070 159.545 120.240 160.145 ;
        RECT 120.410 159.705 120.745 159.955 ;
        RECT 110.355 158.395 115.700 158.830 ;
        RECT 115.875 158.395 119.385 159.485 ;
        RECT 119.555 158.395 119.835 159.535 ;
        RECT 120.005 158.565 120.335 159.545 ;
        RECT 120.505 158.395 120.765 159.535 ;
        RECT 120.935 159.470 121.115 160.270 ;
        RECT 121.390 160.225 122.055 160.395 ;
        RECT 121.390 159.970 121.560 160.225 ;
        RECT 122.315 160.220 122.605 160.945 ;
        RECT 123.695 160.315 124.035 160.775 ;
        RECT 124.205 160.485 124.375 160.945 ;
        RECT 125.005 160.510 125.365 160.775 ;
        RECT 125.010 160.505 125.365 160.510 ;
        RECT 125.015 160.495 125.365 160.505 ;
        RECT 125.020 160.490 125.365 160.495 ;
        RECT 125.025 160.480 125.365 160.490 ;
        RECT 125.605 160.485 125.775 160.945 ;
        RECT 125.030 160.475 125.365 160.480 ;
        RECT 125.040 160.465 125.365 160.475 ;
        RECT 125.050 160.455 125.365 160.465 ;
        RECT 124.545 160.315 124.875 160.395 ;
        RECT 123.695 160.125 124.875 160.315 ;
        RECT 125.065 160.315 125.365 160.455 ;
        RECT 125.065 160.125 125.775 160.315 ;
        RECT 121.285 159.640 121.560 159.970 ;
        RECT 121.785 159.675 122.125 160.045 ;
        RECT 123.695 159.755 124.025 159.955 ;
        RECT 124.335 159.935 124.665 159.955 ;
        RECT 124.215 159.755 124.665 159.935 ;
        RECT 121.390 159.495 121.560 159.640 ;
        RECT 120.935 158.565 121.205 159.470 ;
        RECT 121.390 159.325 122.065 159.495 ;
        RECT 121.375 158.395 121.705 159.155 ;
        RECT 121.885 158.565 122.065 159.325 ;
        RECT 122.315 158.395 122.605 159.560 ;
        RECT 123.695 159.415 123.925 159.755 ;
        RECT 123.705 158.395 124.035 159.115 ;
        RECT 124.215 158.640 124.430 159.755 ;
        RECT 124.835 159.725 125.305 159.955 ;
        RECT 125.490 159.555 125.775 160.125 ;
        RECT 125.945 160.000 126.285 160.775 ;
        RECT 124.625 159.340 125.775 159.555 ;
        RECT 124.625 158.565 124.955 159.340 ;
        RECT 125.125 158.395 125.835 159.170 ;
        RECT 126.005 158.565 126.285 160.000 ;
        RECT 126.455 160.125 127.140 160.765 ;
        RECT 127.310 160.125 127.480 160.945 ;
        RECT 127.650 160.295 127.980 160.760 ;
        RECT 128.150 160.475 128.320 160.945 ;
        RECT 128.580 160.555 129.765 160.725 ;
        RECT 129.935 160.385 130.265 160.775 ;
        RECT 128.965 160.295 129.350 160.385 ;
        RECT 127.650 160.125 129.350 160.295 ;
        RECT 129.755 160.205 130.265 160.385 ;
        RECT 130.685 160.395 130.855 160.775 ;
        RECT 131.035 160.565 131.365 160.945 ;
        RECT 130.685 160.225 131.350 160.395 ;
        RECT 131.545 160.270 131.805 160.775 ;
        RECT 126.455 159.155 126.705 160.125 ;
        RECT 126.875 159.745 127.210 159.955 ;
        RECT 127.380 159.745 127.830 159.955 ;
        RECT 128.020 159.745 128.505 159.955 ;
        RECT 127.040 159.575 127.210 159.745 ;
        RECT 128.130 159.585 128.505 159.745 ;
        RECT 128.695 159.705 129.075 159.955 ;
        RECT 129.255 159.745 129.585 159.955 ;
        RECT 127.040 159.405 127.960 159.575 ;
        RECT 126.455 158.565 127.120 159.155 ;
        RECT 127.290 158.395 127.620 159.235 ;
        RECT 127.790 159.155 127.960 159.405 ;
        RECT 128.130 159.415 128.525 159.585 ;
        RECT 128.130 159.325 128.505 159.415 ;
        RECT 128.695 159.325 129.015 159.705 ;
        RECT 129.755 159.575 129.925 160.205 ;
        RECT 130.095 159.745 130.425 160.035 ;
        RECT 130.615 159.675 130.955 160.045 ;
        RECT 131.180 159.970 131.350 160.225 ;
        RECT 131.180 159.640 131.455 159.970 ;
        RECT 129.185 159.405 130.270 159.575 ;
        RECT 131.180 159.495 131.350 159.640 ;
        RECT 129.185 159.155 129.355 159.405 ;
        RECT 127.790 158.985 129.355 159.155 ;
        RECT 128.130 158.565 128.935 158.985 ;
        RECT 129.525 158.395 129.775 159.235 ;
        RECT 129.970 158.565 130.270 159.405 ;
        RECT 130.675 159.325 131.350 159.495 ;
        RECT 131.625 159.470 131.805 160.270 ;
        RECT 131.975 160.175 134.565 160.945 ;
        RECT 135.355 160.385 135.685 160.775 ;
        RECT 135.855 160.555 137.040 160.725 ;
        RECT 137.300 160.475 137.470 160.945 ;
        RECT 135.355 160.205 135.865 160.385 ;
        RECT 131.975 159.655 133.185 160.175 ;
        RECT 133.355 159.485 134.565 160.005 ;
        RECT 135.195 159.745 135.525 160.035 ;
        RECT 135.695 159.575 135.865 160.205 ;
        RECT 136.270 160.295 136.655 160.385 ;
        RECT 137.640 160.295 137.970 160.760 ;
        RECT 136.270 160.125 137.970 160.295 ;
        RECT 138.140 160.125 138.310 160.945 ;
        RECT 138.480 160.125 139.165 160.765 ;
        RECT 139.495 160.385 139.825 160.775 ;
        RECT 139.995 160.555 141.180 160.725 ;
        RECT 141.440 160.475 141.610 160.945 ;
        RECT 139.495 160.205 140.005 160.385 ;
        RECT 136.035 159.745 136.365 159.955 ;
        RECT 136.545 159.705 136.925 159.955 ;
        RECT 137.115 159.925 137.600 159.955 ;
        RECT 137.095 159.755 137.600 159.925 ;
        RECT 130.675 158.565 130.855 159.325 ;
        RECT 131.035 158.395 131.365 159.155 ;
        RECT 131.535 158.565 131.805 159.470 ;
        RECT 131.975 158.395 134.565 159.485 ;
        RECT 135.350 159.405 136.435 159.575 ;
        RECT 135.350 158.565 135.650 159.405 ;
        RECT 135.845 158.395 136.095 159.235 ;
        RECT 136.265 159.155 136.435 159.405 ;
        RECT 136.605 159.325 136.925 159.705 ;
        RECT 137.115 159.745 137.600 159.755 ;
        RECT 137.790 159.745 138.240 159.955 ;
        RECT 138.410 159.745 138.745 159.955 ;
        RECT 137.115 159.325 137.490 159.745 ;
        RECT 138.410 159.575 138.580 159.745 ;
        RECT 137.660 159.405 138.580 159.575 ;
        RECT 137.660 159.155 137.830 159.405 ;
        RECT 136.265 158.985 137.830 159.155 ;
        RECT 136.685 158.565 137.490 158.985 ;
        RECT 138.000 158.395 138.330 159.235 ;
        RECT 138.915 159.155 139.165 160.125 ;
        RECT 139.335 159.745 139.665 160.035 ;
        RECT 139.835 159.575 140.005 160.205 ;
        RECT 140.410 160.295 140.795 160.385 ;
        RECT 141.780 160.295 142.110 160.760 ;
        RECT 140.410 160.125 142.110 160.295 ;
        RECT 142.280 160.125 142.450 160.945 ;
        RECT 142.620 160.125 143.305 160.765 ;
        RECT 143.935 160.145 144.630 160.775 ;
        RECT 144.835 160.145 145.145 160.945 ;
        RECT 145.480 160.435 145.720 160.945 ;
        RECT 145.900 160.435 146.180 160.765 ;
        RECT 146.410 160.435 146.625 160.945 ;
        RECT 140.175 159.745 140.505 159.955 ;
        RECT 140.685 159.705 141.065 159.955 ;
        RECT 141.255 159.925 141.740 159.955 ;
        RECT 141.235 159.755 141.740 159.925 ;
        RECT 138.500 158.565 139.165 159.155 ;
        RECT 139.490 159.405 140.575 159.575 ;
        RECT 139.490 158.565 139.790 159.405 ;
        RECT 139.985 158.395 140.235 159.235 ;
        RECT 140.405 159.155 140.575 159.405 ;
        RECT 140.745 159.325 141.065 159.705 ;
        RECT 141.255 159.745 141.740 159.755 ;
        RECT 141.930 159.745 142.380 159.955 ;
        RECT 142.550 159.745 142.885 159.955 ;
        RECT 141.255 159.325 141.630 159.745 ;
        RECT 142.550 159.575 142.720 159.745 ;
        RECT 141.800 159.405 142.720 159.575 ;
        RECT 141.800 159.155 141.970 159.405 ;
        RECT 140.405 158.985 141.970 159.155 ;
        RECT 140.825 158.565 141.630 158.985 ;
        RECT 142.140 158.395 142.470 159.235 ;
        RECT 143.055 159.155 143.305 160.125 ;
        RECT 143.955 159.705 144.290 159.955 ;
        RECT 144.460 159.545 144.630 160.145 ;
        RECT 144.800 159.705 145.135 159.975 ;
        RECT 145.375 159.705 145.730 160.265 ;
        RECT 142.640 158.565 143.305 159.155 ;
        RECT 143.935 158.395 144.195 159.535 ;
        RECT 144.365 158.565 144.695 159.545 ;
        RECT 145.900 159.535 146.070 160.435 ;
        RECT 146.240 159.705 146.505 160.265 ;
        RECT 146.795 160.205 147.410 160.775 ;
        RECT 148.075 160.220 148.365 160.945 ;
        RECT 148.535 160.565 149.425 160.735 ;
        RECT 146.755 159.535 146.925 160.035 ;
        RECT 144.865 158.395 145.145 159.535 ;
        RECT 145.500 159.365 146.925 159.535 ;
        RECT 145.500 159.190 145.890 159.365 ;
        RECT 146.375 158.395 146.705 159.195 ;
        RECT 147.095 159.185 147.410 160.205 ;
        RECT 148.535 160.010 149.085 160.395 ;
        RECT 149.255 159.840 149.425 160.565 ;
        RECT 148.535 159.770 149.425 159.840 ;
        RECT 149.595 160.240 149.815 160.725 ;
        RECT 149.985 160.405 150.235 160.945 ;
        RECT 150.405 160.295 150.665 160.775 ;
        RECT 149.595 159.815 149.925 160.240 ;
        RECT 148.535 159.745 149.430 159.770 ;
        RECT 148.535 159.730 149.440 159.745 ;
        RECT 148.535 159.715 149.445 159.730 ;
        RECT 148.535 159.710 149.455 159.715 ;
        RECT 148.535 159.700 149.460 159.710 ;
        RECT 148.535 159.690 149.465 159.700 ;
        RECT 148.535 159.685 149.475 159.690 ;
        RECT 148.535 159.675 149.485 159.685 ;
        RECT 148.535 159.670 149.495 159.675 ;
        RECT 146.875 158.565 147.410 159.185 ;
        RECT 148.075 158.395 148.365 159.560 ;
        RECT 148.535 159.220 148.795 159.670 ;
        RECT 149.160 159.665 149.495 159.670 ;
        RECT 149.160 159.660 149.510 159.665 ;
        RECT 149.160 159.650 149.525 159.660 ;
        RECT 149.160 159.645 149.550 159.650 ;
        RECT 150.095 159.645 150.325 160.040 ;
        RECT 149.160 159.640 150.325 159.645 ;
        RECT 149.190 159.605 150.325 159.640 ;
        RECT 149.225 159.580 150.325 159.605 ;
        RECT 149.255 159.550 150.325 159.580 ;
        RECT 149.275 159.520 150.325 159.550 ;
        RECT 149.295 159.490 150.325 159.520 ;
        RECT 149.365 159.480 150.325 159.490 ;
        RECT 149.390 159.470 150.325 159.480 ;
        RECT 149.410 159.455 150.325 159.470 ;
        RECT 149.430 159.440 150.325 159.455 ;
        RECT 149.435 159.430 150.220 159.440 ;
        RECT 149.450 159.395 150.220 159.430 ;
        RECT 148.965 159.075 149.295 159.320 ;
        RECT 149.465 159.145 150.220 159.395 ;
        RECT 150.495 159.265 150.665 160.295 ;
        RECT 148.965 159.050 149.150 159.075 ;
        RECT 148.535 158.950 149.150 159.050 ;
        RECT 148.535 158.395 149.140 158.950 ;
        RECT 149.315 158.565 149.795 158.905 ;
        RECT 149.965 158.395 150.220 158.940 ;
        RECT 150.390 158.565 150.665 159.265 ;
        RECT 150.835 160.270 151.095 160.775 ;
        RECT 151.275 160.565 151.605 160.945 ;
        RECT 151.785 160.395 151.955 160.775 ;
        RECT 150.835 159.470 151.005 160.270 ;
        RECT 151.290 160.225 151.955 160.395 ;
        RECT 151.290 159.970 151.460 160.225 ;
        RECT 152.215 160.175 154.805 160.945 ;
        RECT 154.975 160.195 156.185 160.945 ;
        RECT 151.175 159.640 151.460 159.970 ;
        RECT 151.695 159.675 152.025 160.045 ;
        RECT 152.215 159.655 153.425 160.175 ;
        RECT 151.290 159.495 151.460 159.640 ;
        RECT 150.835 158.565 151.105 159.470 ;
        RECT 151.290 159.325 151.955 159.495 ;
        RECT 153.595 159.485 154.805 160.005 ;
        RECT 151.275 158.395 151.605 159.155 ;
        RECT 151.785 158.565 151.955 159.325 ;
        RECT 152.215 158.395 154.805 159.485 ;
        RECT 154.975 159.485 155.495 160.025 ;
        RECT 155.665 159.655 156.185 160.195 ;
        RECT 154.975 158.395 156.185 159.485 ;
        RECT 70.710 158.225 156.270 158.395 ;
        RECT 70.795 157.135 72.005 158.225 ;
        RECT 72.175 157.790 77.520 158.225 ;
        RECT 70.795 156.425 71.315 156.965 ;
        RECT 71.485 156.595 72.005 157.135 ;
        RECT 70.795 155.675 72.005 156.425 ;
        RECT 73.760 156.220 74.100 157.050 ;
        RECT 75.580 156.540 75.930 157.790 ;
        RECT 77.695 157.085 77.955 158.225 ;
        RECT 78.125 157.075 78.455 158.055 ;
        RECT 78.625 157.085 78.905 158.225 ;
        RECT 79.075 157.085 79.335 158.225 ;
        RECT 79.505 157.075 79.835 158.055 ;
        RECT 80.005 157.085 80.285 158.225 ;
        RECT 80.655 157.555 80.935 158.225 ;
        RECT 81.105 157.335 81.405 157.885 ;
        RECT 81.605 157.505 81.935 158.225 ;
        RECT 82.125 157.505 82.585 158.055 ;
        RECT 77.715 156.665 78.050 156.915 ;
        RECT 78.220 156.475 78.390 157.075 ;
        RECT 78.560 156.645 78.895 156.915 ;
        RECT 79.095 156.665 79.430 156.915 ;
        RECT 79.600 156.475 79.770 157.075 ;
        RECT 80.470 156.915 80.735 157.275 ;
        RECT 81.105 157.165 82.045 157.335 ;
        RECT 81.875 156.915 82.045 157.165 ;
        RECT 79.940 156.645 80.275 156.915 ;
        RECT 80.470 156.665 81.145 156.915 ;
        RECT 81.365 156.665 81.705 156.915 ;
        RECT 81.875 156.585 82.165 156.915 ;
        RECT 81.875 156.495 82.045 156.585 ;
        RECT 72.175 155.675 77.520 156.220 ;
        RECT 77.695 155.845 78.390 156.475 ;
        RECT 78.595 155.675 78.905 156.475 ;
        RECT 79.075 155.845 79.770 156.475 ;
        RECT 79.975 155.675 80.285 156.475 ;
        RECT 80.655 156.305 82.045 156.495 ;
        RECT 80.655 155.945 80.985 156.305 ;
        RECT 82.335 156.135 82.585 157.505 ;
        RECT 83.675 157.060 83.965 158.225 ;
        RECT 84.135 157.135 85.805 158.225 ;
        RECT 86.445 157.505 86.775 158.225 ;
        RECT 84.135 156.445 84.885 156.965 ;
        RECT 85.055 156.615 85.805 157.135 ;
        RECT 86.435 156.865 86.665 157.205 ;
        RECT 86.955 156.865 87.170 157.980 ;
        RECT 87.365 157.280 87.695 158.055 ;
        RECT 87.865 157.450 88.575 158.225 ;
        RECT 87.365 157.065 88.515 157.280 ;
        RECT 86.435 156.665 86.765 156.865 ;
        RECT 86.955 156.685 87.405 156.865 ;
        RECT 87.075 156.665 87.405 156.685 ;
        RECT 87.575 156.665 88.045 156.895 ;
        RECT 88.230 156.495 88.515 157.065 ;
        RECT 88.745 156.620 89.025 158.055 ;
        RECT 89.200 157.425 89.515 158.225 ;
        RECT 89.780 157.885 90.860 158.040 ;
        RECT 89.715 157.870 90.860 157.885 ;
        RECT 89.715 157.715 89.950 157.870 ;
        RECT 89.780 157.255 89.950 157.715 ;
        RECT 81.605 155.675 81.855 156.135 ;
        RECT 82.025 155.845 82.585 156.135 ;
        RECT 83.675 155.675 83.965 156.400 ;
        RECT 84.135 155.675 85.805 156.445 ;
        RECT 86.435 156.305 87.615 156.495 ;
        RECT 86.435 155.845 86.775 156.305 ;
        RECT 87.285 156.225 87.615 156.305 ;
        RECT 87.805 156.305 88.515 156.495 ;
        RECT 87.805 156.165 88.105 156.305 ;
        RECT 87.790 156.155 88.105 156.165 ;
        RECT 87.780 156.145 88.105 156.155 ;
        RECT 87.770 156.140 88.105 156.145 ;
        RECT 86.945 155.675 87.115 156.135 ;
        RECT 87.765 156.130 88.105 156.140 ;
        RECT 87.760 156.125 88.105 156.130 ;
        RECT 87.755 156.115 88.105 156.125 ;
        RECT 87.750 156.110 88.105 156.115 ;
        RECT 87.745 155.845 88.105 156.110 ;
        RECT 88.345 155.675 88.515 156.135 ;
        RECT 88.685 155.845 89.025 156.620 ;
        RECT 89.195 156.245 89.465 157.255 ;
        RECT 89.635 157.085 89.950 157.255 ;
        RECT 89.635 156.415 89.805 157.085 ;
        RECT 90.120 156.915 90.355 157.595 ;
        RECT 90.525 157.085 90.860 157.870 ;
        RECT 91.045 157.255 91.375 158.040 ;
        RECT 91.045 157.085 91.725 157.255 ;
        RECT 91.905 157.085 92.235 158.225 ;
        RECT 92.955 157.295 93.135 158.055 ;
        RECT 93.315 157.465 93.645 158.225 ;
        RECT 92.955 157.125 93.630 157.295 ;
        RECT 93.815 157.150 94.085 158.055 ;
        RECT 89.975 156.585 90.355 156.915 ;
        RECT 90.525 156.585 90.860 156.915 ;
        RECT 91.035 156.665 91.385 156.915 ;
        RECT 91.555 156.485 91.725 157.085 ;
        RECT 93.460 156.980 93.630 157.125 ;
        RECT 91.895 156.665 92.245 156.915 ;
        RECT 92.895 156.575 93.235 156.945 ;
        RECT 93.460 156.650 93.735 156.980 ;
        RECT 89.635 156.245 90.860 156.415 ;
        RECT 89.265 155.675 89.595 156.075 ;
        RECT 89.765 155.975 89.935 156.245 ;
        RECT 90.105 155.675 90.435 156.075 ;
        RECT 90.605 155.975 90.860 156.245 ;
        RECT 91.055 155.675 91.295 156.485 ;
        RECT 91.465 155.845 91.795 156.485 ;
        RECT 91.965 155.675 92.235 156.485 ;
        RECT 93.460 156.395 93.630 156.650 ;
        RECT 92.965 156.225 93.630 156.395 ;
        RECT 93.905 156.350 94.085 157.150 ;
        RECT 94.795 157.295 94.975 158.055 ;
        RECT 95.155 157.465 95.485 158.225 ;
        RECT 94.795 157.125 95.470 157.295 ;
        RECT 95.655 157.150 95.925 158.055 ;
        RECT 95.300 156.980 95.470 157.125 ;
        RECT 94.735 156.575 95.075 156.945 ;
        RECT 95.300 156.650 95.575 156.980 ;
        RECT 95.300 156.395 95.470 156.650 ;
        RECT 92.965 155.845 93.135 156.225 ;
        RECT 93.315 155.675 93.645 156.055 ;
        RECT 93.825 155.845 94.085 156.350 ;
        RECT 94.805 156.225 95.470 156.395 ;
        RECT 95.745 156.350 95.925 157.150 ;
        RECT 96.175 157.295 96.355 158.055 ;
        RECT 96.535 157.465 96.865 158.225 ;
        RECT 96.175 157.125 96.850 157.295 ;
        RECT 97.035 157.150 97.305 158.055 ;
        RECT 96.680 156.980 96.850 157.125 ;
        RECT 96.115 156.575 96.455 156.945 ;
        RECT 96.680 156.650 96.955 156.980 ;
        RECT 96.680 156.395 96.850 156.650 ;
        RECT 94.805 155.845 94.975 156.225 ;
        RECT 95.155 155.675 95.485 156.055 ;
        RECT 95.665 155.845 95.925 156.350 ;
        RECT 96.185 156.225 96.850 156.395 ;
        RECT 97.125 156.350 97.305 157.150 ;
        RECT 97.555 157.295 97.735 158.055 ;
        RECT 97.915 157.465 98.245 158.225 ;
        RECT 97.555 157.125 98.230 157.295 ;
        RECT 98.415 157.150 98.685 158.055 ;
        RECT 98.060 156.980 98.230 157.125 ;
        RECT 97.495 156.575 97.835 156.945 ;
        RECT 98.060 156.650 98.335 156.980 ;
        RECT 98.060 156.395 98.230 156.650 ;
        RECT 96.185 155.845 96.355 156.225 ;
        RECT 96.535 155.675 96.865 156.055 ;
        RECT 97.045 155.845 97.305 156.350 ;
        RECT 97.565 156.225 98.230 156.395 ;
        RECT 98.505 156.350 98.685 157.150 ;
        RECT 99.855 157.295 100.035 158.055 ;
        RECT 100.215 157.465 100.545 158.225 ;
        RECT 99.855 157.125 100.530 157.295 ;
        RECT 100.715 157.150 100.985 158.055 ;
        RECT 101.155 157.790 106.500 158.225 ;
        RECT 100.360 156.980 100.530 157.125 ;
        RECT 99.795 156.575 100.135 156.945 ;
        RECT 100.360 156.650 100.635 156.980 ;
        RECT 100.360 156.395 100.530 156.650 ;
        RECT 97.565 155.845 97.735 156.225 ;
        RECT 97.915 155.675 98.245 156.055 ;
        RECT 98.425 155.845 98.685 156.350 ;
        RECT 99.865 156.225 100.530 156.395 ;
        RECT 100.805 156.350 100.985 157.150 ;
        RECT 99.865 155.845 100.035 156.225 ;
        RECT 100.215 155.675 100.545 156.055 ;
        RECT 100.725 155.845 100.985 156.350 ;
        RECT 102.740 156.220 103.080 157.050 ;
        RECT 104.560 156.540 104.910 157.790 ;
        RECT 106.675 157.135 109.265 158.225 ;
        RECT 106.675 156.445 107.885 156.965 ;
        RECT 108.055 156.615 109.265 157.135 ;
        RECT 109.435 157.060 109.725 158.225 ;
        RECT 109.895 157.465 110.560 158.055 ;
        RECT 109.895 156.495 110.145 157.465 ;
        RECT 110.730 157.385 111.060 158.225 ;
        RECT 111.570 157.635 112.375 158.055 ;
        RECT 111.230 157.465 112.795 157.635 ;
        RECT 111.230 157.215 111.400 157.465 ;
        RECT 110.480 157.045 111.400 157.215 ;
        RECT 110.480 156.875 110.650 157.045 ;
        RECT 111.570 156.875 111.945 157.295 ;
        RECT 110.315 156.665 110.650 156.875 ;
        RECT 110.820 156.665 111.270 156.875 ;
        RECT 111.460 156.865 111.945 156.875 ;
        RECT 112.135 156.915 112.455 157.295 ;
        RECT 112.625 157.215 112.795 157.465 ;
        RECT 112.965 157.385 113.215 158.225 ;
        RECT 113.410 157.215 113.710 158.055 ;
        RECT 114.045 157.505 114.375 158.225 ;
        RECT 112.625 157.045 113.710 157.215 ;
        RECT 111.460 156.695 111.965 156.865 ;
        RECT 111.460 156.665 111.945 156.695 ;
        RECT 112.135 156.665 112.515 156.915 ;
        RECT 112.695 156.665 113.025 156.875 ;
        RECT 101.155 155.675 106.500 156.220 ;
        RECT 106.675 155.675 109.265 156.445 ;
        RECT 109.435 155.675 109.725 156.400 ;
        RECT 109.895 155.855 110.580 156.495 ;
        RECT 110.750 155.675 110.920 156.495 ;
        RECT 111.090 156.325 112.790 156.495 ;
        RECT 111.090 155.860 111.420 156.325 ;
        RECT 112.405 156.235 112.790 156.325 ;
        RECT 113.195 156.415 113.365 157.045 ;
        RECT 113.535 156.585 113.865 156.875 ;
        RECT 114.035 156.865 114.265 157.205 ;
        RECT 114.555 156.865 114.770 157.980 ;
        RECT 114.965 157.280 115.295 158.055 ;
        RECT 115.465 157.450 116.175 158.225 ;
        RECT 114.965 157.065 116.115 157.280 ;
        RECT 114.035 156.665 114.365 156.865 ;
        RECT 114.555 156.685 115.005 156.865 ;
        RECT 114.675 156.665 115.005 156.685 ;
        RECT 115.175 156.665 115.645 156.895 ;
        RECT 115.830 156.495 116.115 157.065 ;
        RECT 116.345 156.620 116.625 158.055 ;
        RECT 117.795 157.295 117.975 158.055 ;
        RECT 118.155 157.465 118.485 158.225 ;
        RECT 117.795 157.125 118.470 157.295 ;
        RECT 118.655 157.150 118.925 158.055 ;
        RECT 118.300 156.980 118.470 157.125 ;
        RECT 113.195 156.235 113.705 156.415 ;
        RECT 111.590 155.675 111.760 156.145 ;
        RECT 112.020 155.895 113.205 156.065 ;
        RECT 113.375 155.845 113.705 156.235 ;
        RECT 114.035 156.305 115.215 156.495 ;
        RECT 114.035 155.845 114.375 156.305 ;
        RECT 114.885 156.225 115.215 156.305 ;
        RECT 115.405 156.305 116.115 156.495 ;
        RECT 115.405 156.165 115.705 156.305 ;
        RECT 115.390 156.155 115.705 156.165 ;
        RECT 115.380 156.145 115.705 156.155 ;
        RECT 115.370 156.140 115.705 156.145 ;
        RECT 114.545 155.675 114.715 156.135 ;
        RECT 115.365 156.130 115.705 156.140 ;
        RECT 115.360 156.125 115.705 156.130 ;
        RECT 115.355 156.115 115.705 156.125 ;
        RECT 115.350 156.110 115.705 156.115 ;
        RECT 115.345 155.845 115.705 156.110 ;
        RECT 115.945 155.675 116.115 156.135 ;
        RECT 116.285 155.845 116.625 156.620 ;
        RECT 117.735 156.575 118.075 156.945 ;
        RECT 118.300 156.650 118.575 156.980 ;
        RECT 118.300 156.395 118.470 156.650 ;
        RECT 117.805 156.225 118.470 156.395 ;
        RECT 118.745 156.350 118.925 157.150 ;
        RECT 119.095 157.085 119.375 158.225 ;
        RECT 119.545 157.075 119.875 158.055 ;
        RECT 120.045 157.085 120.305 158.225 ;
        RECT 120.555 157.295 120.735 158.055 ;
        RECT 120.915 157.465 121.245 158.225 ;
        RECT 120.555 157.125 121.230 157.295 ;
        RECT 121.415 157.150 121.685 158.055 ;
        RECT 119.105 156.645 119.440 156.915 ;
        RECT 119.610 156.475 119.780 157.075 ;
        RECT 121.060 156.980 121.230 157.125 ;
        RECT 119.950 156.665 120.285 156.915 ;
        RECT 120.495 156.575 120.835 156.945 ;
        RECT 121.060 156.650 121.335 156.980 ;
        RECT 117.805 155.845 117.975 156.225 ;
        RECT 118.155 155.675 118.485 156.055 ;
        RECT 118.665 155.845 118.925 156.350 ;
        RECT 119.095 155.675 119.405 156.475 ;
        RECT 119.610 155.845 120.305 156.475 ;
        RECT 121.060 156.395 121.230 156.650 ;
        RECT 120.565 156.225 121.230 156.395 ;
        RECT 121.505 156.350 121.685 157.150 ;
        RECT 121.855 157.135 123.065 158.225 ;
        RECT 120.565 155.845 120.735 156.225 ;
        RECT 120.915 155.675 121.245 156.055 ;
        RECT 121.425 155.845 121.685 156.350 ;
        RECT 121.855 156.425 122.375 156.965 ;
        RECT 122.545 156.595 123.065 157.135 ;
        RECT 123.245 157.165 123.575 158.015 ;
        RECT 121.855 155.675 123.065 156.425 ;
        RECT 123.245 156.400 123.435 157.165 ;
        RECT 123.745 157.085 123.995 158.225 ;
        RECT 124.185 157.585 124.435 158.005 ;
        RECT 124.665 157.755 124.995 158.225 ;
        RECT 125.225 157.585 125.475 158.005 ;
        RECT 124.185 157.415 125.475 157.585 ;
        RECT 125.655 157.585 125.985 158.015 ;
        RECT 125.655 157.415 126.110 157.585 ;
        RECT 124.175 156.915 124.390 157.245 ;
        RECT 123.605 156.585 123.915 156.915 ;
        RECT 124.085 156.585 124.390 156.915 ;
        RECT 124.565 156.585 124.850 157.245 ;
        RECT 125.045 156.585 125.310 157.245 ;
        RECT 125.525 156.585 125.770 157.245 ;
        RECT 123.745 156.415 123.915 156.585 ;
        RECT 125.940 156.415 126.110 157.415 ;
        RECT 126.455 157.135 128.125 158.225 ;
        RECT 123.245 155.890 123.575 156.400 ;
        RECT 123.745 156.245 126.110 156.415 ;
        RECT 126.455 156.445 127.205 156.965 ;
        RECT 127.375 156.615 128.125 157.135 ;
        RECT 128.295 157.150 128.565 158.055 ;
        RECT 128.735 157.465 129.065 158.225 ;
        RECT 129.245 157.295 129.425 158.055 ;
        RECT 123.745 155.675 124.075 156.075 ;
        RECT 125.125 155.905 125.455 156.245 ;
        RECT 125.625 155.675 125.955 156.075 ;
        RECT 126.455 155.675 128.125 156.445 ;
        RECT 128.295 156.350 128.475 157.150 ;
        RECT 128.750 157.125 129.425 157.295 ;
        RECT 129.675 157.150 129.945 158.055 ;
        RECT 130.115 157.465 130.445 158.225 ;
        RECT 130.625 157.295 130.805 158.055 ;
        RECT 128.750 156.980 128.920 157.125 ;
        RECT 128.645 156.650 128.920 156.980 ;
        RECT 128.750 156.395 128.920 156.650 ;
        RECT 129.145 156.575 129.485 156.945 ;
        RECT 128.295 155.845 128.555 156.350 ;
        RECT 128.750 156.225 129.415 156.395 ;
        RECT 128.735 155.675 129.065 156.055 ;
        RECT 129.245 155.845 129.415 156.225 ;
        RECT 129.675 156.350 129.855 157.150 ;
        RECT 130.130 157.125 130.805 157.295 ;
        RECT 131.055 157.135 134.565 158.225 ;
        RECT 130.130 156.980 130.300 157.125 ;
        RECT 130.025 156.650 130.300 156.980 ;
        RECT 130.130 156.395 130.300 156.650 ;
        RECT 130.525 156.575 130.865 156.945 ;
        RECT 131.055 156.445 132.705 156.965 ;
        RECT 132.875 156.615 134.565 157.135 ;
        RECT 135.195 157.060 135.485 158.225 ;
        RECT 135.655 157.135 137.325 158.225 ;
        RECT 137.505 157.505 137.835 158.225 ;
        RECT 135.655 156.445 136.405 156.965 ;
        RECT 136.575 156.615 137.325 157.135 ;
        RECT 137.495 156.865 137.725 157.205 ;
        RECT 138.015 156.865 138.230 157.980 ;
        RECT 138.425 157.280 138.755 158.055 ;
        RECT 138.925 157.450 139.635 158.225 ;
        RECT 138.425 157.065 139.575 157.280 ;
        RECT 137.495 156.665 137.825 156.865 ;
        RECT 138.015 156.685 138.465 156.865 ;
        RECT 138.135 156.665 138.465 156.685 ;
        RECT 138.635 156.665 139.105 156.895 ;
        RECT 139.290 156.495 139.575 157.065 ;
        RECT 139.805 156.620 140.085 158.055 ;
        RECT 140.265 157.505 140.595 158.225 ;
        RECT 140.255 156.865 140.485 157.205 ;
        RECT 140.775 156.865 140.990 157.980 ;
        RECT 141.185 157.280 141.515 158.055 ;
        RECT 141.685 157.450 142.395 158.225 ;
        RECT 141.185 157.065 142.335 157.280 ;
        RECT 140.255 156.665 140.585 156.865 ;
        RECT 140.775 156.685 141.225 156.865 ;
        RECT 140.895 156.665 141.225 156.685 ;
        RECT 141.395 156.665 141.865 156.895 ;
        RECT 129.675 155.845 129.935 156.350 ;
        RECT 130.130 156.225 130.795 156.395 ;
        RECT 130.115 155.675 130.445 156.055 ;
        RECT 130.625 155.845 130.795 156.225 ;
        RECT 131.055 155.675 134.565 156.445 ;
        RECT 135.195 155.675 135.485 156.400 ;
        RECT 135.655 155.675 137.325 156.445 ;
        RECT 137.495 156.305 138.675 156.495 ;
        RECT 137.495 155.845 137.835 156.305 ;
        RECT 138.345 156.225 138.675 156.305 ;
        RECT 138.865 156.305 139.575 156.495 ;
        RECT 138.865 156.165 139.165 156.305 ;
        RECT 138.850 156.155 139.165 156.165 ;
        RECT 138.840 156.145 139.165 156.155 ;
        RECT 138.830 156.140 139.165 156.145 ;
        RECT 138.005 155.675 138.175 156.135 ;
        RECT 138.825 156.130 139.165 156.140 ;
        RECT 138.820 156.125 139.165 156.130 ;
        RECT 138.815 156.115 139.165 156.125 ;
        RECT 138.810 156.110 139.165 156.115 ;
        RECT 138.805 155.845 139.165 156.110 ;
        RECT 139.405 155.675 139.575 156.135 ;
        RECT 139.745 155.845 140.085 156.620 ;
        RECT 142.050 156.495 142.335 157.065 ;
        RECT 142.565 156.620 142.845 158.055 ;
        RECT 140.255 156.305 141.435 156.495 ;
        RECT 140.255 155.845 140.595 156.305 ;
        RECT 141.105 156.225 141.435 156.305 ;
        RECT 141.625 156.305 142.335 156.495 ;
        RECT 141.625 156.165 141.925 156.305 ;
        RECT 141.610 156.155 141.925 156.165 ;
        RECT 141.600 156.145 141.925 156.155 ;
        RECT 141.590 156.140 141.925 156.145 ;
        RECT 140.765 155.675 140.935 156.135 ;
        RECT 141.585 156.130 141.925 156.140 ;
        RECT 141.580 156.125 141.925 156.130 ;
        RECT 141.575 156.115 141.925 156.125 ;
        RECT 141.570 156.110 141.925 156.115 ;
        RECT 141.565 155.845 141.925 156.110 ;
        RECT 142.165 155.675 142.335 156.135 ;
        RECT 142.505 155.845 142.845 156.620 ;
        RECT 143.015 156.620 143.295 158.055 ;
        RECT 143.465 157.450 144.175 158.225 ;
        RECT 144.345 157.280 144.675 158.055 ;
        RECT 143.525 157.065 144.675 157.280 ;
        RECT 143.015 155.845 143.355 156.620 ;
        RECT 143.525 156.495 143.810 157.065 ;
        RECT 143.995 156.665 144.465 156.895 ;
        RECT 144.870 156.865 145.085 157.980 ;
        RECT 145.265 157.505 145.595 158.225 ;
        RECT 145.775 157.790 151.120 158.225 ;
        RECT 145.375 156.865 145.605 157.205 ;
        RECT 144.635 156.685 145.085 156.865 ;
        RECT 144.635 156.665 144.965 156.685 ;
        RECT 145.275 156.665 145.605 156.865 ;
        RECT 143.525 156.305 144.235 156.495 ;
        RECT 143.935 156.165 144.235 156.305 ;
        RECT 144.425 156.305 145.605 156.495 ;
        RECT 144.425 156.225 144.755 156.305 ;
        RECT 143.935 156.155 144.250 156.165 ;
        RECT 143.935 156.145 144.260 156.155 ;
        RECT 143.935 156.140 144.270 156.145 ;
        RECT 143.525 155.675 143.695 156.135 ;
        RECT 143.935 156.130 144.275 156.140 ;
        RECT 143.935 156.125 144.280 156.130 ;
        RECT 143.935 156.115 144.285 156.125 ;
        RECT 143.935 156.110 144.290 156.115 ;
        RECT 143.935 155.845 144.295 156.110 ;
        RECT 144.925 155.675 145.095 156.135 ;
        RECT 145.265 155.845 145.605 156.305 ;
        RECT 147.360 156.220 147.700 157.050 ;
        RECT 149.180 156.540 149.530 157.790 ;
        RECT 151.295 157.085 151.575 158.225 ;
        RECT 151.745 157.075 152.075 158.055 ;
        RECT 152.245 157.085 152.505 158.225 ;
        RECT 152.675 157.135 154.345 158.225 ;
        RECT 151.305 156.645 151.640 156.915 ;
        RECT 151.810 156.525 151.980 157.075 ;
        RECT 152.150 156.665 152.485 156.915 ;
        RECT 151.810 156.475 151.985 156.525 ;
        RECT 145.775 155.675 151.120 156.220 ;
        RECT 151.295 155.675 151.605 156.475 ;
        RECT 151.810 155.845 152.505 156.475 ;
        RECT 152.675 156.445 153.425 156.965 ;
        RECT 153.595 156.615 154.345 157.135 ;
        RECT 154.975 157.135 156.185 158.225 ;
        RECT 154.975 156.595 155.495 157.135 ;
        RECT 152.675 155.675 154.345 156.445 ;
        RECT 155.665 156.425 156.185 156.965 ;
        RECT 154.975 155.675 156.185 156.425 ;
        RECT 70.710 155.505 156.270 155.675 ;
        RECT 70.795 154.755 72.005 155.505 ;
        RECT 72.265 154.955 72.435 155.245 ;
        RECT 72.605 155.125 72.935 155.505 ;
        RECT 72.265 154.785 72.930 154.955 ;
        RECT 70.795 154.215 71.315 154.755 ;
        RECT 71.485 154.045 72.005 154.585 ;
        RECT 70.795 152.955 72.005 154.045 ;
        RECT 72.180 153.965 72.530 154.615 ;
        RECT 72.700 153.795 72.930 154.785 ;
        RECT 72.265 153.625 72.930 153.795 ;
        RECT 72.265 153.125 72.435 153.625 ;
        RECT 72.605 152.955 72.935 153.455 ;
        RECT 73.105 153.125 73.290 155.245 ;
        RECT 73.545 155.045 73.795 155.505 ;
        RECT 73.965 155.055 74.300 155.225 ;
        RECT 74.495 155.055 75.170 155.225 ;
        RECT 73.965 154.915 74.135 155.055 ;
        RECT 73.460 153.925 73.740 154.875 ;
        RECT 73.910 154.785 74.135 154.915 ;
        RECT 73.910 153.680 74.080 154.785 ;
        RECT 74.305 154.635 74.830 154.855 ;
        RECT 74.250 153.870 74.490 154.465 ;
        RECT 74.660 153.935 74.830 154.635 ;
        RECT 75.000 154.275 75.170 155.055 ;
        RECT 75.490 155.005 75.860 155.505 ;
        RECT 76.040 155.055 76.445 155.225 ;
        RECT 76.615 155.055 77.400 155.225 ;
        RECT 76.040 154.825 76.210 155.055 ;
        RECT 75.380 154.525 76.210 154.825 ;
        RECT 76.595 154.555 77.060 154.885 ;
        RECT 75.380 154.495 75.580 154.525 ;
        RECT 75.700 154.275 75.870 154.345 ;
        RECT 75.000 154.105 75.870 154.275 ;
        RECT 75.360 154.015 75.870 154.105 ;
        RECT 73.910 153.550 74.215 153.680 ;
        RECT 74.660 153.570 75.190 153.935 ;
        RECT 73.530 152.955 73.795 153.415 ;
        RECT 73.965 153.125 74.215 153.550 ;
        RECT 75.360 153.400 75.530 154.015 ;
        RECT 74.425 153.230 75.530 153.400 ;
        RECT 75.700 152.955 75.870 153.755 ;
        RECT 76.040 153.455 76.210 154.525 ;
        RECT 76.380 153.625 76.570 154.345 ;
        RECT 76.740 153.595 77.060 154.555 ;
        RECT 77.230 154.595 77.400 155.055 ;
        RECT 77.675 154.975 77.885 155.505 ;
        RECT 78.145 154.765 78.475 155.290 ;
        RECT 78.645 154.895 78.815 155.505 ;
        RECT 78.985 154.850 79.315 155.285 ;
        RECT 78.985 154.765 79.365 154.850 ;
        RECT 78.275 154.595 78.475 154.765 ;
        RECT 79.140 154.725 79.365 154.765 ;
        RECT 77.230 154.265 78.105 154.595 ;
        RECT 78.275 154.265 79.025 154.595 ;
        RECT 76.040 153.125 76.290 153.455 ;
        RECT 77.230 153.425 77.400 154.265 ;
        RECT 78.275 154.060 78.465 154.265 ;
        RECT 79.195 154.145 79.365 154.725 ;
        RECT 79.535 154.735 81.205 155.505 ;
        RECT 81.465 154.955 81.635 155.335 ;
        RECT 81.815 155.125 82.145 155.505 ;
        RECT 81.465 154.785 82.130 154.955 ;
        RECT 82.325 154.830 82.585 155.335 ;
        RECT 79.535 154.215 80.285 154.735 ;
        RECT 79.150 154.095 79.365 154.145 ;
        RECT 77.570 153.685 78.465 154.060 ;
        RECT 78.975 154.015 79.365 154.095 ;
        RECT 80.455 154.045 81.205 154.565 ;
        RECT 81.395 154.235 81.735 154.605 ;
        RECT 81.960 154.530 82.130 154.785 ;
        RECT 81.960 154.200 82.235 154.530 ;
        RECT 81.960 154.055 82.130 154.200 ;
        RECT 76.515 153.255 77.400 153.425 ;
        RECT 77.580 152.955 77.895 153.455 ;
        RECT 78.125 153.125 78.465 153.685 ;
        RECT 78.635 152.955 78.805 153.965 ;
        RECT 78.975 153.170 79.305 154.015 ;
        RECT 79.535 152.955 81.205 154.045 ;
        RECT 81.455 153.885 82.130 154.055 ;
        RECT 82.405 154.030 82.585 154.830 ;
        RECT 82.755 154.735 85.345 155.505 ;
        RECT 85.985 155.165 87.175 155.335 ;
        RECT 85.985 154.995 86.295 155.165 ;
        RECT 82.755 154.215 83.965 154.735 ;
        RECT 84.135 154.045 85.345 154.565 ;
        RECT 85.980 154.190 86.295 154.825 ;
        RECT 81.455 153.125 81.635 153.885 ;
        RECT 81.815 152.955 82.145 153.715 ;
        RECT 82.315 153.125 82.585 154.030 ;
        RECT 82.755 152.955 85.345 154.045 ;
        RECT 85.985 152.955 86.295 154.020 ;
        RECT 86.465 153.805 86.675 154.995 ;
        RECT 86.845 154.875 87.175 155.165 ;
        RECT 87.415 155.045 87.585 155.505 ;
        RECT 87.815 154.875 88.145 155.335 ;
        RECT 88.325 155.045 88.495 155.505 ;
        RECT 88.675 154.875 89.005 155.335 ;
        RECT 86.845 154.705 89.005 154.875 ;
        RECT 89.210 154.935 89.465 155.285 ;
        RECT 89.635 155.105 89.965 155.505 ;
        RECT 90.135 154.935 90.305 155.285 ;
        RECT 90.475 155.105 90.855 155.505 ;
        RECT 89.210 154.765 90.875 154.935 ;
        RECT 91.045 154.830 91.320 155.175 ;
        RECT 90.705 154.595 90.875 154.765 ;
        RECT 87.015 154.485 87.510 154.515 ;
        RECT 86.955 154.315 87.510 154.485 ;
        RECT 87.690 154.315 88.490 154.515 ;
        RECT 87.015 154.145 87.510 154.315 ;
        RECT 88.660 154.145 88.990 154.535 ;
        RECT 89.195 154.265 89.540 154.595 ;
        RECT 89.710 154.265 90.535 154.595 ;
        RECT 90.705 154.265 90.980 154.595 ;
        RECT 87.015 153.975 88.990 154.145 ;
        RECT 89.215 153.805 89.540 154.095 ;
        RECT 89.710 153.975 89.905 154.265 ;
        RECT 90.705 154.095 90.875 154.265 ;
        RECT 91.150 154.095 91.320 154.830 ;
        RECT 91.515 154.695 91.755 155.505 ;
        RECT 91.925 154.695 92.255 155.335 ;
        RECT 92.425 154.695 92.695 155.505 ;
        RECT 92.875 154.735 96.385 155.505 ;
        RECT 96.555 154.780 96.845 155.505 ;
        RECT 97.015 154.960 102.360 155.505 ;
        RECT 102.865 155.105 103.195 155.505 ;
        RECT 91.495 154.265 91.845 154.515 ;
        RECT 92.015 154.095 92.185 154.695 ;
        RECT 92.355 154.265 92.705 154.515 ;
        RECT 92.875 154.215 94.525 154.735 ;
        RECT 90.215 153.925 90.875 154.095 ;
        RECT 90.215 153.805 90.385 153.925 ;
        RECT 86.465 153.625 88.115 153.805 ;
        RECT 86.465 153.125 86.700 153.625 ;
        RECT 87.815 153.465 88.115 153.625 ;
        RECT 86.870 152.955 87.200 153.415 ;
        RECT 87.395 153.295 87.585 153.455 ;
        RECT 88.285 153.295 88.505 153.805 ;
        RECT 87.395 153.125 88.505 153.295 ;
        RECT 88.675 152.955 89.005 153.805 ;
        RECT 89.215 153.635 90.385 153.805 ;
        RECT 89.195 153.175 90.385 153.465 ;
        RECT 90.555 152.955 90.835 153.755 ;
        RECT 91.045 153.125 91.320 154.095 ;
        RECT 91.505 153.925 92.185 154.095 ;
        RECT 91.505 153.140 91.835 153.925 ;
        RECT 92.365 152.955 92.695 154.095 ;
        RECT 94.695 154.045 96.385 154.565 ;
        RECT 98.600 154.130 98.940 154.960 ;
        RECT 103.365 154.935 103.695 155.275 ;
        RECT 104.745 155.105 105.075 155.505 ;
        RECT 102.710 154.765 105.075 154.935 ;
        RECT 105.245 154.780 105.575 155.290 ;
        RECT 92.875 152.955 96.385 154.045 ;
        RECT 96.555 152.955 96.845 154.120 ;
        RECT 100.420 153.390 100.770 154.640 ;
        RECT 102.710 153.765 102.880 154.765 ;
        RECT 104.905 154.595 105.075 154.765 ;
        RECT 103.050 153.935 103.295 154.595 ;
        RECT 103.510 153.935 103.775 154.595 ;
        RECT 103.970 153.935 104.255 154.595 ;
        RECT 104.430 154.265 104.735 154.595 ;
        RECT 104.905 154.265 105.215 154.595 ;
        RECT 104.430 153.935 104.645 154.265 ;
        RECT 102.710 153.595 103.165 153.765 ;
        RECT 97.015 152.955 102.360 153.390 ;
        RECT 102.835 153.165 103.165 153.595 ;
        RECT 103.345 153.595 104.635 153.765 ;
        RECT 103.345 153.175 103.595 153.595 ;
        RECT 103.825 152.955 104.155 153.425 ;
        RECT 104.385 153.175 104.635 153.595 ;
        RECT 104.825 152.955 105.075 154.095 ;
        RECT 105.385 154.015 105.575 154.780 ;
        RECT 105.755 154.755 106.965 155.505 ;
        RECT 107.295 154.945 107.625 155.335 ;
        RECT 107.795 155.115 108.980 155.285 ;
        RECT 109.240 155.035 109.410 155.505 ;
        RECT 107.295 154.765 107.805 154.945 ;
        RECT 105.755 154.215 106.275 154.755 ;
        RECT 106.445 154.045 106.965 154.585 ;
        RECT 107.135 154.305 107.465 154.595 ;
        RECT 107.635 154.135 107.805 154.765 ;
        RECT 108.210 154.855 108.595 154.945 ;
        RECT 109.580 154.855 109.910 155.320 ;
        RECT 108.210 154.685 109.910 154.855 ;
        RECT 110.080 154.685 110.250 155.505 ;
        RECT 110.420 154.685 111.105 155.325 ;
        RECT 107.975 154.305 108.305 154.515 ;
        RECT 108.485 154.265 108.865 154.515 ;
        RECT 105.245 153.165 105.575 154.015 ;
        RECT 105.755 152.955 106.965 154.045 ;
        RECT 107.290 153.965 108.375 154.135 ;
        RECT 107.290 153.125 107.590 153.965 ;
        RECT 107.785 152.955 108.035 153.795 ;
        RECT 108.205 153.715 108.375 153.965 ;
        RECT 108.545 153.885 108.865 154.265 ;
        RECT 109.055 154.305 109.540 154.515 ;
        RECT 109.730 154.305 110.180 154.515 ;
        RECT 110.350 154.305 110.685 154.515 ;
        RECT 109.055 154.145 109.430 154.305 ;
        RECT 109.035 153.975 109.430 154.145 ;
        RECT 110.350 154.135 110.520 154.305 ;
        RECT 109.055 153.885 109.430 153.975 ;
        RECT 109.600 153.965 110.520 154.135 ;
        RECT 109.600 153.715 109.770 153.965 ;
        RECT 108.205 153.545 109.770 153.715 ;
        RECT 108.625 153.125 109.430 153.545 ;
        RECT 109.940 152.955 110.270 153.795 ;
        RECT 110.855 153.715 111.105 154.685 ;
        RECT 110.440 153.125 111.105 153.715 ;
        RECT 112.195 154.765 112.455 155.335 ;
        RECT 112.625 155.105 113.010 155.505 ;
        RECT 113.180 154.935 113.435 155.335 ;
        RECT 112.625 154.765 113.435 154.935 ;
        RECT 113.625 154.765 113.870 155.335 ;
        RECT 114.040 155.105 114.425 155.505 ;
        RECT 114.595 154.935 114.850 155.335 ;
        RECT 114.040 154.765 114.850 154.935 ;
        RECT 115.040 154.765 115.465 155.335 ;
        RECT 115.635 155.105 116.020 155.505 ;
        RECT 116.190 154.935 116.625 155.335 ;
        RECT 115.635 154.765 116.625 154.935 ;
        RECT 116.885 154.955 117.055 155.335 ;
        RECT 117.235 155.125 117.565 155.505 ;
        RECT 116.885 154.785 117.550 154.955 ;
        RECT 117.745 154.830 118.005 155.335 ;
        RECT 112.195 154.095 112.380 154.765 ;
        RECT 112.625 154.595 112.975 154.765 ;
        RECT 113.625 154.595 113.795 154.765 ;
        RECT 114.040 154.595 114.390 154.765 ;
        RECT 115.040 154.595 115.390 154.765 ;
        RECT 115.635 154.595 115.970 154.765 ;
        RECT 112.550 154.265 112.975 154.595 ;
        RECT 112.195 153.125 112.455 154.095 ;
        RECT 112.625 153.745 112.975 154.265 ;
        RECT 113.145 154.095 113.795 154.595 ;
        RECT 113.965 154.265 114.390 154.595 ;
        RECT 113.145 153.915 113.870 154.095 ;
        RECT 112.625 153.550 113.435 153.745 ;
        RECT 112.625 152.955 113.010 153.380 ;
        RECT 113.180 153.125 113.435 153.550 ;
        RECT 113.625 153.125 113.870 153.915 ;
        RECT 114.040 153.745 114.390 154.265 ;
        RECT 114.560 154.095 115.390 154.595 ;
        RECT 115.560 154.265 115.970 154.595 ;
        RECT 114.560 153.915 115.465 154.095 ;
        RECT 114.040 153.550 114.870 153.745 ;
        RECT 114.040 152.955 114.425 153.380 ;
        RECT 114.595 153.125 114.870 153.550 ;
        RECT 115.040 153.125 115.465 153.915 ;
        RECT 115.635 153.720 115.970 154.265 ;
        RECT 116.140 153.890 116.625 154.595 ;
        RECT 116.815 154.235 117.155 154.605 ;
        RECT 117.380 154.530 117.550 154.785 ;
        RECT 117.380 154.200 117.655 154.530 ;
        RECT 117.380 154.055 117.550 154.200 ;
        RECT 116.875 153.885 117.550 154.055 ;
        RECT 117.825 154.030 118.005 154.830 ;
        RECT 115.635 153.550 116.625 153.720 ;
        RECT 115.635 152.955 116.020 153.380 ;
        RECT 116.190 153.125 116.625 153.550 ;
        RECT 116.875 153.125 117.055 153.885 ;
        RECT 117.235 152.955 117.565 153.715 ;
        RECT 117.735 153.125 118.005 154.030 ;
        RECT 119.105 154.780 119.435 155.290 ;
        RECT 119.605 155.105 119.935 155.505 ;
        RECT 120.985 154.935 121.315 155.275 ;
        RECT 121.485 155.105 121.815 155.505 ;
        RECT 119.105 154.145 119.295 154.780 ;
        RECT 119.605 154.765 121.970 154.935 ;
        RECT 122.315 154.780 122.605 155.505 ;
        RECT 119.605 154.595 119.775 154.765 ;
        RECT 119.465 154.265 119.775 154.595 ;
        RECT 119.945 154.265 120.250 154.595 ;
        RECT 119.105 154.015 119.325 154.145 ;
        RECT 119.105 153.165 119.435 154.015 ;
        RECT 119.605 152.955 119.855 154.095 ;
        RECT 120.035 153.935 120.250 154.265 ;
        RECT 120.425 153.935 120.710 154.595 ;
        RECT 120.905 153.935 121.170 154.595 ;
        RECT 121.385 153.935 121.630 154.595 ;
        RECT 121.800 153.765 121.970 154.765 ;
        RECT 122.775 154.685 123.460 155.325 ;
        RECT 123.630 154.685 123.800 155.505 ;
        RECT 123.970 154.855 124.300 155.320 ;
        RECT 124.470 155.035 124.640 155.505 ;
        RECT 124.900 155.115 126.085 155.285 ;
        RECT 126.255 154.945 126.585 155.335 ;
        RECT 126.915 154.960 132.260 155.505 ;
        RECT 125.285 154.855 125.670 154.945 ;
        RECT 123.970 154.685 125.670 154.855 ;
        RECT 126.075 154.765 126.585 154.945 ;
        RECT 120.045 153.595 121.335 153.765 ;
        RECT 120.045 153.175 120.295 153.595 ;
        RECT 120.525 152.955 120.855 153.425 ;
        RECT 121.085 153.175 121.335 153.595 ;
        RECT 121.515 153.595 121.970 153.765 ;
        RECT 121.515 153.165 121.845 153.595 ;
        RECT 122.315 152.955 122.605 154.120 ;
        RECT 122.775 153.715 123.025 154.685 ;
        RECT 123.195 154.305 123.530 154.515 ;
        RECT 123.700 154.305 124.150 154.515 ;
        RECT 124.340 154.305 124.825 154.515 ;
        RECT 123.360 154.135 123.530 154.305 ;
        RECT 123.360 153.965 124.280 154.135 ;
        RECT 122.775 153.125 123.440 153.715 ;
        RECT 123.610 152.955 123.940 153.795 ;
        RECT 124.110 153.715 124.280 153.965 ;
        RECT 124.450 153.885 124.825 154.305 ;
        RECT 125.015 154.265 125.395 154.515 ;
        RECT 125.575 154.305 125.905 154.515 ;
        RECT 125.015 153.885 125.335 154.265 ;
        RECT 126.075 154.135 126.245 154.765 ;
        RECT 126.415 154.305 126.745 154.595 ;
        RECT 125.505 153.965 126.590 154.135 ;
        RECT 128.500 154.130 128.840 154.960 ;
        RECT 132.435 154.735 135.945 155.505 ;
        RECT 137.125 154.955 137.295 155.335 ;
        RECT 137.475 155.125 137.805 155.505 ;
        RECT 137.125 154.785 137.790 154.955 ;
        RECT 137.985 154.830 138.245 155.335 ;
        RECT 138.415 154.960 143.760 155.505 ;
        RECT 125.505 153.715 125.675 153.965 ;
        RECT 124.110 153.545 125.675 153.715 ;
        RECT 124.450 153.125 125.255 153.545 ;
        RECT 125.845 152.955 126.095 153.795 ;
        RECT 126.290 153.125 126.590 153.965 ;
        RECT 130.320 153.390 130.670 154.640 ;
        RECT 132.435 154.215 134.085 154.735 ;
        RECT 134.255 154.045 135.945 154.565 ;
        RECT 137.055 154.235 137.395 154.605 ;
        RECT 137.620 154.530 137.790 154.785 ;
        RECT 137.620 154.200 137.895 154.530 ;
        RECT 137.620 154.055 137.790 154.200 ;
        RECT 126.915 152.955 132.260 153.390 ;
        RECT 132.435 152.955 135.945 154.045 ;
        RECT 137.115 153.885 137.790 154.055 ;
        RECT 138.065 154.030 138.245 154.830 ;
        RECT 140.000 154.130 140.340 154.960 ;
        RECT 143.935 154.735 147.445 155.505 ;
        RECT 148.075 154.780 148.365 155.505 ;
        RECT 149.030 154.765 149.645 155.335 ;
        RECT 149.815 154.995 150.030 155.505 ;
        RECT 150.260 154.995 150.540 155.325 ;
        RECT 150.720 154.995 150.960 155.505 ;
        RECT 137.115 153.125 137.295 153.885 ;
        RECT 137.475 152.955 137.805 153.715 ;
        RECT 137.975 153.125 138.245 154.030 ;
        RECT 141.820 153.390 142.170 154.640 ;
        RECT 143.935 154.215 145.585 154.735 ;
        RECT 145.755 154.045 147.445 154.565 ;
        RECT 138.415 152.955 143.760 153.390 ;
        RECT 143.935 152.955 147.445 154.045 ;
        RECT 148.075 152.955 148.365 154.120 ;
        RECT 149.030 153.745 149.345 154.765 ;
        RECT 149.515 154.095 149.685 154.595 ;
        RECT 149.935 154.265 150.200 154.825 ;
        RECT 150.370 154.095 150.540 154.995 ;
        RECT 150.710 154.265 151.065 154.825 ;
        RECT 151.295 154.735 154.805 155.505 ;
        RECT 154.975 154.755 156.185 155.505 ;
        RECT 151.295 154.215 152.945 154.735 ;
        RECT 149.515 153.925 150.940 154.095 ;
        RECT 153.115 154.045 154.805 154.565 ;
        RECT 149.030 153.125 149.565 153.745 ;
        RECT 149.735 152.955 150.065 153.755 ;
        RECT 150.550 153.750 150.940 153.925 ;
        RECT 151.295 152.955 154.805 154.045 ;
        RECT 154.975 154.045 155.495 154.585 ;
        RECT 155.665 154.215 156.185 154.755 ;
        RECT 154.975 152.955 156.185 154.045 ;
        RECT 70.710 152.785 156.270 152.955 ;
        RECT 70.795 151.695 72.005 152.785 ;
        RECT 72.175 152.350 77.520 152.785 ;
        RECT 70.795 150.985 71.315 151.525 ;
        RECT 71.485 151.155 72.005 151.695 ;
        RECT 70.795 150.235 72.005 150.985 ;
        RECT 73.760 150.780 74.100 151.610 ;
        RECT 75.580 151.100 75.930 152.350 ;
        RECT 77.695 151.695 80.285 152.785 ;
        RECT 77.695 151.005 78.905 151.525 ;
        RECT 79.075 151.175 80.285 151.695 ;
        RECT 80.915 151.710 81.185 152.615 ;
        RECT 81.355 152.025 81.685 152.785 ;
        RECT 81.865 151.855 82.045 152.615 ;
        RECT 72.175 150.235 77.520 150.780 ;
        RECT 77.695 150.235 80.285 151.005 ;
        RECT 80.915 150.910 81.095 151.710 ;
        RECT 81.370 151.685 82.045 151.855 ;
        RECT 82.295 151.695 83.505 152.785 ;
        RECT 81.370 151.540 81.540 151.685 ;
        RECT 81.265 151.210 81.540 151.540 ;
        RECT 81.370 150.955 81.540 151.210 ;
        RECT 81.765 151.135 82.105 151.505 ;
        RECT 82.295 150.985 82.815 151.525 ;
        RECT 82.985 151.155 83.505 151.695 ;
        RECT 83.675 151.620 83.965 152.785 ;
        RECT 84.135 152.350 89.480 152.785 ;
        RECT 89.655 152.350 95.000 152.785 ;
        RECT 80.915 150.405 81.175 150.910 ;
        RECT 81.370 150.785 82.035 150.955 ;
        RECT 81.355 150.235 81.685 150.615 ;
        RECT 81.865 150.405 82.035 150.785 ;
        RECT 82.295 150.235 83.505 150.985 ;
        RECT 83.675 150.235 83.965 150.960 ;
        RECT 85.720 150.780 86.060 151.610 ;
        RECT 87.540 151.100 87.890 152.350 ;
        RECT 91.240 150.780 91.580 151.610 ;
        RECT 93.060 151.100 93.410 152.350 ;
        RECT 95.175 151.695 96.845 152.785 ;
        RECT 95.175 151.005 95.925 151.525 ;
        RECT 96.095 151.175 96.845 151.695 ;
        RECT 97.015 151.710 97.285 152.615 ;
        RECT 97.455 152.025 97.785 152.785 ;
        RECT 97.965 151.855 98.145 152.615 ;
        RECT 98.395 152.190 98.830 152.615 ;
        RECT 99.000 152.360 99.385 152.785 ;
        RECT 98.395 152.020 99.385 152.190 ;
        RECT 84.135 150.235 89.480 150.780 ;
        RECT 89.655 150.235 95.000 150.780 ;
        RECT 95.175 150.235 96.845 151.005 ;
        RECT 97.015 150.910 97.195 151.710 ;
        RECT 97.470 151.685 98.145 151.855 ;
        RECT 97.470 151.540 97.640 151.685 ;
        RECT 97.365 151.210 97.640 151.540 ;
        RECT 97.470 150.955 97.640 151.210 ;
        RECT 97.865 151.135 98.205 151.505 ;
        RECT 98.395 151.145 98.880 151.850 ;
        RECT 99.050 151.475 99.385 152.020 ;
        RECT 99.555 151.825 99.980 152.615 ;
        RECT 100.150 152.190 100.425 152.615 ;
        RECT 100.595 152.360 100.980 152.785 ;
        RECT 100.150 151.995 100.980 152.190 ;
        RECT 99.555 151.645 100.460 151.825 ;
        RECT 99.050 151.145 99.460 151.475 ;
        RECT 99.630 151.145 100.460 151.645 ;
        RECT 100.630 151.475 100.980 151.995 ;
        RECT 101.150 151.825 101.395 152.615 ;
        RECT 101.585 152.190 101.840 152.615 ;
        RECT 102.010 152.360 102.395 152.785 ;
        RECT 101.585 151.995 102.395 152.190 ;
        RECT 101.150 151.645 101.875 151.825 ;
        RECT 100.630 151.145 101.055 151.475 ;
        RECT 101.225 151.145 101.875 151.645 ;
        RECT 102.045 151.475 102.395 151.995 ;
        RECT 102.565 151.645 102.825 152.615 ;
        RECT 102.045 151.145 102.470 151.475 ;
        RECT 99.050 150.975 99.385 151.145 ;
        RECT 99.630 150.975 99.980 151.145 ;
        RECT 100.630 150.975 100.980 151.145 ;
        RECT 101.225 150.975 101.395 151.145 ;
        RECT 102.045 150.975 102.395 151.145 ;
        RECT 102.640 150.975 102.825 151.645 ;
        RECT 97.015 150.405 97.275 150.910 ;
        RECT 97.470 150.785 98.135 150.955 ;
        RECT 97.455 150.235 97.785 150.615 ;
        RECT 97.965 150.405 98.135 150.785 ;
        RECT 98.395 150.805 99.385 150.975 ;
        RECT 98.395 150.405 98.830 150.805 ;
        RECT 99.000 150.235 99.385 150.635 ;
        RECT 99.555 150.405 99.980 150.975 ;
        RECT 100.170 150.805 100.980 150.975 ;
        RECT 100.170 150.405 100.425 150.805 ;
        RECT 100.595 150.235 100.980 150.635 ;
        RECT 101.150 150.405 101.395 150.975 ;
        RECT 101.585 150.805 102.395 150.975 ;
        RECT 101.585 150.405 101.840 150.805 ;
        RECT 102.010 150.235 102.395 150.635 ;
        RECT 102.565 150.405 102.825 150.975 ;
        RECT 102.995 152.025 103.660 152.615 ;
        RECT 102.995 151.055 103.245 152.025 ;
        RECT 103.830 151.945 104.160 152.785 ;
        RECT 104.670 152.195 105.475 152.615 ;
        RECT 104.330 152.025 105.895 152.195 ;
        RECT 104.330 151.775 104.500 152.025 ;
        RECT 103.580 151.605 104.500 151.775 ;
        RECT 103.580 151.435 103.750 151.605 ;
        RECT 104.670 151.435 105.045 151.855 ;
        RECT 103.415 151.225 103.750 151.435 ;
        RECT 103.920 151.225 104.370 151.435 ;
        RECT 104.560 151.425 105.045 151.435 ;
        RECT 105.235 151.475 105.555 151.855 ;
        RECT 105.725 151.775 105.895 152.025 ;
        RECT 106.065 151.945 106.315 152.785 ;
        RECT 106.510 151.775 106.810 152.615 ;
        RECT 105.725 151.605 106.810 151.775 ;
        RECT 107.135 151.710 107.405 152.615 ;
        RECT 107.575 152.025 107.905 152.785 ;
        RECT 108.085 151.855 108.265 152.615 ;
        RECT 104.560 151.255 105.065 151.425 ;
        RECT 104.560 151.225 105.045 151.255 ;
        RECT 105.235 151.225 105.615 151.475 ;
        RECT 105.795 151.225 106.125 151.435 ;
        RECT 102.995 150.415 103.680 151.055 ;
        RECT 103.850 150.235 104.020 151.055 ;
        RECT 104.190 150.885 105.890 151.055 ;
        RECT 104.190 150.420 104.520 150.885 ;
        RECT 105.505 150.795 105.890 150.885 ;
        RECT 106.295 150.975 106.465 151.605 ;
        RECT 106.635 151.145 106.965 151.435 ;
        RECT 106.295 150.795 106.805 150.975 ;
        RECT 104.690 150.235 104.860 150.705 ;
        RECT 105.120 150.455 106.305 150.625 ;
        RECT 106.475 150.405 106.805 150.795 ;
        RECT 107.135 150.910 107.315 151.710 ;
        RECT 107.590 151.685 108.265 151.855 ;
        RECT 107.590 151.540 107.760 151.685 ;
        RECT 109.435 151.620 109.725 152.785 ;
        RECT 107.485 151.210 107.760 151.540 ;
        RECT 107.590 150.955 107.760 151.210 ;
        RECT 107.985 151.135 108.325 151.505 ;
        RECT 109.895 151.180 110.175 152.615 ;
        RECT 110.345 152.010 111.055 152.785 ;
        RECT 111.225 151.840 111.555 152.615 ;
        RECT 110.405 151.625 111.555 151.840 ;
        RECT 107.135 150.405 107.395 150.910 ;
        RECT 107.590 150.785 108.255 150.955 ;
        RECT 107.575 150.235 107.905 150.615 ;
        RECT 108.085 150.405 108.255 150.785 ;
        RECT 109.435 150.235 109.725 150.960 ;
        RECT 109.895 150.405 110.235 151.180 ;
        RECT 110.405 151.055 110.690 151.625 ;
        RECT 110.875 151.225 111.345 151.455 ;
        RECT 111.750 151.425 111.965 152.540 ;
        RECT 112.145 152.065 112.475 152.785 ;
        RECT 112.735 151.855 112.915 152.615 ;
        RECT 113.095 152.025 113.425 152.785 ;
        RECT 112.255 151.425 112.485 151.765 ;
        RECT 112.735 151.685 113.410 151.855 ;
        RECT 113.595 151.710 113.865 152.615 ;
        RECT 114.035 152.350 119.380 152.785 ;
        RECT 113.240 151.540 113.410 151.685 ;
        RECT 111.515 151.245 111.965 151.425 ;
        RECT 111.515 151.225 111.845 151.245 ;
        RECT 112.155 151.225 112.485 151.425 ;
        RECT 112.675 151.135 113.015 151.505 ;
        RECT 113.240 151.210 113.515 151.540 ;
        RECT 110.405 150.865 111.115 151.055 ;
        RECT 110.815 150.725 111.115 150.865 ;
        RECT 111.305 150.865 112.485 151.055 ;
        RECT 113.240 150.955 113.410 151.210 ;
        RECT 111.305 150.785 111.635 150.865 ;
        RECT 110.815 150.715 111.130 150.725 ;
        RECT 110.815 150.705 111.140 150.715 ;
        RECT 110.815 150.700 111.150 150.705 ;
        RECT 110.405 150.235 110.575 150.695 ;
        RECT 110.815 150.690 111.155 150.700 ;
        RECT 110.815 150.685 111.160 150.690 ;
        RECT 110.815 150.675 111.165 150.685 ;
        RECT 110.815 150.670 111.170 150.675 ;
        RECT 110.815 150.405 111.175 150.670 ;
        RECT 111.805 150.235 111.975 150.695 ;
        RECT 112.145 150.405 112.485 150.865 ;
        RECT 112.745 150.785 113.410 150.955 ;
        RECT 113.685 150.910 113.865 151.710 ;
        RECT 112.745 150.405 112.915 150.785 ;
        RECT 113.095 150.235 113.425 150.615 ;
        RECT 113.605 150.405 113.865 150.910 ;
        RECT 115.620 150.780 115.960 151.610 ;
        RECT 117.440 151.100 117.790 152.350 ;
        RECT 119.555 151.695 123.065 152.785 ;
        RECT 119.555 151.005 121.205 151.525 ;
        RECT 121.375 151.175 123.065 151.695 ;
        RECT 123.235 151.180 123.515 152.615 ;
        RECT 123.685 152.010 124.395 152.785 ;
        RECT 124.565 151.840 124.895 152.615 ;
        RECT 123.745 151.625 124.895 151.840 ;
        RECT 114.035 150.235 119.380 150.780 ;
        RECT 119.555 150.235 123.065 151.005 ;
        RECT 123.235 150.405 123.575 151.180 ;
        RECT 123.745 151.055 124.030 151.625 ;
        RECT 124.215 151.225 124.685 151.455 ;
        RECT 125.090 151.425 125.305 152.540 ;
        RECT 125.485 152.065 125.815 152.785 ;
        RECT 125.595 151.425 125.825 151.765 ;
        RECT 125.995 151.695 127.205 152.785 ;
        RECT 124.855 151.245 125.305 151.425 ;
        RECT 124.855 151.225 125.185 151.245 ;
        RECT 125.495 151.225 125.825 151.425 ;
        RECT 123.745 150.865 124.455 151.055 ;
        RECT 124.155 150.725 124.455 150.865 ;
        RECT 124.645 150.865 125.825 151.055 ;
        RECT 124.645 150.785 124.975 150.865 ;
        RECT 124.155 150.715 124.470 150.725 ;
        RECT 124.155 150.705 124.480 150.715 ;
        RECT 124.155 150.700 124.490 150.705 ;
        RECT 123.745 150.235 123.915 150.695 ;
        RECT 124.155 150.690 124.495 150.700 ;
        RECT 124.155 150.685 124.500 150.690 ;
        RECT 124.155 150.675 124.505 150.685 ;
        RECT 124.155 150.670 124.510 150.675 ;
        RECT 124.155 150.405 124.515 150.670 ;
        RECT 125.145 150.235 125.315 150.695 ;
        RECT 125.485 150.405 125.825 150.865 ;
        RECT 125.995 150.985 126.515 151.525 ;
        RECT 126.685 151.155 127.205 151.695 ;
        RECT 127.455 151.855 127.635 152.615 ;
        RECT 127.815 152.025 128.145 152.785 ;
        RECT 127.455 151.685 128.130 151.855 ;
        RECT 128.315 151.710 128.585 152.615 ;
        RECT 127.960 151.540 128.130 151.685 ;
        RECT 127.395 151.135 127.735 151.505 ;
        RECT 127.960 151.210 128.235 151.540 ;
        RECT 125.995 150.235 127.205 150.985 ;
        RECT 127.960 150.955 128.130 151.210 ;
        RECT 127.465 150.785 128.130 150.955 ;
        RECT 128.405 150.910 128.585 151.710 ;
        RECT 128.755 151.695 130.425 152.785 ;
        RECT 127.465 150.405 127.635 150.785 ;
        RECT 127.815 150.235 128.145 150.615 ;
        RECT 128.325 150.405 128.585 150.910 ;
        RECT 128.755 151.005 129.505 151.525 ;
        RECT 129.675 151.175 130.425 151.695 ;
        RECT 131.055 151.710 131.325 152.615 ;
        RECT 131.495 152.025 131.825 152.785 ;
        RECT 132.005 151.855 132.185 152.615 ;
        RECT 128.755 150.235 130.425 151.005 ;
        RECT 131.055 150.910 131.235 151.710 ;
        RECT 131.510 151.685 132.185 151.855 ;
        RECT 132.435 151.695 135.025 152.785 ;
        RECT 131.510 151.540 131.680 151.685 ;
        RECT 131.405 151.210 131.680 151.540 ;
        RECT 131.510 150.955 131.680 151.210 ;
        RECT 131.905 151.135 132.245 151.505 ;
        RECT 132.435 151.005 133.645 151.525 ;
        RECT 133.815 151.175 135.025 151.695 ;
        RECT 135.195 151.620 135.485 152.785 ;
        RECT 135.810 151.775 136.110 152.615 ;
        RECT 136.305 151.945 136.555 152.785 ;
        RECT 137.145 152.195 137.950 152.615 ;
        RECT 136.725 152.025 138.290 152.195 ;
        RECT 136.725 151.775 136.895 152.025 ;
        RECT 135.810 151.605 136.895 151.775 ;
        RECT 135.655 151.145 135.985 151.435 ;
        RECT 131.055 150.405 131.315 150.910 ;
        RECT 131.510 150.785 132.175 150.955 ;
        RECT 131.495 150.235 131.825 150.615 ;
        RECT 132.005 150.405 132.175 150.785 ;
        RECT 132.435 150.235 135.025 151.005 ;
        RECT 136.155 150.975 136.325 151.605 ;
        RECT 137.065 151.475 137.385 151.855 ;
        RECT 136.495 151.225 136.825 151.435 ;
        RECT 137.005 151.225 137.385 151.475 ;
        RECT 137.575 151.435 137.950 151.855 ;
        RECT 138.120 151.775 138.290 152.025 ;
        RECT 138.460 151.945 138.790 152.785 ;
        RECT 138.960 152.025 139.625 152.615 ;
        RECT 139.805 152.065 140.135 152.785 ;
        RECT 138.120 151.605 139.040 151.775 ;
        RECT 138.870 151.435 139.040 151.605 ;
        RECT 137.575 151.425 138.060 151.435 ;
        RECT 137.555 151.255 138.060 151.425 ;
        RECT 137.575 151.225 138.060 151.255 ;
        RECT 138.250 151.225 138.700 151.435 ;
        RECT 138.870 151.225 139.205 151.435 ;
        RECT 139.375 151.055 139.625 152.025 ;
        RECT 139.795 151.425 140.025 151.765 ;
        RECT 140.315 151.425 140.530 152.540 ;
        RECT 140.725 151.840 141.055 152.615 ;
        RECT 141.225 152.010 141.935 152.785 ;
        RECT 140.725 151.625 141.875 151.840 ;
        RECT 139.795 151.225 140.125 151.425 ;
        RECT 140.315 151.245 140.765 151.425 ;
        RECT 140.435 151.225 140.765 151.245 ;
        RECT 140.935 151.225 141.405 151.455 ;
        RECT 141.590 151.055 141.875 151.625 ;
        RECT 142.105 151.180 142.385 152.615 ;
        RECT 143.475 152.190 143.910 152.615 ;
        RECT 144.080 152.360 144.465 152.785 ;
        RECT 143.475 152.020 144.465 152.190 ;
        RECT 135.195 150.235 135.485 150.960 ;
        RECT 135.815 150.795 136.325 150.975 ;
        RECT 136.730 150.885 138.430 151.055 ;
        RECT 136.730 150.795 137.115 150.885 ;
        RECT 135.815 150.405 136.145 150.795 ;
        RECT 136.315 150.455 137.500 150.625 ;
        RECT 137.760 150.235 137.930 150.705 ;
        RECT 138.100 150.420 138.430 150.885 ;
        RECT 138.600 150.235 138.770 151.055 ;
        RECT 138.940 150.415 139.625 151.055 ;
        RECT 139.795 150.865 140.975 151.055 ;
        RECT 139.795 150.405 140.135 150.865 ;
        RECT 140.645 150.785 140.975 150.865 ;
        RECT 141.165 150.865 141.875 151.055 ;
        RECT 141.165 150.725 141.465 150.865 ;
        RECT 141.150 150.715 141.465 150.725 ;
        RECT 141.140 150.705 141.465 150.715 ;
        RECT 141.130 150.700 141.465 150.705 ;
        RECT 140.305 150.235 140.475 150.695 ;
        RECT 141.125 150.690 141.465 150.700 ;
        RECT 141.120 150.685 141.465 150.690 ;
        RECT 141.115 150.675 141.465 150.685 ;
        RECT 141.110 150.670 141.465 150.675 ;
        RECT 141.105 150.405 141.465 150.670 ;
        RECT 141.705 150.235 141.875 150.695 ;
        RECT 142.045 150.405 142.385 151.180 ;
        RECT 143.475 151.145 143.960 151.850 ;
        RECT 144.130 151.475 144.465 152.020 ;
        RECT 144.635 151.825 145.060 152.615 ;
        RECT 145.230 152.190 145.505 152.615 ;
        RECT 145.675 152.360 146.060 152.785 ;
        RECT 145.230 151.995 146.060 152.190 ;
        RECT 144.635 151.645 145.540 151.825 ;
        RECT 144.130 151.145 144.540 151.475 ;
        RECT 144.710 151.145 145.540 151.645 ;
        RECT 145.710 151.475 146.060 151.995 ;
        RECT 146.230 151.825 146.475 152.615 ;
        RECT 146.665 152.190 146.920 152.615 ;
        RECT 147.090 152.360 147.475 152.785 ;
        RECT 146.665 151.995 147.475 152.190 ;
        RECT 146.230 151.645 146.955 151.825 ;
        RECT 145.710 151.145 146.135 151.475 ;
        RECT 146.305 151.145 146.955 151.645 ;
        RECT 147.125 151.475 147.475 151.995 ;
        RECT 147.645 151.645 147.905 152.615 ;
        RECT 148.075 151.645 148.355 152.785 ;
        RECT 147.125 151.145 147.550 151.475 ;
        RECT 144.130 150.975 144.465 151.145 ;
        RECT 144.710 150.975 145.060 151.145 ;
        RECT 145.710 150.975 146.060 151.145 ;
        RECT 146.305 150.975 146.475 151.145 ;
        RECT 147.125 150.975 147.475 151.145 ;
        RECT 147.720 150.975 147.905 151.645 ;
        RECT 148.525 151.635 148.855 152.615 ;
        RECT 149.025 151.645 149.285 152.785 ;
        RECT 149.455 151.645 149.715 152.785 ;
        RECT 149.885 151.635 150.215 152.615 ;
        RECT 150.385 151.645 150.665 152.785 ;
        RECT 150.875 151.645 151.105 152.785 ;
        RECT 151.275 151.635 151.605 152.615 ;
        RECT 151.775 151.645 151.985 152.785 ;
        RECT 152.215 151.710 152.485 152.615 ;
        RECT 152.655 152.025 152.985 152.785 ;
        RECT 153.165 151.855 153.345 152.615 ;
        RECT 148.085 151.205 148.420 151.475 ;
        RECT 148.590 151.035 148.760 151.635 ;
        RECT 148.930 151.225 149.265 151.475 ;
        RECT 149.475 151.225 149.810 151.475 ;
        RECT 149.980 151.035 150.150 151.635 ;
        RECT 150.320 151.205 150.655 151.475 ;
        RECT 150.855 151.225 151.185 151.475 ;
        RECT 143.475 150.805 144.465 150.975 ;
        RECT 143.475 150.405 143.910 150.805 ;
        RECT 144.080 150.235 144.465 150.635 ;
        RECT 144.635 150.405 145.060 150.975 ;
        RECT 145.250 150.805 146.060 150.975 ;
        RECT 145.250 150.405 145.505 150.805 ;
        RECT 145.675 150.235 146.060 150.635 ;
        RECT 146.230 150.405 146.475 150.975 ;
        RECT 146.665 150.805 147.475 150.975 ;
        RECT 146.665 150.405 146.920 150.805 ;
        RECT 147.090 150.235 147.475 150.635 ;
        RECT 147.645 150.405 147.905 150.975 ;
        RECT 148.075 150.235 148.385 151.035 ;
        RECT 148.590 150.405 149.285 151.035 ;
        RECT 149.455 150.405 150.150 151.035 ;
        RECT 150.355 150.235 150.665 151.035 ;
        RECT 150.875 150.235 151.105 151.055 ;
        RECT 151.355 151.035 151.605 151.635 ;
        RECT 151.275 150.405 151.605 151.035 ;
        RECT 151.775 150.235 151.985 151.055 ;
        RECT 152.215 150.910 152.395 151.710 ;
        RECT 152.670 151.685 153.345 151.855 ;
        RECT 153.595 151.695 154.805 152.785 ;
        RECT 152.670 151.540 152.840 151.685 ;
        RECT 152.565 151.210 152.840 151.540 ;
        RECT 152.670 150.955 152.840 151.210 ;
        RECT 153.065 151.135 153.405 151.505 ;
        RECT 153.595 150.985 154.115 151.525 ;
        RECT 154.285 151.155 154.805 151.695 ;
        RECT 154.975 151.695 156.185 152.785 ;
        RECT 154.975 151.155 155.495 151.695 ;
        RECT 155.665 150.985 156.185 151.525 ;
        RECT 152.215 150.405 152.475 150.910 ;
        RECT 152.670 150.785 153.335 150.955 ;
        RECT 152.655 150.235 152.985 150.615 ;
        RECT 153.165 150.405 153.335 150.785 ;
        RECT 153.595 150.235 154.805 150.985 ;
        RECT 154.975 150.235 156.185 150.985 ;
        RECT 70.710 150.065 156.270 150.235 ;
        RECT 70.795 149.315 72.005 150.065 ;
        RECT 72.265 149.515 72.435 149.805 ;
        RECT 72.605 149.685 72.935 150.065 ;
        RECT 72.265 149.345 72.930 149.515 ;
        RECT 70.795 148.775 71.315 149.315 ;
        RECT 71.485 148.605 72.005 149.145 ;
        RECT 70.795 147.515 72.005 148.605 ;
        RECT 72.180 148.525 72.530 149.175 ;
        RECT 72.700 148.355 72.930 149.345 ;
        RECT 72.265 148.185 72.930 148.355 ;
        RECT 72.265 147.685 72.435 148.185 ;
        RECT 72.605 147.515 72.935 148.015 ;
        RECT 73.105 147.685 73.290 149.805 ;
        RECT 73.545 149.605 73.795 150.065 ;
        RECT 73.965 149.615 74.300 149.785 ;
        RECT 74.495 149.615 75.170 149.785 ;
        RECT 73.965 149.475 74.135 149.615 ;
        RECT 73.460 148.485 73.740 149.435 ;
        RECT 73.910 149.345 74.135 149.475 ;
        RECT 73.910 148.240 74.080 149.345 ;
        RECT 74.305 149.195 74.830 149.415 ;
        RECT 74.250 148.430 74.490 149.025 ;
        RECT 74.660 148.495 74.830 149.195 ;
        RECT 75.000 148.835 75.170 149.615 ;
        RECT 75.490 149.565 75.860 150.065 ;
        RECT 76.040 149.615 76.445 149.785 ;
        RECT 76.615 149.615 77.400 149.785 ;
        RECT 76.040 149.385 76.210 149.615 ;
        RECT 75.380 149.085 76.210 149.385 ;
        RECT 76.595 149.115 77.060 149.445 ;
        RECT 75.380 149.055 75.580 149.085 ;
        RECT 75.700 148.835 75.870 148.905 ;
        RECT 75.000 148.665 75.870 148.835 ;
        RECT 75.360 148.575 75.870 148.665 ;
        RECT 73.910 148.110 74.215 148.240 ;
        RECT 74.660 148.130 75.190 148.495 ;
        RECT 73.530 147.515 73.795 147.975 ;
        RECT 73.965 147.685 74.215 148.110 ;
        RECT 75.360 147.960 75.530 148.575 ;
        RECT 74.425 147.790 75.530 147.960 ;
        RECT 75.700 147.515 75.870 148.315 ;
        RECT 76.040 148.015 76.210 149.085 ;
        RECT 76.380 148.185 76.570 148.905 ;
        RECT 76.740 148.155 77.060 149.115 ;
        RECT 77.230 149.155 77.400 149.615 ;
        RECT 77.675 149.535 77.885 150.065 ;
        RECT 78.145 149.325 78.475 149.850 ;
        RECT 78.645 149.455 78.815 150.065 ;
        RECT 78.985 149.410 79.315 149.845 ;
        RECT 78.985 149.325 79.365 149.410 ;
        RECT 78.275 149.155 78.475 149.325 ;
        RECT 79.140 149.285 79.365 149.325 ;
        RECT 77.230 148.825 78.105 149.155 ;
        RECT 78.275 148.825 79.025 149.155 ;
        RECT 76.040 147.685 76.290 148.015 ;
        RECT 77.230 147.985 77.400 148.825 ;
        RECT 78.275 148.620 78.465 148.825 ;
        RECT 79.195 148.705 79.365 149.285 ;
        RECT 80.465 149.255 80.735 150.065 ;
        RECT 80.905 149.255 81.235 149.895 ;
        RECT 81.405 149.255 81.645 150.065 ;
        RECT 81.845 149.335 82.145 150.065 ;
        RECT 80.455 148.825 80.805 149.075 ;
        RECT 79.150 148.655 79.365 148.705 ;
        RECT 80.975 148.655 81.145 149.255 ;
        RECT 82.325 149.155 82.555 149.775 ;
        RECT 82.755 149.505 82.980 149.885 ;
        RECT 83.150 149.675 83.480 150.065 ;
        RECT 84.135 149.605 84.695 149.895 ;
        RECT 84.865 149.605 85.115 150.065 ;
        RECT 82.755 149.325 83.085 149.505 ;
        RECT 81.315 148.825 81.665 149.075 ;
        RECT 81.850 148.825 82.145 149.155 ;
        RECT 82.325 148.825 82.740 149.155 ;
        RECT 82.910 148.655 83.085 149.325 ;
        RECT 83.255 148.825 83.495 149.475 ;
        RECT 77.570 148.245 78.465 148.620 ;
        RECT 78.975 148.575 79.365 148.655 ;
        RECT 76.515 147.815 77.400 147.985 ;
        RECT 77.580 147.515 77.895 148.015 ;
        RECT 78.125 147.685 78.465 148.245 ;
        RECT 78.635 147.515 78.805 148.525 ;
        RECT 78.975 147.730 79.305 148.575 ;
        RECT 80.465 147.515 80.795 148.655 ;
        RECT 80.975 148.485 81.655 148.655 ;
        RECT 81.325 147.700 81.655 148.485 ;
        RECT 81.845 148.295 82.740 148.625 ;
        RECT 82.910 148.465 83.495 148.655 ;
        RECT 81.845 148.125 83.050 148.295 ;
        RECT 81.845 147.695 82.175 148.125 ;
        RECT 82.355 147.515 82.550 147.955 ;
        RECT 82.720 147.695 83.050 148.125 ;
        RECT 83.220 147.695 83.495 148.465 ;
        RECT 84.135 148.235 84.385 149.605 ;
        RECT 85.735 149.435 86.065 149.795 ;
        RECT 84.675 149.245 86.065 149.435 ;
        RECT 86.525 149.385 86.695 149.760 ;
        RECT 84.675 149.155 84.845 149.245 ;
        RECT 86.495 149.215 86.695 149.385 ;
        RECT 86.885 149.535 87.115 149.840 ;
        RECT 87.285 149.705 87.615 150.065 ;
        RECT 87.810 149.535 88.100 149.885 ;
        RECT 86.885 149.365 88.100 149.535 ;
        RECT 88.275 149.495 88.710 149.895 ;
        RECT 88.880 149.665 89.265 150.065 ;
        RECT 88.275 149.325 89.265 149.495 ;
        RECT 89.435 149.325 89.860 149.895 ;
        RECT 90.050 149.495 90.305 149.895 ;
        RECT 90.475 149.665 90.860 150.065 ;
        RECT 90.050 149.325 90.860 149.495 ;
        RECT 91.030 149.325 91.275 149.895 ;
        RECT 91.465 149.495 91.720 149.895 ;
        RECT 91.890 149.665 92.275 150.065 ;
        RECT 91.465 149.325 92.275 149.495 ;
        RECT 92.445 149.325 92.705 149.895 ;
        RECT 84.555 148.825 84.845 149.155 ;
        RECT 86.525 149.195 86.695 149.215 ;
        RECT 85.015 148.825 85.355 149.075 ;
        RECT 85.575 148.825 86.250 149.075 ;
        RECT 86.525 149.025 87.045 149.195 ;
        RECT 88.930 149.155 89.265 149.325 ;
        RECT 89.510 149.155 89.860 149.325 ;
        RECT 90.510 149.155 90.860 149.325 ;
        RECT 91.105 149.155 91.275 149.325 ;
        RECT 91.925 149.155 92.275 149.325 ;
        RECT 84.675 148.575 84.845 148.825 ;
        RECT 84.675 148.405 85.615 148.575 ;
        RECT 85.985 148.465 86.250 148.825 ;
        RECT 86.440 148.495 86.685 148.855 ;
        RECT 86.875 148.645 87.045 149.025 ;
        RECT 87.215 148.825 87.600 149.155 ;
        RECT 87.780 149.045 88.040 149.155 ;
        RECT 87.780 148.875 88.045 149.045 ;
        RECT 87.780 148.825 88.040 148.875 ;
        RECT 84.135 147.685 84.595 148.235 ;
        RECT 84.785 147.515 85.115 148.235 ;
        RECT 85.315 147.855 85.615 148.405 ;
        RECT 86.875 148.365 87.225 148.645 ;
        RECT 85.785 147.515 86.065 148.185 ;
        RECT 86.440 147.515 86.695 148.315 ;
        RECT 86.895 147.685 87.225 148.365 ;
        RECT 87.405 147.775 87.600 148.825 ;
        RECT 87.780 147.515 88.100 148.655 ;
        RECT 88.275 148.450 88.760 149.155 ;
        RECT 88.930 148.825 89.340 149.155 ;
        RECT 88.930 148.280 89.265 148.825 ;
        RECT 89.510 148.655 90.340 149.155 ;
        RECT 88.275 148.110 89.265 148.280 ;
        RECT 89.435 148.475 90.340 148.655 ;
        RECT 90.510 148.825 90.935 149.155 ;
        RECT 88.275 147.685 88.710 148.110 ;
        RECT 88.880 147.515 89.265 147.940 ;
        RECT 89.435 147.685 89.860 148.475 ;
        RECT 90.510 148.305 90.860 148.825 ;
        RECT 91.105 148.655 91.755 149.155 ;
        RECT 90.030 148.110 90.860 148.305 ;
        RECT 91.030 148.475 91.755 148.655 ;
        RECT 91.925 148.825 92.350 149.155 ;
        RECT 90.030 147.685 90.305 148.110 ;
        RECT 90.475 147.515 90.860 147.940 ;
        RECT 91.030 147.685 91.275 148.475 ;
        RECT 91.925 148.305 92.275 148.825 ;
        RECT 92.520 148.655 92.705 149.325 ;
        RECT 92.875 149.295 96.385 150.065 ;
        RECT 96.555 149.340 96.845 150.065 ;
        RECT 92.875 148.775 94.525 149.295 ;
        RECT 97.015 149.245 97.700 149.885 ;
        RECT 97.870 149.245 98.040 150.065 ;
        RECT 98.210 149.415 98.540 149.880 ;
        RECT 98.710 149.595 98.880 150.065 ;
        RECT 99.140 149.675 100.325 149.845 ;
        RECT 100.495 149.505 100.825 149.895 ;
        RECT 99.525 149.415 99.910 149.505 ;
        RECT 98.210 149.245 99.910 149.415 ;
        RECT 100.315 149.325 100.825 149.505 ;
        RECT 91.465 148.110 92.275 148.305 ;
        RECT 91.465 147.685 91.720 148.110 ;
        RECT 91.890 147.515 92.275 147.940 ;
        RECT 92.445 147.685 92.705 148.655 ;
        RECT 94.695 148.605 96.385 149.125 ;
        RECT 92.875 147.515 96.385 148.605 ;
        RECT 96.555 147.515 96.845 148.680 ;
        RECT 97.015 148.275 97.265 149.245 ;
        RECT 97.435 148.865 97.770 149.075 ;
        RECT 97.940 148.865 98.390 149.075 ;
        RECT 98.580 148.865 99.065 149.075 ;
        RECT 97.600 148.695 97.770 148.865 ;
        RECT 98.690 148.705 99.065 148.865 ;
        RECT 99.255 148.825 99.635 149.075 ;
        RECT 99.815 148.865 100.145 149.075 ;
        RECT 97.600 148.525 98.520 148.695 ;
        RECT 97.015 147.685 97.680 148.275 ;
        RECT 97.850 147.515 98.180 148.355 ;
        RECT 98.350 148.275 98.520 148.525 ;
        RECT 98.690 148.535 99.085 148.705 ;
        RECT 98.690 148.445 99.065 148.535 ;
        RECT 99.255 148.445 99.575 148.825 ;
        RECT 100.315 148.695 100.485 149.325 ;
        RECT 101.155 149.315 102.365 150.065 ;
        RECT 100.655 148.865 100.985 149.155 ;
        RECT 101.155 148.775 101.675 149.315 ;
        RECT 99.745 148.525 100.830 148.695 ;
        RECT 101.845 148.605 102.365 149.145 ;
        RECT 99.745 148.275 99.915 148.525 ;
        RECT 98.350 148.105 99.915 148.275 ;
        RECT 98.690 147.685 99.495 148.105 ;
        RECT 100.085 147.515 100.335 148.355 ;
        RECT 100.530 147.685 100.830 148.525 ;
        RECT 101.155 147.515 102.365 148.605 ;
        RECT 102.535 149.120 102.875 149.895 ;
        RECT 103.045 149.605 103.215 150.065 ;
        RECT 103.455 149.630 103.815 149.895 ;
        RECT 103.455 149.625 103.810 149.630 ;
        RECT 103.455 149.615 103.805 149.625 ;
        RECT 103.455 149.610 103.800 149.615 ;
        RECT 103.455 149.600 103.795 149.610 ;
        RECT 104.445 149.605 104.615 150.065 ;
        RECT 103.455 149.595 103.790 149.600 ;
        RECT 103.455 149.585 103.780 149.595 ;
        RECT 103.455 149.575 103.770 149.585 ;
        RECT 103.455 149.435 103.755 149.575 ;
        RECT 103.045 149.245 103.755 149.435 ;
        RECT 103.945 149.435 104.275 149.515 ;
        RECT 104.785 149.435 105.125 149.895 ;
        RECT 105.295 149.520 110.640 150.065 ;
        RECT 103.945 149.245 105.125 149.435 ;
        RECT 102.535 147.685 102.815 149.120 ;
        RECT 103.045 148.675 103.330 149.245 ;
        RECT 103.515 148.845 103.985 149.075 ;
        RECT 104.155 149.055 104.485 149.075 ;
        RECT 104.155 148.875 104.605 149.055 ;
        RECT 104.795 148.875 105.125 149.075 ;
        RECT 103.045 148.460 104.195 148.675 ;
        RECT 102.985 147.515 103.695 148.290 ;
        RECT 103.865 147.685 104.195 148.460 ;
        RECT 104.390 147.760 104.605 148.875 ;
        RECT 104.895 148.535 105.125 148.875 ;
        RECT 106.880 148.690 107.220 149.520 ;
        RECT 110.815 149.295 113.405 150.065 ;
        RECT 113.575 149.435 113.915 149.895 ;
        RECT 114.085 149.605 114.255 150.065 ;
        RECT 114.885 149.630 115.245 149.895 ;
        RECT 114.890 149.625 115.245 149.630 ;
        RECT 114.895 149.615 115.245 149.625 ;
        RECT 114.900 149.610 115.245 149.615 ;
        RECT 114.905 149.600 115.245 149.610 ;
        RECT 115.485 149.605 115.655 150.065 ;
        RECT 114.910 149.595 115.245 149.600 ;
        RECT 114.920 149.585 115.245 149.595 ;
        RECT 114.930 149.575 115.245 149.585 ;
        RECT 114.425 149.435 114.755 149.515 ;
        RECT 104.785 147.515 105.115 148.235 ;
        RECT 108.700 147.950 109.050 149.200 ;
        RECT 110.815 148.775 112.025 149.295 ;
        RECT 113.575 149.245 114.755 149.435 ;
        RECT 114.945 149.435 115.245 149.575 ;
        RECT 114.945 149.245 115.655 149.435 ;
        RECT 112.195 148.605 113.405 149.125 ;
        RECT 105.295 147.515 110.640 147.950 ;
        RECT 110.815 147.515 113.405 148.605 ;
        RECT 113.575 148.875 113.905 149.075 ;
        RECT 114.215 149.055 114.545 149.075 ;
        RECT 114.095 148.875 114.545 149.055 ;
        RECT 113.575 148.535 113.805 148.875 ;
        RECT 113.585 147.515 113.915 148.235 ;
        RECT 114.095 147.760 114.310 148.875 ;
        RECT 114.715 148.845 115.185 149.075 ;
        RECT 115.370 148.675 115.655 149.245 ;
        RECT 115.825 149.120 116.165 149.895 ;
        RECT 114.505 148.460 115.655 148.675 ;
        RECT 114.505 147.685 114.835 148.460 ;
        RECT 115.005 147.515 115.715 148.290 ;
        RECT 115.885 147.685 116.165 149.120 ;
        RECT 116.370 149.325 116.985 149.895 ;
        RECT 117.155 149.555 117.370 150.065 ;
        RECT 117.600 149.555 117.880 149.885 ;
        RECT 118.060 149.555 118.300 150.065 ;
        RECT 116.370 148.305 116.685 149.325 ;
        RECT 116.855 148.655 117.025 149.155 ;
        RECT 117.275 148.825 117.540 149.385 ;
        RECT 117.710 148.655 117.880 149.555 ;
        RECT 118.635 149.390 118.895 149.895 ;
        RECT 119.075 149.685 119.405 150.065 ;
        RECT 119.585 149.515 119.755 149.895 ;
        RECT 118.050 148.825 118.405 149.385 ;
        RECT 116.855 148.485 118.280 148.655 ;
        RECT 116.370 147.685 116.905 148.305 ;
        RECT 117.075 147.515 117.405 148.315 ;
        RECT 117.890 148.310 118.280 148.485 ;
        RECT 118.635 148.590 118.815 149.390 ;
        RECT 119.090 149.345 119.755 149.515 ;
        RECT 119.090 149.090 119.260 149.345 ;
        RECT 120.015 149.295 121.685 150.065 ;
        RECT 122.315 149.340 122.605 150.065 ;
        RECT 122.775 149.295 126.285 150.065 ;
        RECT 126.455 149.315 127.665 150.065 ;
        RECT 118.985 148.760 119.260 149.090 ;
        RECT 119.485 148.795 119.825 149.165 ;
        RECT 120.015 148.775 120.765 149.295 ;
        RECT 119.090 148.615 119.260 148.760 ;
        RECT 118.635 147.685 118.905 148.590 ;
        RECT 119.090 148.445 119.765 148.615 ;
        RECT 120.935 148.605 121.685 149.125 ;
        RECT 122.775 148.775 124.425 149.295 ;
        RECT 119.075 147.515 119.405 148.275 ;
        RECT 119.585 147.685 119.765 148.445 ;
        RECT 120.015 147.515 121.685 148.605 ;
        RECT 122.315 147.515 122.605 148.680 ;
        RECT 124.595 148.605 126.285 149.125 ;
        RECT 126.455 148.775 126.975 149.315 ;
        RECT 128.040 149.285 128.540 149.895 ;
        RECT 127.145 148.605 127.665 149.145 ;
        RECT 127.835 148.825 128.185 149.075 ;
        RECT 128.370 148.655 128.540 149.285 ;
        RECT 129.170 149.415 129.500 149.895 ;
        RECT 129.670 149.605 129.895 150.065 ;
        RECT 130.065 149.415 130.395 149.895 ;
        RECT 129.170 149.245 130.395 149.415 ;
        RECT 130.585 149.265 130.835 150.065 ;
        RECT 131.005 149.265 131.345 149.895 ;
        RECT 128.710 148.875 129.040 149.075 ;
        RECT 129.210 148.875 129.540 149.075 ;
        RECT 129.710 148.875 130.130 149.075 ;
        RECT 130.305 148.905 131.000 149.075 ;
        RECT 130.305 148.655 130.475 148.905 ;
        RECT 131.170 148.655 131.345 149.265 ;
        RECT 122.775 147.515 126.285 148.605 ;
        RECT 126.455 147.515 127.665 148.605 ;
        RECT 128.040 148.485 130.475 148.655 ;
        RECT 128.040 147.685 128.370 148.485 ;
        RECT 128.540 147.515 128.870 148.315 ;
        RECT 129.170 147.685 129.500 148.485 ;
        RECT 130.145 147.515 130.395 148.315 ;
        RECT 130.665 147.515 130.835 148.655 ;
        RECT 131.005 147.685 131.345 148.655 ;
        RECT 131.515 147.685 131.795 149.785 ;
        RECT 132.025 149.605 132.195 150.065 ;
        RECT 132.465 149.675 133.715 149.855 ;
        RECT 132.850 149.435 133.215 149.505 ;
        RECT 131.965 149.255 133.215 149.435 ;
        RECT 133.385 149.455 133.715 149.675 ;
        RECT 133.885 149.625 134.055 150.065 ;
        RECT 134.225 149.455 134.565 149.870 ;
        RECT 133.385 149.285 134.565 149.455 ;
        RECT 131.965 148.655 132.240 149.255 ;
        RECT 132.410 148.825 132.765 149.075 ;
        RECT 132.960 149.045 133.425 149.075 ;
        RECT 132.955 148.875 133.425 149.045 ;
        RECT 132.960 148.825 133.425 148.875 ;
        RECT 133.595 148.825 133.925 149.075 ;
        RECT 134.100 148.875 134.565 149.075 ;
        RECT 133.745 148.705 133.925 148.825 ;
        RECT 131.965 148.445 133.575 148.655 ;
        RECT 133.745 148.535 134.075 148.705 ;
        RECT 133.165 148.345 133.575 148.445 ;
        RECT 131.985 147.515 132.770 148.275 ;
        RECT 133.165 147.685 133.550 148.345 ;
        RECT 133.875 147.745 134.075 148.535 ;
        RECT 134.245 147.515 134.565 148.695 ;
        RECT 134.735 147.685 135.015 149.785 ;
        RECT 135.245 149.605 135.415 150.065 ;
        RECT 135.685 149.675 136.935 149.855 ;
        RECT 136.070 149.435 136.435 149.505 ;
        RECT 135.185 149.255 136.435 149.435 ;
        RECT 136.605 149.455 136.935 149.675 ;
        RECT 137.105 149.625 137.275 150.065 ;
        RECT 137.445 149.455 137.785 149.870 ;
        RECT 136.605 149.285 137.785 149.455 ;
        RECT 137.955 149.295 140.545 150.065 ;
        RECT 141.175 149.390 141.435 149.895 ;
        RECT 141.615 149.685 141.945 150.065 ;
        RECT 142.125 149.515 142.295 149.895 ;
        RECT 135.185 148.655 135.460 149.255 ;
        RECT 135.630 148.825 135.985 149.075 ;
        RECT 136.180 149.045 136.645 149.075 ;
        RECT 136.175 148.875 136.645 149.045 ;
        RECT 136.180 148.825 136.645 148.875 ;
        RECT 136.815 148.825 137.145 149.075 ;
        RECT 137.320 148.875 137.785 149.075 ;
        RECT 136.965 148.705 137.145 148.825 ;
        RECT 137.955 148.775 139.165 149.295 ;
        RECT 135.185 148.445 136.795 148.655 ;
        RECT 136.965 148.535 137.295 148.705 ;
        RECT 136.385 148.345 136.795 148.445 ;
        RECT 135.205 147.515 135.990 148.275 ;
        RECT 136.385 147.685 136.770 148.345 ;
        RECT 137.095 147.745 137.295 148.535 ;
        RECT 137.465 147.515 137.785 148.695 ;
        RECT 139.335 148.605 140.545 149.125 ;
        RECT 137.955 147.515 140.545 148.605 ;
        RECT 141.175 148.590 141.355 149.390 ;
        RECT 141.630 149.345 142.295 149.515 ;
        RECT 142.555 149.390 142.815 149.895 ;
        RECT 142.995 149.685 143.325 150.065 ;
        RECT 143.505 149.515 143.675 149.895 ;
        RECT 141.630 149.090 141.800 149.345 ;
        RECT 141.525 148.760 141.800 149.090 ;
        RECT 142.025 148.795 142.365 149.165 ;
        RECT 141.630 148.615 141.800 148.760 ;
        RECT 141.175 147.685 141.445 148.590 ;
        RECT 141.630 148.445 142.305 148.615 ;
        RECT 141.615 147.515 141.945 148.275 ;
        RECT 142.125 147.685 142.305 148.445 ;
        RECT 142.555 148.590 142.735 149.390 ;
        RECT 143.010 149.345 143.675 149.515 ;
        RECT 143.010 149.090 143.180 149.345 ;
        RECT 143.935 149.245 144.620 149.885 ;
        RECT 144.790 149.245 144.960 150.065 ;
        RECT 145.130 149.415 145.460 149.880 ;
        RECT 145.630 149.595 145.800 150.065 ;
        RECT 146.060 149.675 147.245 149.845 ;
        RECT 147.415 149.505 147.745 149.895 ;
        RECT 146.445 149.415 146.830 149.505 ;
        RECT 145.130 149.245 146.830 149.415 ;
        RECT 147.235 149.325 147.745 149.505 ;
        RECT 148.075 149.340 148.365 150.065 ;
        RECT 142.905 148.760 143.180 149.090 ;
        RECT 143.405 148.795 143.745 149.165 ;
        RECT 143.010 148.615 143.180 148.760 ;
        RECT 142.555 147.685 142.825 148.590 ;
        RECT 143.010 148.445 143.685 148.615 ;
        RECT 142.995 147.515 143.325 148.275 ;
        RECT 143.505 147.685 143.685 148.445 ;
        RECT 143.935 148.275 144.185 149.245 ;
        RECT 144.355 148.865 144.690 149.075 ;
        RECT 144.860 148.865 145.310 149.075 ;
        RECT 145.500 149.045 145.985 149.075 ;
        RECT 145.500 148.875 146.005 149.045 ;
        RECT 145.500 148.865 145.985 148.875 ;
        RECT 144.520 148.695 144.690 148.865 ;
        RECT 144.520 148.525 145.440 148.695 ;
        RECT 143.935 147.685 144.600 148.275 ;
        RECT 144.770 147.515 145.100 148.355 ;
        RECT 145.270 148.275 145.440 148.525 ;
        RECT 145.610 148.445 145.985 148.865 ;
        RECT 146.175 148.825 146.555 149.075 ;
        RECT 146.735 148.865 147.065 149.075 ;
        RECT 146.175 148.445 146.495 148.825 ;
        RECT 147.235 148.695 147.405 149.325 ;
        RECT 148.595 149.245 148.805 150.065 ;
        RECT 148.975 149.265 149.305 149.895 ;
        RECT 147.575 148.865 147.905 149.155 ;
        RECT 146.665 148.525 147.750 148.695 ;
        RECT 146.665 148.275 146.835 148.525 ;
        RECT 145.270 148.105 146.835 148.275 ;
        RECT 145.610 147.685 146.415 148.105 ;
        RECT 147.005 147.515 147.255 148.355 ;
        RECT 147.450 147.685 147.750 148.525 ;
        RECT 148.075 147.515 148.365 148.680 ;
        RECT 148.975 148.665 149.225 149.265 ;
        RECT 149.475 149.245 149.705 150.065 ;
        RECT 150.380 149.245 150.655 150.065 ;
        RECT 150.825 149.425 151.155 149.895 ;
        RECT 151.325 149.595 151.495 150.065 ;
        RECT 151.665 149.425 151.995 149.895 ;
        RECT 152.165 149.595 152.455 150.065 ;
        RECT 150.825 149.415 151.995 149.425 ;
        RECT 150.825 149.245 152.425 149.415 ;
        RECT 152.695 149.255 152.935 150.065 ;
        RECT 153.105 149.255 153.435 149.895 ;
        RECT 153.605 149.255 153.875 150.065 ;
        RECT 154.975 149.315 156.185 150.065 ;
        RECT 149.395 148.825 149.725 149.075 ;
        RECT 150.380 148.875 151.100 149.075 ;
        RECT 151.270 148.875 152.040 149.075 ;
        RECT 152.210 148.705 152.425 149.245 ;
        RECT 152.675 148.825 153.025 149.075 ;
        RECT 148.595 147.515 148.805 148.655 ;
        RECT 148.975 147.685 149.305 148.665 ;
        RECT 149.475 147.515 149.705 148.655 ;
        RECT 150.380 148.485 151.495 148.695 ;
        RECT 150.380 147.685 150.655 148.485 ;
        RECT 150.825 147.515 151.155 148.315 ;
        RECT 151.325 147.855 151.495 148.485 ;
        RECT 151.665 148.485 152.425 148.705 ;
        RECT 153.195 148.655 153.365 149.255 ;
        RECT 153.535 148.825 153.885 149.075 ;
        RECT 152.685 148.485 153.365 148.655 ;
        RECT 151.665 148.025 151.995 148.485 ;
        RECT 152.165 147.855 152.465 148.315 ;
        RECT 151.325 147.685 152.465 147.855 ;
        RECT 152.685 147.700 153.015 148.485 ;
        RECT 153.545 147.515 153.875 148.655 ;
        RECT 154.975 148.605 155.495 149.145 ;
        RECT 155.665 148.775 156.185 149.315 ;
        RECT 154.975 147.515 156.185 148.605 ;
        RECT 70.710 147.345 156.270 147.515 ;
        RECT 70.795 146.255 72.005 147.345 ;
        RECT 70.795 145.545 71.315 146.085 ;
        RECT 71.485 145.715 72.005 146.255 ;
        RECT 72.175 146.205 72.455 147.345 ;
        RECT 72.625 146.195 72.955 147.175 ;
        RECT 73.125 146.205 73.385 147.345 ;
        RECT 73.615 146.205 73.825 147.345 ;
        RECT 73.995 146.195 74.325 147.175 ;
        RECT 74.495 146.205 74.725 147.345 ;
        RECT 75.120 146.375 75.510 146.550 ;
        RECT 75.995 146.545 76.325 147.345 ;
        RECT 76.495 146.555 77.030 147.175 ;
        RECT 75.120 146.205 76.545 146.375 ;
        RECT 72.185 145.765 72.520 146.035 ;
        RECT 72.690 145.595 72.860 146.195 ;
        RECT 73.030 145.785 73.365 146.035 ;
        RECT 70.795 144.795 72.005 145.545 ;
        RECT 72.175 144.795 72.485 145.595 ;
        RECT 72.690 144.965 73.385 145.595 ;
        RECT 73.615 144.795 73.825 145.615 ;
        RECT 73.995 145.595 74.245 146.195 ;
        RECT 74.415 145.785 74.745 146.035 ;
        RECT 73.995 144.965 74.325 145.595 ;
        RECT 74.495 144.795 74.725 145.615 ;
        RECT 74.995 145.475 75.350 146.035 ;
        RECT 75.520 145.305 75.690 146.205 ;
        RECT 75.860 145.475 76.125 146.035 ;
        RECT 76.375 145.705 76.545 146.205 ;
        RECT 76.715 145.535 77.030 146.555 ;
        RECT 75.100 144.795 75.340 145.305 ;
        RECT 75.520 144.975 75.800 145.305 ;
        RECT 76.030 144.795 76.245 145.305 ;
        RECT 76.415 144.965 77.030 145.535 ;
        RECT 77.235 146.475 77.510 147.175 ;
        RECT 77.680 146.800 77.935 147.345 ;
        RECT 78.105 146.835 78.585 147.175 ;
        RECT 78.760 146.790 79.365 147.345 ;
        RECT 78.750 146.690 79.365 146.790 ;
        RECT 78.750 146.665 78.935 146.690 ;
        RECT 77.235 145.445 77.405 146.475 ;
        RECT 77.680 146.345 78.435 146.595 ;
        RECT 78.605 146.420 78.935 146.665 ;
        RECT 77.680 146.310 78.450 146.345 ;
        RECT 77.680 146.300 78.465 146.310 ;
        RECT 77.575 146.285 78.470 146.300 ;
        RECT 77.575 146.270 78.490 146.285 ;
        RECT 77.575 146.260 78.510 146.270 ;
        RECT 77.575 146.250 78.535 146.260 ;
        RECT 77.575 146.220 78.605 146.250 ;
        RECT 77.575 146.190 78.625 146.220 ;
        RECT 77.575 146.160 78.645 146.190 ;
        RECT 77.575 146.135 78.675 146.160 ;
        RECT 77.575 146.100 78.710 146.135 ;
        RECT 77.575 146.095 78.740 146.100 ;
        RECT 77.575 145.700 77.805 146.095 ;
        RECT 78.350 146.090 78.740 146.095 ;
        RECT 78.375 146.080 78.740 146.090 ;
        RECT 78.390 146.075 78.740 146.080 ;
        RECT 78.405 146.070 78.740 146.075 ;
        RECT 79.105 146.070 79.365 146.520 ;
        RECT 79.540 146.205 79.795 147.345 ;
        RECT 79.965 146.375 80.295 147.175 ;
        RECT 80.465 146.545 80.695 147.345 ;
        RECT 80.865 146.375 81.195 147.175 ;
        RECT 79.965 146.205 81.195 146.375 ;
        RECT 81.375 146.475 81.650 147.175 ;
        RECT 81.820 146.800 82.075 147.345 ;
        RECT 82.245 146.835 82.725 147.175 ;
        RECT 82.900 146.790 83.505 147.345 ;
        RECT 82.890 146.690 83.505 146.790 ;
        RECT 82.890 146.665 83.075 146.690 ;
        RECT 78.405 146.065 79.365 146.070 ;
        RECT 78.415 146.055 79.365 146.065 ;
        RECT 78.425 146.050 79.365 146.055 ;
        RECT 78.435 146.040 79.365 146.050 ;
        RECT 78.440 146.030 79.365 146.040 ;
        RECT 78.445 146.025 79.365 146.030 ;
        RECT 78.455 146.010 79.365 146.025 ;
        RECT 78.460 145.995 79.365 146.010 ;
        RECT 78.470 145.970 79.365 145.995 ;
        RECT 77.975 145.500 78.305 145.925 ;
        RECT 78.055 145.475 78.305 145.500 ;
        RECT 77.235 144.965 77.495 145.445 ;
        RECT 77.665 144.795 77.915 145.335 ;
        RECT 78.085 145.015 78.305 145.475 ;
        RECT 78.475 145.900 79.365 145.970 ;
        RECT 78.475 145.175 78.645 145.900 ;
        RECT 78.815 145.345 79.365 145.730 ;
        RECT 79.560 145.455 79.780 146.035 ;
        RECT 79.965 145.305 80.145 146.205 ;
        RECT 80.315 145.475 80.690 146.035 ;
        RECT 80.895 145.705 81.205 146.035 ;
        RECT 80.865 145.305 81.195 145.535 ;
        RECT 78.475 145.005 79.365 145.175 ;
        RECT 79.540 144.795 79.795 145.285 ;
        RECT 79.965 144.965 81.195 145.305 ;
        RECT 81.375 145.445 81.545 146.475 ;
        RECT 81.820 146.345 82.575 146.595 ;
        RECT 82.745 146.420 83.075 146.665 ;
        RECT 81.820 146.310 82.590 146.345 ;
        RECT 81.820 146.300 82.605 146.310 ;
        RECT 81.715 146.285 82.610 146.300 ;
        RECT 81.715 146.270 82.630 146.285 ;
        RECT 81.715 146.260 82.650 146.270 ;
        RECT 81.715 146.250 82.675 146.260 ;
        RECT 81.715 146.220 82.745 146.250 ;
        RECT 81.715 146.190 82.765 146.220 ;
        RECT 81.715 146.160 82.785 146.190 ;
        RECT 81.715 146.135 82.815 146.160 ;
        RECT 81.715 146.100 82.850 146.135 ;
        RECT 81.715 146.095 82.880 146.100 ;
        RECT 81.715 145.700 81.945 146.095 ;
        RECT 82.490 146.090 82.880 146.095 ;
        RECT 82.515 146.080 82.880 146.090 ;
        RECT 82.530 146.075 82.880 146.080 ;
        RECT 82.545 146.070 82.880 146.075 ;
        RECT 83.245 146.070 83.505 146.520 ;
        RECT 83.675 146.180 83.965 147.345 ;
        RECT 85.065 146.285 85.395 147.135 ;
        RECT 82.545 146.065 83.505 146.070 ;
        RECT 82.555 146.055 83.505 146.065 ;
        RECT 82.565 146.050 83.505 146.055 ;
        RECT 82.575 146.040 83.505 146.050 ;
        RECT 82.580 146.030 83.505 146.040 ;
        RECT 82.585 146.025 83.505 146.030 ;
        RECT 82.595 146.010 83.505 146.025 ;
        RECT 82.600 145.995 83.505 146.010 ;
        RECT 82.610 145.970 83.505 145.995 ;
        RECT 82.115 145.500 82.445 145.925 ;
        RECT 82.195 145.475 82.445 145.500 ;
        RECT 81.375 144.965 81.635 145.445 ;
        RECT 81.805 144.795 82.055 145.335 ;
        RECT 82.225 145.015 82.445 145.475 ;
        RECT 82.615 145.900 83.505 145.970 ;
        RECT 82.615 145.175 82.785 145.900 ;
        RECT 82.955 145.345 83.505 145.730 ;
        RECT 85.065 145.520 85.255 146.285 ;
        RECT 85.565 146.205 85.815 147.345 ;
        RECT 86.005 146.705 86.255 147.125 ;
        RECT 86.485 146.875 86.815 147.345 ;
        RECT 87.045 146.705 87.295 147.125 ;
        RECT 86.005 146.535 87.295 146.705 ;
        RECT 87.475 146.705 87.805 147.135 ;
        RECT 87.475 146.535 87.930 146.705 ;
        RECT 85.995 146.035 86.210 146.365 ;
        RECT 85.425 145.705 85.735 146.035 ;
        RECT 85.905 145.705 86.210 146.035 ;
        RECT 86.385 145.705 86.670 146.365 ;
        RECT 86.865 145.705 87.130 146.365 ;
        RECT 87.345 145.705 87.590 146.365 ;
        RECT 85.565 145.535 85.735 145.705 ;
        RECT 87.760 145.535 87.930 146.535 ;
        RECT 88.355 146.415 88.535 147.175 ;
        RECT 88.715 146.585 89.045 147.345 ;
        RECT 88.355 146.245 89.030 146.415 ;
        RECT 89.215 146.270 89.485 147.175 ;
        RECT 88.860 146.100 89.030 146.245 ;
        RECT 88.295 145.695 88.635 146.065 ;
        RECT 88.860 145.770 89.135 146.100 ;
        RECT 82.615 145.005 83.505 145.175 ;
        RECT 83.675 144.795 83.965 145.520 ;
        RECT 85.065 145.010 85.395 145.520 ;
        RECT 85.565 145.365 87.930 145.535 ;
        RECT 88.860 145.515 89.030 145.770 ;
        RECT 85.565 144.795 85.895 145.195 ;
        RECT 86.945 145.025 87.275 145.365 ;
        RECT 88.365 145.345 89.030 145.515 ;
        RECT 89.305 145.470 89.485 146.270 ;
        RECT 89.655 146.255 92.245 147.345 ;
        RECT 87.445 144.795 87.775 145.195 ;
        RECT 88.365 144.965 88.535 145.345 ;
        RECT 88.715 144.795 89.045 145.175 ;
        RECT 89.225 144.965 89.485 145.470 ;
        RECT 89.655 145.565 90.865 146.085 ;
        RECT 91.035 145.735 92.245 146.255 ;
        RECT 92.570 146.335 92.870 147.175 ;
        RECT 93.065 146.505 93.315 147.345 ;
        RECT 93.905 146.755 94.710 147.175 ;
        RECT 93.485 146.585 95.050 146.755 ;
        RECT 93.485 146.335 93.655 146.585 ;
        RECT 92.570 146.165 93.655 146.335 ;
        RECT 92.415 145.705 92.745 145.995 ;
        RECT 89.655 144.795 92.245 145.565 ;
        RECT 92.915 145.535 93.085 146.165 ;
        RECT 93.825 146.035 94.145 146.415 ;
        RECT 94.335 146.325 94.710 146.415 ;
        RECT 94.315 146.155 94.710 146.325 ;
        RECT 94.880 146.335 95.050 146.585 ;
        RECT 95.220 146.505 95.550 147.345 ;
        RECT 95.720 146.585 96.385 147.175 ;
        RECT 94.880 146.165 95.800 146.335 ;
        RECT 93.255 145.785 93.585 145.995 ;
        RECT 93.765 145.785 94.145 146.035 ;
        RECT 94.335 145.995 94.710 146.155 ;
        RECT 95.630 145.995 95.800 146.165 ;
        RECT 94.335 145.785 94.820 145.995 ;
        RECT 95.010 145.785 95.460 145.995 ;
        RECT 95.630 145.785 95.965 145.995 ;
        RECT 96.135 145.615 96.385 146.585 ;
        RECT 96.555 146.255 98.225 147.345 ;
        RECT 98.855 146.750 99.290 147.175 ;
        RECT 99.460 146.920 99.845 147.345 ;
        RECT 98.855 146.580 99.845 146.750 ;
        RECT 92.575 145.355 93.085 145.535 ;
        RECT 93.490 145.445 95.190 145.615 ;
        RECT 93.490 145.355 93.875 145.445 ;
        RECT 92.575 144.965 92.905 145.355 ;
        RECT 93.075 145.015 94.260 145.185 ;
        RECT 94.520 144.795 94.690 145.265 ;
        RECT 94.860 144.980 95.190 145.445 ;
        RECT 95.360 144.795 95.530 145.615 ;
        RECT 95.700 144.975 96.385 145.615 ;
        RECT 96.555 145.565 97.305 146.085 ;
        RECT 97.475 145.735 98.225 146.255 ;
        RECT 98.855 145.705 99.340 146.410 ;
        RECT 99.510 146.035 99.845 146.580 ;
        RECT 100.015 146.385 100.440 147.175 ;
        RECT 100.610 146.750 100.885 147.175 ;
        RECT 101.055 146.920 101.440 147.345 ;
        RECT 100.610 146.555 101.440 146.750 ;
        RECT 100.015 146.205 100.920 146.385 ;
        RECT 99.510 145.705 99.920 146.035 ;
        RECT 100.090 145.705 100.920 146.205 ;
        RECT 101.090 146.035 101.440 146.555 ;
        RECT 101.610 146.385 101.855 147.175 ;
        RECT 102.045 146.750 102.300 147.175 ;
        RECT 102.470 146.920 102.855 147.345 ;
        RECT 102.045 146.555 102.855 146.750 ;
        RECT 101.610 146.205 102.335 146.385 ;
        RECT 101.090 145.705 101.515 146.035 ;
        RECT 101.685 145.705 102.335 146.205 ;
        RECT 102.505 146.035 102.855 146.555 ;
        RECT 103.025 146.205 103.285 147.175 ;
        RECT 102.505 145.705 102.930 146.035 ;
        RECT 96.555 144.795 98.225 145.565 ;
        RECT 99.510 145.535 99.845 145.705 ;
        RECT 100.090 145.535 100.440 145.705 ;
        RECT 101.090 145.535 101.440 145.705 ;
        RECT 101.685 145.535 101.855 145.705 ;
        RECT 102.505 145.535 102.855 145.705 ;
        RECT 103.100 145.535 103.285 146.205 ;
        RECT 98.855 145.365 99.845 145.535 ;
        RECT 98.855 144.965 99.290 145.365 ;
        RECT 99.460 144.795 99.845 145.195 ;
        RECT 100.015 144.965 100.440 145.535 ;
        RECT 100.630 145.365 101.440 145.535 ;
        RECT 100.630 144.965 100.885 145.365 ;
        RECT 101.055 144.795 101.440 145.195 ;
        RECT 101.610 144.965 101.855 145.535 ;
        RECT 102.045 145.365 102.855 145.535 ;
        RECT 102.045 144.965 102.300 145.365 ;
        RECT 102.470 144.795 102.855 145.195 ;
        RECT 103.025 144.965 103.285 145.535 ;
        RECT 103.455 145.075 103.735 147.175 ;
        RECT 103.925 146.585 104.710 147.345 ;
        RECT 105.105 146.515 105.490 147.175 ;
        RECT 105.105 146.415 105.515 146.515 ;
        RECT 103.905 146.205 105.515 146.415 ;
        RECT 105.815 146.325 106.015 147.115 ;
        RECT 103.905 145.605 104.180 146.205 ;
        RECT 105.685 146.155 106.015 146.325 ;
        RECT 106.185 146.165 106.505 147.345 ;
        RECT 106.675 146.255 109.265 147.345 ;
        RECT 105.685 146.035 105.865 146.155 ;
        RECT 104.350 145.785 104.705 146.035 ;
        RECT 104.900 145.985 105.365 146.035 ;
        RECT 104.895 145.815 105.365 145.985 ;
        RECT 104.900 145.785 105.365 145.815 ;
        RECT 105.535 145.785 105.865 146.035 ;
        RECT 106.040 145.785 106.505 145.985 ;
        RECT 103.905 145.425 105.155 145.605 ;
        RECT 104.790 145.355 105.155 145.425 ;
        RECT 105.325 145.405 106.505 145.575 ;
        RECT 103.965 144.795 104.135 145.255 ;
        RECT 105.325 145.185 105.655 145.405 ;
        RECT 104.405 145.005 105.655 145.185 ;
        RECT 105.825 144.795 105.995 145.235 ;
        RECT 106.165 144.990 106.505 145.405 ;
        RECT 106.675 145.565 107.885 146.085 ;
        RECT 108.055 145.735 109.265 146.255 ;
        RECT 109.435 146.180 109.725 147.345 ;
        RECT 106.675 144.795 109.265 145.565 ;
        RECT 109.435 144.795 109.725 145.520 ;
        RECT 109.895 145.075 110.175 147.175 ;
        RECT 110.365 146.585 111.150 147.345 ;
        RECT 111.545 146.515 111.930 147.175 ;
        RECT 111.545 146.415 111.955 146.515 ;
        RECT 110.345 146.205 111.955 146.415 ;
        RECT 112.255 146.325 112.455 147.115 ;
        RECT 110.345 145.605 110.620 146.205 ;
        RECT 112.125 146.155 112.455 146.325 ;
        RECT 112.625 146.165 112.945 147.345 ;
        RECT 113.195 146.415 113.375 147.175 ;
        RECT 113.555 146.585 113.885 147.345 ;
        RECT 113.195 146.245 113.870 146.415 ;
        RECT 114.055 146.270 114.325 147.175 ;
        RECT 112.125 146.035 112.305 146.155 ;
        RECT 113.700 146.100 113.870 146.245 ;
        RECT 110.790 145.785 111.145 146.035 ;
        RECT 111.340 145.985 111.805 146.035 ;
        RECT 111.335 145.815 111.805 145.985 ;
        RECT 111.340 145.785 111.805 145.815 ;
        RECT 111.975 145.785 112.305 146.035 ;
        RECT 112.480 145.785 112.945 145.985 ;
        RECT 113.135 145.695 113.475 146.065 ;
        RECT 113.700 145.770 113.975 146.100 ;
        RECT 110.345 145.425 111.595 145.605 ;
        RECT 111.230 145.355 111.595 145.425 ;
        RECT 111.765 145.405 112.945 145.575 ;
        RECT 113.700 145.515 113.870 145.770 ;
        RECT 110.405 144.795 110.575 145.255 ;
        RECT 111.765 145.185 112.095 145.405 ;
        RECT 110.845 145.005 112.095 145.185 ;
        RECT 112.265 144.795 112.435 145.235 ;
        RECT 112.605 144.990 112.945 145.405 ;
        RECT 113.205 145.345 113.870 145.515 ;
        RECT 114.145 145.470 114.325 146.270 ;
        RECT 114.495 146.165 114.815 147.345 ;
        RECT 114.985 146.325 115.185 147.115 ;
        RECT 115.510 146.515 115.895 147.175 ;
        RECT 116.290 146.585 117.075 147.345 ;
        RECT 115.485 146.415 115.895 146.515 ;
        RECT 114.985 146.155 115.315 146.325 ;
        RECT 115.485 146.205 117.095 146.415 ;
        RECT 115.135 146.035 115.315 146.155 ;
        RECT 114.495 145.785 114.960 145.985 ;
        RECT 115.135 145.785 115.465 146.035 ;
        RECT 115.635 145.985 116.100 146.035 ;
        RECT 115.635 145.815 116.105 145.985 ;
        RECT 115.635 145.785 116.100 145.815 ;
        RECT 116.295 145.785 116.650 146.035 ;
        RECT 116.820 145.605 117.095 146.205 ;
        RECT 113.205 144.965 113.375 145.345 ;
        RECT 113.555 144.795 113.885 145.175 ;
        RECT 114.065 144.965 114.325 145.470 ;
        RECT 114.495 145.405 115.675 145.575 ;
        RECT 114.495 144.990 114.835 145.405 ;
        RECT 115.005 144.795 115.175 145.235 ;
        RECT 115.345 145.185 115.675 145.405 ;
        RECT 115.845 145.425 117.095 145.605 ;
        RECT 115.845 145.355 116.210 145.425 ;
        RECT 115.345 145.005 116.595 145.185 ;
        RECT 116.865 144.795 117.035 145.255 ;
        RECT 117.265 145.075 117.545 147.175 ;
        RECT 118.635 146.585 119.300 147.175 ;
        RECT 118.635 145.615 118.885 146.585 ;
        RECT 119.470 146.505 119.800 147.345 ;
        RECT 120.310 146.755 121.115 147.175 ;
        RECT 119.970 146.585 121.535 146.755 ;
        RECT 119.970 146.335 120.140 146.585 ;
        RECT 119.220 146.165 120.140 146.335 ;
        RECT 119.220 145.995 119.390 146.165 ;
        RECT 120.310 145.995 120.685 146.415 ;
        RECT 119.055 145.785 119.390 145.995 ;
        RECT 119.560 145.785 120.010 145.995 ;
        RECT 120.200 145.985 120.685 145.995 ;
        RECT 120.875 146.035 121.195 146.415 ;
        RECT 121.365 146.335 121.535 146.585 ;
        RECT 121.705 146.505 121.955 147.345 ;
        RECT 122.150 146.335 122.450 147.175 ;
        RECT 121.365 146.165 122.450 146.335 ;
        RECT 120.200 145.815 120.705 145.985 ;
        RECT 120.200 145.785 120.685 145.815 ;
        RECT 120.875 145.785 121.255 146.035 ;
        RECT 121.435 145.785 121.765 145.995 ;
        RECT 118.635 144.975 119.320 145.615 ;
        RECT 119.490 144.795 119.660 145.615 ;
        RECT 119.830 145.445 121.530 145.615 ;
        RECT 119.830 144.980 120.160 145.445 ;
        RECT 121.145 145.355 121.530 145.445 ;
        RECT 121.935 145.535 122.105 146.165 ;
        RECT 122.275 145.705 122.605 145.995 ;
        RECT 122.775 145.740 123.055 147.175 ;
        RECT 123.225 146.570 123.935 147.345 ;
        RECT 124.105 146.400 124.435 147.175 ;
        RECT 123.285 146.185 124.435 146.400 ;
        RECT 121.935 145.355 122.445 145.535 ;
        RECT 120.330 144.795 120.500 145.265 ;
        RECT 120.760 145.015 121.945 145.185 ;
        RECT 122.115 144.965 122.445 145.355 ;
        RECT 122.775 144.965 123.115 145.740 ;
        RECT 123.285 145.615 123.570 146.185 ;
        RECT 123.755 145.785 124.225 146.015 ;
        RECT 124.630 145.985 124.845 147.100 ;
        RECT 125.025 146.625 125.355 147.345 ;
        RECT 125.135 145.985 125.365 146.325 ;
        RECT 125.535 146.255 127.205 147.345 ;
        RECT 124.395 145.805 124.845 145.985 ;
        RECT 124.395 145.785 124.725 145.805 ;
        RECT 125.035 145.785 125.365 145.985 ;
        RECT 123.285 145.425 123.995 145.615 ;
        RECT 123.695 145.285 123.995 145.425 ;
        RECT 124.185 145.425 125.365 145.615 ;
        RECT 124.185 145.345 124.515 145.425 ;
        RECT 123.695 145.275 124.010 145.285 ;
        RECT 123.695 145.265 124.020 145.275 ;
        RECT 123.695 145.260 124.030 145.265 ;
        RECT 123.285 144.795 123.455 145.255 ;
        RECT 123.695 145.250 124.035 145.260 ;
        RECT 123.695 145.245 124.040 145.250 ;
        RECT 123.695 145.235 124.045 145.245 ;
        RECT 123.695 145.230 124.050 145.235 ;
        RECT 123.695 144.965 124.055 145.230 ;
        RECT 124.685 144.795 124.855 145.255 ;
        RECT 125.025 144.965 125.365 145.425 ;
        RECT 125.535 145.565 126.285 146.085 ;
        RECT 126.455 145.735 127.205 146.255 ;
        RECT 127.530 146.335 127.830 147.175 ;
        RECT 128.025 146.505 128.275 147.345 ;
        RECT 128.865 146.755 129.670 147.175 ;
        RECT 128.445 146.585 130.010 146.755 ;
        RECT 128.445 146.335 128.615 146.585 ;
        RECT 127.530 146.165 128.615 146.335 ;
        RECT 127.375 145.705 127.705 145.995 ;
        RECT 125.535 144.795 127.205 145.565 ;
        RECT 127.875 145.535 128.045 146.165 ;
        RECT 128.785 146.035 129.105 146.415 ;
        RECT 128.215 145.785 128.545 145.995 ;
        RECT 128.725 145.785 129.105 146.035 ;
        RECT 129.295 145.995 129.670 146.415 ;
        RECT 129.840 146.335 130.010 146.585 ;
        RECT 130.180 146.505 130.510 147.345 ;
        RECT 130.680 146.585 131.345 147.175 ;
        RECT 129.840 146.165 130.760 146.335 ;
        RECT 130.590 145.995 130.760 146.165 ;
        RECT 129.295 145.985 129.780 145.995 ;
        RECT 129.275 145.815 129.780 145.985 ;
        RECT 129.295 145.785 129.780 145.815 ;
        RECT 129.970 145.785 130.420 145.995 ;
        RECT 130.590 145.785 130.925 145.995 ;
        RECT 131.095 145.615 131.345 146.585 ;
        RECT 127.535 145.355 128.045 145.535 ;
        RECT 128.450 145.445 130.150 145.615 ;
        RECT 128.450 145.355 128.835 145.445 ;
        RECT 127.535 144.965 127.865 145.355 ;
        RECT 128.035 145.015 129.220 145.185 ;
        RECT 129.480 144.795 129.650 145.265 ;
        RECT 129.820 144.980 130.150 145.445 ;
        RECT 130.320 144.795 130.490 145.615 ;
        RECT 130.660 144.975 131.345 145.615 ;
        RECT 131.515 146.270 131.785 147.175 ;
        RECT 131.955 146.585 132.285 147.345 ;
        RECT 132.465 146.415 132.645 147.175 ;
        RECT 131.515 145.470 131.695 146.270 ;
        RECT 131.970 146.245 132.645 146.415 ;
        RECT 132.895 146.255 134.565 147.345 ;
        RECT 131.970 146.100 132.140 146.245 ;
        RECT 131.865 145.770 132.140 146.100 ;
        RECT 131.970 145.515 132.140 145.770 ;
        RECT 132.365 145.695 132.705 146.065 ;
        RECT 132.895 145.565 133.645 146.085 ;
        RECT 133.815 145.735 134.565 146.255 ;
        RECT 135.195 146.180 135.485 147.345 ;
        RECT 135.655 146.165 135.975 147.345 ;
        RECT 136.145 146.325 136.345 147.115 ;
        RECT 136.670 146.515 137.055 147.175 ;
        RECT 137.450 146.585 138.235 147.345 ;
        RECT 136.645 146.415 137.055 146.515 ;
        RECT 136.145 146.155 136.475 146.325 ;
        RECT 136.645 146.205 138.255 146.415 ;
        RECT 136.295 146.035 136.475 146.155 ;
        RECT 135.655 145.785 136.120 145.985 ;
        RECT 136.295 145.785 136.625 146.035 ;
        RECT 136.795 145.985 137.260 146.035 ;
        RECT 136.795 145.815 137.265 145.985 ;
        RECT 136.795 145.785 137.260 145.815 ;
        RECT 137.455 145.785 137.810 146.035 ;
        RECT 137.980 145.605 138.255 146.205 ;
        RECT 131.515 144.965 131.775 145.470 ;
        RECT 131.970 145.345 132.635 145.515 ;
        RECT 131.955 144.795 132.285 145.175 ;
        RECT 132.465 144.965 132.635 145.345 ;
        RECT 132.895 144.795 134.565 145.565 ;
        RECT 135.195 144.795 135.485 145.520 ;
        RECT 135.655 145.405 136.835 145.575 ;
        RECT 135.655 144.990 135.995 145.405 ;
        RECT 136.165 144.795 136.335 145.235 ;
        RECT 136.505 145.185 136.835 145.405 ;
        RECT 137.005 145.425 138.255 145.605 ;
        RECT 137.005 145.355 137.370 145.425 ;
        RECT 136.505 145.005 137.755 145.185 ;
        RECT 138.025 144.795 138.195 145.255 ;
        RECT 138.425 145.075 138.705 147.175 ;
        RECT 138.875 146.910 144.220 147.345 ;
        RECT 144.395 146.910 149.740 147.345 ;
        RECT 140.460 145.340 140.800 146.170 ;
        RECT 142.280 145.660 142.630 146.910 ;
        RECT 145.980 145.340 146.320 146.170 ;
        RECT 147.800 145.660 148.150 146.910 ;
        RECT 149.915 146.255 153.425 147.345 ;
        RECT 153.595 146.255 154.805 147.345 ;
        RECT 149.915 145.565 151.565 146.085 ;
        RECT 151.735 145.735 153.425 146.255 ;
        RECT 138.875 144.795 144.220 145.340 ;
        RECT 144.395 144.795 149.740 145.340 ;
        RECT 149.915 144.795 153.425 145.565 ;
        RECT 153.595 145.545 154.115 146.085 ;
        RECT 154.285 145.715 154.805 146.255 ;
        RECT 154.975 146.255 156.185 147.345 ;
        RECT 154.975 145.715 155.495 146.255 ;
        RECT 155.665 145.545 156.185 146.085 ;
        RECT 153.595 144.795 154.805 145.545 ;
        RECT 154.975 144.795 156.185 145.545 ;
        RECT 70.710 144.625 156.270 144.795 ;
        RECT 70.795 143.875 72.005 144.625 ;
        RECT 70.795 143.335 71.315 143.875 ;
        RECT 72.175 143.855 73.845 144.625 ;
        RECT 74.015 143.950 74.275 144.455 ;
        RECT 74.455 144.245 74.785 144.625 ;
        RECT 74.965 144.075 75.135 144.455 ;
        RECT 75.860 144.225 76.195 144.625 ;
        RECT 71.485 143.165 72.005 143.705 ;
        RECT 72.175 143.335 72.925 143.855 ;
        RECT 73.095 143.165 73.845 143.685 ;
        RECT 70.795 142.075 72.005 143.165 ;
        RECT 72.175 142.075 73.845 143.165 ;
        RECT 74.015 143.150 74.185 143.950 ;
        RECT 74.470 143.905 75.135 144.075 ;
        RECT 76.365 144.055 76.570 144.455 ;
        RECT 76.780 144.145 77.055 144.625 ;
        RECT 77.265 144.125 77.525 144.455 ;
        RECT 74.470 143.650 74.640 143.905 ;
        RECT 75.885 143.885 76.570 144.055 ;
        RECT 74.355 143.320 74.640 143.650 ;
        RECT 74.875 143.355 75.205 143.725 ;
        RECT 74.470 143.175 74.640 143.320 ;
        RECT 74.015 142.245 74.285 143.150 ;
        RECT 74.470 143.005 75.135 143.175 ;
        RECT 74.455 142.075 74.785 142.835 ;
        RECT 74.965 142.245 75.135 143.005 ;
        RECT 75.885 142.855 76.225 143.885 ;
        RECT 76.395 143.215 76.645 143.715 ;
        RECT 76.825 143.385 77.185 143.965 ;
        RECT 77.355 143.215 77.525 144.125 ;
        RECT 77.695 144.080 83.040 144.625 ;
        RECT 83.305 144.285 83.475 144.320 ;
        RECT 83.275 144.115 83.475 144.285 ;
        RECT 79.280 143.250 79.620 144.080 ;
        RECT 76.395 143.045 77.525 143.215 ;
        RECT 75.885 142.680 76.550 142.855 ;
        RECT 75.860 142.075 76.195 142.500 ;
        RECT 76.365 142.275 76.550 142.680 ;
        RECT 76.755 142.075 77.085 142.855 ;
        RECT 77.255 142.275 77.525 143.045 ;
        RECT 81.100 142.510 81.450 143.760 ;
        RECT 83.305 143.755 83.475 144.115 ;
        RECT 83.665 144.095 83.895 144.400 ;
        RECT 84.065 144.265 84.395 144.625 ;
        RECT 84.590 144.095 84.880 144.445 ;
        RECT 83.665 143.925 84.880 144.095 ;
        RECT 85.145 144.075 85.315 144.455 ;
        RECT 85.495 144.245 85.825 144.625 ;
        RECT 85.145 143.905 85.810 144.075 ;
        RECT 86.005 143.950 86.265 144.455 ;
        RECT 86.435 144.080 91.780 144.625 ;
        RECT 83.305 143.585 83.825 143.755 ;
        RECT 83.220 143.055 83.465 143.415 ;
        RECT 83.655 143.205 83.825 143.585 ;
        RECT 83.995 143.385 84.380 143.715 ;
        RECT 84.560 143.605 84.820 143.715 ;
        RECT 84.560 143.435 84.825 143.605 ;
        RECT 84.560 143.385 84.820 143.435 ;
        RECT 83.655 142.925 84.005 143.205 ;
        RECT 77.695 142.075 83.040 142.510 ;
        RECT 83.220 142.075 83.475 142.875 ;
        RECT 83.675 142.245 84.005 142.925 ;
        RECT 84.185 142.335 84.380 143.385 ;
        RECT 85.075 143.355 85.405 143.725 ;
        RECT 85.640 143.650 85.810 143.905 ;
        RECT 85.640 143.320 85.925 143.650 ;
        RECT 84.560 142.075 84.880 143.215 ;
        RECT 85.640 143.175 85.810 143.320 ;
        RECT 85.145 143.005 85.810 143.175 ;
        RECT 86.095 143.150 86.265 143.950 ;
        RECT 88.020 143.250 88.360 144.080 ;
        RECT 92.575 144.065 92.905 144.455 ;
        RECT 93.075 144.235 94.260 144.405 ;
        RECT 94.520 144.155 94.690 144.625 ;
        RECT 92.575 143.885 93.085 144.065 ;
        RECT 85.145 142.245 85.315 143.005 ;
        RECT 85.495 142.075 85.825 142.835 ;
        RECT 85.995 142.245 86.265 143.150 ;
        RECT 89.840 142.510 90.190 143.760 ;
        RECT 92.415 143.425 92.745 143.715 ;
        RECT 92.915 143.255 93.085 143.885 ;
        RECT 93.490 143.975 93.875 144.065 ;
        RECT 94.860 143.975 95.190 144.440 ;
        RECT 93.490 143.805 95.190 143.975 ;
        RECT 95.360 143.805 95.530 144.625 ;
        RECT 95.700 143.805 96.385 144.445 ;
        RECT 96.555 143.900 96.845 144.625 ;
        RECT 97.175 144.065 97.505 144.455 ;
        RECT 97.675 144.235 98.860 144.405 ;
        RECT 99.120 144.155 99.290 144.625 ;
        RECT 97.175 143.885 97.685 144.065 ;
        RECT 93.255 143.425 93.585 143.635 ;
        RECT 93.765 143.385 94.145 143.635 ;
        RECT 94.335 143.605 94.820 143.635 ;
        RECT 94.315 143.435 94.820 143.605 ;
        RECT 92.570 143.085 93.655 143.255 ;
        RECT 86.435 142.075 91.780 142.510 ;
        RECT 92.570 142.245 92.870 143.085 ;
        RECT 93.065 142.075 93.315 142.915 ;
        RECT 93.485 142.835 93.655 143.085 ;
        RECT 93.825 143.005 94.145 143.385 ;
        RECT 94.335 143.425 94.820 143.435 ;
        RECT 95.010 143.425 95.460 143.635 ;
        RECT 95.630 143.425 95.965 143.635 ;
        RECT 94.335 143.005 94.710 143.425 ;
        RECT 95.630 143.255 95.800 143.425 ;
        RECT 94.880 143.085 95.800 143.255 ;
        RECT 94.880 142.835 95.050 143.085 ;
        RECT 93.485 142.665 95.050 142.835 ;
        RECT 93.905 142.245 94.710 142.665 ;
        RECT 95.220 142.075 95.550 142.915 ;
        RECT 96.135 142.835 96.385 143.805 ;
        RECT 97.015 143.425 97.345 143.715 ;
        RECT 97.515 143.255 97.685 143.885 ;
        RECT 98.090 143.975 98.475 144.065 ;
        RECT 99.460 143.975 99.790 144.440 ;
        RECT 98.090 143.805 99.790 143.975 ;
        RECT 99.960 143.805 100.130 144.625 ;
        RECT 100.300 143.805 100.985 144.445 ;
        RECT 97.855 143.425 98.185 143.635 ;
        RECT 98.365 143.385 98.745 143.635 ;
        RECT 98.935 143.605 99.420 143.635 ;
        RECT 98.915 143.435 99.420 143.605 ;
        RECT 95.720 142.245 96.385 142.835 ;
        RECT 96.555 142.075 96.845 143.240 ;
        RECT 97.170 143.085 98.255 143.255 ;
        RECT 97.170 142.245 97.470 143.085 ;
        RECT 97.665 142.075 97.915 142.915 ;
        RECT 98.085 142.835 98.255 143.085 ;
        RECT 98.425 143.005 98.745 143.385 ;
        RECT 98.935 143.425 99.420 143.435 ;
        RECT 99.610 143.425 100.060 143.635 ;
        RECT 100.230 143.425 100.565 143.635 ;
        RECT 98.935 143.005 99.310 143.425 ;
        RECT 100.230 143.255 100.400 143.425 ;
        RECT 99.480 143.085 100.400 143.255 ;
        RECT 99.480 142.835 99.650 143.085 ;
        RECT 98.085 142.665 99.650 142.835 ;
        RECT 98.505 142.245 99.310 142.665 ;
        RECT 99.820 142.075 100.150 142.915 ;
        RECT 100.735 142.835 100.985 143.805 ;
        RECT 101.155 143.875 102.365 144.625 ;
        RECT 102.535 143.995 102.875 144.455 ;
        RECT 103.045 144.165 103.215 144.625 ;
        RECT 103.845 144.190 104.205 144.455 ;
        RECT 103.850 144.185 104.205 144.190 ;
        RECT 103.855 144.175 104.205 144.185 ;
        RECT 103.860 144.170 104.205 144.175 ;
        RECT 103.865 144.160 104.205 144.170 ;
        RECT 104.445 144.165 104.615 144.625 ;
        RECT 103.870 144.155 104.205 144.160 ;
        RECT 103.880 144.145 104.205 144.155 ;
        RECT 103.890 144.135 104.205 144.145 ;
        RECT 103.385 143.995 103.715 144.075 ;
        RECT 101.155 143.335 101.675 143.875 ;
        RECT 102.535 143.805 103.715 143.995 ;
        RECT 103.905 143.995 104.205 144.135 ;
        RECT 103.905 143.805 104.615 143.995 ;
        RECT 101.845 143.165 102.365 143.705 ;
        RECT 100.320 142.245 100.985 142.835 ;
        RECT 101.155 142.075 102.365 143.165 ;
        RECT 102.535 143.435 102.865 143.635 ;
        RECT 103.175 143.615 103.505 143.635 ;
        RECT 103.055 143.435 103.505 143.615 ;
        RECT 102.535 143.095 102.765 143.435 ;
        RECT 102.545 142.075 102.875 142.795 ;
        RECT 103.055 142.320 103.270 143.435 ;
        RECT 103.675 143.405 104.145 143.635 ;
        RECT 104.330 143.235 104.615 143.805 ;
        RECT 104.785 143.680 105.125 144.455 ;
        RECT 103.465 143.020 104.615 143.235 ;
        RECT 103.465 142.245 103.795 143.020 ;
        RECT 103.965 142.075 104.675 142.850 ;
        RECT 104.845 142.245 105.125 143.680 ;
        RECT 105.295 143.805 105.980 144.445 ;
        RECT 106.150 143.805 106.320 144.625 ;
        RECT 106.490 143.975 106.820 144.440 ;
        RECT 106.990 144.155 107.160 144.625 ;
        RECT 107.420 144.235 108.605 144.405 ;
        RECT 108.775 144.065 109.105 144.455 ;
        RECT 109.435 144.080 114.780 144.625 ;
        RECT 107.805 143.975 108.190 144.065 ;
        RECT 106.490 143.805 108.190 143.975 ;
        RECT 108.595 143.885 109.105 144.065 ;
        RECT 105.295 142.835 105.545 143.805 ;
        RECT 105.715 143.425 106.050 143.635 ;
        RECT 106.220 143.425 106.670 143.635 ;
        RECT 106.860 143.425 107.345 143.635 ;
        RECT 105.880 143.255 106.050 143.425 ;
        RECT 106.970 143.265 107.345 143.425 ;
        RECT 107.535 143.385 107.915 143.635 ;
        RECT 108.095 143.425 108.425 143.635 ;
        RECT 105.880 143.085 106.800 143.255 ;
        RECT 105.295 142.245 105.960 142.835 ;
        RECT 106.130 142.075 106.460 142.915 ;
        RECT 106.630 142.835 106.800 143.085 ;
        RECT 106.970 143.095 107.365 143.265 ;
        RECT 106.970 143.005 107.345 143.095 ;
        RECT 107.535 143.005 107.855 143.385 ;
        RECT 108.595 143.255 108.765 143.885 ;
        RECT 108.935 143.425 109.265 143.715 ;
        RECT 108.025 143.085 109.110 143.255 ;
        RECT 111.020 143.250 111.360 144.080 ;
        RECT 114.955 143.805 115.640 144.445 ;
        RECT 115.810 143.805 115.980 144.625 ;
        RECT 116.150 143.975 116.480 144.440 ;
        RECT 116.650 144.155 116.820 144.625 ;
        RECT 117.080 144.235 118.265 144.405 ;
        RECT 118.435 144.065 118.765 144.455 ;
        RECT 117.465 143.975 117.850 144.065 ;
        RECT 116.150 143.805 117.850 143.975 ;
        RECT 118.255 143.885 118.765 144.065 ;
        RECT 108.025 142.835 108.195 143.085 ;
        RECT 106.630 142.665 108.195 142.835 ;
        RECT 106.970 142.245 107.775 142.665 ;
        RECT 108.365 142.075 108.615 142.915 ;
        RECT 108.810 142.245 109.110 143.085 ;
        RECT 112.840 142.510 113.190 143.760 ;
        RECT 114.955 142.835 115.205 143.805 ;
        RECT 115.375 143.425 115.710 143.635 ;
        RECT 115.880 143.425 116.330 143.635 ;
        RECT 116.520 143.425 117.005 143.635 ;
        RECT 115.540 143.255 115.710 143.425 ;
        RECT 116.630 143.265 117.005 143.425 ;
        RECT 117.195 143.385 117.575 143.635 ;
        RECT 117.755 143.425 118.085 143.635 ;
        RECT 115.540 143.085 116.460 143.255 ;
        RECT 109.435 142.075 114.780 142.510 ;
        RECT 114.955 142.245 115.620 142.835 ;
        RECT 115.790 142.075 116.120 142.915 ;
        RECT 116.290 142.835 116.460 143.085 ;
        RECT 116.630 143.095 117.025 143.265 ;
        RECT 116.630 143.005 117.005 143.095 ;
        RECT 117.195 143.005 117.515 143.385 ;
        RECT 118.255 143.255 118.425 143.885 ;
        RECT 119.095 143.855 121.685 144.625 ;
        RECT 122.315 143.900 122.605 144.625 ;
        RECT 122.775 143.855 124.445 144.625 ;
        RECT 124.615 143.950 124.875 144.455 ;
        RECT 125.055 144.245 125.385 144.625 ;
        RECT 125.565 144.075 125.735 144.455 ;
        RECT 126.160 144.115 126.400 144.625 ;
        RECT 126.580 144.115 126.860 144.445 ;
        RECT 127.090 144.115 127.305 144.625 ;
        RECT 118.595 143.425 118.925 143.715 ;
        RECT 119.095 143.335 120.305 143.855 ;
        RECT 117.685 143.085 118.770 143.255 ;
        RECT 120.475 143.165 121.685 143.685 ;
        RECT 122.775 143.335 123.525 143.855 ;
        RECT 117.685 142.835 117.855 143.085 ;
        RECT 116.290 142.665 117.855 142.835 ;
        RECT 116.630 142.245 117.435 142.665 ;
        RECT 118.025 142.075 118.275 142.915 ;
        RECT 118.470 142.245 118.770 143.085 ;
        RECT 119.095 142.075 121.685 143.165 ;
        RECT 122.315 142.075 122.605 143.240 ;
        RECT 123.695 143.165 124.445 143.685 ;
        RECT 122.775 142.075 124.445 143.165 ;
        RECT 124.615 143.150 124.795 143.950 ;
        RECT 125.070 143.905 125.735 144.075 ;
        RECT 125.070 143.650 125.240 143.905 ;
        RECT 124.965 143.320 125.240 143.650 ;
        RECT 125.465 143.355 125.805 143.725 ;
        RECT 126.055 143.385 126.410 143.945 ;
        RECT 125.070 143.175 125.240 143.320 ;
        RECT 126.580 143.215 126.750 144.115 ;
        RECT 126.920 143.385 127.185 143.945 ;
        RECT 127.475 143.885 128.090 144.455 ;
        RECT 128.295 144.055 128.730 144.455 ;
        RECT 128.900 144.225 129.285 144.625 ;
        RECT 128.295 143.885 129.285 144.055 ;
        RECT 129.455 143.885 129.880 144.455 ;
        RECT 130.070 144.055 130.325 144.455 ;
        RECT 130.495 144.225 130.880 144.625 ;
        RECT 130.070 143.885 130.880 144.055 ;
        RECT 131.050 143.885 131.295 144.455 ;
        RECT 131.485 144.055 131.740 144.455 ;
        RECT 131.910 144.225 132.295 144.625 ;
        RECT 131.485 143.885 132.295 144.055 ;
        RECT 132.465 143.885 132.725 144.455 ;
        RECT 127.435 143.215 127.605 143.715 ;
        RECT 124.615 142.245 124.885 143.150 ;
        RECT 125.070 143.005 125.745 143.175 ;
        RECT 125.055 142.075 125.385 142.835 ;
        RECT 125.565 142.245 125.745 143.005 ;
        RECT 126.180 143.045 127.605 143.215 ;
        RECT 126.180 142.870 126.570 143.045 ;
        RECT 127.055 142.075 127.385 142.875 ;
        RECT 127.775 142.865 128.090 143.885 ;
        RECT 128.950 143.715 129.285 143.885 ;
        RECT 129.530 143.715 129.880 143.885 ;
        RECT 130.530 143.715 130.880 143.885 ;
        RECT 131.125 143.715 131.295 143.885 ;
        RECT 131.945 143.715 132.295 143.885 ;
        RECT 128.295 143.010 128.780 143.715 ;
        RECT 128.950 143.385 129.360 143.715 ;
        RECT 127.555 142.245 128.090 142.865 ;
        RECT 128.950 142.840 129.285 143.385 ;
        RECT 129.530 143.215 130.360 143.715 ;
        RECT 128.295 142.670 129.285 142.840 ;
        RECT 129.455 143.035 130.360 143.215 ;
        RECT 130.530 143.385 130.955 143.715 ;
        RECT 128.295 142.245 128.730 142.670 ;
        RECT 128.900 142.075 129.285 142.500 ;
        RECT 129.455 142.245 129.880 143.035 ;
        RECT 130.530 142.865 130.880 143.385 ;
        RECT 131.125 143.215 131.775 143.715 ;
        RECT 130.050 142.670 130.880 142.865 ;
        RECT 131.050 143.035 131.775 143.215 ;
        RECT 131.945 143.385 132.370 143.715 ;
        RECT 130.050 142.245 130.325 142.670 ;
        RECT 130.495 142.075 130.880 142.500 ;
        RECT 131.050 142.245 131.295 143.035 ;
        RECT 131.945 142.865 132.295 143.385 ;
        RECT 132.540 143.215 132.725 143.885 ;
        RECT 132.895 143.855 135.485 144.625 ;
        RECT 136.445 144.225 136.775 144.625 ;
        RECT 136.945 144.055 137.275 144.395 ;
        RECT 138.325 144.225 138.655 144.625 ;
        RECT 136.290 143.885 138.655 144.055 ;
        RECT 138.825 143.900 139.155 144.410 ;
        RECT 132.895 143.335 134.105 143.855 ;
        RECT 131.485 142.670 132.295 142.865 ;
        RECT 131.485 142.245 131.740 142.670 ;
        RECT 131.910 142.075 132.295 142.500 ;
        RECT 132.465 142.245 132.725 143.215 ;
        RECT 134.275 143.165 135.485 143.685 ;
        RECT 132.895 142.075 135.485 143.165 ;
        RECT 136.290 142.885 136.460 143.885 ;
        RECT 138.485 143.715 138.655 143.885 ;
        RECT 136.630 143.055 136.875 143.715 ;
        RECT 137.090 143.055 137.355 143.715 ;
        RECT 137.550 143.055 137.835 143.715 ;
        RECT 138.010 143.385 138.315 143.715 ;
        RECT 138.485 143.385 138.795 143.715 ;
        RECT 138.010 143.055 138.225 143.385 ;
        RECT 136.290 142.715 136.745 142.885 ;
        RECT 136.415 142.285 136.745 142.715 ;
        RECT 136.925 142.715 138.215 142.885 ;
        RECT 136.925 142.295 137.175 142.715 ;
        RECT 137.405 142.075 137.735 142.545 ;
        RECT 137.965 142.295 138.215 142.715 ;
        RECT 138.405 142.075 138.655 143.215 ;
        RECT 138.965 143.135 139.155 143.900 ;
        RECT 138.825 142.285 139.155 143.135 ;
        RECT 140.290 143.885 140.905 144.455 ;
        RECT 141.075 144.115 141.290 144.625 ;
        RECT 141.520 144.115 141.800 144.445 ;
        RECT 141.980 144.115 142.220 144.625 ;
        RECT 140.290 142.865 140.605 143.885 ;
        RECT 140.775 143.215 140.945 143.715 ;
        RECT 141.195 143.385 141.460 143.945 ;
        RECT 141.630 143.215 141.800 144.115 ;
        RECT 141.970 143.385 142.325 143.945 ;
        RECT 142.555 143.825 143.250 144.455 ;
        RECT 143.455 143.825 143.765 144.625 ;
        RECT 143.935 143.855 147.445 144.625 ;
        RECT 148.075 143.900 148.365 144.625 ;
        RECT 142.575 143.385 142.910 143.635 ;
        RECT 143.080 143.225 143.250 143.825 ;
        RECT 143.420 143.385 143.755 143.655 ;
        RECT 143.935 143.335 145.585 143.855 ;
        RECT 148.995 143.790 149.285 144.625 ;
        RECT 149.455 144.225 150.410 144.395 ;
        RECT 150.825 144.235 151.155 144.625 ;
        RECT 140.775 143.045 142.200 143.215 ;
        RECT 140.290 142.245 140.825 142.865 ;
        RECT 140.995 142.075 141.325 142.875 ;
        RECT 141.810 142.870 142.200 143.045 ;
        RECT 142.555 142.075 142.815 143.215 ;
        RECT 142.985 142.245 143.315 143.225 ;
        RECT 143.485 142.075 143.765 143.215 ;
        RECT 145.755 143.165 147.445 143.685 ;
        RECT 149.455 143.345 149.625 144.225 ;
        RECT 151.325 144.055 151.495 144.375 ;
        RECT 151.665 144.235 151.995 144.625 ;
        RECT 149.795 143.885 152.045 144.055 ;
        RECT 149.795 143.385 150.025 143.885 ;
        RECT 150.195 143.465 150.570 143.635 ;
        RECT 143.935 142.075 147.445 143.165 ;
        RECT 148.075 142.075 148.365 143.240 ;
        RECT 148.995 143.175 149.625 143.345 ;
        RECT 150.400 143.265 150.570 143.465 ;
        RECT 150.740 143.435 151.290 143.635 ;
        RECT 151.460 143.265 151.705 143.715 ;
        RECT 148.995 142.245 149.315 143.175 ;
        RECT 150.400 143.095 151.705 143.265 ;
        RECT 151.875 142.925 152.045 143.885 ;
        RECT 152.215 143.855 154.805 144.625 ;
        RECT 154.975 143.875 156.185 144.625 ;
        RECT 152.215 143.335 153.425 143.855 ;
        RECT 153.595 143.165 154.805 143.685 ;
        RECT 149.495 142.755 150.735 142.925 ;
        RECT 149.495 142.245 149.895 142.755 ;
        RECT 150.065 142.075 150.235 142.585 ;
        RECT 150.405 142.245 150.735 142.755 ;
        RECT 150.905 142.075 151.075 142.925 ;
        RECT 151.665 142.245 152.045 142.925 ;
        RECT 152.215 142.075 154.805 143.165 ;
        RECT 154.975 143.165 155.495 143.705 ;
        RECT 155.665 143.335 156.185 143.875 ;
        RECT 154.975 142.075 156.185 143.165 ;
        RECT 70.710 141.905 156.270 142.075 ;
        RECT 70.795 140.815 72.005 141.905 ;
        RECT 72.265 141.235 72.435 141.735 ;
        RECT 72.605 141.405 72.935 141.905 ;
        RECT 72.265 141.065 72.930 141.235 ;
        RECT 70.795 140.105 71.315 140.645 ;
        RECT 71.485 140.275 72.005 140.815 ;
        RECT 72.180 140.245 72.530 140.895 ;
        RECT 70.795 139.355 72.005 140.105 ;
        RECT 72.700 140.075 72.930 141.065 ;
        RECT 72.265 139.905 72.930 140.075 ;
        RECT 72.265 139.615 72.435 139.905 ;
        RECT 72.605 139.355 72.935 139.735 ;
        RECT 73.105 139.615 73.290 141.735 ;
        RECT 73.530 141.445 73.795 141.905 ;
        RECT 73.965 141.310 74.215 141.735 ;
        RECT 74.425 141.460 75.530 141.630 ;
        RECT 73.910 141.180 74.215 141.310 ;
        RECT 73.460 139.985 73.740 140.935 ;
        RECT 73.910 140.075 74.080 141.180 ;
        RECT 74.250 140.395 74.490 140.990 ;
        RECT 74.660 140.925 75.190 141.290 ;
        RECT 74.660 140.225 74.830 140.925 ;
        RECT 75.360 140.845 75.530 141.460 ;
        RECT 75.700 141.105 75.870 141.905 ;
        RECT 76.040 141.405 76.290 141.735 ;
        RECT 76.515 141.435 77.400 141.605 ;
        RECT 75.360 140.755 75.870 140.845 ;
        RECT 73.910 139.945 74.135 140.075 ;
        RECT 74.305 140.005 74.830 140.225 ;
        RECT 75.000 140.585 75.870 140.755 ;
        RECT 73.545 139.355 73.795 139.815 ;
        RECT 73.965 139.805 74.135 139.945 ;
        RECT 75.000 139.805 75.170 140.585 ;
        RECT 75.700 140.515 75.870 140.585 ;
        RECT 75.380 140.335 75.580 140.365 ;
        RECT 76.040 140.335 76.210 141.405 ;
        RECT 76.380 140.515 76.570 141.235 ;
        RECT 75.380 140.035 76.210 140.335 ;
        RECT 76.740 140.305 77.060 141.265 ;
        RECT 73.965 139.635 74.300 139.805 ;
        RECT 74.495 139.635 75.170 139.805 ;
        RECT 75.490 139.355 75.860 139.855 ;
        RECT 76.040 139.805 76.210 140.035 ;
        RECT 76.595 139.975 77.060 140.305 ;
        RECT 77.230 140.595 77.400 141.435 ;
        RECT 77.580 141.405 77.895 141.905 ;
        RECT 78.125 141.175 78.465 141.735 ;
        RECT 77.570 140.800 78.465 141.175 ;
        RECT 78.635 140.895 78.805 141.905 ;
        RECT 78.275 140.595 78.465 140.800 ;
        RECT 78.975 140.845 79.305 141.690 ;
        RECT 79.535 141.185 79.995 141.735 ;
        RECT 80.185 141.185 80.515 141.905 ;
        RECT 78.975 140.765 79.365 140.845 ;
        RECT 79.150 140.715 79.365 140.765 ;
        RECT 77.230 140.265 78.105 140.595 ;
        RECT 78.275 140.265 79.025 140.595 ;
        RECT 77.230 139.805 77.400 140.265 ;
        RECT 78.275 140.095 78.475 140.265 ;
        RECT 79.195 140.135 79.365 140.715 ;
        RECT 79.140 140.095 79.365 140.135 ;
        RECT 76.040 139.635 76.445 139.805 ;
        RECT 76.615 139.635 77.400 139.805 ;
        RECT 77.675 139.355 77.885 139.885 ;
        RECT 78.145 139.570 78.475 140.095 ;
        RECT 78.985 140.010 79.365 140.095 ;
        RECT 78.645 139.355 78.815 139.965 ;
        RECT 78.985 139.575 79.315 140.010 ;
        RECT 79.535 139.815 79.785 141.185 ;
        RECT 80.715 141.015 81.015 141.565 ;
        RECT 81.185 141.235 81.465 141.905 ;
        RECT 80.075 140.845 81.015 141.015 ;
        RECT 80.075 140.595 80.245 140.845 ;
        RECT 81.385 140.595 81.650 140.955 ;
        RECT 79.955 140.265 80.245 140.595 ;
        RECT 80.415 140.345 80.755 140.595 ;
        RECT 80.975 140.345 81.650 140.595 ;
        RECT 81.835 140.935 82.105 141.705 ;
        RECT 82.275 141.125 82.605 141.905 ;
        RECT 82.810 141.300 82.995 141.705 ;
        RECT 83.165 141.480 83.500 141.905 ;
        RECT 82.810 141.125 83.475 141.300 ;
        RECT 81.835 140.765 82.965 140.935 ;
        RECT 80.075 140.175 80.245 140.265 ;
        RECT 80.075 139.985 81.465 140.175 ;
        RECT 79.535 139.525 80.095 139.815 ;
        RECT 80.265 139.355 80.515 139.815 ;
        RECT 81.135 139.625 81.465 139.985 ;
        RECT 81.835 139.855 82.005 140.765 ;
        RECT 82.175 140.015 82.535 140.595 ;
        RECT 82.715 140.265 82.965 140.765 ;
        RECT 83.135 140.095 83.475 141.125 ;
        RECT 83.675 140.740 83.965 141.905 ;
        RECT 84.225 141.235 84.395 141.735 ;
        RECT 84.565 141.405 84.895 141.905 ;
        RECT 84.225 141.065 84.890 141.235 ;
        RECT 84.140 140.245 84.490 140.895 ;
        RECT 82.790 139.925 83.475 140.095 ;
        RECT 81.835 139.525 82.095 139.855 ;
        RECT 82.305 139.355 82.580 139.835 ;
        RECT 82.790 139.525 82.995 139.925 ;
        RECT 83.165 139.355 83.500 139.755 ;
        RECT 83.675 139.355 83.965 140.080 ;
        RECT 84.660 140.075 84.890 141.065 ;
        RECT 84.225 139.905 84.890 140.075 ;
        RECT 84.225 139.615 84.395 139.905 ;
        RECT 84.565 139.355 84.895 139.735 ;
        RECT 85.065 139.615 85.250 141.735 ;
        RECT 85.490 141.445 85.755 141.905 ;
        RECT 85.925 141.310 86.175 141.735 ;
        RECT 86.385 141.460 87.490 141.630 ;
        RECT 85.870 141.180 86.175 141.310 ;
        RECT 85.420 139.985 85.700 140.935 ;
        RECT 85.870 140.075 86.040 141.180 ;
        RECT 86.210 140.395 86.450 140.990 ;
        RECT 86.620 140.925 87.150 141.290 ;
        RECT 86.620 140.225 86.790 140.925 ;
        RECT 87.320 140.845 87.490 141.460 ;
        RECT 87.660 141.105 87.830 141.905 ;
        RECT 88.000 141.405 88.250 141.735 ;
        RECT 88.475 141.435 89.360 141.605 ;
        RECT 87.320 140.755 87.830 140.845 ;
        RECT 85.870 139.945 86.095 140.075 ;
        RECT 86.265 140.005 86.790 140.225 ;
        RECT 86.960 140.585 87.830 140.755 ;
        RECT 85.505 139.355 85.755 139.815 ;
        RECT 85.925 139.805 86.095 139.945 ;
        RECT 86.960 139.805 87.130 140.585 ;
        RECT 87.660 140.515 87.830 140.585 ;
        RECT 87.340 140.335 87.540 140.365 ;
        RECT 88.000 140.335 88.170 141.405 ;
        RECT 88.340 140.515 88.530 141.235 ;
        RECT 87.340 140.035 88.170 140.335 ;
        RECT 88.700 140.305 89.020 141.265 ;
        RECT 85.925 139.635 86.260 139.805 ;
        RECT 86.455 139.635 87.130 139.805 ;
        RECT 87.450 139.355 87.820 139.855 ;
        RECT 88.000 139.805 88.170 140.035 ;
        RECT 88.555 139.975 89.020 140.305 ;
        RECT 89.190 140.595 89.360 141.435 ;
        RECT 89.540 141.405 89.855 141.905 ;
        RECT 90.085 141.175 90.425 141.735 ;
        RECT 89.530 140.800 90.425 141.175 ;
        RECT 90.595 140.895 90.765 141.905 ;
        RECT 90.235 140.595 90.425 140.800 ;
        RECT 90.935 140.845 91.265 141.690 ;
        RECT 90.935 140.765 91.325 140.845 ;
        RECT 91.495 140.815 94.085 141.905 ;
        RECT 91.110 140.715 91.325 140.765 ;
        RECT 89.190 140.265 90.065 140.595 ;
        RECT 90.235 140.265 90.985 140.595 ;
        RECT 89.190 139.805 89.360 140.265 ;
        RECT 90.235 140.095 90.435 140.265 ;
        RECT 91.155 140.135 91.325 140.715 ;
        RECT 91.100 140.095 91.325 140.135 ;
        RECT 88.000 139.635 88.405 139.805 ;
        RECT 88.575 139.635 89.360 139.805 ;
        RECT 89.635 139.355 89.845 139.885 ;
        RECT 90.105 139.570 90.435 140.095 ;
        RECT 90.945 140.010 91.325 140.095 ;
        RECT 91.495 140.125 92.705 140.645 ;
        RECT 92.875 140.295 94.085 140.815 ;
        RECT 94.715 140.765 95.055 141.735 ;
        RECT 95.225 140.765 95.395 141.905 ;
        RECT 95.665 141.105 95.915 141.905 ;
        RECT 96.560 140.935 96.890 141.735 ;
        RECT 97.190 141.105 97.520 141.905 ;
        RECT 97.690 140.935 98.020 141.735 ;
        RECT 98.405 141.185 98.735 141.905 ;
        RECT 95.585 140.765 98.020 140.935 ;
        RECT 94.715 140.155 94.890 140.765 ;
        RECT 95.585 140.515 95.755 140.765 ;
        RECT 95.060 140.345 95.755 140.515 ;
        RECT 95.930 140.345 96.350 140.545 ;
        RECT 96.520 140.345 96.850 140.545 ;
        RECT 97.020 140.345 97.350 140.545 ;
        RECT 90.605 139.355 90.775 139.965 ;
        RECT 90.945 139.575 91.275 140.010 ;
        RECT 91.495 139.355 94.085 140.125 ;
        RECT 94.715 139.525 95.055 140.155 ;
        RECT 95.225 139.355 95.475 140.155 ;
        RECT 95.665 140.005 96.890 140.175 ;
        RECT 95.665 139.525 95.995 140.005 ;
        RECT 96.165 139.355 96.390 139.815 ;
        RECT 96.560 139.525 96.890 140.005 ;
        RECT 97.520 140.135 97.690 140.765 ;
        RECT 97.875 140.345 98.225 140.595 ;
        RECT 98.395 140.545 98.625 140.885 ;
        RECT 98.915 140.545 99.130 141.660 ;
        RECT 99.325 140.960 99.655 141.735 ;
        RECT 99.825 141.130 100.535 141.905 ;
        RECT 99.325 140.745 100.475 140.960 ;
        RECT 98.395 140.345 98.725 140.545 ;
        RECT 98.915 140.365 99.365 140.545 ;
        RECT 99.035 140.345 99.365 140.365 ;
        RECT 99.535 140.345 100.005 140.575 ;
        RECT 100.190 140.175 100.475 140.745 ;
        RECT 100.705 140.300 100.985 141.735 ;
        RECT 101.155 140.815 103.745 141.905 ;
        RECT 97.520 139.525 98.020 140.135 ;
        RECT 98.395 139.985 99.575 140.175 ;
        RECT 98.395 139.525 98.735 139.985 ;
        RECT 99.245 139.905 99.575 139.985 ;
        RECT 99.765 139.985 100.475 140.175 ;
        RECT 99.765 139.845 100.065 139.985 ;
        RECT 99.750 139.835 100.065 139.845 ;
        RECT 99.740 139.825 100.065 139.835 ;
        RECT 99.730 139.820 100.065 139.825 ;
        RECT 98.905 139.355 99.075 139.815 ;
        RECT 99.725 139.810 100.065 139.820 ;
        RECT 99.720 139.805 100.065 139.810 ;
        RECT 99.715 139.795 100.065 139.805 ;
        RECT 99.710 139.790 100.065 139.795 ;
        RECT 99.705 139.525 100.065 139.790 ;
        RECT 100.305 139.355 100.475 139.815 ;
        RECT 100.645 139.525 100.985 140.300 ;
        RECT 101.155 140.125 102.365 140.645 ;
        RECT 102.535 140.295 103.745 140.815 ;
        RECT 103.915 140.300 104.195 141.735 ;
        RECT 104.365 141.130 105.075 141.905 ;
        RECT 105.245 140.960 105.575 141.735 ;
        RECT 104.425 140.745 105.575 140.960 ;
        RECT 101.155 139.355 103.745 140.125 ;
        RECT 103.915 139.525 104.255 140.300 ;
        RECT 104.425 140.175 104.710 140.745 ;
        RECT 104.895 140.345 105.365 140.575 ;
        RECT 105.770 140.545 105.985 141.660 ;
        RECT 106.165 141.185 106.495 141.905 ;
        RECT 106.275 140.545 106.505 140.885 ;
        RECT 106.675 140.815 109.265 141.905 ;
        RECT 105.535 140.365 105.985 140.545 ;
        RECT 105.535 140.345 105.865 140.365 ;
        RECT 106.175 140.345 106.505 140.545 ;
        RECT 104.425 139.985 105.135 140.175 ;
        RECT 104.835 139.845 105.135 139.985 ;
        RECT 105.325 139.985 106.505 140.175 ;
        RECT 105.325 139.905 105.655 139.985 ;
        RECT 104.835 139.835 105.150 139.845 ;
        RECT 104.835 139.825 105.160 139.835 ;
        RECT 104.835 139.820 105.170 139.825 ;
        RECT 104.425 139.355 104.595 139.815 ;
        RECT 104.835 139.810 105.175 139.820 ;
        RECT 104.835 139.805 105.180 139.810 ;
        RECT 104.835 139.795 105.185 139.805 ;
        RECT 104.835 139.790 105.190 139.795 ;
        RECT 104.835 139.525 105.195 139.790 ;
        RECT 105.825 139.355 105.995 139.815 ;
        RECT 106.165 139.525 106.505 139.985 ;
        RECT 106.675 140.125 107.885 140.645 ;
        RECT 108.055 140.295 109.265 140.815 ;
        RECT 109.435 140.740 109.725 141.905 ;
        RECT 109.895 141.470 115.240 141.905 ;
        RECT 106.675 139.355 109.265 140.125 ;
        RECT 109.435 139.355 109.725 140.080 ;
        RECT 111.480 139.900 111.820 140.730 ;
        RECT 113.300 140.220 113.650 141.470 ;
        RECT 115.875 140.765 116.155 141.905 ;
        RECT 116.325 140.755 116.655 141.735 ;
        RECT 116.825 140.765 117.085 141.905 ;
        RECT 117.255 140.815 119.845 141.905 ;
        RECT 115.885 140.325 116.220 140.595 ;
        RECT 116.390 140.155 116.560 140.755 ;
        RECT 116.730 140.345 117.065 140.595 ;
        RECT 109.895 139.355 115.240 139.900 ;
        RECT 115.875 139.355 116.185 140.155 ;
        RECT 116.390 139.525 117.085 140.155 ;
        RECT 117.255 140.125 118.465 140.645 ;
        RECT 118.635 140.295 119.845 140.815 ;
        RECT 120.475 140.765 120.735 141.735 ;
        RECT 120.905 141.480 121.290 141.905 ;
        RECT 121.460 141.310 121.715 141.735 ;
        RECT 120.905 141.115 121.715 141.310 ;
        RECT 117.255 139.355 119.845 140.125 ;
        RECT 120.475 140.095 120.660 140.765 ;
        RECT 120.905 140.595 121.255 141.115 ;
        RECT 121.905 140.945 122.150 141.735 ;
        RECT 122.320 141.480 122.705 141.905 ;
        RECT 122.875 141.310 123.150 141.735 ;
        RECT 120.830 140.265 121.255 140.595 ;
        RECT 121.425 140.765 122.150 140.945 ;
        RECT 122.320 141.115 123.150 141.310 ;
        RECT 121.425 140.265 122.075 140.765 ;
        RECT 122.320 140.595 122.670 141.115 ;
        RECT 123.320 140.945 123.745 141.735 ;
        RECT 123.915 141.480 124.300 141.905 ;
        RECT 124.470 141.310 124.905 141.735 ;
        RECT 122.245 140.265 122.670 140.595 ;
        RECT 122.840 140.765 123.745 140.945 ;
        RECT 123.915 141.140 124.905 141.310 ;
        RECT 122.840 140.265 123.670 140.765 ;
        RECT 123.915 140.595 124.250 141.140 ;
        RECT 123.840 140.265 124.250 140.595 ;
        RECT 124.420 140.265 124.905 140.970 ;
        RECT 125.075 140.830 125.345 141.735 ;
        RECT 125.515 141.145 125.845 141.905 ;
        RECT 126.025 140.975 126.205 141.735 ;
        RECT 120.905 140.095 121.255 140.265 ;
        RECT 121.905 140.095 122.075 140.265 ;
        RECT 122.320 140.095 122.670 140.265 ;
        RECT 123.320 140.095 123.670 140.265 ;
        RECT 123.915 140.095 124.250 140.265 ;
        RECT 120.475 139.525 120.735 140.095 ;
        RECT 120.905 139.925 121.715 140.095 ;
        RECT 120.905 139.355 121.290 139.755 ;
        RECT 121.460 139.525 121.715 139.925 ;
        RECT 121.905 139.525 122.150 140.095 ;
        RECT 122.320 139.925 123.130 140.095 ;
        RECT 122.320 139.355 122.705 139.755 ;
        RECT 122.875 139.525 123.130 139.925 ;
        RECT 123.320 139.525 123.745 140.095 ;
        RECT 123.915 139.925 124.905 140.095 ;
        RECT 123.915 139.355 124.300 139.755 ;
        RECT 124.470 139.525 124.905 139.925 ;
        RECT 125.075 140.030 125.255 140.830 ;
        RECT 125.530 140.805 126.205 140.975 ;
        RECT 125.530 140.660 125.700 140.805 ;
        RECT 125.425 140.330 125.700 140.660 ;
        RECT 126.915 140.765 127.175 141.735 ;
        RECT 127.345 141.480 127.730 141.905 ;
        RECT 127.900 141.310 128.155 141.735 ;
        RECT 127.345 141.115 128.155 141.310 ;
        RECT 125.530 140.075 125.700 140.330 ;
        RECT 125.925 140.255 126.265 140.625 ;
        RECT 126.915 140.095 127.100 140.765 ;
        RECT 127.345 140.595 127.695 141.115 ;
        RECT 128.345 140.945 128.590 141.735 ;
        RECT 128.760 141.480 129.145 141.905 ;
        RECT 129.315 141.310 129.590 141.735 ;
        RECT 127.270 140.265 127.695 140.595 ;
        RECT 127.865 140.765 128.590 140.945 ;
        RECT 128.760 141.115 129.590 141.310 ;
        RECT 127.865 140.265 128.515 140.765 ;
        RECT 128.760 140.595 129.110 141.115 ;
        RECT 129.760 140.945 130.185 141.735 ;
        RECT 130.355 141.480 130.740 141.905 ;
        RECT 130.910 141.310 131.345 141.735 ;
        RECT 128.685 140.265 129.110 140.595 ;
        RECT 129.280 140.765 130.185 140.945 ;
        RECT 130.355 141.140 131.345 141.310 ;
        RECT 132.275 141.265 132.605 141.695 ;
        RECT 129.280 140.265 130.110 140.765 ;
        RECT 130.355 140.595 130.690 141.140 ;
        RECT 132.150 141.095 132.605 141.265 ;
        RECT 132.785 141.265 133.035 141.685 ;
        RECT 133.265 141.435 133.595 141.905 ;
        RECT 133.825 141.265 134.075 141.685 ;
        RECT 132.785 141.095 134.075 141.265 ;
        RECT 130.280 140.265 130.690 140.595 ;
        RECT 130.860 140.265 131.345 140.970 ;
        RECT 127.345 140.095 127.695 140.265 ;
        RECT 128.345 140.095 128.515 140.265 ;
        RECT 128.760 140.095 129.110 140.265 ;
        RECT 129.760 140.095 130.110 140.265 ;
        RECT 130.355 140.095 130.690 140.265 ;
        RECT 132.150 140.095 132.320 141.095 ;
        RECT 132.490 140.265 132.735 140.925 ;
        RECT 132.950 140.265 133.215 140.925 ;
        RECT 133.410 140.265 133.695 140.925 ;
        RECT 133.870 140.595 134.085 140.925 ;
        RECT 134.265 140.765 134.515 141.905 ;
        RECT 134.685 140.845 135.015 141.695 ;
        RECT 133.870 140.265 134.175 140.595 ;
        RECT 134.345 140.265 134.655 140.595 ;
        RECT 134.345 140.095 134.515 140.265 ;
        RECT 125.075 139.525 125.335 140.030 ;
        RECT 125.530 139.905 126.195 140.075 ;
        RECT 125.515 139.355 125.845 139.735 ;
        RECT 126.025 139.525 126.195 139.905 ;
        RECT 126.915 139.525 127.175 140.095 ;
        RECT 127.345 139.925 128.155 140.095 ;
        RECT 127.345 139.355 127.730 139.755 ;
        RECT 127.900 139.525 128.155 139.925 ;
        RECT 128.345 139.525 128.590 140.095 ;
        RECT 128.760 139.925 129.570 140.095 ;
        RECT 128.760 139.355 129.145 139.755 ;
        RECT 129.315 139.525 129.570 139.925 ;
        RECT 129.760 139.525 130.185 140.095 ;
        RECT 130.355 139.925 131.345 140.095 ;
        RECT 132.150 139.925 134.515 140.095 ;
        RECT 134.825 140.080 135.015 140.845 ;
        RECT 135.195 140.740 135.485 141.905 ;
        RECT 135.655 140.765 135.995 141.735 ;
        RECT 136.165 140.765 136.335 141.905 ;
        RECT 136.605 141.105 136.855 141.905 ;
        RECT 137.500 140.935 137.830 141.735 ;
        RECT 138.130 141.105 138.460 141.905 ;
        RECT 138.630 140.935 138.960 141.735 ;
        RECT 136.525 140.765 138.960 140.935 ;
        RECT 139.345 140.845 139.675 141.695 ;
        RECT 135.655 140.155 135.830 140.765 ;
        RECT 136.525 140.515 136.695 140.765 ;
        RECT 136.000 140.345 136.695 140.515 ;
        RECT 136.870 140.345 137.290 140.545 ;
        RECT 137.460 140.345 137.790 140.545 ;
        RECT 137.960 140.345 138.290 140.545 ;
        RECT 130.355 139.355 130.740 139.755 ;
        RECT 130.910 139.525 131.345 139.925 ;
        RECT 132.305 139.355 132.635 139.755 ;
        RECT 132.805 139.585 133.135 139.925 ;
        RECT 134.185 139.355 134.515 139.755 ;
        RECT 134.685 139.570 135.015 140.080 ;
        RECT 135.195 139.355 135.485 140.080 ;
        RECT 135.655 139.525 135.995 140.155 ;
        RECT 136.165 139.355 136.415 140.155 ;
        RECT 136.605 140.005 137.830 140.175 ;
        RECT 136.605 139.525 136.935 140.005 ;
        RECT 137.105 139.355 137.330 139.815 ;
        RECT 137.500 139.525 137.830 140.005 ;
        RECT 138.460 140.135 138.630 140.765 ;
        RECT 138.815 140.345 139.165 140.595 ;
        RECT 138.460 139.525 138.960 140.135 ;
        RECT 139.345 140.080 139.535 140.845 ;
        RECT 139.845 140.765 140.095 141.905 ;
        RECT 140.285 141.265 140.535 141.685 ;
        RECT 140.765 141.435 141.095 141.905 ;
        RECT 141.325 141.265 141.575 141.685 ;
        RECT 140.285 141.095 141.575 141.265 ;
        RECT 141.755 141.265 142.085 141.695 ;
        RECT 141.755 141.095 142.210 141.265 ;
        RECT 140.275 140.595 140.490 140.925 ;
        RECT 139.705 140.265 140.015 140.595 ;
        RECT 140.185 140.265 140.490 140.595 ;
        RECT 140.665 140.265 140.950 140.925 ;
        RECT 141.145 140.265 141.410 140.925 ;
        RECT 141.625 140.265 141.870 140.925 ;
        RECT 139.845 140.095 140.015 140.265 ;
        RECT 142.040 140.095 142.210 141.095 ;
        RECT 139.345 139.570 139.675 140.080 ;
        RECT 139.845 139.925 142.210 140.095 ;
        RECT 143.475 140.795 143.735 141.735 ;
        RECT 143.905 141.505 144.235 141.905 ;
        RECT 145.380 141.640 145.635 141.735 ;
        RECT 144.495 141.470 145.635 141.640 ;
        RECT 145.805 141.525 146.135 141.695 ;
        RECT 144.495 141.245 144.665 141.470 ;
        RECT 143.905 141.075 144.665 141.245 ;
        RECT 145.380 141.335 145.635 141.470 ;
        RECT 143.475 140.080 143.650 140.795 ;
        RECT 143.905 140.595 144.075 141.075 ;
        RECT 144.930 140.985 145.100 141.175 ;
        RECT 145.380 141.165 145.790 141.335 ;
        RECT 143.820 140.265 144.075 140.595 ;
        RECT 144.300 140.265 144.630 140.885 ;
        RECT 144.930 140.815 145.450 140.985 ;
        RECT 144.800 140.265 145.090 140.645 ;
        RECT 145.280 140.095 145.450 140.815 ;
        RECT 139.845 139.355 140.175 139.755 ;
        RECT 141.225 139.585 141.555 139.925 ;
        RECT 141.725 139.355 142.055 139.755 ;
        RECT 143.475 139.525 143.735 140.080 ;
        RECT 144.570 139.925 145.450 140.095 ;
        RECT 145.620 140.140 145.790 141.165 ;
        RECT 145.965 141.275 146.135 141.525 ;
        RECT 146.305 141.445 146.555 141.905 ;
        RECT 146.725 141.275 146.905 141.735 ;
        RECT 145.965 141.105 146.905 141.275 ;
        RECT 147.155 141.105 147.595 141.735 ;
        RECT 145.990 140.625 146.470 140.925 ;
        RECT 145.620 139.970 145.970 140.140 ;
        RECT 146.210 140.035 146.470 140.625 ;
        RECT 146.670 140.035 146.930 140.925 ;
        RECT 147.155 140.095 147.465 141.105 ;
        RECT 147.770 141.055 148.085 141.905 ;
        RECT 148.255 141.565 149.685 141.735 ;
        RECT 148.255 140.885 148.425 141.565 ;
        RECT 147.635 140.715 148.425 140.885 ;
        RECT 147.635 140.265 147.805 140.715 ;
        RECT 148.595 140.595 148.795 141.395 ;
        RECT 147.975 140.265 148.365 140.545 ;
        RECT 148.550 140.265 148.795 140.595 ;
        RECT 148.995 140.265 149.245 141.395 ;
        RECT 149.435 140.935 149.685 141.565 ;
        RECT 149.865 141.105 150.195 141.905 ;
        RECT 149.435 140.765 150.205 140.935 ;
        RECT 150.375 140.815 151.585 141.905 ;
        RECT 151.775 141.055 152.105 141.905 ;
        RECT 152.275 141.565 153.385 141.735 ;
        RECT 152.275 141.055 152.495 141.565 ;
        RECT 153.195 141.405 153.385 141.565 ;
        RECT 153.580 141.445 153.910 141.905 ;
        RECT 152.665 141.235 152.965 141.395 ;
        RECT 154.080 141.235 154.315 141.735 ;
        RECT 152.665 141.055 154.315 141.235 ;
        RECT 149.460 140.265 149.865 140.595 ;
        RECT 150.035 140.095 150.205 140.765 ;
        RECT 143.905 139.355 144.335 139.800 ;
        RECT 144.570 139.525 144.740 139.925 ;
        RECT 144.910 139.355 145.630 139.755 ;
        RECT 145.800 139.525 145.970 139.970 ;
        RECT 146.545 139.355 146.945 139.865 ;
        RECT 147.155 139.535 147.595 140.095 ;
        RECT 147.765 139.355 148.215 140.095 ;
        RECT 148.385 139.925 149.545 140.095 ;
        RECT 148.385 139.525 148.555 139.925 ;
        RECT 148.725 139.355 149.145 139.755 ;
        RECT 149.315 139.525 149.545 139.925 ;
        RECT 149.715 139.525 150.205 140.095 ;
        RECT 150.375 140.105 150.895 140.645 ;
        RECT 151.065 140.275 151.585 140.815 ;
        RECT 151.790 140.715 153.765 140.885 ;
        RECT 151.790 140.325 152.120 140.715 ;
        RECT 152.290 140.345 153.090 140.545 ;
        RECT 153.270 140.345 153.765 140.715 ;
        RECT 150.375 139.355 151.585 140.105 ;
        RECT 151.775 139.985 153.935 140.155 ;
        RECT 151.775 139.525 152.105 139.985 ;
        RECT 152.285 139.355 152.455 139.815 ;
        RECT 152.635 139.525 152.965 139.985 ;
        RECT 153.195 139.355 153.365 139.815 ;
        RECT 153.605 139.695 153.935 139.985 ;
        RECT 154.105 139.865 154.315 141.055 ;
        RECT 154.485 140.840 154.795 141.905 ;
        RECT 154.975 140.815 156.185 141.905 ;
        RECT 154.485 140.035 154.800 140.670 ;
        RECT 154.975 140.275 155.495 140.815 ;
        RECT 155.665 140.105 156.185 140.645 ;
        RECT 154.485 139.695 154.795 139.865 ;
        RECT 153.605 139.525 154.795 139.695 ;
        RECT 154.975 139.355 156.185 140.105 ;
        RECT 70.710 139.185 156.270 139.355 ;
        RECT 70.795 138.435 72.005 139.185 ;
        RECT 70.795 137.895 71.315 138.435 ;
        RECT 72.175 138.415 75.685 139.185 ;
        RECT 75.855 138.435 77.065 139.185 ;
        RECT 71.485 137.725 72.005 138.265 ;
        RECT 72.175 137.895 73.825 138.415 ;
        RECT 73.995 137.725 75.685 138.245 ;
        RECT 75.855 137.895 76.375 138.435 ;
        RECT 76.545 137.725 77.065 138.265 ;
        RECT 70.795 136.635 72.005 137.725 ;
        RECT 72.175 136.635 75.685 137.725 ;
        RECT 75.855 136.635 77.065 137.725 ;
        RECT 77.245 136.815 77.505 139.005 ;
        RECT 77.765 138.815 78.435 139.185 ;
        RECT 78.615 138.635 78.925 139.005 ;
        RECT 77.695 138.435 78.925 138.635 ;
        RECT 77.695 137.765 77.985 138.435 ;
        RECT 79.105 138.255 79.335 138.895 ;
        RECT 79.515 138.455 79.805 139.185 ;
        RECT 80.015 138.375 80.255 139.185 ;
        RECT 80.425 138.375 80.755 139.015 ;
        RECT 80.925 138.375 81.195 139.185 ;
        RECT 78.165 137.945 78.630 138.255 ;
        RECT 78.810 137.945 79.335 138.255 ;
        RECT 79.515 137.945 79.815 138.275 ;
        RECT 79.995 137.945 80.345 138.195 ;
        RECT 80.515 137.775 80.685 138.375 ;
        RECT 81.435 138.365 81.645 139.185 ;
        RECT 81.815 138.385 82.145 139.015 ;
        RECT 80.855 137.945 81.205 138.195 ;
        RECT 81.815 137.785 82.065 138.385 ;
        RECT 82.315 138.365 82.545 139.185 ;
        RECT 82.755 138.445 83.015 139.015 ;
        RECT 83.185 138.785 83.570 139.185 ;
        RECT 83.740 138.615 83.995 139.015 ;
        RECT 83.185 138.445 83.995 138.615 ;
        RECT 84.185 138.445 84.430 139.015 ;
        RECT 84.600 138.785 84.985 139.185 ;
        RECT 85.155 138.615 85.410 139.015 ;
        RECT 84.600 138.445 85.410 138.615 ;
        RECT 85.600 138.445 86.025 139.015 ;
        RECT 86.195 138.785 86.580 139.185 ;
        RECT 86.750 138.615 87.185 139.015 ;
        RECT 87.355 138.640 92.700 139.185 ;
        RECT 86.195 138.445 87.185 138.615 ;
        RECT 82.235 137.945 82.565 138.195 ;
        RECT 77.695 137.545 78.465 137.765 ;
        RECT 77.675 136.635 78.015 137.365 ;
        RECT 78.195 136.815 78.465 137.545 ;
        RECT 78.645 137.525 79.805 137.765 ;
        RECT 78.645 136.815 78.875 137.525 ;
        RECT 79.045 136.635 79.375 137.345 ;
        RECT 79.545 136.815 79.805 137.525 ;
        RECT 80.005 137.605 80.685 137.775 ;
        RECT 80.005 136.820 80.335 137.605 ;
        RECT 80.865 136.635 81.195 137.775 ;
        RECT 81.435 136.635 81.645 137.775 ;
        RECT 81.815 136.805 82.145 137.785 ;
        RECT 82.755 137.775 82.940 138.445 ;
        RECT 83.185 138.275 83.535 138.445 ;
        RECT 84.185 138.275 84.355 138.445 ;
        RECT 84.600 138.275 84.950 138.445 ;
        RECT 85.600 138.275 85.950 138.445 ;
        RECT 86.195 138.275 86.530 138.445 ;
        RECT 83.110 137.945 83.535 138.275 ;
        RECT 82.315 136.635 82.545 137.775 ;
        RECT 82.755 136.805 83.015 137.775 ;
        RECT 83.185 137.425 83.535 137.945 ;
        RECT 83.705 137.775 84.355 138.275 ;
        RECT 84.525 137.945 84.950 138.275 ;
        RECT 83.705 137.595 84.430 137.775 ;
        RECT 83.185 137.230 83.995 137.425 ;
        RECT 83.185 136.635 83.570 137.060 ;
        RECT 83.740 136.805 83.995 137.230 ;
        RECT 84.185 136.805 84.430 137.595 ;
        RECT 84.600 137.425 84.950 137.945 ;
        RECT 85.120 137.775 85.950 138.275 ;
        RECT 86.120 137.945 86.530 138.275 ;
        RECT 85.120 137.595 86.025 137.775 ;
        RECT 84.600 137.230 85.430 137.425 ;
        RECT 84.600 136.635 84.985 137.060 ;
        RECT 85.155 136.805 85.430 137.230 ;
        RECT 85.600 136.805 86.025 137.595 ;
        RECT 86.195 137.400 86.530 137.945 ;
        RECT 86.700 137.570 87.185 138.275 ;
        RECT 88.940 137.810 89.280 138.640 ;
        RECT 92.875 138.435 94.085 139.185 ;
        RECT 94.420 138.675 94.660 139.185 ;
        RECT 94.840 138.675 95.120 139.005 ;
        RECT 95.350 138.675 95.565 139.185 ;
        RECT 86.195 137.230 87.185 137.400 ;
        RECT 86.195 136.635 86.580 137.060 ;
        RECT 86.750 136.805 87.185 137.230 ;
        RECT 90.760 137.070 91.110 138.320 ;
        RECT 92.875 137.895 93.395 138.435 ;
        RECT 93.565 137.725 94.085 138.265 ;
        RECT 94.315 137.945 94.670 138.505 ;
        RECT 94.840 137.775 95.010 138.675 ;
        RECT 95.180 137.945 95.445 138.505 ;
        RECT 95.735 138.445 96.350 139.015 ;
        RECT 96.555 138.460 96.845 139.185 ;
        RECT 95.695 137.775 95.865 138.275 ;
        RECT 87.355 136.635 92.700 137.070 ;
        RECT 92.875 136.635 94.085 137.725 ;
        RECT 94.440 137.605 95.865 137.775 ;
        RECT 94.440 137.430 94.830 137.605 ;
        RECT 95.315 136.635 95.645 137.435 ;
        RECT 96.035 137.425 96.350 138.445 ;
        RECT 97.510 138.445 98.125 139.015 ;
        RECT 98.295 138.675 98.510 139.185 ;
        RECT 98.740 138.675 99.020 139.005 ;
        RECT 99.200 138.675 99.440 139.185 ;
        RECT 95.815 136.805 96.350 137.425 ;
        RECT 96.555 136.635 96.845 137.800 ;
        RECT 97.510 137.425 97.825 138.445 ;
        RECT 97.995 137.775 98.165 138.275 ;
        RECT 98.415 137.945 98.680 138.505 ;
        RECT 98.850 137.775 99.020 138.675 ;
        RECT 99.865 138.635 100.035 139.015 ;
        RECT 100.215 138.805 100.545 139.185 ;
        RECT 99.190 137.945 99.545 138.505 ;
        RECT 99.865 138.465 100.530 138.635 ;
        RECT 100.725 138.510 100.985 139.015 ;
        RECT 99.795 137.915 100.135 138.285 ;
        RECT 100.360 138.210 100.530 138.465 ;
        RECT 100.360 137.880 100.635 138.210 ;
        RECT 97.995 137.605 99.420 137.775 ;
        RECT 100.360 137.735 100.530 137.880 ;
        RECT 97.510 136.805 98.045 137.425 ;
        RECT 98.215 136.635 98.545 137.435 ;
        RECT 99.030 137.430 99.420 137.605 ;
        RECT 99.855 137.565 100.530 137.735 ;
        RECT 100.805 137.710 100.985 138.510 ;
        RECT 101.155 138.415 104.665 139.185 ;
        RECT 101.155 137.895 102.805 138.415 ;
        RECT 105.755 138.385 106.095 139.015 ;
        RECT 106.265 138.385 106.515 139.185 ;
        RECT 106.705 138.535 107.035 139.015 ;
        RECT 107.205 138.725 107.430 139.185 ;
        RECT 107.600 138.535 107.930 139.015 ;
        RECT 102.975 137.725 104.665 138.245 ;
        RECT 99.855 136.805 100.035 137.565 ;
        RECT 100.215 136.635 100.545 137.395 ;
        RECT 100.715 136.805 100.985 137.710 ;
        RECT 101.155 136.635 104.665 137.725 ;
        RECT 105.755 137.775 105.930 138.385 ;
        RECT 106.705 138.365 107.930 138.535 ;
        RECT 108.560 138.405 109.060 139.015 ;
        RECT 109.435 138.415 112.025 139.185 ;
        RECT 112.820 138.675 113.060 139.185 ;
        RECT 113.240 138.675 113.520 139.005 ;
        RECT 113.750 138.675 113.965 139.185 ;
        RECT 106.100 138.025 106.795 138.195 ;
        RECT 106.625 137.775 106.795 138.025 ;
        RECT 106.970 137.995 107.390 138.195 ;
        RECT 107.560 137.995 107.890 138.195 ;
        RECT 108.060 137.995 108.390 138.195 ;
        RECT 108.560 137.775 108.730 138.405 ;
        RECT 108.915 137.945 109.265 138.195 ;
        RECT 109.435 137.895 110.645 138.415 ;
        RECT 105.755 136.805 106.095 137.775 ;
        RECT 106.265 136.635 106.435 137.775 ;
        RECT 106.625 137.605 109.060 137.775 ;
        RECT 110.815 137.725 112.025 138.245 ;
        RECT 112.715 137.945 113.070 138.505 ;
        RECT 113.240 137.775 113.410 138.675 ;
        RECT 113.580 137.945 113.845 138.505 ;
        RECT 114.135 138.445 114.750 139.015 ;
        RECT 114.095 137.775 114.265 138.275 ;
        RECT 106.705 136.635 106.955 137.435 ;
        RECT 107.600 136.805 107.930 137.605 ;
        RECT 108.230 136.635 108.560 137.435 ;
        RECT 108.730 136.805 109.060 137.605 ;
        RECT 109.435 136.635 112.025 137.725 ;
        RECT 112.840 137.605 114.265 137.775 ;
        RECT 112.840 137.430 113.230 137.605 ;
        RECT 113.715 136.635 114.045 137.435 ;
        RECT 114.435 137.425 114.750 138.445 ;
        RECT 114.215 136.805 114.750 137.425 ;
        RECT 115.415 138.385 115.755 139.015 ;
        RECT 115.925 138.385 116.175 139.185 ;
        RECT 116.365 138.535 116.695 139.015 ;
        RECT 116.865 138.725 117.090 139.185 ;
        RECT 117.260 138.535 117.590 139.015 ;
        RECT 115.415 138.335 115.645 138.385 ;
        RECT 116.365 138.365 117.590 138.535 ;
        RECT 118.220 138.405 118.720 139.015 ;
        RECT 119.425 138.785 119.755 139.185 ;
        RECT 119.925 138.615 120.255 138.955 ;
        RECT 121.305 138.785 121.635 139.185 ;
        RECT 119.270 138.445 121.635 138.615 ;
        RECT 121.805 138.460 122.135 138.970 ;
        RECT 122.315 138.460 122.605 139.185 ;
        RECT 115.415 137.775 115.590 138.335 ;
        RECT 115.760 138.025 116.455 138.195 ;
        RECT 116.285 137.775 116.455 138.025 ;
        RECT 116.630 137.995 117.050 138.195 ;
        RECT 117.220 137.995 117.550 138.195 ;
        RECT 117.720 137.995 118.050 138.195 ;
        RECT 118.220 137.775 118.390 138.405 ;
        RECT 118.575 137.945 118.925 138.195 ;
        RECT 115.415 136.805 115.755 137.775 ;
        RECT 115.925 136.635 116.095 137.775 ;
        RECT 116.285 137.605 118.720 137.775 ;
        RECT 116.365 136.635 116.615 137.435 ;
        RECT 117.260 136.805 117.590 137.605 ;
        RECT 117.890 136.635 118.220 137.435 ;
        RECT 118.390 136.805 118.720 137.605 ;
        RECT 119.270 137.445 119.440 138.445 ;
        RECT 121.465 138.275 121.635 138.445 ;
        RECT 119.610 137.615 119.855 138.275 ;
        RECT 120.070 137.615 120.335 138.275 ;
        RECT 120.530 137.615 120.815 138.275 ;
        RECT 120.990 137.945 121.295 138.275 ;
        RECT 121.465 137.945 121.775 138.275 ;
        RECT 120.990 137.615 121.205 137.945 ;
        RECT 121.945 137.825 122.135 138.460 ;
        RECT 122.775 138.415 125.365 139.185 ;
        RECT 126.015 138.495 126.255 139.015 ;
        RECT 126.425 138.690 126.820 139.185 ;
        RECT 127.385 138.855 127.555 139.000 ;
        RECT 127.180 138.660 127.555 138.855 ;
        RECT 122.775 137.895 123.985 138.415 ;
        RECT 119.270 137.275 119.725 137.445 ;
        RECT 119.395 136.845 119.725 137.275 ;
        RECT 119.905 137.275 121.195 137.445 ;
        RECT 119.905 136.855 120.155 137.275 ;
        RECT 120.385 136.635 120.715 137.105 ;
        RECT 120.945 136.855 121.195 137.275 ;
        RECT 121.385 136.635 121.635 137.775 ;
        RECT 121.915 137.695 122.135 137.825 ;
        RECT 121.805 136.845 122.135 137.695 ;
        RECT 122.315 136.635 122.605 137.800 ;
        RECT 124.155 137.725 125.365 138.245 ;
        RECT 122.775 136.635 125.365 137.725 ;
        RECT 126.015 137.690 126.190 138.495 ;
        RECT 127.180 138.325 127.350 138.660 ;
        RECT 127.835 138.615 128.075 138.990 ;
        RECT 128.245 138.680 128.580 139.185 ;
        RECT 128.845 138.635 129.015 139.015 ;
        RECT 129.195 138.805 129.525 139.185 ;
        RECT 127.835 138.465 128.055 138.615 ;
        RECT 126.365 137.965 127.350 138.325 ;
        RECT 127.520 138.135 128.055 138.465 ;
        RECT 126.365 137.945 127.650 137.965 ;
        RECT 126.790 137.795 127.650 137.945 ;
        RECT 126.015 136.905 126.320 137.690 ;
        RECT 126.495 137.315 127.190 137.625 ;
        RECT 126.500 136.635 127.185 137.105 ;
        RECT 127.365 136.850 127.650 137.795 ;
        RECT 127.820 137.485 128.055 138.135 ;
        RECT 128.225 137.655 128.525 138.505 ;
        RECT 128.845 138.465 129.510 138.635 ;
        RECT 129.705 138.510 129.965 139.015 ;
        RECT 128.775 137.915 129.115 138.285 ;
        RECT 129.340 138.210 129.510 138.465 ;
        RECT 129.340 137.880 129.615 138.210 ;
        RECT 129.340 137.735 129.510 137.880 ;
        RECT 128.835 137.565 129.510 137.735 ;
        RECT 129.785 137.710 129.965 138.510 ;
        RECT 130.135 138.385 130.830 139.015 ;
        RECT 131.035 138.385 131.345 139.185 ;
        RECT 131.515 138.415 133.185 139.185 ;
        RECT 130.155 137.945 130.490 138.195 ;
        RECT 130.660 137.785 130.830 138.385 ;
        RECT 131.000 137.945 131.335 138.215 ;
        RECT 131.515 137.895 132.265 138.415 ;
        RECT 133.560 138.405 134.060 139.015 ;
        RECT 127.820 137.255 128.495 137.485 ;
        RECT 127.825 136.635 128.155 137.085 ;
        RECT 128.325 136.825 128.495 137.255 ;
        RECT 128.835 136.805 129.015 137.565 ;
        RECT 129.195 136.635 129.525 137.395 ;
        RECT 129.695 136.805 129.965 137.710 ;
        RECT 130.135 136.635 130.395 137.775 ;
        RECT 130.565 136.805 130.895 137.785 ;
        RECT 131.065 136.635 131.345 137.775 ;
        RECT 132.435 137.725 133.185 138.245 ;
        RECT 133.355 137.945 133.705 138.195 ;
        RECT 133.890 137.775 134.060 138.405 ;
        RECT 134.690 138.535 135.020 139.015 ;
        RECT 135.190 138.725 135.415 139.185 ;
        RECT 135.585 138.535 135.915 139.015 ;
        RECT 134.690 138.365 135.915 138.535 ;
        RECT 136.105 138.385 136.355 139.185 ;
        RECT 136.525 138.385 136.865 139.015 ;
        RECT 137.035 138.385 137.730 139.015 ;
        RECT 137.935 138.385 138.245 139.185 ;
        RECT 138.745 138.785 139.075 139.185 ;
        RECT 139.245 138.615 139.575 138.955 ;
        RECT 140.625 138.785 140.955 139.185 ;
        RECT 138.590 138.445 140.955 138.615 ;
        RECT 141.125 138.460 141.455 138.970 ;
        RECT 134.230 137.995 134.560 138.195 ;
        RECT 134.730 137.995 135.060 138.195 ;
        RECT 135.230 137.995 135.650 138.195 ;
        RECT 135.825 138.025 136.520 138.195 ;
        RECT 135.825 137.775 135.995 138.025 ;
        RECT 136.690 137.775 136.865 138.385 ;
        RECT 137.055 137.945 137.390 138.195 ;
        RECT 137.560 137.785 137.730 138.385 ;
        RECT 137.900 137.945 138.235 138.215 ;
        RECT 131.515 136.635 133.185 137.725 ;
        RECT 133.560 137.605 135.995 137.775 ;
        RECT 133.560 136.805 133.890 137.605 ;
        RECT 134.060 136.635 134.390 137.435 ;
        RECT 134.690 136.805 135.020 137.605 ;
        RECT 135.665 136.635 135.915 137.435 ;
        RECT 136.185 136.635 136.355 137.775 ;
        RECT 136.525 136.805 136.865 137.775 ;
        RECT 137.035 136.635 137.295 137.775 ;
        RECT 137.465 136.805 137.795 137.785 ;
        RECT 137.965 136.635 138.245 137.775 ;
        RECT 138.590 137.445 138.760 138.445 ;
        RECT 140.785 138.275 140.955 138.445 ;
        RECT 138.930 137.615 139.175 138.275 ;
        RECT 139.390 137.615 139.655 138.275 ;
        RECT 139.850 137.615 140.135 138.275 ;
        RECT 140.310 137.945 140.615 138.275 ;
        RECT 140.785 137.945 141.095 138.275 ;
        RECT 140.310 137.615 140.525 137.945 ;
        RECT 138.590 137.275 139.045 137.445 ;
        RECT 138.715 136.845 139.045 137.275 ;
        RECT 139.225 137.275 140.515 137.445 ;
        RECT 139.225 136.855 139.475 137.275 ;
        RECT 139.705 136.635 140.035 137.105 ;
        RECT 140.265 136.855 140.515 137.275 ;
        RECT 140.705 136.635 140.955 137.775 ;
        RECT 141.265 137.695 141.455 138.460 ;
        RECT 141.635 138.615 142.070 139.015 ;
        RECT 142.240 138.785 142.625 139.185 ;
        RECT 141.635 138.445 142.625 138.615 ;
        RECT 142.795 138.445 143.220 139.015 ;
        RECT 143.410 138.615 143.665 139.015 ;
        RECT 143.835 138.785 144.220 139.185 ;
        RECT 143.410 138.445 144.220 138.615 ;
        RECT 144.390 138.445 144.635 139.015 ;
        RECT 144.825 138.615 145.080 139.015 ;
        RECT 145.250 138.785 145.635 139.185 ;
        RECT 144.825 138.445 145.635 138.615 ;
        RECT 145.805 138.445 146.065 139.015 ;
        RECT 142.290 138.275 142.625 138.445 ;
        RECT 142.870 138.275 143.220 138.445 ;
        RECT 143.870 138.275 144.220 138.445 ;
        RECT 144.465 138.275 144.635 138.445 ;
        RECT 145.285 138.275 145.635 138.445 ;
        RECT 141.125 136.845 141.455 137.695 ;
        RECT 141.635 137.570 142.120 138.275 ;
        RECT 142.290 137.945 142.700 138.275 ;
        RECT 142.290 137.400 142.625 137.945 ;
        RECT 142.870 137.775 143.700 138.275 ;
        RECT 141.635 137.230 142.625 137.400 ;
        RECT 142.795 137.595 143.700 137.775 ;
        RECT 143.870 137.945 144.295 138.275 ;
        RECT 141.635 136.805 142.070 137.230 ;
        RECT 142.240 136.635 142.625 137.060 ;
        RECT 142.795 136.805 143.220 137.595 ;
        RECT 143.870 137.425 144.220 137.945 ;
        RECT 144.465 137.775 145.115 138.275 ;
        RECT 143.390 137.230 144.220 137.425 ;
        RECT 144.390 137.595 145.115 137.775 ;
        RECT 145.285 137.945 145.710 138.275 ;
        RECT 143.390 136.805 143.665 137.230 ;
        RECT 143.835 136.635 144.220 137.060 ;
        RECT 144.390 136.805 144.635 137.595 ;
        RECT 145.285 137.425 145.635 137.945 ;
        RECT 145.880 137.775 146.065 138.445 ;
        RECT 146.235 138.415 147.905 139.185 ;
        RECT 148.075 138.460 148.365 139.185 ;
        RECT 146.235 137.895 146.985 138.415 ;
        RECT 148.535 138.350 148.825 139.185 ;
        RECT 148.995 138.785 149.950 138.955 ;
        RECT 150.365 138.795 150.695 139.185 ;
        RECT 144.825 137.230 145.635 137.425 ;
        RECT 144.825 136.805 145.080 137.230 ;
        RECT 145.250 136.635 145.635 137.060 ;
        RECT 145.805 136.805 146.065 137.775 ;
        RECT 147.155 137.725 147.905 138.245 ;
        RECT 148.995 137.905 149.165 138.785 ;
        RECT 150.865 138.615 151.035 138.935 ;
        RECT 151.205 138.795 151.535 139.185 ;
        RECT 149.335 138.445 151.585 138.615 ;
        RECT 149.335 137.945 149.565 138.445 ;
        RECT 149.735 138.025 150.110 138.195 ;
        RECT 146.235 136.635 147.905 137.725 ;
        RECT 148.075 136.635 148.365 137.800 ;
        RECT 148.535 137.735 149.165 137.905 ;
        RECT 149.940 137.825 150.110 138.025 ;
        RECT 150.280 137.995 150.830 138.195 ;
        RECT 151.000 137.825 151.245 138.275 ;
        RECT 148.535 136.805 148.855 137.735 ;
        RECT 149.940 137.655 151.245 137.825 ;
        RECT 151.415 137.485 151.585 138.445 ;
        RECT 151.780 138.535 152.090 139.005 ;
        RECT 152.260 138.705 152.995 139.185 ;
        RECT 153.165 138.615 153.335 138.965 ;
        RECT 153.505 138.785 153.885 139.185 ;
        RECT 151.780 138.365 152.515 138.535 ;
        RECT 153.165 138.445 153.905 138.615 ;
        RECT 154.075 138.510 154.345 138.855 ;
        RECT 152.265 138.275 152.515 138.365 ;
        RECT 153.735 138.275 153.905 138.445 ;
        RECT 151.760 137.945 152.095 138.195 ;
        RECT 152.265 137.945 153.005 138.275 ;
        RECT 153.735 137.945 153.965 138.275 ;
        RECT 149.035 137.315 150.275 137.485 ;
        RECT 149.035 136.805 149.435 137.315 ;
        RECT 149.605 136.635 149.775 137.145 ;
        RECT 149.945 136.805 150.275 137.315 ;
        RECT 150.445 136.635 150.615 137.485 ;
        RECT 151.205 136.805 151.585 137.485 ;
        RECT 151.760 136.635 152.015 137.775 ;
        RECT 152.265 137.385 152.435 137.945 ;
        RECT 153.735 137.775 153.905 137.945 ;
        RECT 154.175 137.775 154.345 138.510 ;
        RECT 154.975 138.435 156.185 139.185 ;
        RECT 152.660 137.605 153.905 137.775 ;
        RECT 152.660 137.355 153.080 137.605 ;
        RECT 152.210 136.855 153.405 137.185 ;
        RECT 153.585 136.635 153.865 137.435 ;
        RECT 154.075 136.805 154.345 137.775 ;
        RECT 154.975 137.725 155.495 138.265 ;
        RECT 155.665 137.895 156.185 138.435 ;
        RECT 154.975 136.635 156.185 137.725 ;
        RECT 70.710 136.465 156.270 136.635 ;
        RECT 70.795 135.375 72.005 136.465 ;
        RECT 72.175 135.375 74.765 136.465 ;
        RECT 75.395 135.955 75.695 136.465 ;
        RECT 75.865 135.785 76.195 136.295 ;
        RECT 76.365 135.955 76.995 136.465 ;
        RECT 77.575 135.955 77.955 136.125 ;
        RECT 78.125 135.955 78.425 136.465 ;
        RECT 77.785 135.785 77.955 135.955 ;
        RECT 70.795 134.665 71.315 135.205 ;
        RECT 71.485 134.835 72.005 135.375 ;
        RECT 72.175 134.685 73.385 135.205 ;
        RECT 73.555 134.855 74.765 135.375 ;
        RECT 75.395 135.615 77.615 135.785 ;
        RECT 70.795 133.915 72.005 134.665 ;
        RECT 72.175 133.915 74.765 134.685 ;
        RECT 75.395 134.655 75.565 135.615 ;
        RECT 75.735 135.275 77.275 135.445 ;
        RECT 75.735 134.825 75.980 135.275 ;
        RECT 76.240 134.905 76.935 135.105 ;
        RECT 77.105 135.075 77.275 135.275 ;
        RECT 77.445 135.415 77.615 135.615 ;
        RECT 77.785 135.585 78.445 135.785 ;
        RECT 77.445 135.245 78.105 135.415 ;
        RECT 77.105 134.905 77.705 135.075 ;
        RECT 77.935 134.825 78.105 135.245 ;
        RECT 75.395 134.110 75.860 134.655 ;
        RECT 76.365 133.915 76.535 134.735 ;
        RECT 76.705 134.655 77.615 134.735 ;
        RECT 78.275 134.655 78.445 135.585 ;
        RECT 78.625 135.495 78.955 136.280 ;
        RECT 78.625 135.325 79.305 135.495 ;
        RECT 79.485 135.325 79.815 136.465 ;
        RECT 79.995 135.375 83.505 136.465 ;
        RECT 78.615 134.905 78.965 135.155 ;
        RECT 79.135 134.725 79.305 135.325 ;
        RECT 79.475 134.905 79.825 135.155 ;
        RECT 76.705 134.565 77.955 134.655 ;
        RECT 76.705 134.085 77.035 134.565 ;
        RECT 77.445 134.485 77.955 134.565 ;
        RECT 77.205 133.915 77.555 134.305 ;
        RECT 77.725 134.085 77.955 134.485 ;
        RECT 78.125 134.175 78.445 134.655 ;
        RECT 78.635 133.915 78.875 134.725 ;
        RECT 79.045 134.085 79.375 134.725 ;
        RECT 79.545 133.915 79.815 134.725 ;
        RECT 79.995 134.685 81.645 135.205 ;
        RECT 81.815 134.855 83.505 135.375 ;
        RECT 83.675 135.300 83.965 136.465 ;
        RECT 84.135 135.375 85.805 136.465 ;
        RECT 84.135 134.685 84.885 135.205 ;
        RECT 85.055 134.855 85.805 135.375 ;
        RECT 86.445 135.325 86.775 136.465 ;
        RECT 87.305 135.495 87.635 136.280 ;
        RECT 88.015 135.795 88.295 136.465 ;
        RECT 88.465 135.575 88.765 136.125 ;
        RECT 88.965 135.745 89.295 136.465 ;
        RECT 89.485 135.745 89.945 136.295 ;
        RECT 86.955 135.325 87.635 135.495 ;
        RECT 86.435 134.905 86.785 135.155 ;
        RECT 86.955 134.725 87.125 135.325 ;
        RECT 87.830 135.155 88.095 135.515 ;
        RECT 88.465 135.405 89.405 135.575 ;
        RECT 89.235 135.155 89.405 135.405 ;
        RECT 87.295 134.905 87.645 135.155 ;
        RECT 87.830 134.905 88.505 135.155 ;
        RECT 88.725 134.905 89.065 135.155 ;
        RECT 89.235 134.825 89.525 135.155 ;
        RECT 89.235 134.735 89.405 134.825 ;
        RECT 79.995 133.915 83.505 134.685 ;
        RECT 83.675 133.915 83.965 134.640 ;
        RECT 84.135 133.915 85.805 134.685 ;
        RECT 86.445 133.915 86.715 134.725 ;
        RECT 86.885 134.085 87.215 134.725 ;
        RECT 87.385 133.915 87.625 134.725 ;
        RECT 88.015 134.545 89.405 134.735 ;
        RECT 88.015 134.185 88.345 134.545 ;
        RECT 89.695 134.375 89.945 135.745 ;
        RECT 88.965 133.915 89.215 134.375 ;
        RECT 89.385 134.085 89.945 134.375 ;
        RECT 90.115 135.745 90.575 136.295 ;
        RECT 90.765 135.745 91.095 136.465 ;
        RECT 90.115 134.375 90.365 135.745 ;
        RECT 91.295 135.575 91.595 136.125 ;
        RECT 91.765 135.795 92.045 136.465 ;
        RECT 90.655 135.405 91.595 135.575 ;
        RECT 90.655 135.155 90.825 135.405 ;
        RECT 91.965 135.155 92.230 135.515 ;
        RECT 92.415 135.375 94.085 136.465 ;
        RECT 90.535 134.825 90.825 135.155 ;
        RECT 90.995 134.905 91.335 135.155 ;
        RECT 91.555 134.905 92.230 135.155 ;
        RECT 90.655 134.735 90.825 134.825 ;
        RECT 90.655 134.545 92.045 134.735 ;
        RECT 90.115 134.085 90.675 134.375 ;
        RECT 90.845 133.915 91.095 134.375 ;
        RECT 91.715 134.185 92.045 134.545 ;
        RECT 92.415 134.685 93.165 135.205 ;
        RECT 93.335 134.855 94.085 135.375 ;
        RECT 94.255 135.325 94.535 136.465 ;
        RECT 94.705 135.315 95.035 136.295 ;
        RECT 95.205 135.325 95.465 136.465 ;
        RECT 95.640 135.745 95.975 136.255 ;
        RECT 94.265 134.885 94.600 135.155 ;
        RECT 94.770 134.765 94.940 135.315 ;
        RECT 95.110 134.905 95.445 135.155 ;
        RECT 94.770 134.715 94.945 134.765 ;
        RECT 92.415 133.915 94.085 134.685 ;
        RECT 94.255 133.915 94.565 134.715 ;
        RECT 94.770 134.085 95.465 134.715 ;
        RECT 95.640 134.390 95.895 135.745 ;
        RECT 96.225 135.665 96.555 136.465 ;
        RECT 96.800 135.875 97.085 136.295 ;
        RECT 97.340 136.045 97.670 136.465 ;
        RECT 97.895 136.125 99.055 136.295 ;
        RECT 97.895 135.875 98.225 136.125 ;
        RECT 96.800 135.705 98.225 135.875 ;
        RECT 98.455 135.495 98.625 135.955 ;
        RECT 98.885 135.625 99.055 136.125 ;
        RECT 99.615 135.825 99.945 136.255 ;
        RECT 99.490 135.655 99.945 135.825 ;
        RECT 100.125 135.825 100.375 136.245 ;
        RECT 100.605 135.995 100.935 136.465 ;
        RECT 101.165 135.825 101.415 136.245 ;
        RECT 100.125 135.655 101.415 135.825 ;
        RECT 96.255 135.325 98.625 135.495 ;
        RECT 96.255 135.155 96.425 135.325 ;
        RECT 98.875 135.155 99.080 135.445 ;
        RECT 96.120 134.825 96.425 135.155 ;
        RECT 96.620 135.105 96.870 135.155 ;
        RECT 97.080 135.105 97.350 135.155 ;
        RECT 97.540 135.105 97.830 135.155 ;
        RECT 96.615 134.935 96.870 135.105 ;
        RECT 97.075 134.935 97.350 135.105 ;
        RECT 97.535 134.935 97.830 135.105 ;
        RECT 96.620 134.825 96.870 134.935 ;
        RECT 96.255 134.655 96.425 134.825 ;
        RECT 96.255 134.485 96.815 134.655 ;
        RECT 97.080 134.495 97.350 134.935 ;
        RECT 97.540 134.495 97.830 134.935 ;
        RECT 98.000 134.490 98.420 135.155 ;
        RECT 98.730 135.105 99.080 135.155 ;
        RECT 98.730 134.935 99.085 135.105 ;
        RECT 98.730 134.825 99.080 134.935 ;
        RECT 99.490 134.655 99.660 135.655 ;
        RECT 99.830 134.825 100.075 135.485 ;
        RECT 100.290 134.825 100.555 135.485 ;
        RECT 100.750 134.825 101.035 135.485 ;
        RECT 101.210 135.155 101.425 135.485 ;
        RECT 101.605 135.325 101.855 136.465 ;
        RECT 102.025 135.405 102.355 136.255 ;
        RECT 101.210 134.825 101.515 135.155 ;
        RECT 101.685 134.825 101.995 135.155 ;
        RECT 101.685 134.655 101.855 134.825 ;
        RECT 95.640 134.130 95.975 134.390 ;
        RECT 96.645 134.315 96.815 134.485 ;
        RECT 96.145 133.915 96.475 134.315 ;
        RECT 96.645 134.145 98.260 134.315 ;
        RECT 98.805 133.915 99.135 134.635 ;
        RECT 99.490 134.485 101.855 134.655 ;
        RECT 102.165 134.640 102.355 135.405 ;
        RECT 103.075 135.535 103.255 136.295 ;
        RECT 103.435 135.705 103.765 136.465 ;
        RECT 103.075 135.365 103.750 135.535 ;
        RECT 103.935 135.390 104.205 136.295 ;
        RECT 103.580 135.220 103.750 135.365 ;
        RECT 103.015 134.815 103.355 135.185 ;
        RECT 103.580 134.890 103.855 135.220 ;
        RECT 99.645 133.915 99.975 134.315 ;
        RECT 100.145 134.145 100.475 134.485 ;
        RECT 101.525 133.915 101.855 134.315 ;
        RECT 102.025 134.130 102.355 134.640 ;
        RECT 103.580 134.635 103.750 134.890 ;
        RECT 103.085 134.465 103.750 134.635 ;
        RECT 104.025 134.590 104.205 135.390 ;
        RECT 104.455 135.535 104.635 136.295 ;
        RECT 104.815 135.705 105.145 136.465 ;
        RECT 104.455 135.365 105.130 135.535 ;
        RECT 105.315 135.390 105.585 136.295 ;
        RECT 106.055 135.825 106.385 136.255 ;
        RECT 104.960 135.220 105.130 135.365 ;
        RECT 104.395 134.815 104.735 135.185 ;
        RECT 104.960 134.890 105.235 135.220 ;
        RECT 104.960 134.635 105.130 134.890 ;
        RECT 103.085 134.085 103.255 134.465 ;
        RECT 103.435 133.915 103.765 134.295 ;
        RECT 103.945 134.085 104.205 134.590 ;
        RECT 104.465 134.465 105.130 134.635 ;
        RECT 105.405 134.590 105.585 135.390 ;
        RECT 104.465 134.085 104.635 134.465 ;
        RECT 104.815 133.915 105.145 134.295 ;
        RECT 105.325 134.085 105.585 134.590 ;
        RECT 105.930 135.655 106.385 135.825 ;
        RECT 106.565 135.825 106.815 136.245 ;
        RECT 107.045 135.995 107.375 136.465 ;
        RECT 107.605 135.825 107.855 136.245 ;
        RECT 106.565 135.655 107.855 135.825 ;
        RECT 105.930 134.655 106.100 135.655 ;
        RECT 106.270 134.825 106.515 135.485 ;
        RECT 106.730 134.825 106.995 135.485 ;
        RECT 107.190 134.825 107.475 135.485 ;
        RECT 107.650 135.155 107.865 135.485 ;
        RECT 108.045 135.325 108.295 136.465 ;
        RECT 108.465 135.405 108.795 136.255 ;
        RECT 107.650 134.825 107.955 135.155 ;
        RECT 108.125 134.825 108.435 135.155 ;
        RECT 108.125 134.655 108.295 134.825 ;
        RECT 105.930 134.485 108.295 134.655 ;
        RECT 108.605 134.640 108.795 135.405 ;
        RECT 109.435 135.300 109.725 136.465 ;
        RECT 109.895 135.375 113.405 136.465 ;
        RECT 113.575 135.375 114.785 136.465 ;
        RECT 109.895 134.685 111.545 135.205 ;
        RECT 111.715 134.855 113.405 135.375 ;
        RECT 106.085 133.915 106.415 134.315 ;
        RECT 106.585 134.145 106.915 134.485 ;
        RECT 107.965 133.915 108.295 134.315 ;
        RECT 108.465 134.130 108.795 134.640 ;
        RECT 109.435 133.915 109.725 134.640 ;
        RECT 109.895 133.915 113.405 134.685 ;
        RECT 113.575 134.665 114.095 135.205 ;
        RECT 114.265 134.835 114.785 135.375 ;
        RECT 114.965 135.405 115.295 136.255 ;
        RECT 113.575 133.915 114.785 134.665 ;
        RECT 114.965 134.640 115.155 135.405 ;
        RECT 115.465 135.325 115.715 136.465 ;
        RECT 115.905 135.825 116.155 136.245 ;
        RECT 116.385 135.995 116.715 136.465 ;
        RECT 116.945 135.825 117.195 136.245 ;
        RECT 115.905 135.655 117.195 135.825 ;
        RECT 117.375 135.825 117.705 136.255 ;
        RECT 118.175 136.030 123.520 136.465 ;
        RECT 117.375 135.655 117.830 135.825 ;
        RECT 115.895 135.155 116.110 135.485 ;
        RECT 115.325 134.825 115.635 135.155 ;
        RECT 115.805 134.825 116.110 135.155 ;
        RECT 116.285 134.825 116.570 135.485 ;
        RECT 116.765 134.825 117.030 135.485 ;
        RECT 117.245 134.825 117.490 135.485 ;
        RECT 115.465 134.655 115.635 134.825 ;
        RECT 117.660 134.655 117.830 135.655 ;
        RECT 114.965 134.130 115.295 134.640 ;
        RECT 115.465 134.485 117.830 134.655 ;
        RECT 115.465 133.915 115.795 134.315 ;
        RECT 116.845 134.145 117.175 134.485 ;
        RECT 119.760 134.460 120.100 135.290 ;
        RECT 121.580 134.780 121.930 136.030 ;
        RECT 123.695 135.375 126.285 136.465 ;
        RECT 123.695 134.685 124.905 135.205 ;
        RECT 125.075 134.855 126.285 135.375 ;
        RECT 126.920 135.515 127.185 136.285 ;
        RECT 127.355 135.745 127.685 136.465 ;
        RECT 127.875 135.925 128.135 136.285 ;
        RECT 128.305 136.095 128.635 136.465 ;
        RECT 128.805 135.925 129.065 136.285 ;
        RECT 127.875 135.695 129.065 135.925 ;
        RECT 129.635 135.515 129.925 136.285 ;
        RECT 117.345 133.915 117.675 134.315 ;
        RECT 118.175 133.915 123.520 134.460 ;
        RECT 123.695 133.915 126.285 134.685 ;
        RECT 126.920 134.095 127.255 135.515 ;
        RECT 127.430 135.335 129.925 135.515 ;
        RECT 130.135 135.375 133.645 136.465 ;
        RECT 127.430 134.645 127.655 135.335 ;
        RECT 127.855 134.825 128.135 135.155 ;
        RECT 128.315 134.825 128.890 135.155 ;
        RECT 129.070 134.825 129.505 135.155 ;
        RECT 129.685 134.825 129.955 135.155 ;
        RECT 130.135 134.685 131.785 135.205 ;
        RECT 131.955 134.855 133.645 135.375 ;
        RECT 133.895 135.535 134.075 136.295 ;
        RECT 134.255 135.705 134.585 136.465 ;
        RECT 133.895 135.365 134.570 135.535 ;
        RECT 134.755 135.390 135.025 136.295 ;
        RECT 134.400 135.220 134.570 135.365 ;
        RECT 133.835 134.815 134.175 135.185 ;
        RECT 134.400 134.890 134.675 135.220 ;
        RECT 127.430 134.455 129.915 134.645 ;
        RECT 127.435 133.915 128.180 134.285 ;
        RECT 128.745 134.095 129.000 134.455 ;
        RECT 129.180 133.915 129.510 134.285 ;
        RECT 129.690 134.095 129.915 134.455 ;
        RECT 130.135 133.915 133.645 134.685 ;
        RECT 134.400 134.635 134.570 134.890 ;
        RECT 133.905 134.465 134.570 134.635 ;
        RECT 134.845 134.590 135.025 135.390 ;
        RECT 135.195 135.300 135.485 136.465 ;
        RECT 135.665 135.405 135.995 136.255 ;
        RECT 135.665 135.275 135.885 135.405 ;
        RECT 136.165 135.325 136.415 136.465 ;
        RECT 136.605 135.825 136.855 136.245 ;
        RECT 137.085 135.995 137.415 136.465 ;
        RECT 137.645 135.825 137.895 136.245 ;
        RECT 136.605 135.655 137.895 135.825 ;
        RECT 138.075 135.825 138.405 136.255 ;
        RECT 138.075 135.655 138.530 135.825 ;
        RECT 135.665 134.640 135.855 135.275 ;
        RECT 136.595 135.155 136.810 135.485 ;
        RECT 136.025 134.825 136.335 135.155 ;
        RECT 136.505 134.825 136.810 135.155 ;
        RECT 136.985 134.825 137.270 135.485 ;
        RECT 137.465 134.825 137.730 135.485 ;
        RECT 137.945 134.825 138.190 135.485 ;
        RECT 136.165 134.655 136.335 134.825 ;
        RECT 138.360 134.655 138.530 135.655 ;
        RECT 133.905 134.085 134.075 134.465 ;
        RECT 134.255 133.915 134.585 134.295 ;
        RECT 134.765 134.085 135.025 134.590 ;
        RECT 135.195 133.915 135.485 134.640 ;
        RECT 135.665 134.130 135.995 134.640 ;
        RECT 136.165 134.485 138.530 134.655 ;
        RECT 138.910 135.675 139.445 136.295 ;
        RECT 138.910 134.655 139.225 135.675 ;
        RECT 139.615 135.665 139.945 136.465 ;
        RECT 140.430 135.495 140.820 135.670 ;
        RECT 139.395 135.325 140.820 135.495 ;
        RECT 141.175 135.375 143.765 136.465 ;
        RECT 144.395 135.870 144.830 136.295 ;
        RECT 145.000 136.040 145.385 136.465 ;
        RECT 144.395 135.700 145.385 135.870 ;
        RECT 139.395 134.825 139.565 135.325 ;
        RECT 136.165 133.915 136.495 134.315 ;
        RECT 137.545 134.145 137.875 134.485 ;
        RECT 138.045 133.915 138.375 134.315 ;
        RECT 138.910 134.085 139.525 134.655 ;
        RECT 139.815 134.595 140.080 135.155 ;
        RECT 140.250 134.425 140.420 135.325 ;
        RECT 140.590 134.595 140.945 135.155 ;
        RECT 141.175 134.685 142.385 135.205 ;
        RECT 142.555 134.855 143.765 135.375 ;
        RECT 144.395 134.825 144.880 135.530 ;
        RECT 145.050 135.155 145.385 135.700 ;
        RECT 145.555 135.505 145.980 136.295 ;
        RECT 146.150 135.870 146.425 136.295 ;
        RECT 146.595 136.040 146.980 136.465 ;
        RECT 146.150 135.675 146.980 135.870 ;
        RECT 145.555 135.325 146.460 135.505 ;
        RECT 145.050 134.825 145.460 135.155 ;
        RECT 145.630 134.825 146.460 135.325 ;
        RECT 146.630 135.155 146.980 135.675 ;
        RECT 147.150 135.505 147.395 136.295 ;
        RECT 147.585 135.870 147.840 136.295 ;
        RECT 148.010 136.040 148.395 136.465 ;
        RECT 147.585 135.675 148.395 135.870 ;
        RECT 147.150 135.325 147.875 135.505 ;
        RECT 146.630 134.825 147.055 135.155 ;
        RECT 147.225 134.825 147.875 135.325 ;
        RECT 148.045 135.155 148.395 135.675 ;
        RECT 148.565 135.325 148.825 136.295 ;
        RECT 150.005 135.535 150.175 136.295 ;
        RECT 150.390 135.705 150.720 136.465 ;
        RECT 150.005 135.365 150.720 135.535 ;
        RECT 150.890 135.390 151.145 136.295 ;
        RECT 148.045 134.825 148.470 135.155 ;
        RECT 139.695 133.915 139.910 134.425 ;
        RECT 140.140 134.095 140.420 134.425 ;
        RECT 140.600 133.915 140.840 134.425 ;
        RECT 141.175 133.915 143.765 134.685 ;
        RECT 145.050 134.655 145.385 134.825 ;
        RECT 145.630 134.655 145.980 134.825 ;
        RECT 146.630 134.655 146.980 134.825 ;
        RECT 147.225 134.655 147.395 134.825 ;
        RECT 148.045 134.655 148.395 134.825 ;
        RECT 148.640 134.655 148.825 135.325 ;
        RECT 149.915 134.815 150.270 135.185 ;
        RECT 150.550 135.155 150.720 135.365 ;
        RECT 150.550 134.825 150.805 135.155 ;
        RECT 144.395 134.485 145.385 134.655 ;
        RECT 144.395 134.085 144.830 134.485 ;
        RECT 145.000 133.915 145.385 134.315 ;
        RECT 145.555 134.085 145.980 134.655 ;
        RECT 146.170 134.485 146.980 134.655 ;
        RECT 146.170 134.085 146.425 134.485 ;
        RECT 146.595 133.915 146.980 134.315 ;
        RECT 147.150 134.085 147.395 134.655 ;
        RECT 147.585 134.485 148.395 134.655 ;
        RECT 147.585 134.085 147.840 134.485 ;
        RECT 148.010 133.915 148.395 134.315 ;
        RECT 148.565 134.085 148.825 134.655 ;
        RECT 150.550 134.635 150.720 134.825 ;
        RECT 150.975 134.660 151.145 135.390 ;
        RECT 151.320 135.315 151.580 136.465 ;
        RECT 151.760 135.325 152.080 136.465 ;
        RECT 152.260 135.155 152.455 136.205 ;
        RECT 152.635 135.615 152.965 136.295 ;
        RECT 153.165 135.665 153.420 136.465 ;
        RECT 152.635 135.335 152.985 135.615 ;
        RECT 151.820 135.105 152.080 135.155 ;
        RECT 151.815 134.935 152.080 135.105 ;
        RECT 151.820 134.825 152.080 134.935 ;
        RECT 152.260 134.825 152.645 135.155 ;
        RECT 152.815 134.955 152.985 135.335 ;
        RECT 153.175 135.125 153.420 135.485 ;
        RECT 153.595 135.325 153.875 136.465 ;
        RECT 154.045 135.315 154.375 136.295 ;
        RECT 154.545 135.325 154.805 136.465 ;
        RECT 154.975 135.375 156.185 136.465 ;
        RECT 152.815 134.785 153.335 134.955 ;
        RECT 153.605 134.885 153.940 135.155 ;
        RECT 153.165 134.765 153.335 134.785 ;
        RECT 150.005 134.465 150.720 134.635 ;
        RECT 150.005 134.085 150.175 134.465 ;
        RECT 150.390 133.915 150.720 134.295 ;
        RECT 150.890 134.085 151.145 134.660 ;
        RECT 151.320 133.915 151.580 134.755 ;
        RECT 151.760 134.445 152.975 134.615 ;
        RECT 151.760 134.095 152.050 134.445 ;
        RECT 152.245 133.915 152.575 134.275 ;
        RECT 152.745 134.140 152.975 134.445 ;
        RECT 153.165 134.595 153.365 134.765 ;
        RECT 154.110 134.715 154.280 135.315 ;
        RECT 154.450 134.905 154.785 135.155 ;
        RECT 154.975 134.835 155.495 135.375 ;
        RECT 153.165 134.220 153.335 134.595 ;
        RECT 153.595 133.915 153.905 134.715 ;
        RECT 154.110 134.085 154.805 134.715 ;
        RECT 155.665 134.665 156.185 135.205 ;
        RECT 154.975 133.915 156.185 134.665 ;
        RECT 70.710 133.745 156.270 133.915 ;
        RECT 70.795 132.995 72.005 133.745 ;
        RECT 72.175 133.005 72.640 133.550 ;
        RECT 70.795 132.455 71.315 132.995 ;
        RECT 71.485 132.285 72.005 132.825 ;
        RECT 70.795 131.195 72.005 132.285 ;
        RECT 72.175 132.045 72.345 133.005 ;
        RECT 73.145 132.925 73.315 133.745 ;
        RECT 73.485 133.095 73.815 133.575 ;
        RECT 73.985 133.355 74.335 133.745 ;
        RECT 74.505 133.175 74.735 133.575 ;
        RECT 74.225 133.095 74.735 133.175 ;
        RECT 73.485 133.005 74.735 133.095 ;
        RECT 74.905 133.005 75.225 133.485 ;
        RECT 75.395 133.200 80.740 133.745 ;
        RECT 73.485 132.925 74.395 133.005 ;
        RECT 72.515 132.385 72.760 132.835 ;
        RECT 73.020 132.555 73.715 132.755 ;
        RECT 73.885 132.585 74.485 132.755 ;
        RECT 73.885 132.385 74.055 132.585 ;
        RECT 74.715 132.415 74.885 132.835 ;
        RECT 72.515 132.215 74.055 132.385 ;
        RECT 74.225 132.245 74.885 132.415 ;
        RECT 74.225 132.045 74.395 132.245 ;
        RECT 75.055 132.075 75.225 133.005 ;
        RECT 76.980 132.370 77.320 133.200 ;
        RECT 80.915 132.975 82.585 133.745 ;
        RECT 83.220 133.005 83.555 133.745 ;
        RECT 72.175 131.875 74.395 132.045 ;
        RECT 74.565 131.875 75.225 132.075 ;
        RECT 72.175 131.195 72.475 131.705 ;
        RECT 72.645 131.365 72.975 131.875 ;
        RECT 74.565 131.705 74.735 131.875 ;
        RECT 73.145 131.195 73.775 131.705 ;
        RECT 74.355 131.535 74.735 131.705 ;
        RECT 74.905 131.195 75.205 131.705 ;
        RECT 78.800 131.630 79.150 132.880 ;
        RECT 80.915 132.455 81.665 132.975 ;
        RECT 83.725 132.835 83.940 133.530 ;
        RECT 84.130 133.005 84.480 133.530 ;
        RECT 84.650 133.005 85.345 133.575 ;
        RECT 84.275 132.835 84.480 133.005 ;
        RECT 81.835 132.285 82.585 132.805 ;
        RECT 83.240 132.505 83.525 132.835 ;
        RECT 83.725 132.505 84.105 132.835 ;
        RECT 84.275 132.505 84.585 132.835 ;
        RECT 84.755 132.335 84.925 133.005 ;
        RECT 85.515 132.975 88.105 133.745 ;
        RECT 75.395 131.195 80.740 131.630 ;
        RECT 80.915 131.195 82.585 132.285 ;
        RECT 83.215 131.195 83.475 132.335 ;
        RECT 83.645 132.165 84.925 132.335 ;
        RECT 85.105 132.165 85.345 132.835 ;
        RECT 85.515 132.455 86.725 132.975 ;
        RECT 88.295 132.935 88.535 133.745 ;
        RECT 88.705 132.935 89.035 133.575 ;
        RECT 89.205 132.935 89.475 133.745 ;
        RECT 89.655 133.200 95.000 133.745 ;
        RECT 86.895 132.285 88.105 132.805 ;
        RECT 88.275 132.505 88.625 132.755 ;
        RECT 88.795 132.335 88.965 132.935 ;
        RECT 89.135 132.505 89.485 132.755 ;
        RECT 91.240 132.370 91.580 133.200 ;
        RECT 95.175 132.995 96.385 133.745 ;
        RECT 96.555 133.020 96.845 133.745 ;
        RECT 83.645 131.365 83.975 132.165 ;
        RECT 84.145 131.195 84.315 131.995 ;
        RECT 84.515 131.365 84.845 132.165 ;
        RECT 85.045 131.195 85.325 131.995 ;
        RECT 85.515 131.195 88.105 132.285 ;
        RECT 88.285 132.165 88.965 132.335 ;
        RECT 88.285 131.380 88.615 132.165 ;
        RECT 89.145 131.195 89.475 132.335 ;
        RECT 93.060 131.630 93.410 132.880 ;
        RECT 95.175 132.455 95.695 132.995 ;
        RECT 95.865 132.285 96.385 132.825 ;
        RECT 97.015 132.800 97.355 133.575 ;
        RECT 97.525 133.285 97.695 133.745 ;
        RECT 97.935 133.310 98.295 133.575 ;
        RECT 97.935 133.305 98.290 133.310 ;
        RECT 97.935 133.295 98.285 133.305 ;
        RECT 97.935 133.290 98.280 133.295 ;
        RECT 97.935 133.280 98.275 133.290 ;
        RECT 98.925 133.285 99.095 133.745 ;
        RECT 97.935 133.275 98.270 133.280 ;
        RECT 97.935 133.265 98.260 133.275 ;
        RECT 97.935 133.255 98.250 133.265 ;
        RECT 97.935 133.115 98.235 133.255 ;
        RECT 97.525 132.925 98.235 133.115 ;
        RECT 98.425 133.115 98.755 133.195 ;
        RECT 99.265 133.115 99.605 133.575 ;
        RECT 98.425 132.925 99.605 133.115 ;
        RECT 99.775 133.070 100.035 133.575 ;
        RECT 100.215 133.365 100.545 133.745 ;
        RECT 100.725 133.195 100.895 133.575 ;
        RECT 89.655 131.195 95.000 131.630 ;
        RECT 95.175 131.195 96.385 132.285 ;
        RECT 96.555 131.195 96.845 132.360 ;
        RECT 97.015 131.365 97.295 132.800 ;
        RECT 97.525 132.355 97.810 132.925 ;
        RECT 97.995 132.525 98.465 132.755 ;
        RECT 98.635 132.735 98.965 132.755 ;
        RECT 98.635 132.555 99.085 132.735 ;
        RECT 99.275 132.555 99.605 132.755 ;
        RECT 97.525 132.140 98.675 132.355 ;
        RECT 97.465 131.195 98.175 131.970 ;
        RECT 98.345 131.365 98.675 132.140 ;
        RECT 98.870 131.440 99.085 132.555 ;
        RECT 99.375 132.215 99.605 132.555 ;
        RECT 99.775 132.270 99.955 133.070 ;
        RECT 100.230 133.025 100.895 133.195 ;
        RECT 100.230 132.770 100.400 133.025 ;
        RECT 101.155 132.975 103.745 133.745 ;
        RECT 104.410 133.005 105.025 133.575 ;
        RECT 105.195 133.235 105.410 133.745 ;
        RECT 105.640 133.235 105.920 133.565 ;
        RECT 106.100 133.235 106.340 133.745 ;
        RECT 100.125 132.440 100.400 132.770 ;
        RECT 100.625 132.475 100.965 132.845 ;
        RECT 101.155 132.455 102.365 132.975 ;
        RECT 100.230 132.295 100.400 132.440 ;
        RECT 99.265 131.195 99.595 131.915 ;
        RECT 99.775 131.365 100.045 132.270 ;
        RECT 100.230 132.125 100.905 132.295 ;
        RECT 102.535 132.285 103.745 132.805 ;
        RECT 100.215 131.195 100.545 131.955 ;
        RECT 100.725 131.365 100.905 132.125 ;
        RECT 101.155 131.195 103.745 132.285 ;
        RECT 104.410 131.985 104.725 133.005 ;
        RECT 104.895 132.335 105.065 132.835 ;
        RECT 105.315 132.505 105.580 133.065 ;
        RECT 105.750 132.335 105.920 133.235 ;
        RECT 106.675 133.200 112.020 133.745 ;
        RECT 106.090 132.505 106.445 133.065 ;
        RECT 108.260 132.370 108.600 133.200 ;
        RECT 104.895 132.165 106.320 132.335 ;
        RECT 104.410 131.365 104.945 131.985 ;
        RECT 105.115 131.195 105.445 131.995 ;
        RECT 105.930 131.990 106.320 132.165 ;
        RECT 110.080 131.630 110.430 132.880 ;
        RECT 112.200 132.145 112.535 133.565 ;
        RECT 112.715 133.375 113.460 133.745 ;
        RECT 114.025 133.205 114.280 133.565 ;
        RECT 114.460 133.375 114.790 133.745 ;
        RECT 114.970 133.205 115.195 133.565 ;
        RECT 112.710 133.015 115.195 133.205 ;
        RECT 115.415 133.200 120.760 133.745 ;
        RECT 112.710 132.325 112.935 133.015 ;
        RECT 113.135 132.505 113.415 132.835 ;
        RECT 113.595 132.505 114.170 132.835 ;
        RECT 114.350 132.505 114.785 132.835 ;
        RECT 114.965 132.505 115.235 132.835 ;
        RECT 117.000 132.370 117.340 133.200 ;
        RECT 120.935 132.995 122.145 133.745 ;
        RECT 122.315 133.020 122.605 133.745 ;
        RECT 122.775 133.245 123.035 133.575 ;
        RECT 123.245 133.265 123.520 133.745 ;
        RECT 112.710 132.145 115.205 132.325 ;
        RECT 106.675 131.195 112.020 131.630 ;
        RECT 112.200 131.375 112.465 132.145 ;
        RECT 112.635 131.195 112.965 131.915 ;
        RECT 113.155 131.735 114.345 131.965 ;
        RECT 113.155 131.375 113.415 131.735 ;
        RECT 113.585 131.195 113.915 131.565 ;
        RECT 114.085 131.375 114.345 131.735 ;
        RECT 114.915 131.375 115.205 132.145 ;
        RECT 118.820 131.630 119.170 132.880 ;
        RECT 120.935 132.455 121.455 132.995 ;
        RECT 121.625 132.285 122.145 132.825 ;
        RECT 115.415 131.195 120.760 131.630 ;
        RECT 120.935 131.195 122.145 132.285 ;
        RECT 122.315 131.195 122.605 132.360 ;
        RECT 122.775 132.335 122.945 133.245 ;
        RECT 123.730 133.175 123.935 133.575 ;
        RECT 124.105 133.345 124.440 133.745 ;
        RECT 124.705 133.195 124.875 133.575 ;
        RECT 125.055 133.365 125.385 133.745 ;
        RECT 123.115 132.505 123.475 133.085 ;
        RECT 123.730 133.005 124.415 133.175 ;
        RECT 124.705 133.025 125.370 133.195 ;
        RECT 125.565 133.070 125.825 133.575 ;
        RECT 123.655 132.335 123.905 132.835 ;
        RECT 122.775 132.165 123.905 132.335 ;
        RECT 122.775 131.395 123.045 132.165 ;
        RECT 124.075 131.975 124.415 133.005 ;
        RECT 124.635 132.475 124.975 132.845 ;
        RECT 125.200 132.770 125.370 133.025 ;
        RECT 125.200 132.440 125.475 132.770 ;
        RECT 125.200 132.295 125.370 132.440 ;
        RECT 123.215 131.195 123.545 131.975 ;
        RECT 123.750 131.800 124.415 131.975 ;
        RECT 124.695 132.125 125.370 132.295 ;
        RECT 125.645 132.270 125.825 133.070 ;
        RECT 125.995 132.975 128.585 133.745 ;
        RECT 129.215 133.070 129.475 133.575 ;
        RECT 129.655 133.365 129.985 133.745 ;
        RECT 130.165 133.195 130.335 133.575 ;
        RECT 125.995 132.455 127.205 132.975 ;
        RECT 127.375 132.285 128.585 132.805 ;
        RECT 123.750 131.395 123.935 131.800 ;
        RECT 124.105 131.195 124.440 131.620 ;
        RECT 124.695 131.365 124.875 132.125 ;
        RECT 125.055 131.195 125.385 131.955 ;
        RECT 125.555 131.365 125.825 132.270 ;
        RECT 125.995 131.195 128.585 132.285 ;
        RECT 129.215 132.270 129.395 133.070 ;
        RECT 129.670 133.025 130.335 133.195 ;
        RECT 130.685 133.195 130.855 133.575 ;
        RECT 131.035 133.365 131.365 133.745 ;
        RECT 130.685 133.025 131.350 133.195 ;
        RECT 131.545 133.070 131.805 133.575 ;
        RECT 129.670 132.770 129.840 133.025 ;
        RECT 129.565 132.440 129.840 132.770 ;
        RECT 130.065 132.475 130.405 132.845 ;
        RECT 130.615 132.475 130.945 132.845 ;
        RECT 131.180 132.770 131.350 133.025 ;
        RECT 129.670 132.295 129.840 132.440 ;
        RECT 131.180 132.440 131.465 132.770 ;
        RECT 131.180 132.295 131.350 132.440 ;
        RECT 129.215 131.365 129.485 132.270 ;
        RECT 129.670 132.125 130.345 132.295 ;
        RECT 129.655 131.195 129.985 131.955 ;
        RECT 130.165 131.365 130.345 132.125 ;
        RECT 130.685 132.125 131.350 132.295 ;
        RECT 131.635 132.270 131.805 133.070 ;
        RECT 132.065 133.195 132.235 133.575 ;
        RECT 132.415 133.365 132.745 133.745 ;
        RECT 132.065 133.025 132.730 133.195 ;
        RECT 132.925 133.070 133.185 133.575 ;
        RECT 131.995 132.475 132.335 132.845 ;
        RECT 132.560 132.770 132.730 133.025 ;
        RECT 132.560 132.440 132.835 132.770 ;
        RECT 132.560 132.295 132.730 132.440 ;
        RECT 130.685 131.365 130.855 132.125 ;
        RECT 131.035 131.195 131.365 131.955 ;
        RECT 131.535 131.365 131.805 132.270 ;
        RECT 132.055 132.125 132.730 132.295 ;
        RECT 133.005 132.270 133.185 133.070 ;
        RECT 133.355 132.975 136.865 133.745 ;
        RECT 137.035 132.995 138.245 133.745 ;
        RECT 138.425 133.020 138.755 133.530 ;
        RECT 138.925 133.345 139.255 133.745 ;
        RECT 140.305 133.175 140.635 133.515 ;
        RECT 140.805 133.345 141.135 133.745 ;
        RECT 133.355 132.455 135.005 132.975 ;
        RECT 135.175 132.285 136.865 132.805 ;
        RECT 137.035 132.455 137.555 132.995 ;
        RECT 137.725 132.285 138.245 132.825 ;
        RECT 132.055 131.365 132.235 132.125 ;
        RECT 132.415 131.195 132.745 131.955 ;
        RECT 132.915 131.365 133.185 132.270 ;
        RECT 133.355 131.195 136.865 132.285 ;
        RECT 137.035 131.195 138.245 132.285 ;
        RECT 138.425 132.255 138.615 133.020 ;
        RECT 138.925 133.005 141.290 133.175 ;
        RECT 138.925 132.835 139.095 133.005 ;
        RECT 138.785 132.505 139.095 132.835 ;
        RECT 139.265 132.505 139.570 132.835 ;
        RECT 138.425 131.405 138.755 132.255 ;
        RECT 138.925 131.195 139.175 132.335 ;
        RECT 139.355 132.175 139.570 132.505 ;
        RECT 139.745 132.175 140.030 132.835 ;
        RECT 140.225 132.175 140.490 132.835 ;
        RECT 140.705 132.175 140.950 132.835 ;
        RECT 141.120 132.005 141.290 133.005 ;
        RECT 141.635 132.945 142.330 133.575 ;
        RECT 142.535 132.945 142.845 133.745 ;
        RECT 141.655 132.505 141.990 132.755 ;
        RECT 142.160 132.385 142.330 132.945 ;
        RECT 143.485 132.935 143.755 133.745 ;
        RECT 143.925 132.935 144.255 133.575 ;
        RECT 144.425 132.935 144.665 133.745 ;
        RECT 144.875 132.935 145.115 133.745 ;
        RECT 145.285 132.935 145.615 133.575 ;
        RECT 145.785 132.935 146.055 133.745 ;
        RECT 146.325 133.195 146.495 133.575 ;
        RECT 146.710 133.365 147.040 133.745 ;
        RECT 146.325 133.025 147.040 133.195 ;
        RECT 142.500 132.505 142.835 132.775 ;
        RECT 143.475 132.505 143.825 132.755 ;
        RECT 142.155 132.345 142.330 132.385 ;
        RECT 139.365 131.835 140.655 132.005 ;
        RECT 139.365 131.415 139.615 131.835 ;
        RECT 139.845 131.195 140.175 131.665 ;
        RECT 140.405 131.415 140.655 131.835 ;
        RECT 140.835 131.835 141.290 132.005 ;
        RECT 140.835 131.405 141.165 131.835 ;
        RECT 141.635 131.195 141.895 132.335 ;
        RECT 142.065 131.365 142.395 132.345 ;
        RECT 143.995 132.335 144.165 132.935 ;
        RECT 144.335 132.505 144.685 132.755 ;
        RECT 144.855 132.505 145.205 132.755 ;
        RECT 145.375 132.335 145.545 132.935 ;
        RECT 145.715 132.505 146.065 132.755 ;
        RECT 146.235 132.475 146.590 132.845 ;
        RECT 146.870 132.835 147.040 133.025 ;
        RECT 147.210 133.000 147.465 133.575 ;
        RECT 146.870 132.505 147.125 132.835 ;
        RECT 142.565 131.195 142.845 132.335 ;
        RECT 143.485 131.195 143.815 132.335 ;
        RECT 143.995 132.165 144.675 132.335 ;
        RECT 144.345 131.380 144.675 132.165 ;
        RECT 144.865 132.165 145.545 132.335 ;
        RECT 144.865 131.380 145.195 132.165 ;
        RECT 145.725 131.195 146.055 132.335 ;
        RECT 146.870 132.295 147.040 132.505 ;
        RECT 146.325 132.125 147.040 132.295 ;
        RECT 147.295 132.270 147.465 133.000 ;
        RECT 147.640 132.905 147.900 133.745 ;
        RECT 148.075 133.020 148.365 133.745 ;
        RECT 148.535 133.365 149.425 133.535 ;
        RECT 148.535 132.810 149.085 133.195 ;
        RECT 149.255 132.640 149.425 133.365 ;
        RECT 148.535 132.570 149.425 132.640 ;
        RECT 149.595 133.040 149.815 133.525 ;
        RECT 149.985 133.205 150.235 133.745 ;
        RECT 150.405 133.095 150.665 133.575 ;
        RECT 149.595 132.615 149.925 133.040 ;
        RECT 148.535 132.545 149.430 132.570 ;
        RECT 148.535 132.530 149.440 132.545 ;
        RECT 148.535 132.515 149.445 132.530 ;
        RECT 148.535 132.510 149.455 132.515 ;
        RECT 148.535 132.500 149.460 132.510 ;
        RECT 148.535 132.490 149.465 132.500 ;
        RECT 148.535 132.485 149.475 132.490 ;
        RECT 148.535 132.475 149.485 132.485 ;
        RECT 148.535 132.470 149.495 132.475 ;
        RECT 146.325 131.365 146.495 132.125 ;
        RECT 146.710 131.195 147.040 131.955 ;
        RECT 147.210 131.365 147.465 132.270 ;
        RECT 147.640 131.195 147.900 132.345 ;
        RECT 148.075 131.195 148.365 132.360 ;
        RECT 148.535 132.020 148.795 132.470 ;
        RECT 149.160 132.465 149.495 132.470 ;
        RECT 149.160 132.460 149.510 132.465 ;
        RECT 149.160 132.450 149.525 132.460 ;
        RECT 149.160 132.445 149.550 132.450 ;
        RECT 150.095 132.445 150.325 132.840 ;
        RECT 149.160 132.440 150.325 132.445 ;
        RECT 149.190 132.405 150.325 132.440 ;
        RECT 149.225 132.380 150.325 132.405 ;
        RECT 149.255 132.350 150.325 132.380 ;
        RECT 149.275 132.320 150.325 132.350 ;
        RECT 149.295 132.290 150.325 132.320 ;
        RECT 149.365 132.280 150.325 132.290 ;
        RECT 149.390 132.270 150.325 132.280 ;
        RECT 149.410 132.255 150.325 132.270 ;
        RECT 149.430 132.240 150.325 132.255 ;
        RECT 149.435 132.230 150.220 132.240 ;
        RECT 149.450 132.195 150.220 132.230 ;
        RECT 148.965 131.875 149.295 132.120 ;
        RECT 149.465 131.945 150.220 132.195 ;
        RECT 150.495 132.065 150.665 133.095 ;
        RECT 148.965 131.850 149.150 131.875 ;
        RECT 148.535 131.750 149.150 131.850 ;
        RECT 148.535 131.195 149.140 131.750 ;
        RECT 149.315 131.365 149.795 131.705 ;
        RECT 149.965 131.195 150.220 131.740 ;
        RECT 150.390 131.365 150.665 132.065 ;
        RECT 151.330 133.005 151.945 133.575 ;
        RECT 152.115 133.235 152.330 133.745 ;
        RECT 152.560 133.235 152.840 133.565 ;
        RECT 153.020 133.235 153.260 133.745 ;
        RECT 151.330 131.985 151.645 133.005 ;
        RECT 151.815 132.335 151.985 132.835 ;
        RECT 152.235 132.505 152.500 133.065 ;
        RECT 152.670 132.335 152.840 133.235 ;
        RECT 153.010 132.505 153.365 133.065 ;
        RECT 153.595 132.945 154.290 133.575 ;
        RECT 154.495 132.945 154.805 133.745 ;
        RECT 154.975 132.995 156.185 133.745 ;
        RECT 153.615 132.505 153.950 132.755 ;
        RECT 154.120 132.345 154.290 132.945 ;
        RECT 154.460 132.505 154.795 132.775 ;
        RECT 151.815 132.165 153.240 132.335 ;
        RECT 151.330 131.365 151.865 131.985 ;
        RECT 152.035 131.195 152.365 131.995 ;
        RECT 152.850 131.990 153.240 132.165 ;
        RECT 153.595 131.195 153.855 132.335 ;
        RECT 154.025 131.365 154.355 132.345 ;
        RECT 154.525 131.195 154.805 132.335 ;
        RECT 154.975 132.285 155.495 132.825 ;
        RECT 155.665 132.455 156.185 132.995 ;
        RECT 154.975 131.195 156.185 132.285 ;
        RECT 70.710 131.025 156.270 131.195 ;
        RECT 70.795 129.935 72.005 131.025 ;
        RECT 72.175 129.935 73.845 131.025 ;
        RECT 74.015 130.515 74.315 131.025 ;
        RECT 74.485 130.345 74.815 130.855 ;
        RECT 74.985 130.515 75.615 131.025 ;
        RECT 76.195 130.515 76.575 130.685 ;
        RECT 76.745 130.515 77.045 131.025 ;
        RECT 76.405 130.345 76.575 130.515 ;
        RECT 70.795 129.225 71.315 129.765 ;
        RECT 71.485 129.395 72.005 129.935 ;
        RECT 72.175 129.245 72.925 129.765 ;
        RECT 73.095 129.415 73.845 129.935 ;
        RECT 74.015 130.175 76.235 130.345 ;
        RECT 70.795 128.475 72.005 129.225 ;
        RECT 72.175 128.475 73.845 129.245 ;
        RECT 74.015 129.215 74.185 130.175 ;
        RECT 74.355 129.835 75.895 130.005 ;
        RECT 74.355 129.385 74.600 129.835 ;
        RECT 74.860 129.465 75.555 129.665 ;
        RECT 75.725 129.635 75.895 129.835 ;
        RECT 76.065 129.975 76.235 130.175 ;
        RECT 76.405 130.145 77.065 130.345 ;
        RECT 76.065 129.805 76.725 129.975 ;
        RECT 75.725 129.465 76.325 129.635 ;
        RECT 76.555 129.385 76.725 129.805 ;
        RECT 74.015 128.670 74.480 129.215 ;
        RECT 74.985 128.475 75.155 129.295 ;
        RECT 75.325 129.215 76.235 129.295 ;
        RECT 76.895 129.215 77.065 130.145 ;
        RECT 77.695 129.885 77.975 131.025 ;
        RECT 78.145 129.875 78.475 130.855 ;
        RECT 78.645 129.885 78.905 131.025 ;
        RECT 79.095 130.135 79.355 130.845 ;
        RECT 79.525 130.315 79.855 131.025 ;
        RECT 80.025 130.135 80.255 130.845 ;
        RECT 79.095 129.895 80.255 130.135 ;
        RECT 80.435 130.115 80.705 130.845 ;
        RECT 80.885 130.295 81.225 131.025 ;
        RECT 80.435 129.895 81.205 130.115 ;
        RECT 77.705 129.445 78.040 129.715 ;
        RECT 78.210 129.275 78.380 129.875 ;
        RECT 78.550 129.465 78.885 129.715 ;
        RECT 79.085 129.385 79.385 129.715 ;
        RECT 79.565 129.405 80.090 129.715 ;
        RECT 80.270 129.405 80.735 129.715 ;
        RECT 75.325 129.125 76.575 129.215 ;
        RECT 75.325 128.645 75.655 129.125 ;
        RECT 76.065 129.045 76.575 129.125 ;
        RECT 75.825 128.475 76.175 128.865 ;
        RECT 76.345 128.645 76.575 129.045 ;
        RECT 76.745 128.735 77.065 129.215 ;
        RECT 77.695 128.475 78.005 129.275 ;
        RECT 78.210 128.645 78.905 129.275 ;
        RECT 79.095 128.475 79.385 129.205 ;
        RECT 79.565 128.765 79.795 129.405 ;
        RECT 80.915 129.225 81.205 129.895 ;
        RECT 79.975 129.025 81.205 129.225 ;
        RECT 79.975 128.655 80.285 129.025 ;
        RECT 80.465 128.475 81.135 128.845 ;
        RECT 81.395 128.655 81.655 130.845 ;
        RECT 81.835 129.885 82.115 131.025 ;
        RECT 82.285 129.875 82.615 130.855 ;
        RECT 82.785 129.885 83.045 131.025 ;
        RECT 81.845 129.445 82.180 129.715 ;
        RECT 82.350 129.275 82.520 129.875 ;
        RECT 83.675 129.860 83.965 131.025 ;
        RECT 84.135 130.470 84.740 131.025 ;
        RECT 84.915 130.515 85.395 130.855 ;
        RECT 85.565 130.480 85.820 131.025 ;
        RECT 84.135 130.370 84.750 130.470 ;
        RECT 84.565 130.345 84.750 130.370 ;
        RECT 84.135 129.750 84.395 130.200 ;
        RECT 84.565 130.100 84.895 130.345 ;
        RECT 85.065 130.025 85.820 130.275 ;
        RECT 85.990 130.155 86.265 130.855 ;
        RECT 85.050 129.990 85.820 130.025 ;
        RECT 85.035 129.980 85.820 129.990 ;
        RECT 85.030 129.965 85.925 129.980 ;
        RECT 85.010 129.950 85.925 129.965 ;
        RECT 84.990 129.940 85.925 129.950 ;
        RECT 84.965 129.930 85.925 129.940 ;
        RECT 84.895 129.900 85.925 129.930 ;
        RECT 84.875 129.870 85.925 129.900 ;
        RECT 84.855 129.840 85.925 129.870 ;
        RECT 84.825 129.815 85.925 129.840 ;
        RECT 84.790 129.780 85.925 129.815 ;
        RECT 84.760 129.775 85.925 129.780 ;
        RECT 84.760 129.770 85.150 129.775 ;
        RECT 84.760 129.760 85.125 129.770 ;
        RECT 84.760 129.755 85.110 129.760 ;
        RECT 84.760 129.750 85.095 129.755 ;
        RECT 84.135 129.745 85.095 129.750 ;
        RECT 84.135 129.735 85.085 129.745 ;
        RECT 84.135 129.730 85.075 129.735 ;
        RECT 84.135 129.720 85.065 129.730 ;
        RECT 82.690 129.465 83.025 129.715 ;
        RECT 84.135 129.710 85.060 129.720 ;
        RECT 84.135 129.705 85.055 129.710 ;
        RECT 84.135 129.690 85.045 129.705 ;
        RECT 84.135 129.675 85.040 129.690 ;
        RECT 84.135 129.650 85.030 129.675 ;
        RECT 84.135 129.580 85.025 129.650 ;
        RECT 81.835 128.475 82.145 129.275 ;
        RECT 82.350 128.645 83.045 129.275 ;
        RECT 83.675 128.475 83.965 129.200 ;
        RECT 84.135 129.025 84.685 129.410 ;
        RECT 84.855 128.855 85.025 129.580 ;
        RECT 84.135 128.685 85.025 128.855 ;
        RECT 85.195 129.180 85.525 129.605 ;
        RECT 85.695 129.380 85.925 129.775 ;
        RECT 85.195 128.695 85.415 129.180 ;
        RECT 86.095 129.125 86.265 130.155 ;
        RECT 86.475 130.075 86.765 130.845 ;
        RECT 87.335 130.485 87.595 130.845 ;
        RECT 87.765 130.655 88.095 131.025 ;
        RECT 88.265 130.485 88.525 130.845 ;
        RECT 87.335 130.255 88.525 130.485 ;
        RECT 88.715 130.305 89.045 131.025 ;
        RECT 89.215 130.075 89.480 130.845 ;
        RECT 89.660 130.645 89.995 131.025 ;
        RECT 86.475 129.895 88.970 130.075 ;
        RECT 86.445 129.385 86.715 129.715 ;
        RECT 86.895 129.385 87.330 129.715 ;
        RECT 87.510 129.385 88.085 129.715 ;
        RECT 88.265 129.385 88.545 129.715 ;
        RECT 88.745 129.205 88.970 129.895 ;
        RECT 85.585 128.475 85.835 129.015 ;
        RECT 86.005 128.645 86.265 129.125 ;
        RECT 86.485 129.015 88.970 129.205 ;
        RECT 86.485 128.655 86.710 129.015 ;
        RECT 86.890 128.475 87.220 128.845 ;
        RECT 87.400 128.655 87.655 129.015 ;
        RECT 88.220 128.475 88.965 128.845 ;
        RECT 89.145 128.655 89.480 130.075 ;
        RECT 89.655 129.155 89.895 130.465 ;
        RECT 90.165 130.055 90.415 130.855 ;
        RECT 90.635 130.305 90.965 131.025 ;
        RECT 91.150 130.055 91.400 130.855 ;
        RECT 91.865 130.225 92.195 131.025 ;
        RECT 92.365 130.595 92.705 130.855 ;
        RECT 90.065 129.885 92.255 130.055 ;
        RECT 90.065 128.975 90.235 129.885 ;
        RECT 91.940 129.715 92.255 129.885 ;
        RECT 89.740 128.645 90.235 128.975 ;
        RECT 90.455 128.750 90.805 129.715 ;
        RECT 90.985 128.745 91.285 129.715 ;
        RECT 91.465 128.745 91.745 129.715 ;
        RECT 91.940 129.465 92.270 129.715 ;
        RECT 91.925 128.475 92.195 129.275 ;
        RECT 92.445 129.195 92.705 130.595 ;
        RECT 92.365 128.685 92.705 129.195 ;
        RECT 92.875 130.225 93.315 130.855 ;
        RECT 92.875 129.215 93.185 130.225 ;
        RECT 93.490 130.175 93.805 131.025 ;
        RECT 93.975 130.685 95.405 130.855 ;
        RECT 93.975 130.005 94.145 130.685 ;
        RECT 93.355 129.835 94.145 130.005 ;
        RECT 93.355 129.385 93.525 129.835 ;
        RECT 94.315 129.715 94.515 130.515 ;
        RECT 93.695 129.385 94.085 129.665 ;
        RECT 94.270 129.385 94.515 129.715 ;
        RECT 94.715 129.385 94.965 130.515 ;
        RECT 95.155 130.055 95.405 130.685 ;
        RECT 95.585 130.225 95.915 131.025 ;
        RECT 95.155 129.885 95.925 130.055 ;
        RECT 96.095 129.935 97.765 131.025 ;
        RECT 95.180 129.385 95.585 129.715 ;
        RECT 95.755 129.215 95.925 129.885 ;
        RECT 92.875 128.655 93.315 129.215 ;
        RECT 93.485 128.475 93.935 129.215 ;
        RECT 94.105 129.045 95.265 129.215 ;
        RECT 94.105 128.645 94.275 129.045 ;
        RECT 94.445 128.475 94.865 128.875 ;
        RECT 95.035 128.645 95.265 129.045 ;
        RECT 95.435 128.645 95.925 129.215 ;
        RECT 96.095 129.245 96.845 129.765 ;
        RECT 97.015 129.415 97.765 129.935 ;
        RECT 98.395 130.225 98.835 130.855 ;
        RECT 96.095 128.475 97.765 129.245 ;
        RECT 98.395 129.215 98.705 130.225 ;
        RECT 99.010 130.175 99.325 131.025 ;
        RECT 99.495 130.685 100.925 130.855 ;
        RECT 99.495 130.005 99.665 130.685 ;
        RECT 98.875 129.835 99.665 130.005 ;
        RECT 98.875 129.385 99.045 129.835 ;
        RECT 99.835 129.715 100.035 130.515 ;
        RECT 99.215 129.385 99.605 129.665 ;
        RECT 99.790 129.385 100.035 129.715 ;
        RECT 100.235 129.385 100.485 130.515 ;
        RECT 100.675 130.055 100.925 130.685 ;
        RECT 101.105 130.225 101.435 131.025 ;
        RECT 101.915 130.385 102.245 130.815 ;
        RECT 101.790 130.215 102.245 130.385 ;
        RECT 102.425 130.385 102.675 130.805 ;
        RECT 102.905 130.555 103.235 131.025 ;
        RECT 103.465 130.385 103.715 130.805 ;
        RECT 102.425 130.215 103.715 130.385 ;
        RECT 100.675 129.885 101.445 130.055 ;
        RECT 100.700 129.385 101.105 129.715 ;
        RECT 101.275 129.215 101.445 129.885 ;
        RECT 98.395 128.655 98.835 129.215 ;
        RECT 99.005 128.475 99.455 129.215 ;
        RECT 99.625 129.045 100.785 129.215 ;
        RECT 99.625 128.645 99.795 129.045 ;
        RECT 99.965 128.475 100.385 128.875 ;
        RECT 100.555 128.645 100.785 129.045 ;
        RECT 100.955 128.645 101.445 129.215 ;
        RECT 101.790 129.215 101.960 130.215 ;
        RECT 102.130 129.385 102.375 130.045 ;
        RECT 102.590 129.385 102.855 130.045 ;
        RECT 103.050 129.385 103.335 130.045 ;
        RECT 103.510 129.715 103.725 130.045 ;
        RECT 103.905 129.885 104.155 131.025 ;
        RECT 104.325 129.965 104.655 130.815 ;
        RECT 104.835 130.430 105.270 130.855 ;
        RECT 105.440 130.600 105.825 131.025 ;
        RECT 104.835 130.260 105.825 130.430 ;
        RECT 103.510 129.385 103.815 129.715 ;
        RECT 103.985 129.385 104.295 129.715 ;
        RECT 103.985 129.215 104.155 129.385 ;
        RECT 101.790 129.045 104.155 129.215 ;
        RECT 104.465 129.200 104.655 129.965 ;
        RECT 104.835 129.385 105.320 130.090 ;
        RECT 105.490 129.715 105.825 130.260 ;
        RECT 105.995 130.065 106.420 130.855 ;
        RECT 106.590 130.430 106.865 130.855 ;
        RECT 107.035 130.600 107.420 131.025 ;
        RECT 106.590 130.235 107.420 130.430 ;
        RECT 105.995 129.885 106.900 130.065 ;
        RECT 105.490 129.385 105.900 129.715 ;
        RECT 106.070 129.385 106.900 129.885 ;
        RECT 107.070 129.715 107.420 130.235 ;
        RECT 107.590 130.065 107.835 130.855 ;
        RECT 108.025 130.430 108.280 130.855 ;
        RECT 108.450 130.600 108.835 131.025 ;
        RECT 108.025 130.235 108.835 130.430 ;
        RECT 107.590 129.885 108.315 130.065 ;
        RECT 107.070 129.385 107.495 129.715 ;
        RECT 107.665 129.385 108.315 129.885 ;
        RECT 108.485 129.715 108.835 130.235 ;
        RECT 109.005 129.885 109.265 130.855 ;
        RECT 108.485 129.385 108.910 129.715 ;
        RECT 105.490 129.215 105.825 129.385 ;
        RECT 106.070 129.215 106.420 129.385 ;
        RECT 107.070 129.215 107.420 129.385 ;
        RECT 107.665 129.215 107.835 129.385 ;
        RECT 108.485 129.215 108.835 129.385 ;
        RECT 109.080 129.215 109.265 129.885 ;
        RECT 109.435 129.860 109.725 131.025 ;
        RECT 109.975 130.095 110.155 130.855 ;
        RECT 110.335 130.265 110.665 131.025 ;
        RECT 109.975 129.925 110.650 130.095 ;
        RECT 110.835 129.950 111.105 130.855 ;
        RECT 110.480 129.780 110.650 129.925 ;
        RECT 109.915 129.375 110.255 129.745 ;
        RECT 110.480 129.450 110.755 129.780 ;
        RECT 101.945 128.475 102.275 128.875 ;
        RECT 102.445 128.705 102.775 129.045 ;
        RECT 103.825 128.475 104.155 128.875 ;
        RECT 104.325 128.690 104.655 129.200 ;
        RECT 104.835 129.045 105.825 129.215 ;
        RECT 104.835 128.645 105.270 129.045 ;
        RECT 105.440 128.475 105.825 128.875 ;
        RECT 105.995 128.645 106.420 129.215 ;
        RECT 106.610 129.045 107.420 129.215 ;
        RECT 106.610 128.645 106.865 129.045 ;
        RECT 107.035 128.475 107.420 128.875 ;
        RECT 107.590 128.645 107.835 129.215 ;
        RECT 108.025 129.045 108.835 129.215 ;
        RECT 108.025 128.645 108.280 129.045 ;
        RECT 108.450 128.475 108.835 128.875 ;
        RECT 109.005 128.645 109.265 129.215 ;
        RECT 109.435 128.475 109.725 129.200 ;
        RECT 110.480 129.195 110.650 129.450 ;
        RECT 109.985 129.025 110.650 129.195 ;
        RECT 110.925 129.150 111.105 129.950 ;
        RECT 109.985 128.645 110.155 129.025 ;
        RECT 110.335 128.475 110.665 128.855 ;
        RECT 110.845 128.645 111.105 129.150 ;
        RECT 111.275 130.305 111.735 130.855 ;
        RECT 111.925 130.305 112.255 131.025 ;
        RECT 111.275 128.935 111.525 130.305 ;
        RECT 112.455 130.135 112.755 130.685 ;
        RECT 112.925 130.355 113.205 131.025 ;
        RECT 111.815 129.965 112.755 130.135 ;
        RECT 111.815 129.715 111.985 129.965 ;
        RECT 113.125 129.715 113.390 130.075 ;
        RECT 111.695 129.385 111.985 129.715 ;
        RECT 112.155 129.465 112.495 129.715 ;
        RECT 112.715 129.465 113.390 129.715 ;
        RECT 111.815 129.295 111.985 129.385 ;
        RECT 113.575 129.420 113.855 130.855 ;
        RECT 114.025 130.250 114.735 131.025 ;
        RECT 114.905 130.080 115.235 130.855 ;
        RECT 114.085 129.865 115.235 130.080 ;
        RECT 111.815 129.105 113.205 129.295 ;
        RECT 111.275 128.645 111.835 128.935 ;
        RECT 112.005 128.475 112.255 128.935 ;
        RECT 112.875 128.745 113.205 129.105 ;
        RECT 113.575 128.645 113.915 129.420 ;
        RECT 114.085 129.295 114.370 129.865 ;
        RECT 114.555 129.465 115.025 129.695 ;
        RECT 115.430 129.665 115.645 130.780 ;
        RECT 115.825 130.305 116.155 131.025 ;
        RECT 116.355 130.135 116.615 130.845 ;
        RECT 116.785 130.315 117.115 131.025 ;
        RECT 117.285 130.135 117.515 130.845 ;
        RECT 115.935 129.665 116.165 130.005 ;
        RECT 116.355 129.895 117.515 130.135 ;
        RECT 117.695 130.115 117.965 130.845 ;
        RECT 118.145 130.295 118.485 131.025 ;
        RECT 117.695 129.895 118.465 130.115 ;
        RECT 115.195 129.485 115.645 129.665 ;
        RECT 115.195 129.465 115.525 129.485 ;
        RECT 115.835 129.465 116.165 129.665 ;
        RECT 116.345 129.385 116.645 129.715 ;
        RECT 116.825 129.405 117.350 129.715 ;
        RECT 117.530 129.405 117.995 129.715 ;
        RECT 114.085 129.105 114.795 129.295 ;
        RECT 114.495 128.965 114.795 129.105 ;
        RECT 114.985 129.105 116.165 129.295 ;
        RECT 114.985 129.025 115.315 129.105 ;
        RECT 114.495 128.955 114.810 128.965 ;
        RECT 114.495 128.945 114.820 128.955 ;
        RECT 114.495 128.940 114.830 128.945 ;
        RECT 114.085 128.475 114.255 128.935 ;
        RECT 114.495 128.930 114.835 128.940 ;
        RECT 114.495 128.925 114.840 128.930 ;
        RECT 114.495 128.915 114.845 128.925 ;
        RECT 114.495 128.910 114.850 128.915 ;
        RECT 114.495 128.645 114.855 128.910 ;
        RECT 115.485 128.475 115.655 128.935 ;
        RECT 115.825 128.645 116.165 129.105 ;
        RECT 116.355 128.475 116.645 129.205 ;
        RECT 116.825 128.765 117.055 129.405 ;
        RECT 118.175 129.225 118.465 129.895 ;
        RECT 117.235 129.025 118.465 129.225 ;
        RECT 117.235 128.655 117.545 129.025 ;
        RECT 117.725 128.475 118.395 128.845 ;
        RECT 118.655 128.655 118.915 130.845 ;
        RECT 119.095 129.950 119.365 130.855 ;
        RECT 119.535 130.265 119.865 131.025 ;
        RECT 120.045 130.095 120.225 130.855 ;
        RECT 119.095 129.150 119.275 129.950 ;
        RECT 119.550 129.925 120.225 130.095 ;
        RECT 120.475 129.950 120.745 130.855 ;
        RECT 120.915 130.265 121.245 131.025 ;
        RECT 121.425 130.095 121.605 130.855 ;
        RECT 119.550 129.780 119.720 129.925 ;
        RECT 119.445 129.450 119.720 129.780 ;
        RECT 119.550 129.195 119.720 129.450 ;
        RECT 119.945 129.375 120.285 129.745 ;
        RECT 119.095 128.645 119.355 129.150 ;
        RECT 119.550 129.025 120.215 129.195 ;
        RECT 119.535 128.475 119.865 128.855 ;
        RECT 120.045 128.645 120.215 129.025 ;
        RECT 120.475 129.150 120.655 129.950 ;
        RECT 120.930 129.925 121.605 130.095 ;
        RECT 121.855 129.950 122.125 130.855 ;
        RECT 122.295 130.265 122.625 131.025 ;
        RECT 122.805 130.095 122.985 130.855 ;
        RECT 120.930 129.780 121.100 129.925 ;
        RECT 120.825 129.450 121.100 129.780 ;
        RECT 120.930 129.195 121.100 129.450 ;
        RECT 121.325 129.375 121.665 129.745 ;
        RECT 120.475 128.645 120.735 129.150 ;
        RECT 120.930 129.025 121.595 129.195 ;
        RECT 120.915 128.475 121.245 128.855 ;
        RECT 121.425 128.645 121.595 129.025 ;
        RECT 121.855 129.150 122.035 129.950 ;
        RECT 122.310 129.925 122.985 130.095 ;
        RECT 123.695 129.950 123.965 130.855 ;
        RECT 124.135 130.265 124.465 131.025 ;
        RECT 124.645 130.095 124.825 130.855 ;
        RECT 122.310 129.780 122.480 129.925 ;
        RECT 122.205 129.450 122.480 129.780 ;
        RECT 122.310 129.195 122.480 129.450 ;
        RECT 122.705 129.375 123.045 129.745 ;
        RECT 121.855 128.645 122.115 129.150 ;
        RECT 122.310 129.025 122.975 129.195 ;
        RECT 122.295 128.475 122.625 128.855 ;
        RECT 122.805 128.645 122.975 129.025 ;
        RECT 123.695 129.150 123.875 129.950 ;
        RECT 124.150 129.925 124.825 130.095 ;
        RECT 124.150 129.780 124.320 129.925 ;
        RECT 124.045 129.450 124.320 129.780 ;
        RECT 125.075 129.885 125.335 130.855 ;
        RECT 125.505 130.600 125.890 131.025 ;
        RECT 126.060 130.430 126.315 130.855 ;
        RECT 125.505 130.235 126.315 130.430 ;
        RECT 124.150 129.195 124.320 129.450 ;
        RECT 124.545 129.375 124.885 129.745 ;
        RECT 125.075 129.215 125.260 129.885 ;
        RECT 125.505 129.715 125.855 130.235 ;
        RECT 126.505 130.065 126.750 130.855 ;
        RECT 126.920 130.600 127.305 131.025 ;
        RECT 127.475 130.430 127.750 130.855 ;
        RECT 125.430 129.385 125.855 129.715 ;
        RECT 126.025 129.885 126.750 130.065 ;
        RECT 126.920 130.235 127.750 130.430 ;
        RECT 126.025 129.385 126.675 129.885 ;
        RECT 126.920 129.715 127.270 130.235 ;
        RECT 127.920 130.065 128.345 130.855 ;
        RECT 128.515 130.600 128.900 131.025 ;
        RECT 129.070 130.430 129.505 130.855 ;
        RECT 126.845 129.385 127.270 129.715 ;
        RECT 127.440 129.885 128.345 130.065 ;
        RECT 128.515 130.260 129.505 130.430 ;
        RECT 127.440 129.385 128.270 129.885 ;
        RECT 128.515 129.715 128.850 130.260 ;
        RECT 129.765 130.095 129.935 130.855 ;
        RECT 130.115 130.265 130.445 131.025 ;
        RECT 128.440 129.385 128.850 129.715 ;
        RECT 129.020 129.385 129.505 130.090 ;
        RECT 129.765 129.925 130.430 130.095 ;
        RECT 130.615 129.950 130.885 130.855 ;
        RECT 130.260 129.780 130.430 129.925 ;
        RECT 125.505 129.215 125.855 129.385 ;
        RECT 126.505 129.215 126.675 129.385 ;
        RECT 126.920 129.215 127.270 129.385 ;
        RECT 127.920 129.215 128.270 129.385 ;
        RECT 128.515 129.215 128.850 129.385 ;
        RECT 129.695 129.375 130.025 129.745 ;
        RECT 130.260 129.450 130.545 129.780 ;
        RECT 123.695 128.645 123.955 129.150 ;
        RECT 124.150 129.025 124.815 129.195 ;
        RECT 124.135 128.475 124.465 128.855 ;
        RECT 124.645 128.645 124.815 129.025 ;
        RECT 125.075 128.645 125.335 129.215 ;
        RECT 125.505 129.045 126.315 129.215 ;
        RECT 125.505 128.475 125.890 128.875 ;
        RECT 126.060 128.645 126.315 129.045 ;
        RECT 126.505 128.645 126.750 129.215 ;
        RECT 126.920 129.045 127.730 129.215 ;
        RECT 126.920 128.475 127.305 128.875 ;
        RECT 127.475 128.645 127.730 129.045 ;
        RECT 127.920 128.645 128.345 129.215 ;
        RECT 128.515 129.045 129.505 129.215 ;
        RECT 130.260 129.195 130.430 129.450 ;
        RECT 128.515 128.475 128.900 128.875 ;
        RECT 129.070 128.645 129.505 129.045 ;
        RECT 129.765 129.025 130.430 129.195 ;
        RECT 130.715 129.150 130.885 129.950 ;
        RECT 129.765 128.645 129.935 129.025 ;
        RECT 130.115 128.475 130.445 128.855 ;
        RECT 130.625 128.645 130.885 129.150 ;
        RECT 131.055 129.885 131.395 130.855 ;
        RECT 131.565 129.885 131.735 131.025 ;
        RECT 132.005 130.225 132.255 131.025 ;
        RECT 132.900 130.055 133.230 130.855 ;
        RECT 133.530 130.225 133.860 131.025 ;
        RECT 134.030 130.055 134.360 130.855 ;
        RECT 131.925 129.885 134.360 130.055 ;
        RECT 131.055 129.275 131.230 129.885 ;
        RECT 131.925 129.635 132.095 129.885 ;
        RECT 131.400 129.465 132.095 129.635 ;
        RECT 132.270 129.465 132.690 129.665 ;
        RECT 132.860 129.465 133.190 129.665 ;
        RECT 133.360 129.465 133.690 129.665 ;
        RECT 131.055 128.645 131.395 129.275 ;
        RECT 131.565 128.475 131.815 129.275 ;
        RECT 132.005 129.125 133.230 129.295 ;
        RECT 132.005 128.645 132.335 129.125 ;
        RECT 132.505 128.475 132.730 128.935 ;
        RECT 132.900 128.645 133.230 129.125 ;
        RECT 133.860 129.255 134.030 129.885 ;
        RECT 135.195 129.860 135.485 131.025 ;
        RECT 135.955 130.385 136.285 130.815 ;
        RECT 135.830 130.215 136.285 130.385 ;
        RECT 136.465 130.385 136.715 130.805 ;
        RECT 136.945 130.555 137.275 131.025 ;
        RECT 137.505 130.385 137.755 130.805 ;
        RECT 136.465 130.215 137.755 130.385 ;
        RECT 134.215 129.465 134.565 129.715 ;
        RECT 133.860 128.645 134.360 129.255 ;
        RECT 135.830 129.215 136.000 130.215 ;
        RECT 136.170 129.385 136.415 130.045 ;
        RECT 136.630 129.385 136.895 130.045 ;
        RECT 137.090 129.385 137.375 130.045 ;
        RECT 137.550 129.715 137.765 130.045 ;
        RECT 137.945 129.885 138.195 131.025 ;
        RECT 138.365 129.965 138.695 130.815 ;
        RECT 137.550 129.385 137.855 129.715 ;
        RECT 138.025 129.385 138.335 129.715 ;
        RECT 138.025 129.215 138.195 129.385 ;
        RECT 135.195 128.475 135.485 129.200 ;
        RECT 135.830 129.045 138.195 129.215 ;
        RECT 138.505 129.200 138.695 129.965 ;
        RECT 138.935 129.885 139.145 131.025 ;
        RECT 139.315 129.875 139.645 130.855 ;
        RECT 139.815 129.885 140.045 131.025 ;
        RECT 140.265 129.885 140.595 131.025 ;
        RECT 141.125 130.055 141.455 130.840 ;
        RECT 140.775 129.885 141.455 130.055 ;
        RECT 135.985 128.475 136.315 128.875 ;
        RECT 136.485 128.705 136.815 129.045 ;
        RECT 137.865 128.475 138.195 128.875 ;
        RECT 138.365 128.690 138.695 129.200 ;
        RECT 138.935 128.475 139.145 129.295 ;
        RECT 139.315 129.275 139.565 129.875 ;
        RECT 139.735 129.465 140.065 129.715 ;
        RECT 140.255 129.465 140.605 129.715 ;
        RECT 139.315 128.645 139.645 129.275 ;
        RECT 139.815 128.475 140.045 129.295 ;
        RECT 140.775 129.285 140.945 129.885 ;
        RECT 141.640 129.875 141.900 131.025 ;
        RECT 142.075 129.950 142.330 130.855 ;
        RECT 142.500 130.265 142.830 131.025 ;
        RECT 143.045 130.095 143.215 130.855 ;
        RECT 143.675 130.355 143.955 131.025 ;
        RECT 141.115 129.465 141.465 129.715 ;
        RECT 140.265 128.475 140.535 129.285 ;
        RECT 140.705 128.645 141.035 129.285 ;
        RECT 141.205 128.475 141.445 129.285 ;
        RECT 141.640 128.475 141.900 129.315 ;
        RECT 142.075 129.220 142.245 129.950 ;
        RECT 142.500 129.925 143.215 130.095 ;
        RECT 144.125 130.135 144.425 130.685 ;
        RECT 144.625 130.305 144.955 131.025 ;
        RECT 145.145 130.305 145.605 130.855 ;
        RECT 142.500 129.715 142.670 129.925 ;
        RECT 142.415 129.385 142.670 129.715 ;
        RECT 142.075 128.645 142.330 129.220 ;
        RECT 142.500 129.195 142.670 129.385 ;
        RECT 142.950 129.375 143.305 129.745 ;
        RECT 143.490 129.715 143.755 130.075 ;
        RECT 144.125 129.965 145.065 130.135 ;
        RECT 144.895 129.715 145.065 129.965 ;
        RECT 143.490 129.465 144.165 129.715 ;
        RECT 144.385 129.465 144.725 129.715 ;
        RECT 144.895 129.385 145.185 129.715 ;
        RECT 144.895 129.295 145.065 129.385 ;
        RECT 142.500 129.025 143.215 129.195 ;
        RECT 142.500 128.475 142.830 128.855 ;
        RECT 143.045 128.645 143.215 129.025 ;
        RECT 143.675 129.105 145.065 129.295 ;
        RECT 143.675 128.745 144.005 129.105 ;
        RECT 145.355 128.935 145.605 130.305 ;
        RECT 145.780 129.885 146.035 131.025 ;
        RECT 144.625 128.475 144.875 128.935 ;
        RECT 145.045 128.645 145.605 128.935 ;
        RECT 145.780 128.475 146.035 129.275 ;
        RECT 146.205 128.685 146.535 130.815 ;
        RECT 146.850 130.225 147.070 131.025 ;
        RECT 147.280 130.395 147.530 130.855 ;
        RECT 147.815 130.645 148.145 131.025 ;
        RECT 148.405 130.395 148.715 130.855 ;
        RECT 147.280 130.225 148.715 130.395 ;
        RECT 149.485 130.055 149.655 130.855 ;
        RECT 146.705 129.885 149.655 130.055 ;
        RECT 149.915 129.885 150.190 130.855 ;
        RECT 150.400 130.225 150.680 131.025 ;
        RECT 150.850 130.685 152.900 130.805 ;
        RECT 150.850 130.515 152.905 130.685 ;
        RECT 150.850 130.175 152.480 130.345 ;
        RECT 150.850 130.055 151.020 130.175 ;
        RECT 150.360 129.885 151.020 130.055 ;
        RECT 146.705 129.215 146.875 129.885 ;
        RECT 147.185 129.385 147.400 129.715 ;
        RECT 146.705 129.045 147.385 129.215 ;
        RECT 146.705 128.475 147.035 128.855 ;
        RECT 147.215 128.815 147.385 129.045 ;
        RECT 147.585 128.995 147.855 129.715 ;
        RECT 148.130 129.385 148.365 129.715 ;
        RECT 148.585 129.385 148.925 129.715 ;
        RECT 149.385 129.385 149.695 129.715 ;
        RECT 148.130 128.995 148.310 129.385 ;
        RECT 148.480 129.045 149.655 129.215 ;
        RECT 148.480 128.815 148.650 129.045 ;
        RECT 147.215 128.645 148.650 128.815 ;
        RECT 148.910 128.475 149.240 128.875 ;
        RECT 149.485 128.645 149.655 129.045 ;
        RECT 149.915 129.150 150.085 129.885 ;
        RECT 150.360 129.715 150.530 129.885 ;
        RECT 150.255 129.385 150.530 129.715 ;
        RECT 150.700 129.385 151.080 129.715 ;
        RECT 151.250 129.385 151.990 130.005 ;
        RECT 152.160 129.885 152.480 130.175 ;
        RECT 152.675 129.715 152.915 130.310 ;
        RECT 153.085 129.950 153.425 131.025 ;
        RECT 153.605 130.055 153.935 130.840 ;
        RECT 153.605 129.885 154.285 130.055 ;
        RECT 154.465 129.885 154.795 131.025 ;
        RECT 154.975 129.935 156.185 131.025 ;
        RECT 152.260 129.385 152.915 129.715 ;
        RECT 150.360 129.215 150.530 129.385 ;
        RECT 149.915 128.805 150.190 129.150 ;
        RECT 150.360 129.045 151.945 129.215 ;
        RECT 150.380 128.475 150.760 128.875 ;
        RECT 150.930 128.695 151.100 129.045 ;
        RECT 151.270 128.475 151.600 128.875 ;
        RECT 151.775 128.695 151.945 129.045 ;
        RECT 152.145 128.475 152.475 128.975 ;
        RECT 152.670 128.695 152.915 129.385 ;
        RECT 153.085 129.145 153.425 129.715 ;
        RECT 153.595 129.465 153.945 129.715 ;
        RECT 154.115 129.285 154.285 129.885 ;
        RECT 154.455 129.465 154.805 129.715 ;
        RECT 154.975 129.395 155.495 129.935 ;
        RECT 153.085 128.475 153.425 128.975 ;
        RECT 153.615 128.475 153.855 129.285 ;
        RECT 154.025 128.645 154.355 129.285 ;
        RECT 154.525 128.475 154.795 129.285 ;
        RECT 155.665 129.225 156.185 129.765 ;
        RECT 154.975 128.475 156.185 129.225 ;
        RECT 70.710 128.305 156.270 128.475 ;
        RECT 70.795 127.555 72.005 128.305 ;
        RECT 72.175 127.555 73.385 128.305 ;
        RECT 73.555 127.630 73.815 128.135 ;
        RECT 73.995 127.925 74.325 128.305 ;
        RECT 74.505 127.755 74.675 128.135 ;
        RECT 70.795 127.015 71.315 127.555 ;
        RECT 71.485 126.845 72.005 127.385 ;
        RECT 72.175 127.015 72.695 127.555 ;
        RECT 72.865 126.845 73.385 127.385 ;
        RECT 70.795 125.755 72.005 126.845 ;
        RECT 72.175 125.755 73.385 126.845 ;
        RECT 73.555 126.830 73.725 127.630 ;
        RECT 74.010 127.585 74.675 127.755 ;
        RECT 75.395 127.630 75.655 128.135 ;
        RECT 75.835 127.925 76.165 128.305 ;
        RECT 76.345 127.755 76.515 128.135 ;
        RECT 74.010 127.330 74.180 127.585 ;
        RECT 73.895 127.000 74.180 127.330 ;
        RECT 74.415 127.035 74.745 127.405 ;
        RECT 74.010 126.855 74.180 127.000 ;
        RECT 73.555 125.925 73.825 126.830 ;
        RECT 74.010 126.685 74.675 126.855 ;
        RECT 73.995 125.755 74.325 126.515 ;
        RECT 74.505 125.925 74.675 126.685 ;
        RECT 75.395 126.830 75.565 127.630 ;
        RECT 75.850 127.585 76.515 127.755 ;
        RECT 75.850 127.330 76.020 127.585 ;
        RECT 76.775 127.555 77.985 128.305 ;
        RECT 78.320 127.795 78.560 128.305 ;
        RECT 78.740 127.795 79.020 128.125 ;
        RECT 79.250 127.795 79.465 128.305 ;
        RECT 75.735 127.000 76.020 127.330 ;
        RECT 76.255 127.035 76.585 127.405 ;
        RECT 76.775 127.015 77.295 127.555 ;
        RECT 75.850 126.855 76.020 127.000 ;
        RECT 75.395 125.925 75.665 126.830 ;
        RECT 75.850 126.685 76.515 126.855 ;
        RECT 77.465 126.845 77.985 127.385 ;
        RECT 78.215 127.065 78.570 127.625 ;
        RECT 78.740 126.895 78.910 127.795 ;
        RECT 79.080 127.065 79.345 127.625 ;
        RECT 79.635 127.565 80.250 128.135 ;
        RECT 80.915 127.925 81.805 128.095 ;
        RECT 79.595 126.895 79.765 127.395 ;
        RECT 75.835 125.755 76.165 126.515 ;
        RECT 76.345 125.925 76.515 126.685 ;
        RECT 76.775 125.755 77.985 126.845 ;
        RECT 78.340 126.725 79.765 126.895 ;
        RECT 78.340 126.550 78.730 126.725 ;
        RECT 79.215 125.755 79.545 126.555 ;
        RECT 79.935 126.545 80.250 127.565 ;
        RECT 80.915 127.370 81.465 127.755 ;
        RECT 81.635 127.200 81.805 127.925 ;
        RECT 80.915 127.130 81.805 127.200 ;
        RECT 81.975 127.600 82.195 128.085 ;
        RECT 82.365 127.765 82.615 128.305 ;
        RECT 82.785 127.655 83.045 128.135 ;
        RECT 84.005 127.905 84.335 128.305 ;
        RECT 84.505 127.735 84.835 128.075 ;
        RECT 85.885 127.905 86.215 128.305 ;
        RECT 81.975 127.175 82.305 127.600 ;
        RECT 80.915 127.105 81.810 127.130 ;
        RECT 80.915 127.090 81.820 127.105 ;
        RECT 80.915 127.075 81.825 127.090 ;
        RECT 80.915 127.070 81.835 127.075 ;
        RECT 80.915 127.060 81.840 127.070 ;
        RECT 80.915 127.050 81.845 127.060 ;
        RECT 80.915 127.045 81.855 127.050 ;
        RECT 80.915 127.035 81.865 127.045 ;
        RECT 80.915 127.030 81.875 127.035 ;
        RECT 80.915 126.580 81.175 127.030 ;
        RECT 81.540 127.025 81.875 127.030 ;
        RECT 81.540 127.020 81.890 127.025 ;
        RECT 81.540 127.010 81.905 127.020 ;
        RECT 81.540 127.005 81.930 127.010 ;
        RECT 82.475 127.005 82.705 127.400 ;
        RECT 81.540 127.000 82.705 127.005 ;
        RECT 81.570 126.965 82.705 127.000 ;
        RECT 81.605 126.940 82.705 126.965 ;
        RECT 81.635 126.910 82.705 126.940 ;
        RECT 81.655 126.880 82.705 126.910 ;
        RECT 81.675 126.850 82.705 126.880 ;
        RECT 81.745 126.840 82.705 126.850 ;
        RECT 81.770 126.830 82.705 126.840 ;
        RECT 81.790 126.815 82.705 126.830 ;
        RECT 81.810 126.800 82.705 126.815 ;
        RECT 81.815 126.790 82.600 126.800 ;
        RECT 81.830 126.755 82.600 126.790 ;
        RECT 79.715 125.925 80.250 126.545 ;
        RECT 81.345 126.435 81.675 126.680 ;
        RECT 81.845 126.505 82.600 126.755 ;
        RECT 82.875 126.625 83.045 127.655 ;
        RECT 81.345 126.410 81.530 126.435 ;
        RECT 80.915 126.310 81.530 126.410 ;
        RECT 80.915 125.755 81.520 126.310 ;
        RECT 81.695 125.925 82.175 126.265 ;
        RECT 82.345 125.755 82.600 126.300 ;
        RECT 82.770 125.925 83.045 126.625 ;
        RECT 83.850 127.565 86.215 127.735 ;
        RECT 86.385 127.580 86.715 128.090 ;
        RECT 86.900 127.815 87.155 128.305 ;
        RECT 87.325 127.795 88.555 128.135 ;
        RECT 83.850 126.565 84.020 127.565 ;
        RECT 86.045 127.395 86.215 127.565 ;
        RECT 84.190 126.735 84.435 127.395 ;
        RECT 84.650 126.735 84.915 127.395 ;
        RECT 85.110 126.735 85.395 127.395 ;
        RECT 85.570 127.065 85.875 127.395 ;
        RECT 86.045 127.065 86.355 127.395 ;
        RECT 85.570 126.735 85.785 127.065 ;
        RECT 83.850 126.395 84.305 126.565 ;
        RECT 83.975 125.965 84.305 126.395 ;
        RECT 84.485 126.395 85.775 126.565 ;
        RECT 84.485 125.975 84.735 126.395 ;
        RECT 84.965 125.755 85.295 126.225 ;
        RECT 85.525 125.975 85.775 126.395 ;
        RECT 85.965 125.755 86.215 126.895 ;
        RECT 86.525 126.815 86.715 127.580 ;
        RECT 86.920 127.065 87.140 127.645 ;
        RECT 87.325 126.895 87.505 127.795 ;
        RECT 87.675 127.065 88.050 127.625 ;
        RECT 88.225 127.565 88.555 127.795 ;
        RECT 88.735 127.505 89.430 128.135 ;
        RECT 89.635 127.505 89.945 128.305 ;
        RECT 91.085 127.915 91.415 128.305 ;
        RECT 91.585 127.735 91.755 128.055 ;
        RECT 91.925 127.915 92.255 128.305 ;
        RECT 92.670 127.905 93.625 128.075 ;
        RECT 91.035 127.565 93.285 127.735 ;
        RECT 88.255 127.065 88.565 127.395 ;
        RECT 88.755 127.065 89.090 127.315 ;
        RECT 89.260 126.905 89.430 127.505 ;
        RECT 89.600 127.065 89.935 127.335 ;
        RECT 86.385 125.965 86.715 126.815 ;
        RECT 86.900 125.755 87.155 126.895 ;
        RECT 87.325 126.725 88.555 126.895 ;
        RECT 87.325 125.925 87.655 126.725 ;
        RECT 87.825 125.755 88.055 126.555 ;
        RECT 88.225 125.925 88.555 126.725 ;
        RECT 88.735 125.755 88.995 126.895 ;
        RECT 89.165 125.925 89.495 126.905 ;
        RECT 89.665 125.755 89.945 126.895 ;
        RECT 91.035 126.605 91.205 127.565 ;
        RECT 91.375 126.945 91.620 127.395 ;
        RECT 91.790 127.115 92.340 127.315 ;
        RECT 92.510 127.145 92.885 127.315 ;
        RECT 92.510 126.945 92.680 127.145 ;
        RECT 93.055 127.065 93.285 127.565 ;
        RECT 91.375 126.775 92.680 126.945 ;
        RECT 93.455 127.025 93.625 127.905 ;
        RECT 93.795 127.470 94.085 128.305 ;
        RECT 94.715 127.630 94.975 128.135 ;
        RECT 95.155 127.925 95.485 128.305 ;
        RECT 95.665 127.755 95.835 128.135 ;
        RECT 93.455 126.855 94.085 127.025 ;
        RECT 91.035 125.925 91.415 126.605 ;
        RECT 92.005 125.755 92.175 126.605 ;
        RECT 92.345 126.435 93.585 126.605 ;
        RECT 92.345 125.925 92.675 126.435 ;
        RECT 92.845 125.755 93.015 126.265 ;
        RECT 93.185 125.925 93.585 126.435 ;
        RECT 93.765 125.925 94.085 126.855 ;
        RECT 94.715 126.830 94.885 127.630 ;
        RECT 95.170 127.585 95.835 127.755 ;
        RECT 95.170 127.330 95.340 127.585 ;
        RECT 96.555 127.580 96.845 128.305 ;
        RECT 97.015 127.565 97.455 128.125 ;
        RECT 97.625 127.565 98.075 128.305 ;
        RECT 98.245 127.735 98.415 128.135 ;
        RECT 98.585 127.905 99.005 128.305 ;
        RECT 99.175 127.735 99.405 128.135 ;
        RECT 98.245 127.565 99.405 127.735 ;
        RECT 99.575 127.565 100.065 128.135 ;
        RECT 100.325 127.755 100.495 128.135 ;
        RECT 100.675 127.925 101.005 128.305 ;
        RECT 100.325 127.585 100.990 127.755 ;
        RECT 101.185 127.630 101.445 128.135 ;
        RECT 95.055 127.000 95.340 127.330 ;
        RECT 95.575 127.035 95.905 127.405 ;
        RECT 95.170 126.855 95.340 127.000 ;
        RECT 94.715 125.925 94.985 126.830 ;
        RECT 95.170 126.685 95.835 126.855 ;
        RECT 95.155 125.755 95.485 126.515 ;
        RECT 95.665 125.925 95.835 126.685 ;
        RECT 96.555 125.755 96.845 126.920 ;
        RECT 97.015 126.555 97.325 127.565 ;
        RECT 97.495 126.945 97.665 127.395 ;
        RECT 97.835 127.115 98.225 127.395 ;
        RECT 98.410 127.065 98.655 127.395 ;
        RECT 97.495 126.775 98.285 126.945 ;
        RECT 97.015 125.925 97.455 126.555 ;
        RECT 97.630 125.755 97.945 126.605 ;
        RECT 98.115 126.095 98.285 126.775 ;
        RECT 98.455 126.265 98.655 127.065 ;
        RECT 98.855 126.265 99.105 127.395 ;
        RECT 99.320 127.065 99.725 127.395 ;
        RECT 99.895 126.895 100.065 127.565 ;
        RECT 100.255 127.035 100.585 127.405 ;
        RECT 100.820 127.330 100.990 127.585 ;
        RECT 99.295 126.725 100.065 126.895 ;
        RECT 100.820 127.000 101.105 127.330 ;
        RECT 100.820 126.855 100.990 127.000 ;
        RECT 99.295 126.095 99.545 126.725 ;
        RECT 100.325 126.685 100.990 126.855 ;
        RECT 101.275 126.830 101.445 127.630 ;
        RECT 98.115 125.925 99.545 126.095 ;
        RECT 99.725 125.755 100.055 126.555 ;
        RECT 100.325 125.925 100.495 126.685 ;
        RECT 100.675 125.755 101.005 126.515 ;
        RECT 101.175 125.925 101.445 126.830 ;
        RECT 101.615 127.630 101.875 128.135 ;
        RECT 102.055 127.925 102.385 128.305 ;
        RECT 102.565 127.755 102.735 128.135 ;
        RECT 101.615 126.830 101.785 127.630 ;
        RECT 102.070 127.585 102.735 127.755 ;
        RECT 102.070 127.330 102.240 127.585 ;
        RECT 102.995 127.505 103.690 128.135 ;
        RECT 103.895 127.505 104.205 128.305 ;
        RECT 101.955 127.000 102.240 127.330 ;
        RECT 102.475 127.035 102.805 127.405 ;
        RECT 103.015 127.065 103.350 127.315 ;
        RECT 102.070 126.855 102.240 127.000 ;
        RECT 103.520 126.905 103.690 127.505 ;
        RECT 104.375 127.360 104.715 128.135 ;
        RECT 104.885 127.845 105.055 128.305 ;
        RECT 105.295 127.870 105.655 128.135 ;
        RECT 105.295 127.865 105.650 127.870 ;
        RECT 105.295 127.855 105.645 127.865 ;
        RECT 105.295 127.850 105.640 127.855 ;
        RECT 105.295 127.840 105.635 127.850 ;
        RECT 106.285 127.845 106.455 128.305 ;
        RECT 105.295 127.835 105.630 127.840 ;
        RECT 105.295 127.825 105.620 127.835 ;
        RECT 105.295 127.815 105.610 127.825 ;
        RECT 105.295 127.675 105.595 127.815 ;
        RECT 104.885 127.485 105.595 127.675 ;
        RECT 105.785 127.675 106.115 127.755 ;
        RECT 106.625 127.675 106.965 128.135 ;
        RECT 105.785 127.485 106.965 127.675 ;
        RECT 107.135 127.675 107.475 128.135 ;
        RECT 107.645 127.845 107.815 128.305 ;
        RECT 108.445 127.870 108.805 128.135 ;
        RECT 108.450 127.865 108.805 127.870 ;
        RECT 108.455 127.855 108.805 127.865 ;
        RECT 108.460 127.850 108.805 127.855 ;
        RECT 108.465 127.840 108.805 127.850 ;
        RECT 109.045 127.845 109.215 128.305 ;
        RECT 108.470 127.835 108.805 127.840 ;
        RECT 108.480 127.825 108.805 127.835 ;
        RECT 108.490 127.815 108.805 127.825 ;
        RECT 107.985 127.675 108.315 127.755 ;
        RECT 107.135 127.485 108.315 127.675 ;
        RECT 108.505 127.675 108.805 127.815 ;
        RECT 108.505 127.485 109.215 127.675 ;
        RECT 103.860 127.065 104.195 127.335 ;
        RECT 101.615 125.925 101.885 126.830 ;
        RECT 102.070 126.685 102.735 126.855 ;
        RECT 102.055 125.755 102.385 126.515 ;
        RECT 102.565 125.925 102.735 126.685 ;
        RECT 102.995 125.755 103.255 126.895 ;
        RECT 103.425 125.925 103.755 126.905 ;
        RECT 103.925 125.755 104.205 126.895 ;
        RECT 104.375 125.925 104.655 127.360 ;
        RECT 104.885 126.915 105.170 127.485 ;
        RECT 105.355 127.085 105.825 127.315 ;
        RECT 105.995 127.295 106.325 127.315 ;
        RECT 105.995 127.115 106.445 127.295 ;
        RECT 106.635 127.115 106.965 127.315 ;
        RECT 104.885 126.700 106.035 126.915 ;
        RECT 104.825 125.755 105.535 126.530 ;
        RECT 105.705 125.925 106.035 126.700 ;
        RECT 106.230 126.000 106.445 127.115 ;
        RECT 106.735 126.775 106.965 127.115 ;
        RECT 107.135 127.115 107.465 127.315 ;
        RECT 107.775 127.295 108.105 127.315 ;
        RECT 107.655 127.115 108.105 127.295 ;
        RECT 107.135 126.775 107.365 127.115 ;
        RECT 106.625 125.755 106.955 126.475 ;
        RECT 107.145 125.755 107.475 126.475 ;
        RECT 107.655 126.000 107.870 127.115 ;
        RECT 108.275 127.085 108.745 127.315 ;
        RECT 108.930 126.915 109.215 127.485 ;
        RECT 109.385 127.360 109.725 128.135 ;
        RECT 108.065 126.700 109.215 126.915 ;
        RECT 108.065 125.925 108.395 126.700 ;
        RECT 108.565 125.755 109.275 126.530 ;
        RECT 109.445 125.925 109.725 127.360 ;
        RECT 109.895 127.535 111.565 128.305 ;
        RECT 109.895 127.015 110.645 127.535 ;
        RECT 110.815 126.845 111.565 127.365 ;
        RECT 109.895 125.755 111.565 126.845 ;
        RECT 112.195 127.360 112.535 128.135 ;
        RECT 112.705 127.845 112.875 128.305 ;
        RECT 113.115 127.870 113.475 128.135 ;
        RECT 113.115 127.865 113.470 127.870 ;
        RECT 113.115 127.855 113.465 127.865 ;
        RECT 113.115 127.850 113.460 127.855 ;
        RECT 113.115 127.840 113.455 127.850 ;
        RECT 114.105 127.845 114.275 128.305 ;
        RECT 113.115 127.835 113.450 127.840 ;
        RECT 113.115 127.825 113.440 127.835 ;
        RECT 113.115 127.815 113.430 127.825 ;
        RECT 113.115 127.675 113.415 127.815 ;
        RECT 112.705 127.485 113.415 127.675 ;
        RECT 113.605 127.675 113.935 127.755 ;
        RECT 114.445 127.675 114.785 128.135 ;
        RECT 113.605 127.485 114.785 127.675 ;
        RECT 114.955 127.505 115.295 128.135 ;
        RECT 115.465 127.505 115.715 128.305 ;
        RECT 115.905 127.655 116.235 128.135 ;
        RECT 116.405 127.845 116.630 128.305 ;
        RECT 116.800 127.655 117.130 128.135 ;
        RECT 112.195 125.925 112.475 127.360 ;
        RECT 112.705 126.915 112.990 127.485 ;
        RECT 113.175 127.085 113.645 127.315 ;
        RECT 113.815 127.295 114.145 127.315 ;
        RECT 113.815 127.115 114.265 127.295 ;
        RECT 114.455 127.115 114.785 127.315 ;
        RECT 112.705 126.700 113.855 126.915 ;
        RECT 112.645 125.755 113.355 126.530 ;
        RECT 113.525 125.925 113.855 126.700 ;
        RECT 114.050 126.000 114.265 127.115 ;
        RECT 114.555 126.775 114.785 127.115 ;
        RECT 114.955 126.895 115.130 127.505 ;
        RECT 115.905 127.485 117.130 127.655 ;
        RECT 117.760 127.525 118.260 128.135 ;
        RECT 118.635 127.565 119.075 128.125 ;
        RECT 119.245 127.565 119.695 128.305 ;
        RECT 119.865 127.735 120.035 128.135 ;
        RECT 120.205 127.905 120.625 128.305 ;
        RECT 120.795 127.735 121.025 128.135 ;
        RECT 119.865 127.565 121.025 127.735 ;
        RECT 121.195 127.565 121.685 128.135 ;
        RECT 122.315 127.580 122.605 128.305 ;
        RECT 122.775 127.675 123.115 128.135 ;
        RECT 123.285 127.845 123.455 128.305 ;
        RECT 124.085 127.870 124.445 128.135 ;
        RECT 124.090 127.865 124.445 127.870 ;
        RECT 124.095 127.855 124.445 127.865 ;
        RECT 124.100 127.850 124.445 127.855 ;
        RECT 124.105 127.840 124.445 127.850 ;
        RECT 124.685 127.845 124.855 128.305 ;
        RECT 124.110 127.835 124.445 127.840 ;
        RECT 124.120 127.825 124.445 127.835 ;
        RECT 124.130 127.815 124.445 127.825 ;
        RECT 123.625 127.675 123.955 127.755 ;
        RECT 115.300 127.145 115.995 127.315 ;
        RECT 115.825 126.895 115.995 127.145 ;
        RECT 116.170 127.115 116.590 127.315 ;
        RECT 116.760 127.115 117.090 127.315 ;
        RECT 117.260 127.115 117.590 127.315 ;
        RECT 117.760 126.895 117.930 127.525 ;
        RECT 118.115 127.065 118.465 127.315 ;
        RECT 114.445 125.755 114.775 126.475 ;
        RECT 114.955 125.925 115.295 126.895 ;
        RECT 115.465 125.755 115.635 126.895 ;
        RECT 115.825 126.725 118.260 126.895 ;
        RECT 115.905 125.755 116.155 126.555 ;
        RECT 116.800 125.925 117.130 126.725 ;
        RECT 117.430 125.755 117.760 126.555 ;
        RECT 117.930 125.925 118.260 126.725 ;
        RECT 118.635 126.555 118.945 127.565 ;
        RECT 119.115 126.945 119.285 127.395 ;
        RECT 119.455 127.115 119.845 127.395 ;
        RECT 120.030 127.065 120.275 127.395 ;
        RECT 119.115 126.775 119.905 126.945 ;
        RECT 118.635 125.925 119.075 126.555 ;
        RECT 119.250 125.755 119.565 126.605 ;
        RECT 119.735 126.095 119.905 126.775 ;
        RECT 120.075 126.265 120.275 127.065 ;
        RECT 120.475 126.265 120.725 127.395 ;
        RECT 120.940 127.065 121.345 127.395 ;
        RECT 121.515 126.895 121.685 127.565 ;
        RECT 122.775 127.485 123.955 127.675 ;
        RECT 124.145 127.675 124.445 127.815 ;
        RECT 124.145 127.485 124.855 127.675 ;
        RECT 122.775 127.115 123.105 127.315 ;
        RECT 123.415 127.295 123.745 127.315 ;
        RECT 123.295 127.115 123.745 127.295 ;
        RECT 120.915 126.725 121.685 126.895 ;
        RECT 120.915 126.095 121.165 126.725 ;
        RECT 119.735 125.925 121.165 126.095 ;
        RECT 121.345 125.755 121.675 126.555 ;
        RECT 122.315 125.755 122.605 126.920 ;
        RECT 122.775 126.775 123.005 127.115 ;
        RECT 122.785 125.755 123.115 126.475 ;
        RECT 123.295 126.000 123.510 127.115 ;
        RECT 123.915 127.085 124.385 127.315 ;
        RECT 124.570 126.915 124.855 127.485 ;
        RECT 125.025 127.360 125.365 128.135 ;
        RECT 125.595 127.825 125.875 128.305 ;
        RECT 126.045 127.655 126.305 128.045 ;
        RECT 126.480 127.825 126.735 128.305 ;
        RECT 126.905 127.655 127.200 128.045 ;
        RECT 127.380 127.825 127.655 128.305 ;
        RECT 127.825 127.805 128.125 128.135 ;
        RECT 123.705 126.700 124.855 126.915 ;
        RECT 123.705 125.925 124.035 126.700 ;
        RECT 124.205 125.755 124.915 126.530 ;
        RECT 125.085 125.925 125.365 127.360 ;
        RECT 125.550 127.485 127.200 127.655 ;
        RECT 125.550 126.975 125.955 127.485 ;
        RECT 126.125 127.145 127.265 127.315 ;
        RECT 125.550 126.805 126.305 126.975 ;
        RECT 125.590 125.755 125.875 126.625 ;
        RECT 126.045 126.555 126.305 126.805 ;
        RECT 127.095 126.895 127.265 127.145 ;
        RECT 127.435 127.065 127.785 127.635 ;
        RECT 127.955 126.895 128.125 127.805 ;
        RECT 128.295 127.675 128.635 128.135 ;
        RECT 128.805 127.845 128.975 128.305 ;
        RECT 129.605 127.870 129.965 128.135 ;
        RECT 129.610 127.865 129.965 127.870 ;
        RECT 129.615 127.855 129.965 127.865 ;
        RECT 129.620 127.850 129.965 127.855 ;
        RECT 129.625 127.840 129.965 127.850 ;
        RECT 130.205 127.845 130.375 128.305 ;
        RECT 129.630 127.835 129.965 127.840 ;
        RECT 129.640 127.825 129.965 127.835 ;
        RECT 129.650 127.815 129.965 127.825 ;
        RECT 129.145 127.675 129.475 127.755 ;
        RECT 128.295 127.485 129.475 127.675 ;
        RECT 129.665 127.675 129.965 127.815 ;
        RECT 129.665 127.485 130.375 127.675 ;
        RECT 127.095 126.725 128.125 126.895 ;
        RECT 128.295 127.115 128.625 127.315 ;
        RECT 128.935 127.295 129.265 127.315 ;
        RECT 128.815 127.115 129.265 127.295 ;
        RECT 128.295 126.775 128.525 127.115 ;
        RECT 126.045 126.385 127.165 126.555 ;
        RECT 126.045 125.925 126.305 126.385 ;
        RECT 126.480 125.755 126.735 126.215 ;
        RECT 126.905 125.925 127.165 126.385 ;
        RECT 127.335 125.755 127.645 126.555 ;
        RECT 127.815 125.925 128.125 126.725 ;
        RECT 128.305 125.755 128.635 126.475 ;
        RECT 128.815 126.000 129.030 127.115 ;
        RECT 129.435 127.085 129.905 127.315 ;
        RECT 130.090 126.915 130.375 127.485 ;
        RECT 130.545 127.360 130.885 128.135 ;
        RECT 129.225 126.700 130.375 126.915 ;
        RECT 129.225 125.925 129.555 126.700 ;
        RECT 129.725 125.755 130.435 126.530 ;
        RECT 130.605 125.925 130.885 127.360 ;
        RECT 131.055 127.360 131.395 128.135 ;
        RECT 131.565 127.845 131.735 128.305 ;
        RECT 131.975 127.870 132.335 128.135 ;
        RECT 131.975 127.865 132.330 127.870 ;
        RECT 131.975 127.855 132.325 127.865 ;
        RECT 131.975 127.850 132.320 127.855 ;
        RECT 131.975 127.840 132.315 127.850 ;
        RECT 132.965 127.845 133.135 128.305 ;
        RECT 131.975 127.835 132.310 127.840 ;
        RECT 131.975 127.825 132.300 127.835 ;
        RECT 131.975 127.815 132.290 127.825 ;
        RECT 131.975 127.675 132.275 127.815 ;
        RECT 131.565 127.485 132.275 127.675 ;
        RECT 132.465 127.675 132.795 127.755 ;
        RECT 133.305 127.675 133.645 128.135 ;
        RECT 132.465 127.485 133.645 127.675 ;
        RECT 131.055 125.925 131.335 127.360 ;
        RECT 131.565 126.915 131.850 127.485 ;
        RECT 133.815 127.360 134.155 128.135 ;
        RECT 134.325 127.845 134.495 128.305 ;
        RECT 134.735 127.870 135.095 128.135 ;
        RECT 134.735 127.865 135.090 127.870 ;
        RECT 134.735 127.855 135.085 127.865 ;
        RECT 134.735 127.850 135.080 127.855 ;
        RECT 134.735 127.840 135.075 127.850 ;
        RECT 135.725 127.845 135.895 128.305 ;
        RECT 134.735 127.835 135.070 127.840 ;
        RECT 134.735 127.825 135.060 127.835 ;
        RECT 134.735 127.815 135.050 127.825 ;
        RECT 134.735 127.675 135.035 127.815 ;
        RECT 134.325 127.485 135.035 127.675 ;
        RECT 135.225 127.675 135.555 127.755 ;
        RECT 136.065 127.675 136.405 128.135 ;
        RECT 135.225 127.485 136.405 127.675 ;
        RECT 132.035 127.085 132.505 127.315 ;
        RECT 132.675 127.295 133.005 127.315 ;
        RECT 132.675 127.115 133.125 127.295 ;
        RECT 133.315 127.115 133.645 127.315 ;
        RECT 131.565 126.700 132.715 126.915 ;
        RECT 131.505 125.755 132.215 126.530 ;
        RECT 132.385 125.925 132.715 126.700 ;
        RECT 132.910 126.000 133.125 127.115 ;
        RECT 133.415 126.775 133.645 127.115 ;
        RECT 133.305 125.755 133.635 126.475 ;
        RECT 133.815 125.925 134.095 127.360 ;
        RECT 134.325 126.915 134.610 127.485 ;
        RECT 136.575 127.360 136.915 128.135 ;
        RECT 137.085 127.845 137.255 128.305 ;
        RECT 137.495 127.870 137.855 128.135 ;
        RECT 137.495 127.865 137.850 127.870 ;
        RECT 137.495 127.855 137.845 127.865 ;
        RECT 137.495 127.850 137.840 127.855 ;
        RECT 137.495 127.840 137.835 127.850 ;
        RECT 138.485 127.845 138.655 128.305 ;
        RECT 137.495 127.835 137.830 127.840 ;
        RECT 137.495 127.825 137.820 127.835 ;
        RECT 137.495 127.815 137.810 127.825 ;
        RECT 137.495 127.675 137.795 127.815 ;
        RECT 137.085 127.485 137.795 127.675 ;
        RECT 137.985 127.675 138.315 127.755 ;
        RECT 138.825 127.675 139.165 128.135 ;
        RECT 137.985 127.485 139.165 127.675 ;
        RECT 139.335 127.675 139.675 128.135 ;
        RECT 139.845 127.845 140.015 128.305 ;
        RECT 140.645 127.870 141.005 128.135 ;
        RECT 140.650 127.865 141.005 127.870 ;
        RECT 140.655 127.855 141.005 127.865 ;
        RECT 140.660 127.850 141.005 127.855 ;
        RECT 140.665 127.840 141.005 127.850 ;
        RECT 141.245 127.845 141.415 128.305 ;
        RECT 140.670 127.835 141.005 127.840 ;
        RECT 140.680 127.825 141.005 127.835 ;
        RECT 140.690 127.815 141.005 127.825 ;
        RECT 140.185 127.675 140.515 127.755 ;
        RECT 139.335 127.485 140.515 127.675 ;
        RECT 140.705 127.675 141.005 127.815 ;
        RECT 140.705 127.485 141.415 127.675 ;
        RECT 134.795 127.085 135.265 127.315 ;
        RECT 135.435 127.295 135.765 127.315 ;
        RECT 135.435 127.115 135.885 127.295 ;
        RECT 136.075 127.115 136.405 127.315 ;
        RECT 134.325 126.700 135.475 126.915 ;
        RECT 134.265 125.755 134.975 126.530 ;
        RECT 135.145 125.925 135.475 126.700 ;
        RECT 135.670 126.000 135.885 127.115 ;
        RECT 136.175 126.775 136.405 127.115 ;
        RECT 136.065 125.755 136.395 126.475 ;
        RECT 136.575 125.925 136.855 127.360 ;
        RECT 137.085 126.915 137.370 127.485 ;
        RECT 137.555 127.085 138.025 127.315 ;
        RECT 138.195 127.295 138.525 127.315 ;
        RECT 138.195 127.115 138.645 127.295 ;
        RECT 138.835 127.115 139.165 127.315 ;
        RECT 137.085 126.700 138.235 126.915 ;
        RECT 137.025 125.755 137.735 126.530 ;
        RECT 137.905 125.925 138.235 126.700 ;
        RECT 138.430 126.000 138.645 127.115 ;
        RECT 138.935 126.775 139.165 127.115 ;
        RECT 139.335 127.115 139.665 127.315 ;
        RECT 139.975 127.295 140.305 127.315 ;
        RECT 139.855 127.115 140.305 127.295 ;
        RECT 139.335 126.775 139.565 127.115 ;
        RECT 138.825 125.755 139.155 126.475 ;
        RECT 139.345 125.755 139.675 126.475 ;
        RECT 139.855 126.000 140.070 127.115 ;
        RECT 140.475 127.085 140.945 127.315 ;
        RECT 141.130 126.915 141.415 127.485 ;
        RECT 141.585 127.360 141.925 128.135 ;
        RECT 142.185 127.755 142.355 128.135 ;
        RECT 142.570 127.925 142.900 128.305 ;
        RECT 142.185 127.585 142.900 127.755 ;
        RECT 140.265 126.700 141.415 126.915 ;
        RECT 140.265 125.925 140.595 126.700 ;
        RECT 140.765 125.755 141.475 126.530 ;
        RECT 141.645 125.925 141.925 127.360 ;
        RECT 142.095 127.035 142.450 127.405 ;
        RECT 142.730 127.395 142.900 127.585 ;
        RECT 143.070 127.560 143.325 128.135 ;
        RECT 142.730 127.065 142.985 127.395 ;
        RECT 142.730 126.855 142.900 127.065 ;
        RECT 142.185 126.685 142.900 126.855 ;
        RECT 143.155 126.830 143.325 127.560 ;
        RECT 143.500 127.465 143.760 128.305 ;
        RECT 143.935 127.565 144.400 128.110 ;
        RECT 142.185 125.925 142.355 126.685 ;
        RECT 142.570 125.755 142.900 126.515 ;
        RECT 143.070 125.925 143.325 126.830 ;
        RECT 143.500 125.755 143.760 126.905 ;
        RECT 143.935 126.605 144.105 127.565 ;
        RECT 144.905 127.485 145.075 128.305 ;
        RECT 145.245 127.655 145.575 128.135 ;
        RECT 145.745 127.915 146.095 128.305 ;
        RECT 146.265 127.735 146.495 128.135 ;
        RECT 145.985 127.655 146.495 127.735 ;
        RECT 145.245 127.565 146.495 127.655 ;
        RECT 146.665 127.565 146.985 128.045 ;
        RECT 148.075 127.580 148.365 128.305 ;
        RECT 148.535 127.805 148.835 128.135 ;
        RECT 149.005 127.825 149.280 128.305 ;
        RECT 145.245 127.485 146.155 127.565 ;
        RECT 144.275 126.945 144.520 127.395 ;
        RECT 144.780 127.115 145.475 127.315 ;
        RECT 145.645 127.145 146.245 127.315 ;
        RECT 145.645 126.945 145.815 127.145 ;
        RECT 146.475 126.975 146.645 127.395 ;
        RECT 144.275 126.775 145.815 126.945 ;
        RECT 145.985 126.805 146.645 126.975 ;
        RECT 145.985 126.605 146.155 126.805 ;
        RECT 146.815 126.635 146.985 127.565 ;
        RECT 143.935 126.435 146.155 126.605 ;
        RECT 146.325 126.435 146.985 126.635 ;
        RECT 143.935 125.755 144.235 126.265 ;
        RECT 144.405 125.925 144.735 126.435 ;
        RECT 146.325 126.265 146.495 126.435 ;
        RECT 144.905 125.755 145.535 126.265 ;
        RECT 146.115 126.095 146.495 126.265 ;
        RECT 146.665 125.755 146.965 126.265 ;
        RECT 148.075 125.755 148.365 126.920 ;
        RECT 148.535 126.895 148.705 127.805 ;
        RECT 149.460 127.655 149.755 128.045 ;
        RECT 149.925 127.825 150.180 128.305 ;
        RECT 150.355 127.655 150.615 128.045 ;
        RECT 150.785 127.825 151.065 128.305 ;
        RECT 148.875 127.065 149.225 127.635 ;
        RECT 149.460 127.485 151.110 127.655 ;
        RECT 149.395 127.145 150.535 127.315 ;
        RECT 149.395 126.895 149.565 127.145 ;
        RECT 150.705 126.975 151.110 127.485 ;
        RECT 148.535 126.725 149.565 126.895 ;
        RECT 150.355 126.805 151.110 126.975 ;
        RECT 151.330 127.565 151.945 128.135 ;
        RECT 152.115 127.795 152.330 128.305 ;
        RECT 152.560 127.795 152.840 128.125 ;
        RECT 153.020 127.795 153.260 128.305 ;
        RECT 148.535 125.925 148.845 126.725 ;
        RECT 150.355 126.555 150.615 126.805 ;
        RECT 149.015 125.755 149.325 126.555 ;
        RECT 149.495 126.385 150.615 126.555 ;
        RECT 149.495 125.925 149.755 126.385 ;
        RECT 149.925 125.755 150.180 126.215 ;
        RECT 150.355 125.925 150.615 126.385 ;
        RECT 150.785 125.755 151.070 126.625 ;
        RECT 151.330 126.545 151.645 127.565 ;
        RECT 151.815 126.895 151.985 127.395 ;
        RECT 152.235 127.065 152.500 127.625 ;
        RECT 152.670 126.895 152.840 127.795 ;
        RECT 153.010 127.065 153.365 127.625 ;
        RECT 153.595 127.555 154.805 128.305 ;
        RECT 154.975 127.555 156.185 128.305 ;
        RECT 153.595 127.015 154.115 127.555 ;
        RECT 151.815 126.725 153.240 126.895 ;
        RECT 154.285 126.845 154.805 127.385 ;
        RECT 151.330 125.925 151.865 126.545 ;
        RECT 152.035 125.755 152.365 126.555 ;
        RECT 152.850 126.550 153.240 126.725 ;
        RECT 153.595 125.755 154.805 126.845 ;
        RECT 154.975 126.845 155.495 127.385 ;
        RECT 155.665 127.015 156.185 127.555 ;
        RECT 154.975 125.755 156.185 126.845 ;
        RECT 70.710 125.585 156.270 125.755 ;
        RECT 70.795 124.495 72.005 125.585 ;
        RECT 70.795 123.785 71.315 124.325 ;
        RECT 71.485 123.955 72.005 124.495 ;
        RECT 72.180 124.435 72.440 125.585 ;
        RECT 72.615 124.510 72.870 125.415 ;
        RECT 73.040 124.825 73.370 125.585 ;
        RECT 73.585 124.655 73.755 125.415 ;
        RECT 74.070 124.715 74.355 125.585 ;
        RECT 74.525 124.955 74.785 125.415 ;
        RECT 74.960 125.125 75.215 125.585 ;
        RECT 75.385 124.955 75.645 125.415 ;
        RECT 74.525 124.785 75.645 124.955 ;
        RECT 75.815 124.785 76.125 125.585 ;
        RECT 70.795 123.035 72.005 123.785 ;
        RECT 72.180 123.035 72.440 123.875 ;
        RECT 72.615 123.780 72.785 124.510 ;
        RECT 73.040 124.485 73.755 124.655 ;
        RECT 74.525 124.535 74.785 124.785 ;
        RECT 76.295 124.615 76.605 125.415 ;
        RECT 73.040 124.275 73.210 124.485 ;
        RECT 74.030 124.365 74.785 124.535 ;
        RECT 75.575 124.445 76.605 124.615 ;
        RECT 76.775 124.495 78.445 125.585 ;
        RECT 72.955 123.945 73.210 124.275 ;
        RECT 72.615 123.205 72.870 123.780 ;
        RECT 73.040 123.755 73.210 123.945 ;
        RECT 73.490 123.935 73.845 124.305 ;
        RECT 74.030 123.855 74.435 124.365 ;
        RECT 75.575 124.195 75.745 124.445 ;
        RECT 74.605 124.025 75.745 124.195 ;
        RECT 73.040 123.585 73.755 123.755 ;
        RECT 74.030 123.685 75.680 123.855 ;
        RECT 75.915 123.705 76.265 124.275 ;
        RECT 73.040 123.035 73.370 123.415 ;
        RECT 73.585 123.205 73.755 123.585 ;
        RECT 74.075 123.035 74.355 123.515 ;
        RECT 74.525 123.295 74.785 123.685 ;
        RECT 74.960 123.035 75.215 123.515 ;
        RECT 75.385 123.295 75.680 123.685 ;
        RECT 76.435 123.535 76.605 124.445 ;
        RECT 75.860 123.035 76.135 123.515 ;
        RECT 76.305 123.205 76.605 123.535 ;
        RECT 76.775 123.805 77.525 124.325 ;
        RECT 77.695 123.975 78.445 124.495 ;
        RECT 79.080 124.445 79.335 125.585 ;
        RECT 79.505 124.615 79.835 125.415 ;
        RECT 80.005 124.785 80.235 125.585 ;
        RECT 80.405 124.615 80.735 125.415 ;
        RECT 79.505 124.445 80.735 124.615 ;
        RECT 76.775 123.035 78.445 123.805 ;
        RECT 79.100 123.695 79.320 124.275 ;
        RECT 79.505 123.545 79.685 124.445 ;
        RECT 80.920 124.435 81.180 125.585 ;
        RECT 81.355 124.510 81.610 125.415 ;
        RECT 81.780 124.825 82.110 125.585 ;
        RECT 82.325 124.655 82.495 125.415 ;
        RECT 79.855 123.715 80.230 124.275 ;
        RECT 80.435 123.945 80.745 124.275 ;
        RECT 80.405 123.545 80.735 123.775 ;
        RECT 79.080 123.035 79.335 123.525 ;
        RECT 79.505 123.205 80.735 123.545 ;
        RECT 80.920 123.035 81.180 123.875 ;
        RECT 81.355 123.780 81.525 124.510 ;
        RECT 81.780 124.485 82.495 124.655 ;
        RECT 81.780 124.275 81.950 124.485 ;
        RECT 83.675 124.420 83.965 125.585 ;
        RECT 84.140 124.435 84.400 125.585 ;
        RECT 84.575 124.510 84.830 125.415 ;
        RECT 85.000 124.825 85.330 125.585 ;
        RECT 85.545 124.655 85.715 125.415 ;
        RECT 81.695 123.945 81.950 124.275 ;
        RECT 81.355 123.205 81.610 123.780 ;
        RECT 81.780 123.755 81.950 123.945 ;
        RECT 82.230 123.935 82.585 124.305 ;
        RECT 81.780 123.585 82.495 123.755 ;
        RECT 81.780 123.035 82.110 123.415 ;
        RECT 82.325 123.205 82.495 123.585 ;
        RECT 83.675 123.035 83.965 123.760 ;
        RECT 84.140 123.035 84.400 123.875 ;
        RECT 84.575 123.780 84.745 124.510 ;
        RECT 85.000 124.485 85.715 124.655 ;
        RECT 85.000 124.275 85.170 124.485 ;
        RECT 85.980 124.435 86.240 125.585 ;
        RECT 86.415 124.510 86.670 125.415 ;
        RECT 86.840 124.825 87.170 125.585 ;
        RECT 87.385 124.655 87.555 125.415 ;
        RECT 84.915 123.945 85.170 124.275 ;
        RECT 84.575 123.205 84.830 123.780 ;
        RECT 85.000 123.755 85.170 123.945 ;
        RECT 85.450 123.935 85.805 124.305 ;
        RECT 85.000 123.585 85.715 123.755 ;
        RECT 85.000 123.035 85.330 123.415 ;
        RECT 85.545 123.205 85.715 123.585 ;
        RECT 85.980 123.035 86.240 123.875 ;
        RECT 86.415 123.780 86.585 124.510 ;
        RECT 86.840 124.485 87.555 124.655 ;
        RECT 87.815 124.495 89.485 125.585 ;
        RECT 86.840 124.275 87.010 124.485 ;
        RECT 86.755 123.945 87.010 124.275 ;
        RECT 86.415 123.205 86.670 123.780 ;
        RECT 86.840 123.755 87.010 123.945 ;
        RECT 87.290 123.935 87.645 124.305 ;
        RECT 87.815 123.805 88.565 124.325 ;
        RECT 88.735 123.975 89.485 124.495 ;
        RECT 89.660 124.435 89.920 125.585 ;
        RECT 90.095 124.510 90.350 125.415 ;
        RECT 90.520 124.825 90.850 125.585 ;
        RECT 91.065 124.655 91.235 125.415 ;
        RECT 86.840 123.585 87.555 123.755 ;
        RECT 86.840 123.035 87.170 123.415 ;
        RECT 87.385 123.205 87.555 123.585 ;
        RECT 87.815 123.035 89.485 123.805 ;
        RECT 89.660 123.035 89.920 123.875 ;
        RECT 90.095 123.780 90.265 124.510 ;
        RECT 90.520 124.485 91.235 124.655 ;
        RECT 91.495 124.495 93.165 125.585 ;
        RECT 90.520 124.275 90.690 124.485 ;
        RECT 90.435 123.945 90.690 124.275 ;
        RECT 90.095 123.205 90.350 123.780 ;
        RECT 90.520 123.755 90.690 123.945 ;
        RECT 90.970 123.935 91.325 124.305 ;
        RECT 91.495 123.805 92.245 124.325 ;
        RECT 92.415 123.975 93.165 124.495 ;
        RECT 93.340 124.435 93.600 125.585 ;
        RECT 93.775 124.510 94.030 125.415 ;
        RECT 94.200 124.825 94.530 125.585 ;
        RECT 94.745 124.655 94.915 125.415 ;
        RECT 90.520 123.585 91.235 123.755 ;
        RECT 90.520 123.035 90.850 123.415 ;
        RECT 91.065 123.205 91.235 123.585 ;
        RECT 91.495 123.035 93.165 123.805 ;
        RECT 93.340 123.035 93.600 123.875 ;
        RECT 93.775 123.780 93.945 124.510 ;
        RECT 94.200 124.485 94.915 124.655 ;
        RECT 95.175 124.495 96.385 125.585 ;
        RECT 94.200 124.275 94.370 124.485 ;
        RECT 94.115 123.945 94.370 124.275 ;
        RECT 93.775 123.205 94.030 123.780 ;
        RECT 94.200 123.755 94.370 123.945 ;
        RECT 94.650 123.935 95.005 124.305 ;
        RECT 95.175 123.785 95.695 124.325 ;
        RECT 95.865 123.955 96.385 124.495 ;
        RECT 96.555 124.420 96.845 125.585 ;
        RECT 97.020 124.435 97.280 125.585 ;
        RECT 97.455 124.510 97.710 125.415 ;
        RECT 97.880 124.825 98.210 125.585 ;
        RECT 98.425 124.655 98.595 125.415 ;
        RECT 94.200 123.585 94.915 123.755 ;
        RECT 94.200 123.035 94.530 123.415 ;
        RECT 94.745 123.205 94.915 123.585 ;
        RECT 95.175 123.035 96.385 123.785 ;
        RECT 96.555 123.035 96.845 123.760 ;
        RECT 97.020 123.035 97.280 123.875 ;
        RECT 97.455 123.780 97.625 124.510 ;
        RECT 97.880 124.485 98.595 124.655 ;
        RECT 98.855 124.495 100.525 125.585 ;
        RECT 97.880 124.275 98.050 124.485 ;
        RECT 97.795 123.945 98.050 124.275 ;
        RECT 97.455 123.205 97.710 123.780 ;
        RECT 97.880 123.755 98.050 123.945 ;
        RECT 98.330 123.935 98.685 124.305 ;
        RECT 98.855 123.805 99.605 124.325 ;
        RECT 99.775 123.975 100.525 124.495 ;
        RECT 100.700 124.435 100.960 125.585 ;
        RECT 101.135 124.510 101.390 125.415 ;
        RECT 101.560 124.825 101.890 125.585 ;
        RECT 102.105 124.655 102.275 125.415 ;
        RECT 97.880 123.585 98.595 123.755 ;
        RECT 97.880 123.035 98.210 123.415 ;
        RECT 98.425 123.205 98.595 123.585 ;
        RECT 98.855 123.035 100.525 123.805 ;
        RECT 100.700 123.035 100.960 123.875 ;
        RECT 101.135 123.780 101.305 124.510 ;
        RECT 101.560 124.485 102.275 124.655 ;
        RECT 102.535 124.495 104.205 125.585 ;
        RECT 101.560 124.275 101.730 124.485 ;
        RECT 101.475 123.945 101.730 124.275 ;
        RECT 101.135 123.205 101.390 123.780 ;
        RECT 101.560 123.755 101.730 123.945 ;
        RECT 102.010 123.935 102.365 124.305 ;
        RECT 102.535 123.805 103.285 124.325 ;
        RECT 103.455 123.975 104.205 124.495 ;
        RECT 104.465 124.655 104.635 125.415 ;
        RECT 104.850 124.825 105.180 125.585 ;
        RECT 104.465 124.485 105.180 124.655 ;
        RECT 105.350 124.510 105.605 125.415 ;
        RECT 104.375 123.935 104.730 124.305 ;
        RECT 105.010 124.275 105.180 124.485 ;
        RECT 105.010 123.945 105.265 124.275 ;
        RECT 101.560 123.585 102.275 123.755 ;
        RECT 101.560 123.035 101.890 123.415 ;
        RECT 102.105 123.205 102.275 123.585 ;
        RECT 102.535 123.035 104.205 123.805 ;
        RECT 105.010 123.755 105.180 123.945 ;
        RECT 105.435 123.780 105.605 124.510 ;
        RECT 105.780 124.435 106.040 125.585 ;
        RECT 106.215 124.495 107.425 125.585 ;
        RECT 104.465 123.585 105.180 123.755 ;
        RECT 104.465 123.205 104.635 123.585 ;
        RECT 104.850 123.035 105.180 123.415 ;
        RECT 105.350 123.205 105.605 123.780 ;
        RECT 105.780 123.035 106.040 123.875 ;
        RECT 106.215 123.785 106.735 124.325 ;
        RECT 106.905 123.955 107.425 124.495 ;
        RECT 107.600 124.435 107.860 125.585 ;
        RECT 108.035 124.510 108.290 125.415 ;
        RECT 108.460 124.825 108.790 125.585 ;
        RECT 109.005 124.655 109.175 125.415 ;
        RECT 106.215 123.035 107.425 123.785 ;
        RECT 107.600 123.035 107.860 123.875 ;
        RECT 108.035 123.780 108.205 124.510 ;
        RECT 108.460 124.485 109.175 124.655 ;
        RECT 108.460 124.275 108.630 124.485 ;
        RECT 109.435 124.420 109.725 125.585 ;
        RECT 109.895 124.615 110.205 125.415 ;
        RECT 110.375 124.785 110.685 125.585 ;
        RECT 110.855 124.955 111.115 125.415 ;
        RECT 111.285 125.125 111.540 125.585 ;
        RECT 111.715 124.955 111.975 125.415 ;
        RECT 110.855 124.785 111.975 124.955 ;
        RECT 109.895 124.445 110.925 124.615 ;
        RECT 108.375 123.945 108.630 124.275 ;
        RECT 108.035 123.205 108.290 123.780 ;
        RECT 108.460 123.755 108.630 123.945 ;
        RECT 108.910 123.935 109.265 124.305 ;
        RECT 108.460 123.585 109.175 123.755 ;
        RECT 108.460 123.035 108.790 123.415 ;
        RECT 109.005 123.205 109.175 123.585 ;
        RECT 109.435 123.035 109.725 123.760 ;
        RECT 109.895 123.535 110.065 124.445 ;
        RECT 110.235 123.705 110.585 124.275 ;
        RECT 110.755 124.195 110.925 124.445 ;
        RECT 111.715 124.535 111.975 124.785 ;
        RECT 112.145 124.715 112.430 125.585 ;
        RECT 111.715 124.365 112.470 124.535 ;
        RECT 112.655 124.495 113.865 125.585 ;
        RECT 114.090 124.715 114.375 125.585 ;
        RECT 114.545 124.955 114.805 125.415 ;
        RECT 114.980 125.125 115.235 125.585 ;
        RECT 115.405 124.955 115.665 125.415 ;
        RECT 114.545 124.785 115.665 124.955 ;
        RECT 115.835 124.785 116.145 125.585 ;
        RECT 114.545 124.535 114.805 124.785 ;
        RECT 116.315 124.615 116.625 125.415 ;
        RECT 116.805 124.865 117.135 125.585 ;
        RECT 110.755 124.025 111.895 124.195 ;
        RECT 112.065 123.855 112.470 124.365 ;
        RECT 110.820 123.685 112.470 123.855 ;
        RECT 112.655 123.785 113.175 124.325 ;
        RECT 113.345 123.955 113.865 124.495 ;
        RECT 114.050 124.365 114.805 124.535 ;
        RECT 115.595 124.445 116.625 124.615 ;
        RECT 114.050 123.855 114.455 124.365 ;
        RECT 115.595 124.195 115.765 124.445 ;
        RECT 114.625 124.025 115.765 124.195 ;
        RECT 109.895 123.205 110.195 123.535 ;
        RECT 110.365 123.035 110.640 123.515 ;
        RECT 110.820 123.295 111.115 123.685 ;
        RECT 111.285 123.035 111.540 123.515 ;
        RECT 111.715 123.295 111.975 123.685 ;
        RECT 112.145 123.035 112.425 123.515 ;
        RECT 112.655 123.035 113.865 123.785 ;
        RECT 114.050 123.685 115.700 123.855 ;
        RECT 115.935 123.705 116.285 124.275 ;
        RECT 114.095 123.035 114.375 123.515 ;
        RECT 114.545 123.295 114.805 123.685 ;
        RECT 114.980 123.035 115.235 123.515 ;
        RECT 115.405 123.295 115.700 123.685 ;
        RECT 116.455 123.535 116.625 124.445 ;
        RECT 116.795 124.225 117.025 124.565 ;
        RECT 117.315 124.225 117.530 125.340 ;
        RECT 117.725 124.640 118.055 125.415 ;
        RECT 118.225 124.810 118.935 125.585 ;
        RECT 117.725 124.425 118.875 124.640 ;
        RECT 116.795 124.025 117.125 124.225 ;
        RECT 117.315 124.045 117.765 124.225 ;
        RECT 117.435 124.025 117.765 124.045 ;
        RECT 117.935 124.025 118.405 124.255 ;
        RECT 118.590 123.855 118.875 124.425 ;
        RECT 119.105 123.980 119.385 125.415 ;
        RECT 115.880 123.035 116.155 123.515 ;
        RECT 116.325 123.205 116.625 123.535 ;
        RECT 116.795 123.665 117.975 123.855 ;
        RECT 116.795 123.205 117.135 123.665 ;
        RECT 117.645 123.585 117.975 123.665 ;
        RECT 118.165 123.665 118.875 123.855 ;
        RECT 118.165 123.525 118.465 123.665 ;
        RECT 118.150 123.515 118.465 123.525 ;
        RECT 118.140 123.505 118.465 123.515 ;
        RECT 118.130 123.500 118.465 123.505 ;
        RECT 117.305 123.035 117.475 123.495 ;
        RECT 118.125 123.490 118.465 123.500 ;
        RECT 118.120 123.485 118.465 123.490 ;
        RECT 118.115 123.475 118.465 123.485 ;
        RECT 118.110 123.470 118.465 123.475 ;
        RECT 118.105 123.205 118.465 123.470 ;
        RECT 118.705 123.035 118.875 123.495 ;
        RECT 119.045 123.205 119.385 123.980 ;
        RECT 119.555 124.615 119.865 125.415 ;
        RECT 120.035 124.785 120.345 125.585 ;
        RECT 120.515 124.955 120.775 125.415 ;
        RECT 120.945 125.125 121.200 125.585 ;
        RECT 121.375 124.955 121.635 125.415 ;
        RECT 120.515 124.785 121.635 124.955 ;
        RECT 119.555 124.445 120.585 124.615 ;
        RECT 119.555 123.535 119.725 124.445 ;
        RECT 119.895 123.705 120.245 124.275 ;
        RECT 120.415 124.195 120.585 124.445 ;
        RECT 121.375 124.535 121.635 124.785 ;
        RECT 121.805 124.715 122.090 125.585 ;
        RECT 121.375 124.365 122.130 124.535 ;
        RECT 122.315 124.420 122.605 125.585 ;
        RECT 122.785 124.865 123.115 125.585 ;
        RECT 120.415 124.025 121.555 124.195 ;
        RECT 121.725 123.855 122.130 124.365 ;
        RECT 122.775 124.225 123.005 124.565 ;
        RECT 123.295 124.225 123.510 125.340 ;
        RECT 123.705 124.640 124.035 125.415 ;
        RECT 124.205 124.810 124.915 125.585 ;
        RECT 123.705 124.425 124.855 124.640 ;
        RECT 122.775 124.025 123.105 124.225 ;
        RECT 123.295 124.045 123.745 124.225 ;
        RECT 123.415 124.025 123.745 124.045 ;
        RECT 123.915 124.025 124.385 124.255 ;
        RECT 124.570 123.855 124.855 124.425 ;
        RECT 125.085 123.980 125.365 125.415 ;
        RECT 120.480 123.685 122.130 123.855 ;
        RECT 119.555 123.205 119.855 123.535 ;
        RECT 120.025 123.035 120.300 123.515 ;
        RECT 120.480 123.295 120.775 123.685 ;
        RECT 120.945 123.035 121.200 123.515 ;
        RECT 121.375 123.295 121.635 123.685 ;
        RECT 121.805 123.035 122.085 123.515 ;
        RECT 122.315 123.035 122.605 123.760 ;
        RECT 122.775 123.665 123.955 123.855 ;
        RECT 122.775 123.205 123.115 123.665 ;
        RECT 123.625 123.585 123.955 123.665 ;
        RECT 124.145 123.665 124.855 123.855 ;
        RECT 124.145 123.525 124.445 123.665 ;
        RECT 124.130 123.515 124.445 123.525 ;
        RECT 124.120 123.505 124.445 123.515 ;
        RECT 124.110 123.500 124.445 123.505 ;
        RECT 123.285 123.035 123.455 123.495 ;
        RECT 124.105 123.490 124.445 123.500 ;
        RECT 124.100 123.485 124.445 123.490 ;
        RECT 124.095 123.475 124.445 123.485 ;
        RECT 124.090 123.470 124.445 123.475 ;
        RECT 124.085 123.205 124.445 123.470 ;
        RECT 124.685 123.035 124.855 123.495 ;
        RECT 125.025 123.205 125.365 123.980 ;
        RECT 125.995 124.865 126.455 125.415 ;
        RECT 126.645 124.865 126.975 125.585 ;
        RECT 125.995 123.495 126.245 124.865 ;
        RECT 127.175 124.695 127.475 125.245 ;
        RECT 127.645 124.915 127.925 125.585 ;
        RECT 128.350 124.715 128.635 125.585 ;
        RECT 128.805 124.955 129.065 125.415 ;
        RECT 129.240 125.125 129.495 125.585 ;
        RECT 129.665 124.955 129.925 125.415 ;
        RECT 128.805 124.785 129.925 124.955 ;
        RECT 130.095 124.785 130.405 125.585 ;
        RECT 126.535 124.525 127.475 124.695 ;
        RECT 126.535 124.275 126.705 124.525 ;
        RECT 127.845 124.275 128.110 124.635 ;
        RECT 128.805 124.535 129.065 124.785 ;
        RECT 130.575 124.615 130.885 125.415 ;
        RECT 126.415 123.945 126.705 124.275 ;
        RECT 126.875 124.025 127.215 124.275 ;
        RECT 127.435 124.025 128.110 124.275 ;
        RECT 128.310 124.365 129.065 124.535 ;
        RECT 129.855 124.445 130.885 124.615 ;
        RECT 126.535 123.855 126.705 123.945 ;
        RECT 128.310 123.855 128.715 124.365 ;
        RECT 129.855 124.195 130.025 124.445 ;
        RECT 128.885 124.025 130.025 124.195 ;
        RECT 126.535 123.665 127.925 123.855 ;
        RECT 128.310 123.685 129.960 123.855 ;
        RECT 130.195 123.705 130.545 124.275 ;
        RECT 125.995 123.205 126.555 123.495 ;
        RECT 126.725 123.035 126.975 123.495 ;
        RECT 127.595 123.305 127.925 123.665 ;
        RECT 128.355 123.035 128.635 123.515 ;
        RECT 128.805 123.295 129.065 123.685 ;
        RECT 129.240 123.035 129.495 123.515 ;
        RECT 129.665 123.295 129.960 123.685 ;
        RECT 130.715 123.535 130.885 124.445 ;
        RECT 130.140 123.035 130.415 123.515 ;
        RECT 130.585 123.205 130.885 123.535 ;
        RECT 131.515 123.980 131.795 125.415 ;
        RECT 131.965 124.810 132.675 125.585 ;
        RECT 132.845 124.640 133.175 125.415 ;
        RECT 132.025 124.425 133.175 124.640 ;
        RECT 131.515 123.205 131.855 123.980 ;
        RECT 132.025 123.855 132.310 124.425 ;
        RECT 132.495 124.025 132.965 124.255 ;
        RECT 133.370 124.225 133.585 125.340 ;
        RECT 133.765 124.865 134.095 125.585 ;
        RECT 133.875 124.225 134.105 124.565 ;
        RECT 135.195 124.420 135.485 125.585 ;
        RECT 135.655 124.615 135.965 125.415 ;
        RECT 136.135 124.785 136.445 125.585 ;
        RECT 136.615 124.955 136.875 125.415 ;
        RECT 137.045 125.125 137.300 125.585 ;
        RECT 137.475 124.955 137.735 125.415 ;
        RECT 136.615 124.785 137.735 124.955 ;
        RECT 135.655 124.445 136.685 124.615 ;
        RECT 133.135 124.045 133.585 124.225 ;
        RECT 133.135 124.025 133.465 124.045 ;
        RECT 133.775 124.025 134.105 124.225 ;
        RECT 132.025 123.665 132.735 123.855 ;
        RECT 132.435 123.525 132.735 123.665 ;
        RECT 132.925 123.665 134.105 123.855 ;
        RECT 132.925 123.585 133.255 123.665 ;
        RECT 132.435 123.515 132.750 123.525 ;
        RECT 132.435 123.505 132.760 123.515 ;
        RECT 132.435 123.500 132.770 123.505 ;
        RECT 132.025 123.035 132.195 123.495 ;
        RECT 132.435 123.490 132.775 123.500 ;
        RECT 132.435 123.485 132.780 123.490 ;
        RECT 132.435 123.475 132.785 123.485 ;
        RECT 132.435 123.470 132.790 123.475 ;
        RECT 132.435 123.205 132.795 123.470 ;
        RECT 133.425 123.035 133.595 123.495 ;
        RECT 133.765 123.205 134.105 123.665 ;
        RECT 135.195 123.035 135.485 123.760 ;
        RECT 135.655 123.535 135.825 124.445 ;
        RECT 135.995 123.705 136.345 124.275 ;
        RECT 136.515 124.195 136.685 124.445 ;
        RECT 137.475 124.535 137.735 124.785 ;
        RECT 137.905 124.715 138.190 125.585 ;
        RECT 139.345 124.865 139.675 125.585 ;
        RECT 137.475 124.365 138.230 124.535 ;
        RECT 136.515 124.025 137.655 124.195 ;
        RECT 137.825 123.855 138.230 124.365 ;
        RECT 139.335 124.225 139.565 124.565 ;
        RECT 139.855 124.225 140.070 125.340 ;
        RECT 140.265 124.640 140.595 125.415 ;
        RECT 140.765 124.810 141.475 125.585 ;
        RECT 140.265 124.425 141.415 124.640 ;
        RECT 139.335 124.025 139.665 124.225 ;
        RECT 139.855 124.045 140.305 124.225 ;
        RECT 139.975 124.025 140.305 124.045 ;
        RECT 140.475 124.025 140.945 124.255 ;
        RECT 141.130 123.855 141.415 124.425 ;
        RECT 141.645 123.980 141.925 125.415 ;
        RECT 142.105 124.865 142.435 125.585 ;
        RECT 142.095 124.225 142.325 124.565 ;
        RECT 142.615 124.225 142.830 125.340 ;
        RECT 143.025 124.640 143.355 125.415 ;
        RECT 143.525 124.810 144.235 125.585 ;
        RECT 143.025 124.425 144.175 124.640 ;
        RECT 142.095 124.025 142.425 124.225 ;
        RECT 142.615 124.045 143.065 124.225 ;
        RECT 142.735 124.025 143.065 124.045 ;
        RECT 143.235 124.025 143.705 124.255 ;
        RECT 136.580 123.685 138.230 123.855 ;
        RECT 135.655 123.205 135.955 123.535 ;
        RECT 136.125 123.035 136.400 123.515 ;
        RECT 136.580 123.295 136.875 123.685 ;
        RECT 137.045 123.035 137.300 123.515 ;
        RECT 137.475 123.295 137.735 123.685 ;
        RECT 139.335 123.665 140.515 123.855 ;
        RECT 137.905 123.035 138.185 123.515 ;
        RECT 139.335 123.205 139.675 123.665 ;
        RECT 140.185 123.585 140.515 123.665 ;
        RECT 140.705 123.665 141.415 123.855 ;
        RECT 140.705 123.525 141.005 123.665 ;
        RECT 140.690 123.515 141.005 123.525 ;
        RECT 140.680 123.505 141.005 123.515 ;
        RECT 140.670 123.500 141.005 123.505 ;
        RECT 139.845 123.035 140.015 123.495 ;
        RECT 140.665 123.490 141.005 123.500 ;
        RECT 140.660 123.485 141.005 123.490 ;
        RECT 140.655 123.475 141.005 123.485 ;
        RECT 140.650 123.470 141.005 123.475 ;
        RECT 140.645 123.205 141.005 123.470 ;
        RECT 141.245 123.035 141.415 123.495 ;
        RECT 141.585 123.205 141.925 123.980 ;
        RECT 143.890 123.855 144.175 124.425 ;
        RECT 144.405 123.980 144.685 125.415 ;
        RECT 142.095 123.665 143.275 123.855 ;
        RECT 142.095 123.205 142.435 123.665 ;
        RECT 142.945 123.585 143.275 123.665 ;
        RECT 143.465 123.665 144.175 123.855 ;
        RECT 143.465 123.525 143.765 123.665 ;
        RECT 143.450 123.515 143.765 123.525 ;
        RECT 143.440 123.505 143.765 123.515 ;
        RECT 143.430 123.500 143.765 123.505 ;
        RECT 142.605 123.035 142.775 123.495 ;
        RECT 143.425 123.490 143.765 123.500 ;
        RECT 143.420 123.485 143.765 123.490 ;
        RECT 143.415 123.475 143.765 123.485 ;
        RECT 143.410 123.470 143.765 123.475 ;
        RECT 143.405 123.205 143.765 123.470 ;
        RECT 144.005 123.035 144.175 123.495 ;
        RECT 144.345 123.205 144.685 123.980 ;
        RECT 144.855 124.615 145.165 125.415 ;
        RECT 145.335 124.785 145.645 125.585 ;
        RECT 145.815 124.955 146.075 125.415 ;
        RECT 146.245 125.125 146.500 125.585 ;
        RECT 146.675 124.955 146.935 125.415 ;
        RECT 145.815 124.785 146.935 124.955 ;
        RECT 144.855 124.445 145.885 124.615 ;
        RECT 144.855 123.535 145.025 124.445 ;
        RECT 145.195 123.705 145.545 124.275 ;
        RECT 145.715 124.195 145.885 124.445 ;
        RECT 146.675 124.535 146.935 124.785 ;
        RECT 147.105 124.715 147.390 125.585 ;
        RECT 146.675 124.365 147.430 124.535 ;
        RECT 148.075 124.420 148.365 125.585 ;
        RECT 148.535 124.615 148.845 125.415 ;
        RECT 149.015 124.785 149.325 125.585 ;
        RECT 149.495 124.955 149.755 125.415 ;
        RECT 149.925 125.125 150.180 125.585 ;
        RECT 150.355 124.955 150.615 125.415 ;
        RECT 149.495 124.785 150.615 124.955 ;
        RECT 148.535 124.445 149.565 124.615 ;
        RECT 145.715 124.025 146.855 124.195 ;
        RECT 147.025 123.855 147.430 124.365 ;
        RECT 145.780 123.685 147.430 123.855 ;
        RECT 144.855 123.205 145.155 123.535 ;
        RECT 145.325 123.035 145.600 123.515 ;
        RECT 145.780 123.295 146.075 123.685 ;
        RECT 146.245 123.035 146.500 123.515 ;
        RECT 146.675 123.295 146.935 123.685 ;
        RECT 147.105 123.035 147.385 123.515 ;
        RECT 148.075 123.035 148.365 123.760 ;
        RECT 148.535 123.535 148.705 124.445 ;
        RECT 148.875 123.705 149.225 124.275 ;
        RECT 149.395 124.195 149.565 124.445 ;
        RECT 150.355 124.535 150.615 124.785 ;
        RECT 150.785 124.715 151.070 125.585 ;
        RECT 151.495 124.915 151.775 125.585 ;
        RECT 151.945 124.695 152.245 125.245 ;
        RECT 152.445 124.865 152.775 125.585 ;
        RECT 152.965 124.865 153.425 125.415 ;
        RECT 150.355 124.365 151.110 124.535 ;
        RECT 149.395 124.025 150.535 124.195 ;
        RECT 150.705 123.855 151.110 124.365 ;
        RECT 151.310 124.275 151.575 124.635 ;
        RECT 151.945 124.525 152.885 124.695 ;
        RECT 152.715 124.275 152.885 124.525 ;
        RECT 151.310 124.025 151.985 124.275 ;
        RECT 152.205 124.025 152.545 124.275 ;
        RECT 152.715 123.945 153.005 124.275 ;
        RECT 152.715 123.855 152.885 123.945 ;
        RECT 149.460 123.685 151.110 123.855 ;
        RECT 148.535 123.205 148.835 123.535 ;
        RECT 149.005 123.035 149.280 123.515 ;
        RECT 149.460 123.295 149.755 123.685 ;
        RECT 149.925 123.035 150.180 123.515 ;
        RECT 150.355 123.295 150.615 123.685 ;
        RECT 151.495 123.665 152.885 123.855 ;
        RECT 150.785 123.035 151.065 123.515 ;
        RECT 151.495 123.305 151.825 123.665 ;
        RECT 153.175 123.495 153.425 124.865 ;
        RECT 153.595 124.495 154.805 125.585 ;
        RECT 152.445 123.035 152.695 123.495 ;
        RECT 152.865 123.205 153.425 123.495 ;
        RECT 153.595 123.785 154.115 124.325 ;
        RECT 154.285 123.955 154.805 124.495 ;
        RECT 154.975 124.495 156.185 125.585 ;
        RECT 154.975 123.955 155.495 124.495 ;
        RECT 155.665 123.785 156.185 124.325 ;
        RECT 153.595 123.035 154.805 123.785 ;
        RECT 154.975 123.035 156.185 123.785 ;
        RECT 70.710 122.865 156.270 123.035 ;
        RECT 51.110 103.480 53.100 103.650 ;
        RECT 51.110 79.970 51.280 103.480 ;
        RECT 51.760 100.840 52.450 103.000 ;
        RECT 52.930 79.970 53.100 103.480 ;
        RECT 55.110 103.480 57.100 103.650 ;
        RECT 55.110 79.970 55.280 103.480 ;
        RECT 55.760 100.840 56.450 103.000 ;
        RECT 56.930 79.970 57.100 103.480 ;
        RECT 59.110 103.480 61.100 103.650 ;
        RECT 59.110 79.970 59.280 103.480 ;
        RECT 59.760 100.840 60.450 103.000 ;
        RECT 60.930 79.970 61.100 103.480 ;
        RECT 63.110 103.480 65.100 103.650 ;
        RECT 63.110 79.970 63.280 103.480 ;
        RECT 63.760 100.840 64.450 103.000 ;
        RECT 64.930 79.970 65.100 103.480 ;
        RECT 67.110 103.480 69.100 103.650 ;
        RECT 67.110 79.970 67.280 103.480 ;
        RECT 67.760 100.840 68.450 103.000 ;
        RECT 68.930 79.970 69.100 103.480 ;
        RECT 71.110 103.480 73.100 103.650 ;
        RECT 71.110 79.970 71.280 103.480 ;
        RECT 71.760 100.840 72.450 103.000 ;
        RECT 72.930 79.970 73.100 103.480 ;
        RECT 75.110 103.480 77.100 103.650 ;
        RECT 75.110 79.970 75.280 103.480 ;
        RECT 75.760 100.840 76.450 103.000 ;
        RECT 76.930 79.970 77.100 103.480 ;
        RECT 79.110 103.480 81.100 103.650 ;
        RECT 79.110 79.970 79.280 103.480 ;
        RECT 79.760 100.840 80.450 103.000 ;
        RECT 80.930 79.970 81.100 103.480 ;
        RECT 88.110 103.480 90.100 103.650 ;
        RECT 88.110 79.970 88.280 103.480 ;
        RECT 88.760 100.840 89.450 103.000 ;
        RECT 89.930 79.970 90.100 103.480 ;
        RECT 92.110 103.480 94.100 103.650 ;
        RECT 92.110 79.970 92.280 103.480 ;
        RECT 92.760 100.840 93.450 103.000 ;
        RECT 93.930 79.970 94.100 103.480 ;
        RECT 96.110 103.480 98.100 103.650 ;
        RECT 96.110 79.970 96.280 103.480 ;
        RECT 96.760 100.840 97.450 103.000 ;
        RECT 97.930 79.970 98.100 103.480 ;
        RECT 100.110 103.480 102.100 103.650 ;
        RECT 100.110 79.970 100.280 103.480 ;
        RECT 100.760 100.840 101.450 103.000 ;
        RECT 101.930 79.970 102.100 103.480 ;
        RECT 104.110 103.480 106.100 103.650 ;
        RECT 104.110 79.970 104.280 103.480 ;
        RECT 104.760 100.840 105.450 103.000 ;
        RECT 105.930 79.970 106.100 103.480 ;
        RECT 108.110 103.480 110.100 103.650 ;
        RECT 108.110 79.970 108.280 103.480 ;
        RECT 108.760 100.840 109.450 103.000 ;
        RECT 109.930 79.970 110.100 103.480 ;
        RECT 112.110 103.480 114.100 103.650 ;
        RECT 112.110 79.970 112.280 103.480 ;
        RECT 112.760 100.840 113.450 103.000 ;
        RECT 113.930 79.970 114.100 103.480 ;
        RECT 116.110 103.480 118.100 103.650 ;
        RECT 116.110 79.970 116.280 103.480 ;
        RECT 116.760 100.840 117.450 103.000 ;
        RECT 117.930 79.970 118.100 103.480 ;
        RECT 125.110 103.480 127.100 103.650 ;
        RECT 125.110 79.970 125.280 103.480 ;
        RECT 125.760 100.840 126.450 103.000 ;
        RECT 126.930 79.970 127.100 103.480 ;
        RECT 129.110 103.480 131.100 103.650 ;
        RECT 129.110 79.970 129.280 103.480 ;
        RECT 129.760 100.840 130.450 103.000 ;
        RECT 130.930 79.970 131.100 103.480 ;
        RECT 133.110 103.480 135.100 103.650 ;
        RECT 133.110 79.970 133.280 103.480 ;
        RECT 133.760 100.840 134.450 103.000 ;
        RECT 134.930 79.970 135.100 103.480 ;
        RECT 137.110 103.480 139.100 103.650 ;
        RECT 137.110 79.970 137.280 103.480 ;
        RECT 137.760 100.840 138.450 103.000 ;
        RECT 138.930 79.970 139.100 103.480 ;
        RECT 141.110 103.480 143.100 103.650 ;
        RECT 141.110 79.970 141.280 103.480 ;
        RECT 141.760 100.840 142.450 103.000 ;
        RECT 142.930 79.970 143.100 103.480 ;
        RECT 145.110 103.480 147.100 103.650 ;
        RECT 145.110 79.970 145.280 103.480 ;
        RECT 145.760 100.840 146.450 103.000 ;
        RECT 146.930 79.970 147.100 103.480 ;
        RECT 149.110 103.480 151.100 103.650 ;
        RECT 149.110 79.970 149.280 103.480 ;
        RECT 149.760 100.840 150.450 103.000 ;
        RECT 150.930 79.970 151.100 103.480 ;
        RECT 153.110 103.480 155.100 103.650 ;
        RECT 153.110 79.970 153.280 103.480 ;
        RECT 153.760 100.840 154.450 103.000 ;
        RECT 154.930 79.970 155.100 103.480 ;
        RECT 51.030 79.170 51.370 79.970 ;
        RECT 52.830 79.170 53.170 79.970 ;
        RECT 55.030 79.170 55.370 79.970 ;
        RECT 56.830 79.170 57.170 79.970 ;
        RECT 59.030 79.170 59.370 79.970 ;
        RECT 60.830 79.170 61.170 79.970 ;
        RECT 63.030 79.170 63.370 79.970 ;
        RECT 64.830 79.170 65.170 79.970 ;
        RECT 67.030 79.170 67.370 79.970 ;
        RECT 68.830 79.170 69.170 79.970 ;
        RECT 71.030 79.170 71.370 79.970 ;
        RECT 72.830 79.170 73.170 79.970 ;
        RECT 75.030 79.170 75.370 79.970 ;
        RECT 76.830 79.170 77.170 79.970 ;
        RECT 79.030 79.170 79.370 79.970 ;
        RECT 80.830 79.170 81.170 79.970 ;
        RECT 88.030 79.170 88.370 79.970 ;
        RECT 89.830 79.170 90.170 79.970 ;
        RECT 92.030 79.170 92.370 79.970 ;
        RECT 93.830 79.170 94.170 79.970 ;
        RECT 96.030 79.170 96.370 79.970 ;
        RECT 97.830 79.170 98.170 79.970 ;
        RECT 100.030 79.170 100.370 79.970 ;
        RECT 101.830 79.170 102.170 79.970 ;
        RECT 104.030 79.170 104.370 79.970 ;
        RECT 105.830 79.170 106.170 79.970 ;
        RECT 108.030 79.170 108.370 79.970 ;
        RECT 109.830 79.170 110.170 79.970 ;
        RECT 112.030 79.170 112.370 79.970 ;
        RECT 113.830 79.170 114.170 79.970 ;
        RECT 116.030 79.170 116.370 79.970 ;
        RECT 117.830 79.170 118.170 79.970 ;
        RECT 125.030 79.170 125.370 79.970 ;
        RECT 126.830 79.170 127.170 79.970 ;
        RECT 129.030 79.170 129.370 79.970 ;
        RECT 130.830 79.170 131.170 79.970 ;
        RECT 133.030 79.170 133.370 79.970 ;
        RECT 134.830 79.170 135.170 79.970 ;
        RECT 137.030 79.170 137.370 79.970 ;
        RECT 138.830 79.170 139.170 79.970 ;
        RECT 141.030 79.170 141.370 79.970 ;
        RECT 142.830 79.170 143.170 79.970 ;
        RECT 145.030 79.170 145.370 79.970 ;
        RECT 146.830 79.170 147.170 79.970 ;
        RECT 149.030 79.170 149.370 79.970 ;
        RECT 150.830 79.170 151.170 79.970 ;
        RECT 153.030 79.170 153.370 79.970 ;
        RECT 154.830 79.170 155.170 79.970 ;
        RECT 51.110 58.460 51.280 79.170 ;
        RECT 51.760 58.940 52.450 61.100 ;
        RECT 52.930 58.460 53.100 79.170 ;
        RECT 51.110 58.290 53.100 58.460 ;
        RECT 55.110 58.460 55.280 79.170 ;
        RECT 55.760 58.940 56.450 61.100 ;
        RECT 56.930 58.460 57.100 79.170 ;
        RECT 55.110 58.290 57.100 58.460 ;
        RECT 59.110 58.460 59.280 79.170 ;
        RECT 59.760 58.940 60.450 61.100 ;
        RECT 60.930 58.460 61.100 79.170 ;
        RECT 59.110 58.290 61.100 58.460 ;
        RECT 63.110 58.460 63.280 79.170 ;
        RECT 63.760 58.940 64.450 61.100 ;
        RECT 64.930 58.460 65.100 79.170 ;
        RECT 63.110 58.290 65.100 58.460 ;
        RECT 67.110 58.460 67.280 79.170 ;
        RECT 67.760 58.940 68.450 61.100 ;
        RECT 68.930 58.460 69.100 79.170 ;
        RECT 67.110 58.290 69.100 58.460 ;
        RECT 71.110 58.460 71.280 79.170 ;
        RECT 71.760 58.940 72.450 61.100 ;
        RECT 72.930 58.460 73.100 79.170 ;
        RECT 71.110 58.290 73.100 58.460 ;
        RECT 75.110 58.460 75.280 79.170 ;
        RECT 75.760 58.940 76.450 61.100 ;
        RECT 76.930 58.460 77.100 79.170 ;
        RECT 75.110 58.290 77.100 58.460 ;
        RECT 79.110 58.460 79.280 79.170 ;
        RECT 79.760 58.940 80.450 61.100 ;
        RECT 80.930 58.460 81.100 79.170 ;
        RECT 79.110 58.290 81.100 58.460 ;
        RECT 88.110 58.460 88.280 79.170 ;
        RECT 88.760 58.940 89.450 61.100 ;
        RECT 89.930 58.460 90.100 79.170 ;
        RECT 88.110 58.290 90.100 58.460 ;
        RECT 92.110 58.460 92.280 79.170 ;
        RECT 92.760 58.940 93.450 61.100 ;
        RECT 93.930 58.460 94.100 79.170 ;
        RECT 92.110 58.290 94.100 58.460 ;
        RECT 96.110 58.460 96.280 79.170 ;
        RECT 96.760 58.940 97.450 61.100 ;
        RECT 97.930 58.460 98.100 79.170 ;
        RECT 96.110 58.290 98.100 58.460 ;
        RECT 100.110 58.460 100.280 79.170 ;
        RECT 100.760 58.940 101.450 61.100 ;
        RECT 101.930 58.460 102.100 79.170 ;
        RECT 100.110 58.290 102.100 58.460 ;
        RECT 104.110 58.460 104.280 79.170 ;
        RECT 104.760 58.940 105.450 61.100 ;
        RECT 105.930 58.460 106.100 79.170 ;
        RECT 104.110 58.290 106.100 58.460 ;
        RECT 108.110 58.460 108.280 79.170 ;
        RECT 108.760 58.940 109.450 61.100 ;
        RECT 109.930 58.460 110.100 79.170 ;
        RECT 108.110 58.290 110.100 58.460 ;
        RECT 112.110 58.460 112.280 79.170 ;
        RECT 112.760 58.940 113.450 61.100 ;
        RECT 113.930 58.460 114.100 79.170 ;
        RECT 112.110 58.290 114.100 58.460 ;
        RECT 116.110 58.460 116.280 79.170 ;
        RECT 116.760 58.940 117.450 61.100 ;
        RECT 117.930 58.460 118.100 79.170 ;
        RECT 116.110 58.290 118.100 58.460 ;
        RECT 125.110 58.460 125.280 79.170 ;
        RECT 125.760 58.940 126.450 61.100 ;
        RECT 126.930 58.460 127.100 79.170 ;
        RECT 125.110 58.290 127.100 58.460 ;
        RECT 129.110 58.460 129.280 79.170 ;
        RECT 129.760 58.940 130.450 61.100 ;
        RECT 130.930 58.460 131.100 79.170 ;
        RECT 129.110 58.290 131.100 58.460 ;
        RECT 133.110 58.460 133.280 79.170 ;
        RECT 133.760 58.940 134.450 61.100 ;
        RECT 134.930 58.460 135.100 79.170 ;
        RECT 133.110 58.290 135.100 58.460 ;
        RECT 137.110 58.460 137.280 79.170 ;
        RECT 137.760 58.940 138.450 61.100 ;
        RECT 138.930 58.460 139.100 79.170 ;
        RECT 137.110 58.290 139.100 58.460 ;
        RECT 141.110 58.460 141.280 79.170 ;
        RECT 141.760 58.940 142.450 61.100 ;
        RECT 142.930 58.460 143.100 79.170 ;
        RECT 141.110 58.290 143.100 58.460 ;
        RECT 145.110 58.460 145.280 79.170 ;
        RECT 145.760 58.940 146.450 61.100 ;
        RECT 146.930 58.460 147.100 79.170 ;
        RECT 145.110 58.290 147.100 58.460 ;
        RECT 149.110 58.460 149.280 79.170 ;
        RECT 149.760 58.940 150.450 61.100 ;
        RECT 150.930 58.460 151.100 79.170 ;
        RECT 149.110 58.290 151.100 58.460 ;
        RECT 153.110 58.460 153.280 79.170 ;
        RECT 153.760 58.940 154.450 61.100 ;
        RECT 154.930 58.460 155.100 79.170 ;
        RECT 153.110 58.290 155.100 58.460 ;
        RECT 51.110 55.480 53.100 55.650 ;
        RECT 51.110 30.810 51.280 55.480 ;
        RECT 51.760 52.840 52.450 55.000 ;
        RECT 51.760 31.290 52.450 33.450 ;
        RECT 51.480 30.810 52.740 30.900 ;
        RECT 52.930 30.810 53.100 55.480 ;
        RECT 51.110 30.640 53.100 30.810 ;
        RECT 55.110 55.480 57.100 55.650 ;
        RECT 55.110 30.810 55.280 55.480 ;
        RECT 55.760 52.840 56.450 55.000 ;
        RECT 55.760 31.290 56.450 33.450 ;
        RECT 55.480 30.810 56.740 30.900 ;
        RECT 56.930 30.810 57.100 55.480 ;
        RECT 55.110 30.640 57.100 30.810 ;
        RECT 59.110 55.480 61.100 55.650 ;
        RECT 59.110 30.810 59.280 55.480 ;
        RECT 59.760 52.840 60.450 55.000 ;
        RECT 59.760 31.290 60.450 33.450 ;
        RECT 59.480 30.810 60.740 30.900 ;
        RECT 60.930 30.810 61.100 55.480 ;
        RECT 59.110 30.640 61.100 30.810 ;
        RECT 63.110 55.480 65.100 55.650 ;
        RECT 63.110 30.810 63.280 55.480 ;
        RECT 63.760 52.840 64.450 55.000 ;
        RECT 63.760 31.290 64.450 33.450 ;
        RECT 63.480 30.810 64.740 30.900 ;
        RECT 64.930 30.810 65.100 55.480 ;
        RECT 63.110 30.640 65.100 30.810 ;
        RECT 67.110 55.480 69.100 55.650 ;
        RECT 67.110 30.810 67.280 55.480 ;
        RECT 67.760 52.840 68.450 55.000 ;
        RECT 67.760 31.290 68.450 33.450 ;
        RECT 67.480 30.810 68.740 30.900 ;
        RECT 68.930 30.810 69.100 55.480 ;
        RECT 67.110 30.640 69.100 30.810 ;
        RECT 71.110 55.480 73.100 55.650 ;
        RECT 71.110 30.810 71.280 55.480 ;
        RECT 71.760 52.840 72.450 55.000 ;
        RECT 71.760 31.290 72.450 33.450 ;
        RECT 71.480 30.810 72.740 30.900 ;
        RECT 72.930 30.810 73.100 55.480 ;
        RECT 71.110 30.640 73.100 30.810 ;
        RECT 75.110 55.480 77.100 55.650 ;
        RECT 75.110 30.810 75.280 55.480 ;
        RECT 75.760 52.840 76.450 55.000 ;
        RECT 75.760 31.290 76.450 33.450 ;
        RECT 75.480 30.810 76.740 30.900 ;
        RECT 76.930 30.810 77.100 55.480 ;
        RECT 75.110 30.640 77.100 30.810 ;
        RECT 79.110 55.480 81.100 55.650 ;
        RECT 79.110 30.810 79.280 55.480 ;
        RECT 79.760 52.840 80.450 55.000 ;
        RECT 79.760 31.290 80.450 33.450 ;
        RECT 79.480 30.810 80.740 30.900 ;
        RECT 80.930 30.810 81.100 55.480 ;
        RECT 79.110 30.640 81.100 30.810 ;
        RECT 88.110 55.480 90.100 55.650 ;
        RECT 88.110 30.810 88.280 55.480 ;
        RECT 88.760 52.840 89.450 55.000 ;
        RECT 88.760 31.290 89.450 33.450 ;
        RECT 88.480 30.810 89.740 30.900 ;
        RECT 89.930 30.810 90.100 55.480 ;
        RECT 88.110 30.640 90.100 30.810 ;
        RECT 92.110 55.480 94.100 55.650 ;
        RECT 92.110 30.810 92.280 55.480 ;
        RECT 92.760 52.840 93.450 55.000 ;
        RECT 92.760 31.290 93.450 33.450 ;
        RECT 92.480 30.810 93.740 30.900 ;
        RECT 93.930 30.810 94.100 55.480 ;
        RECT 92.110 30.640 94.100 30.810 ;
        RECT 96.110 55.480 98.100 55.650 ;
        RECT 96.110 30.810 96.280 55.480 ;
        RECT 96.760 52.840 97.450 55.000 ;
        RECT 96.760 31.290 97.450 33.450 ;
        RECT 96.480 30.810 97.740 30.900 ;
        RECT 97.930 30.810 98.100 55.480 ;
        RECT 96.110 30.640 98.100 30.810 ;
        RECT 100.110 55.480 102.100 55.650 ;
        RECT 100.110 30.810 100.280 55.480 ;
        RECT 100.760 52.840 101.450 55.000 ;
        RECT 100.760 31.290 101.450 33.450 ;
        RECT 100.480 30.810 101.740 30.900 ;
        RECT 101.930 30.810 102.100 55.480 ;
        RECT 100.110 30.640 102.100 30.810 ;
        RECT 104.110 55.480 106.100 55.650 ;
        RECT 104.110 30.810 104.280 55.480 ;
        RECT 104.760 52.840 105.450 55.000 ;
        RECT 104.760 31.290 105.450 33.450 ;
        RECT 104.480 30.810 105.740 30.900 ;
        RECT 105.930 30.810 106.100 55.480 ;
        RECT 104.110 30.640 106.100 30.810 ;
        RECT 108.110 55.480 110.100 55.650 ;
        RECT 108.110 30.810 108.280 55.480 ;
        RECT 108.760 52.840 109.450 55.000 ;
        RECT 108.760 31.290 109.450 33.450 ;
        RECT 108.480 30.810 109.740 30.900 ;
        RECT 109.930 30.810 110.100 55.480 ;
        RECT 108.110 30.640 110.100 30.810 ;
        RECT 112.110 55.480 114.100 55.650 ;
        RECT 112.110 30.810 112.280 55.480 ;
        RECT 112.760 52.840 113.450 55.000 ;
        RECT 112.760 31.290 113.450 33.450 ;
        RECT 112.480 30.810 113.740 30.900 ;
        RECT 113.930 30.810 114.100 55.480 ;
        RECT 112.110 30.640 114.100 30.810 ;
        RECT 116.110 55.480 118.100 55.650 ;
        RECT 116.110 30.810 116.280 55.480 ;
        RECT 116.760 52.840 117.450 55.000 ;
        RECT 116.760 31.290 117.450 33.450 ;
        RECT 116.480 30.810 117.740 30.900 ;
        RECT 117.930 30.810 118.100 55.480 ;
        RECT 116.110 30.640 118.100 30.810 ;
        RECT 125.110 55.480 127.100 55.650 ;
        RECT 125.110 30.810 125.280 55.480 ;
        RECT 125.760 52.840 126.450 55.000 ;
        RECT 125.760 31.290 126.450 33.450 ;
        RECT 125.480 30.810 126.740 30.900 ;
        RECT 126.930 30.810 127.100 55.480 ;
        RECT 125.110 30.640 127.100 30.810 ;
        RECT 129.110 55.480 131.100 55.650 ;
        RECT 129.110 30.810 129.280 55.480 ;
        RECT 129.760 52.840 130.450 55.000 ;
        RECT 129.760 31.290 130.450 33.450 ;
        RECT 129.480 30.810 130.740 30.900 ;
        RECT 130.930 30.810 131.100 55.480 ;
        RECT 129.110 30.640 131.100 30.810 ;
        RECT 133.110 55.480 135.100 55.650 ;
        RECT 133.110 30.810 133.280 55.480 ;
        RECT 133.760 52.840 134.450 55.000 ;
        RECT 133.760 31.290 134.450 33.450 ;
        RECT 133.480 30.810 134.740 30.900 ;
        RECT 134.930 30.810 135.100 55.480 ;
        RECT 133.110 30.640 135.100 30.810 ;
        RECT 137.110 55.480 139.100 55.650 ;
        RECT 137.110 30.810 137.280 55.480 ;
        RECT 137.760 52.840 138.450 55.000 ;
        RECT 137.760 31.290 138.450 33.450 ;
        RECT 137.480 30.810 138.740 30.900 ;
        RECT 138.930 30.810 139.100 55.480 ;
        RECT 137.110 30.640 139.100 30.810 ;
        RECT 141.110 55.480 143.100 55.650 ;
        RECT 141.110 30.810 141.280 55.480 ;
        RECT 141.760 52.840 142.450 55.000 ;
        RECT 141.760 31.290 142.450 33.450 ;
        RECT 141.480 30.810 142.740 30.900 ;
        RECT 142.930 30.810 143.100 55.480 ;
        RECT 141.110 30.640 143.100 30.810 ;
        RECT 145.110 55.480 147.100 55.650 ;
        RECT 145.110 30.810 145.280 55.480 ;
        RECT 145.760 52.840 146.450 55.000 ;
        RECT 145.760 31.290 146.450 33.450 ;
        RECT 145.480 30.810 146.740 30.900 ;
        RECT 146.930 30.810 147.100 55.480 ;
        RECT 145.110 30.640 147.100 30.810 ;
        RECT 149.110 55.480 151.100 55.650 ;
        RECT 149.110 30.810 149.280 55.480 ;
        RECT 149.760 52.840 150.450 55.000 ;
        RECT 149.760 31.290 150.450 33.450 ;
        RECT 149.480 30.810 150.740 30.900 ;
        RECT 150.930 30.810 151.100 55.480 ;
        RECT 149.110 30.640 151.100 30.810 ;
        RECT 153.110 55.480 155.100 55.650 ;
        RECT 153.110 30.810 153.280 55.480 ;
        RECT 153.760 52.840 154.450 55.000 ;
        RECT 153.760 31.290 154.450 33.450 ;
        RECT 153.480 30.810 154.740 30.900 ;
        RECT 154.930 30.810 155.100 55.480 ;
        RECT 153.110 30.640 155.100 30.810 ;
        RECT 51.480 30.540 52.740 30.640 ;
        RECT 55.480 30.540 56.740 30.640 ;
        RECT 59.480 30.540 60.740 30.640 ;
        RECT 63.480 30.540 64.740 30.640 ;
        RECT 67.480 30.540 68.740 30.640 ;
        RECT 71.480 30.540 72.740 30.640 ;
        RECT 75.480 30.540 76.740 30.640 ;
        RECT 79.480 30.540 80.740 30.640 ;
        RECT 88.480 30.540 89.740 30.640 ;
        RECT 92.480 30.540 93.740 30.640 ;
        RECT 96.480 30.540 97.740 30.640 ;
        RECT 100.480 30.540 101.740 30.640 ;
        RECT 104.480 30.540 105.740 30.640 ;
        RECT 108.480 30.540 109.740 30.640 ;
        RECT 112.480 30.540 113.740 30.640 ;
        RECT 116.480 30.540 117.740 30.640 ;
        RECT 125.480 30.540 126.740 30.640 ;
        RECT 129.480 30.540 130.740 30.640 ;
        RECT 133.480 30.540 134.740 30.640 ;
        RECT 137.480 30.540 138.740 30.640 ;
        RECT 141.480 30.540 142.740 30.640 ;
        RECT 145.480 30.540 146.740 30.640 ;
        RECT 149.480 30.540 150.740 30.640 ;
        RECT 153.480 30.540 154.740 30.640 ;
        RECT 31.285 26.620 33.035 26.790 ;
        RECT 31.285 22.445 31.455 26.620 ;
        RECT 31.995 26.110 32.325 26.280 ;
        RECT 31.220 21.745 31.520 22.445 ;
        RECT 31.285 17.130 31.455 21.745 ;
        RECT 31.855 17.855 32.025 25.895 ;
        RECT 32.295 17.855 32.465 25.895 ;
        RECT 31.995 17.470 32.325 17.640 ;
        RECT 32.865 17.130 33.035 26.620 ;
        RECT 34.100 24.595 35.850 24.765 ;
        RECT 34.100 19.195 34.270 24.595 ;
        RECT 34.810 24.085 35.140 24.255 ;
        RECT 34.670 19.875 34.840 23.915 ;
        RECT 35.110 19.875 35.280 23.915 ;
        RECT 35.680 23.645 35.850 24.595 ;
        RECT 35.620 22.845 35.920 23.645 ;
        RECT 34.810 19.535 35.140 19.705 ;
        RECT 35.680 19.195 35.850 22.845 ;
        RECT 34.100 19.025 35.850 19.195 ;
        RECT 31.285 16.960 33.035 17.130 ;
      LAYER mcon ;
        RECT 70.855 207.185 71.025 207.355 ;
        RECT 71.315 207.185 71.485 207.355 ;
        RECT 71.775 207.185 71.945 207.355 ;
        RECT 72.235 207.185 72.405 207.355 ;
        RECT 72.695 207.185 72.865 207.355 ;
        RECT 73.155 207.185 73.325 207.355 ;
        RECT 73.615 207.185 73.785 207.355 ;
        RECT 74.075 207.185 74.245 207.355 ;
        RECT 74.535 207.185 74.705 207.355 ;
        RECT 74.995 207.185 75.165 207.355 ;
        RECT 75.455 207.185 75.625 207.355 ;
        RECT 75.915 207.185 76.085 207.355 ;
        RECT 76.375 207.185 76.545 207.355 ;
        RECT 76.835 207.185 77.005 207.355 ;
        RECT 77.295 207.185 77.465 207.355 ;
        RECT 77.755 207.185 77.925 207.355 ;
        RECT 78.215 207.185 78.385 207.355 ;
        RECT 78.675 207.185 78.845 207.355 ;
        RECT 79.135 207.185 79.305 207.355 ;
        RECT 79.595 207.185 79.765 207.355 ;
        RECT 80.055 207.185 80.225 207.355 ;
        RECT 80.515 207.185 80.685 207.355 ;
        RECT 80.975 207.185 81.145 207.355 ;
        RECT 81.435 207.185 81.605 207.355 ;
        RECT 81.895 207.185 82.065 207.355 ;
        RECT 82.355 207.185 82.525 207.355 ;
        RECT 82.815 207.185 82.985 207.355 ;
        RECT 83.275 207.185 83.445 207.355 ;
        RECT 83.735 207.185 83.905 207.355 ;
        RECT 84.195 207.185 84.365 207.355 ;
        RECT 84.655 207.185 84.825 207.355 ;
        RECT 85.115 207.185 85.285 207.355 ;
        RECT 85.575 207.185 85.745 207.355 ;
        RECT 86.035 207.185 86.205 207.355 ;
        RECT 86.495 207.185 86.665 207.355 ;
        RECT 86.955 207.185 87.125 207.355 ;
        RECT 87.415 207.185 87.585 207.355 ;
        RECT 87.875 207.185 88.045 207.355 ;
        RECT 88.335 207.185 88.505 207.355 ;
        RECT 88.795 207.185 88.965 207.355 ;
        RECT 89.255 207.185 89.425 207.355 ;
        RECT 89.715 207.185 89.885 207.355 ;
        RECT 90.175 207.185 90.345 207.355 ;
        RECT 90.635 207.185 90.805 207.355 ;
        RECT 91.095 207.185 91.265 207.355 ;
        RECT 91.555 207.185 91.725 207.355 ;
        RECT 92.015 207.185 92.185 207.355 ;
        RECT 92.475 207.185 92.645 207.355 ;
        RECT 92.935 207.185 93.105 207.355 ;
        RECT 93.395 207.185 93.565 207.355 ;
        RECT 93.855 207.185 94.025 207.355 ;
        RECT 94.315 207.185 94.485 207.355 ;
        RECT 94.775 207.185 94.945 207.355 ;
        RECT 95.235 207.185 95.405 207.355 ;
        RECT 95.695 207.185 95.865 207.355 ;
        RECT 96.155 207.185 96.325 207.355 ;
        RECT 96.615 207.185 96.785 207.355 ;
        RECT 97.075 207.185 97.245 207.355 ;
        RECT 97.535 207.185 97.705 207.355 ;
        RECT 97.995 207.185 98.165 207.355 ;
        RECT 98.455 207.185 98.625 207.355 ;
        RECT 98.915 207.185 99.085 207.355 ;
        RECT 99.375 207.185 99.545 207.355 ;
        RECT 99.835 207.185 100.005 207.355 ;
        RECT 100.295 207.185 100.465 207.355 ;
        RECT 100.755 207.185 100.925 207.355 ;
        RECT 101.215 207.185 101.385 207.355 ;
        RECT 101.675 207.185 101.845 207.355 ;
        RECT 102.135 207.185 102.305 207.355 ;
        RECT 102.595 207.185 102.765 207.355 ;
        RECT 103.055 207.185 103.225 207.355 ;
        RECT 103.515 207.185 103.685 207.355 ;
        RECT 103.975 207.185 104.145 207.355 ;
        RECT 104.435 207.185 104.605 207.355 ;
        RECT 104.895 207.185 105.065 207.355 ;
        RECT 105.355 207.185 105.525 207.355 ;
        RECT 105.815 207.185 105.985 207.355 ;
        RECT 106.275 207.185 106.445 207.355 ;
        RECT 106.735 207.185 106.905 207.355 ;
        RECT 107.195 207.185 107.365 207.355 ;
        RECT 107.655 207.185 107.825 207.355 ;
        RECT 108.115 207.185 108.285 207.355 ;
        RECT 108.575 207.185 108.745 207.355 ;
        RECT 109.035 207.185 109.205 207.355 ;
        RECT 109.495 207.185 109.665 207.355 ;
        RECT 109.955 207.185 110.125 207.355 ;
        RECT 110.415 207.185 110.585 207.355 ;
        RECT 110.875 207.185 111.045 207.355 ;
        RECT 111.335 207.185 111.505 207.355 ;
        RECT 111.795 207.185 111.965 207.355 ;
        RECT 112.255 207.185 112.425 207.355 ;
        RECT 112.715 207.185 112.885 207.355 ;
        RECT 113.175 207.185 113.345 207.355 ;
        RECT 113.635 207.185 113.805 207.355 ;
        RECT 114.095 207.185 114.265 207.355 ;
        RECT 114.555 207.185 114.725 207.355 ;
        RECT 115.015 207.185 115.185 207.355 ;
        RECT 115.475 207.185 115.645 207.355 ;
        RECT 115.935 207.185 116.105 207.355 ;
        RECT 116.395 207.185 116.565 207.355 ;
        RECT 116.855 207.185 117.025 207.355 ;
        RECT 117.315 207.185 117.485 207.355 ;
        RECT 117.775 207.185 117.945 207.355 ;
        RECT 118.235 207.185 118.405 207.355 ;
        RECT 118.695 207.185 118.865 207.355 ;
        RECT 119.155 207.185 119.325 207.355 ;
        RECT 119.615 207.185 119.785 207.355 ;
        RECT 120.075 207.185 120.245 207.355 ;
        RECT 120.535 207.185 120.705 207.355 ;
        RECT 120.995 207.185 121.165 207.355 ;
        RECT 121.455 207.185 121.625 207.355 ;
        RECT 121.915 207.185 122.085 207.355 ;
        RECT 122.375 207.185 122.545 207.355 ;
        RECT 122.835 207.185 123.005 207.355 ;
        RECT 123.295 207.185 123.465 207.355 ;
        RECT 123.755 207.185 123.925 207.355 ;
        RECT 124.215 207.185 124.385 207.355 ;
        RECT 124.675 207.185 124.845 207.355 ;
        RECT 125.135 207.185 125.305 207.355 ;
        RECT 125.595 207.185 125.765 207.355 ;
        RECT 126.055 207.185 126.225 207.355 ;
        RECT 126.515 207.185 126.685 207.355 ;
        RECT 126.975 207.185 127.145 207.355 ;
        RECT 127.435 207.185 127.605 207.355 ;
        RECT 127.895 207.185 128.065 207.355 ;
        RECT 128.355 207.185 128.525 207.355 ;
        RECT 128.815 207.185 128.985 207.355 ;
        RECT 129.275 207.185 129.445 207.355 ;
        RECT 129.735 207.185 129.905 207.355 ;
        RECT 130.195 207.185 130.365 207.355 ;
        RECT 130.655 207.185 130.825 207.355 ;
        RECT 131.115 207.185 131.285 207.355 ;
        RECT 131.575 207.185 131.745 207.355 ;
        RECT 132.035 207.185 132.205 207.355 ;
        RECT 132.495 207.185 132.665 207.355 ;
        RECT 132.955 207.185 133.125 207.355 ;
        RECT 133.415 207.185 133.585 207.355 ;
        RECT 133.875 207.185 134.045 207.355 ;
        RECT 134.335 207.185 134.505 207.355 ;
        RECT 134.795 207.185 134.965 207.355 ;
        RECT 135.255 207.185 135.425 207.355 ;
        RECT 135.715 207.185 135.885 207.355 ;
        RECT 136.175 207.185 136.345 207.355 ;
        RECT 136.635 207.185 136.805 207.355 ;
        RECT 137.095 207.185 137.265 207.355 ;
        RECT 137.555 207.185 137.725 207.355 ;
        RECT 138.015 207.185 138.185 207.355 ;
        RECT 138.475 207.185 138.645 207.355 ;
        RECT 138.935 207.185 139.105 207.355 ;
        RECT 139.395 207.185 139.565 207.355 ;
        RECT 139.855 207.185 140.025 207.355 ;
        RECT 140.315 207.185 140.485 207.355 ;
        RECT 140.775 207.185 140.945 207.355 ;
        RECT 141.235 207.185 141.405 207.355 ;
        RECT 141.695 207.185 141.865 207.355 ;
        RECT 142.155 207.185 142.325 207.355 ;
        RECT 142.615 207.185 142.785 207.355 ;
        RECT 143.075 207.185 143.245 207.355 ;
        RECT 143.535 207.185 143.705 207.355 ;
        RECT 143.995 207.185 144.165 207.355 ;
        RECT 144.455 207.185 144.625 207.355 ;
        RECT 144.915 207.185 145.085 207.355 ;
        RECT 145.375 207.185 145.545 207.355 ;
        RECT 145.835 207.185 146.005 207.355 ;
        RECT 146.295 207.185 146.465 207.355 ;
        RECT 146.755 207.185 146.925 207.355 ;
        RECT 147.215 207.185 147.385 207.355 ;
        RECT 147.675 207.185 147.845 207.355 ;
        RECT 148.135 207.185 148.305 207.355 ;
        RECT 148.595 207.185 148.765 207.355 ;
        RECT 149.055 207.185 149.225 207.355 ;
        RECT 149.515 207.185 149.685 207.355 ;
        RECT 149.975 207.185 150.145 207.355 ;
        RECT 150.435 207.185 150.605 207.355 ;
        RECT 150.895 207.185 151.065 207.355 ;
        RECT 151.355 207.185 151.525 207.355 ;
        RECT 151.815 207.185 151.985 207.355 ;
        RECT 152.275 207.185 152.445 207.355 ;
        RECT 152.735 207.185 152.905 207.355 ;
        RECT 153.195 207.185 153.365 207.355 ;
        RECT 153.655 207.185 153.825 207.355 ;
        RECT 154.115 207.185 154.285 207.355 ;
        RECT 154.575 207.185 154.745 207.355 ;
        RECT 155.035 207.185 155.205 207.355 ;
        RECT 155.495 207.185 155.665 207.355 ;
        RECT 155.955 207.185 156.125 207.355 ;
        RECT 74.075 206.675 74.245 206.845 ;
        RECT 75.455 205.655 75.625 205.825 ;
        RECT 78.215 206.675 78.385 206.845 ;
        RECT 77.295 205.655 77.465 205.825 ;
        RECT 76.375 204.975 76.545 205.145 ;
        RECT 79.135 205.655 79.305 205.825 ;
        RECT 79.595 204.975 79.765 205.145 ;
        RECT 82.815 205.995 82.985 206.165 ;
        RECT 81.895 204.975 82.065 205.145 ;
        RECT 84.195 205.315 84.365 205.485 ;
        RECT 88.335 206.675 88.505 206.845 ;
        RECT 86.955 205.655 87.125 205.825 ;
        RECT 89.255 205.655 89.425 205.825 ;
        RECT 91.555 206.675 91.725 206.845 ;
        RECT 92.475 205.655 92.645 205.825 ;
        RECT 97.535 206.675 97.705 206.845 ;
        RECT 93.395 205.315 93.565 205.485 ;
        RECT 100.755 206.335 100.925 206.505 ;
        RECT 104.435 206.675 104.605 206.845 ;
        RECT 98.915 205.315 99.085 205.485 ;
        RECT 100.755 205.315 100.925 205.485 ;
        RECT 102.135 205.655 102.305 205.825 ;
        RECT 103.515 205.655 103.685 205.825 ;
        RECT 101.675 205.315 101.845 205.485 ;
        RECT 106.275 206.335 106.445 206.505 ;
        RECT 105.355 205.655 105.525 205.825 ;
        RECT 108.575 206.675 108.745 206.845 ;
        RECT 107.655 205.655 107.825 205.825 ;
        RECT 110.415 205.995 110.585 206.165 ;
        RECT 112.255 206.675 112.425 206.845 ;
        RECT 110.875 205.655 111.045 205.825 ;
        RECT 113.175 205.655 113.345 205.825 ;
        RECT 113.635 205.655 113.805 205.825 ;
        RECT 114.555 204.975 114.725 205.145 ;
        RECT 116.855 205.655 117.025 205.825 ;
        RECT 117.315 205.655 117.485 205.825 ;
        RECT 115.935 204.975 116.105 205.145 ;
        RECT 118.235 204.975 118.405 205.145 ;
        RECT 118.695 204.975 118.865 205.145 ;
        RECT 121.915 205.655 122.085 205.825 ;
        RECT 125.595 205.995 125.765 206.165 ;
        RECT 123.295 204.975 123.465 205.145 ;
        RECT 126.055 205.995 126.225 206.165 ;
        RECT 127.435 204.975 127.605 205.145 ;
        RECT 130.195 205.995 130.365 206.165 ;
        RECT 131.575 206.335 131.745 206.505 ;
        RECT 129.735 204.975 129.905 205.145 ;
        RECT 135.715 206.335 135.885 206.505 ;
        RECT 134.795 205.655 134.965 205.825 ;
        RECT 137.095 206.335 137.265 206.505 ;
        RECT 136.635 205.655 136.805 205.825 ;
        RECT 138.015 205.655 138.185 205.825 ;
        RECT 141.260 206.335 141.430 206.505 ;
        RECT 139.395 205.655 139.565 205.825 ;
        RECT 140.775 205.655 140.945 205.825 ;
        RECT 138.475 204.975 138.645 205.145 ;
        RECT 141.655 205.995 141.825 206.165 ;
        RECT 142.110 205.315 142.280 205.485 ;
        RECT 143.360 206.335 143.530 206.505 ;
        RECT 142.845 205.995 143.015 206.165 ;
        RECT 144.930 206.335 145.100 206.505 ;
        RECT 145.365 205.995 145.535 206.165 ;
        RECT 149.055 205.995 149.225 206.165 ;
        RECT 150.435 205.655 150.605 205.825 ;
        RECT 147.675 204.975 147.845 205.145 ;
        RECT 70.855 204.465 71.025 204.635 ;
        RECT 71.315 204.465 71.485 204.635 ;
        RECT 71.775 204.465 71.945 204.635 ;
        RECT 72.235 204.465 72.405 204.635 ;
        RECT 72.695 204.465 72.865 204.635 ;
        RECT 73.155 204.465 73.325 204.635 ;
        RECT 73.615 204.465 73.785 204.635 ;
        RECT 74.075 204.465 74.245 204.635 ;
        RECT 74.535 204.465 74.705 204.635 ;
        RECT 74.995 204.465 75.165 204.635 ;
        RECT 75.455 204.465 75.625 204.635 ;
        RECT 75.915 204.465 76.085 204.635 ;
        RECT 76.375 204.465 76.545 204.635 ;
        RECT 76.835 204.465 77.005 204.635 ;
        RECT 77.295 204.465 77.465 204.635 ;
        RECT 77.755 204.465 77.925 204.635 ;
        RECT 78.215 204.465 78.385 204.635 ;
        RECT 78.675 204.465 78.845 204.635 ;
        RECT 79.135 204.465 79.305 204.635 ;
        RECT 79.595 204.465 79.765 204.635 ;
        RECT 80.055 204.465 80.225 204.635 ;
        RECT 80.515 204.465 80.685 204.635 ;
        RECT 80.975 204.465 81.145 204.635 ;
        RECT 81.435 204.465 81.605 204.635 ;
        RECT 81.895 204.465 82.065 204.635 ;
        RECT 82.355 204.465 82.525 204.635 ;
        RECT 82.815 204.465 82.985 204.635 ;
        RECT 83.275 204.465 83.445 204.635 ;
        RECT 83.735 204.465 83.905 204.635 ;
        RECT 84.195 204.465 84.365 204.635 ;
        RECT 84.655 204.465 84.825 204.635 ;
        RECT 85.115 204.465 85.285 204.635 ;
        RECT 85.575 204.465 85.745 204.635 ;
        RECT 86.035 204.465 86.205 204.635 ;
        RECT 86.495 204.465 86.665 204.635 ;
        RECT 86.955 204.465 87.125 204.635 ;
        RECT 87.415 204.465 87.585 204.635 ;
        RECT 87.875 204.465 88.045 204.635 ;
        RECT 88.335 204.465 88.505 204.635 ;
        RECT 88.795 204.465 88.965 204.635 ;
        RECT 89.255 204.465 89.425 204.635 ;
        RECT 89.715 204.465 89.885 204.635 ;
        RECT 90.175 204.465 90.345 204.635 ;
        RECT 90.635 204.465 90.805 204.635 ;
        RECT 91.095 204.465 91.265 204.635 ;
        RECT 91.555 204.465 91.725 204.635 ;
        RECT 92.015 204.465 92.185 204.635 ;
        RECT 92.475 204.465 92.645 204.635 ;
        RECT 92.935 204.465 93.105 204.635 ;
        RECT 93.395 204.465 93.565 204.635 ;
        RECT 93.855 204.465 94.025 204.635 ;
        RECT 94.315 204.465 94.485 204.635 ;
        RECT 94.775 204.465 94.945 204.635 ;
        RECT 95.235 204.465 95.405 204.635 ;
        RECT 95.695 204.465 95.865 204.635 ;
        RECT 96.155 204.465 96.325 204.635 ;
        RECT 96.615 204.465 96.785 204.635 ;
        RECT 97.075 204.465 97.245 204.635 ;
        RECT 97.535 204.465 97.705 204.635 ;
        RECT 97.995 204.465 98.165 204.635 ;
        RECT 98.455 204.465 98.625 204.635 ;
        RECT 98.915 204.465 99.085 204.635 ;
        RECT 99.375 204.465 99.545 204.635 ;
        RECT 99.835 204.465 100.005 204.635 ;
        RECT 100.295 204.465 100.465 204.635 ;
        RECT 100.755 204.465 100.925 204.635 ;
        RECT 101.215 204.465 101.385 204.635 ;
        RECT 101.675 204.465 101.845 204.635 ;
        RECT 102.135 204.465 102.305 204.635 ;
        RECT 102.595 204.465 102.765 204.635 ;
        RECT 103.055 204.465 103.225 204.635 ;
        RECT 103.515 204.465 103.685 204.635 ;
        RECT 103.975 204.465 104.145 204.635 ;
        RECT 104.435 204.465 104.605 204.635 ;
        RECT 104.895 204.465 105.065 204.635 ;
        RECT 105.355 204.465 105.525 204.635 ;
        RECT 105.815 204.465 105.985 204.635 ;
        RECT 106.275 204.465 106.445 204.635 ;
        RECT 106.735 204.465 106.905 204.635 ;
        RECT 107.195 204.465 107.365 204.635 ;
        RECT 107.655 204.465 107.825 204.635 ;
        RECT 108.115 204.465 108.285 204.635 ;
        RECT 108.575 204.465 108.745 204.635 ;
        RECT 109.035 204.465 109.205 204.635 ;
        RECT 109.495 204.465 109.665 204.635 ;
        RECT 109.955 204.465 110.125 204.635 ;
        RECT 110.415 204.465 110.585 204.635 ;
        RECT 110.875 204.465 111.045 204.635 ;
        RECT 111.335 204.465 111.505 204.635 ;
        RECT 111.795 204.465 111.965 204.635 ;
        RECT 112.255 204.465 112.425 204.635 ;
        RECT 112.715 204.465 112.885 204.635 ;
        RECT 113.175 204.465 113.345 204.635 ;
        RECT 113.635 204.465 113.805 204.635 ;
        RECT 114.095 204.465 114.265 204.635 ;
        RECT 114.555 204.465 114.725 204.635 ;
        RECT 115.015 204.465 115.185 204.635 ;
        RECT 115.475 204.465 115.645 204.635 ;
        RECT 115.935 204.465 116.105 204.635 ;
        RECT 116.395 204.465 116.565 204.635 ;
        RECT 116.855 204.465 117.025 204.635 ;
        RECT 117.315 204.465 117.485 204.635 ;
        RECT 117.775 204.465 117.945 204.635 ;
        RECT 118.235 204.465 118.405 204.635 ;
        RECT 118.695 204.465 118.865 204.635 ;
        RECT 119.155 204.465 119.325 204.635 ;
        RECT 119.615 204.465 119.785 204.635 ;
        RECT 120.075 204.465 120.245 204.635 ;
        RECT 120.535 204.465 120.705 204.635 ;
        RECT 120.995 204.465 121.165 204.635 ;
        RECT 121.455 204.465 121.625 204.635 ;
        RECT 121.915 204.465 122.085 204.635 ;
        RECT 122.375 204.465 122.545 204.635 ;
        RECT 122.835 204.465 123.005 204.635 ;
        RECT 123.295 204.465 123.465 204.635 ;
        RECT 123.755 204.465 123.925 204.635 ;
        RECT 124.215 204.465 124.385 204.635 ;
        RECT 124.675 204.465 124.845 204.635 ;
        RECT 125.135 204.465 125.305 204.635 ;
        RECT 125.595 204.465 125.765 204.635 ;
        RECT 126.055 204.465 126.225 204.635 ;
        RECT 126.515 204.465 126.685 204.635 ;
        RECT 126.975 204.465 127.145 204.635 ;
        RECT 127.435 204.465 127.605 204.635 ;
        RECT 127.895 204.465 128.065 204.635 ;
        RECT 128.355 204.465 128.525 204.635 ;
        RECT 128.815 204.465 128.985 204.635 ;
        RECT 129.275 204.465 129.445 204.635 ;
        RECT 129.735 204.465 129.905 204.635 ;
        RECT 130.195 204.465 130.365 204.635 ;
        RECT 130.655 204.465 130.825 204.635 ;
        RECT 131.115 204.465 131.285 204.635 ;
        RECT 131.575 204.465 131.745 204.635 ;
        RECT 132.035 204.465 132.205 204.635 ;
        RECT 132.495 204.465 132.665 204.635 ;
        RECT 132.955 204.465 133.125 204.635 ;
        RECT 133.415 204.465 133.585 204.635 ;
        RECT 133.875 204.465 134.045 204.635 ;
        RECT 134.335 204.465 134.505 204.635 ;
        RECT 134.795 204.465 134.965 204.635 ;
        RECT 135.255 204.465 135.425 204.635 ;
        RECT 135.715 204.465 135.885 204.635 ;
        RECT 136.175 204.465 136.345 204.635 ;
        RECT 136.635 204.465 136.805 204.635 ;
        RECT 137.095 204.465 137.265 204.635 ;
        RECT 137.555 204.465 137.725 204.635 ;
        RECT 138.015 204.465 138.185 204.635 ;
        RECT 138.475 204.465 138.645 204.635 ;
        RECT 138.935 204.465 139.105 204.635 ;
        RECT 139.395 204.465 139.565 204.635 ;
        RECT 139.855 204.465 140.025 204.635 ;
        RECT 140.315 204.465 140.485 204.635 ;
        RECT 140.775 204.465 140.945 204.635 ;
        RECT 141.235 204.465 141.405 204.635 ;
        RECT 141.695 204.465 141.865 204.635 ;
        RECT 142.155 204.465 142.325 204.635 ;
        RECT 142.615 204.465 142.785 204.635 ;
        RECT 143.075 204.465 143.245 204.635 ;
        RECT 143.535 204.465 143.705 204.635 ;
        RECT 143.995 204.465 144.165 204.635 ;
        RECT 144.455 204.465 144.625 204.635 ;
        RECT 144.915 204.465 145.085 204.635 ;
        RECT 145.375 204.465 145.545 204.635 ;
        RECT 145.835 204.465 146.005 204.635 ;
        RECT 146.295 204.465 146.465 204.635 ;
        RECT 146.755 204.465 146.925 204.635 ;
        RECT 147.215 204.465 147.385 204.635 ;
        RECT 147.675 204.465 147.845 204.635 ;
        RECT 148.135 204.465 148.305 204.635 ;
        RECT 148.595 204.465 148.765 204.635 ;
        RECT 149.055 204.465 149.225 204.635 ;
        RECT 149.515 204.465 149.685 204.635 ;
        RECT 149.975 204.465 150.145 204.635 ;
        RECT 150.435 204.465 150.605 204.635 ;
        RECT 150.895 204.465 151.065 204.635 ;
        RECT 151.355 204.465 151.525 204.635 ;
        RECT 151.815 204.465 151.985 204.635 ;
        RECT 152.275 204.465 152.445 204.635 ;
        RECT 152.735 204.465 152.905 204.635 ;
        RECT 153.195 204.465 153.365 204.635 ;
        RECT 153.655 204.465 153.825 204.635 ;
        RECT 154.115 204.465 154.285 204.635 ;
        RECT 154.575 204.465 154.745 204.635 ;
        RECT 155.035 204.465 155.205 204.635 ;
        RECT 155.495 204.465 155.665 204.635 ;
        RECT 155.955 204.465 156.125 204.635 ;
        RECT 73.155 202.935 73.325 203.105 ;
        RECT 73.640 202.595 73.810 202.765 ;
        RECT 74.035 202.935 74.205 203.105 ;
        RECT 74.490 203.615 74.660 203.785 ;
        RECT 75.225 202.935 75.395 203.105 ;
        RECT 75.740 202.595 75.910 202.765 ;
        RECT 77.310 202.595 77.480 202.765 ;
        RECT 77.745 202.935 77.915 203.105 ;
        RECT 80.055 203.955 80.225 204.125 ;
        RECT 82.355 203.275 82.525 203.445 ;
        RECT 83.275 203.275 83.445 203.445 ;
        RECT 83.735 202.935 83.905 203.105 ;
        RECT 83.275 202.255 83.445 202.425 ;
        RECT 84.220 202.595 84.390 202.765 ;
        RECT 84.615 202.935 84.785 203.105 ;
        RECT 85.015 203.275 85.185 203.445 ;
        RECT 85.805 202.935 85.975 203.105 ;
        RECT 86.320 202.595 86.490 202.765 ;
        RECT 87.890 202.595 88.060 202.765 ;
        RECT 88.325 202.935 88.495 203.105 ;
        RECT 94.315 203.955 94.485 204.125 ;
        RECT 92.015 203.275 92.185 203.445 ;
        RECT 93.395 203.275 93.565 203.445 ;
        RECT 90.635 202.255 90.805 202.425 ;
        RECT 91.095 202.255 91.265 202.425 ;
        RECT 95.695 203.275 95.865 203.445 ;
        RECT 94.775 202.255 94.945 202.425 ;
        RECT 99.835 203.955 100.005 204.125 ;
        RECT 97.995 203.275 98.165 203.445 ;
        RECT 98.455 202.935 98.625 203.105 ;
        RECT 100.755 203.955 100.925 204.125 ;
        RECT 101.675 203.615 101.845 203.785 ;
        RECT 104.895 203.955 105.065 204.125 ;
        RECT 101.675 202.255 101.845 202.425 ;
        RECT 103.515 202.595 103.685 202.765 ;
        RECT 106.735 203.615 106.905 203.785 ;
        RECT 107.195 202.935 107.365 203.105 ;
        RECT 107.655 202.935 107.825 203.105 ;
        RECT 109.035 202.255 109.205 202.425 ;
        RECT 111.345 202.935 111.515 203.105 ;
        RECT 111.780 202.595 111.950 202.765 ;
        RECT 113.865 202.935 114.035 203.105 ;
        RECT 113.350 202.595 113.520 202.765 ;
        RECT 114.600 203.275 114.770 203.445 ;
        RECT 115.055 202.935 115.225 203.105 ;
        RECT 115.935 203.275 116.105 203.445 ;
        RECT 117.315 203.275 117.485 203.445 ;
        RECT 115.450 202.595 115.620 202.765 ;
        RECT 116.395 202.255 116.565 202.425 ;
        RECT 117.775 202.595 117.945 202.765 ;
        RECT 120.075 203.955 120.245 204.125 ;
        RECT 120.995 202.935 121.165 203.105 ;
        RECT 124.215 203.275 124.385 203.445 ;
        RECT 125.595 203.275 125.765 203.445 ;
        RECT 125.135 202.595 125.305 202.765 ;
        RECT 126.080 202.595 126.250 202.765 ;
        RECT 126.475 202.935 126.645 203.105 ;
        RECT 126.875 203.275 127.045 203.445 ;
        RECT 127.665 202.935 127.835 203.105 ;
        RECT 128.180 202.595 128.350 202.765 ;
        RECT 129.750 202.595 129.920 202.765 ;
        RECT 130.185 202.935 130.355 203.105 ;
        RECT 134.335 203.275 134.505 203.445 ;
        RECT 135.715 203.275 135.885 203.445 ;
        RECT 132.495 202.595 132.665 202.765 ;
        RECT 133.415 202.255 133.585 202.425 ;
        RECT 137.095 203.275 137.265 203.445 ;
        RECT 136.635 202.595 136.805 202.765 ;
        RECT 137.580 202.595 137.750 202.765 ;
        RECT 137.975 202.935 138.145 203.105 ;
        RECT 138.375 203.275 138.545 203.445 ;
        RECT 139.165 202.935 139.335 203.105 ;
        RECT 139.680 202.595 139.850 202.765 ;
        RECT 141.250 202.595 141.420 202.765 ;
        RECT 141.685 202.935 141.855 203.105 ;
        RECT 145.375 203.275 145.545 203.445 ;
        RECT 143.995 202.255 144.165 202.425 ;
        RECT 144.455 202.255 144.625 202.425 ;
        RECT 146.755 203.275 146.925 203.445 ;
        RECT 145.835 202.255 146.005 202.425 ;
        RECT 148.595 202.255 148.765 202.425 ;
        RECT 150.895 202.935 151.065 203.105 ;
        RECT 151.355 202.935 151.525 203.105 ;
        RECT 153.655 203.275 153.825 203.445 ;
        RECT 152.735 202.595 152.905 202.765 ;
        RECT 70.855 201.745 71.025 201.915 ;
        RECT 71.315 201.745 71.485 201.915 ;
        RECT 71.775 201.745 71.945 201.915 ;
        RECT 72.235 201.745 72.405 201.915 ;
        RECT 72.695 201.745 72.865 201.915 ;
        RECT 73.155 201.745 73.325 201.915 ;
        RECT 73.615 201.745 73.785 201.915 ;
        RECT 74.075 201.745 74.245 201.915 ;
        RECT 74.535 201.745 74.705 201.915 ;
        RECT 74.995 201.745 75.165 201.915 ;
        RECT 75.455 201.745 75.625 201.915 ;
        RECT 75.915 201.745 76.085 201.915 ;
        RECT 76.375 201.745 76.545 201.915 ;
        RECT 76.835 201.745 77.005 201.915 ;
        RECT 77.295 201.745 77.465 201.915 ;
        RECT 77.755 201.745 77.925 201.915 ;
        RECT 78.215 201.745 78.385 201.915 ;
        RECT 78.675 201.745 78.845 201.915 ;
        RECT 79.135 201.745 79.305 201.915 ;
        RECT 79.595 201.745 79.765 201.915 ;
        RECT 80.055 201.745 80.225 201.915 ;
        RECT 80.515 201.745 80.685 201.915 ;
        RECT 80.975 201.745 81.145 201.915 ;
        RECT 81.435 201.745 81.605 201.915 ;
        RECT 81.895 201.745 82.065 201.915 ;
        RECT 82.355 201.745 82.525 201.915 ;
        RECT 82.815 201.745 82.985 201.915 ;
        RECT 83.275 201.745 83.445 201.915 ;
        RECT 83.735 201.745 83.905 201.915 ;
        RECT 84.195 201.745 84.365 201.915 ;
        RECT 84.655 201.745 84.825 201.915 ;
        RECT 85.115 201.745 85.285 201.915 ;
        RECT 85.575 201.745 85.745 201.915 ;
        RECT 86.035 201.745 86.205 201.915 ;
        RECT 86.495 201.745 86.665 201.915 ;
        RECT 86.955 201.745 87.125 201.915 ;
        RECT 87.415 201.745 87.585 201.915 ;
        RECT 87.875 201.745 88.045 201.915 ;
        RECT 88.335 201.745 88.505 201.915 ;
        RECT 88.795 201.745 88.965 201.915 ;
        RECT 89.255 201.745 89.425 201.915 ;
        RECT 89.715 201.745 89.885 201.915 ;
        RECT 90.175 201.745 90.345 201.915 ;
        RECT 90.635 201.745 90.805 201.915 ;
        RECT 91.095 201.745 91.265 201.915 ;
        RECT 91.555 201.745 91.725 201.915 ;
        RECT 92.015 201.745 92.185 201.915 ;
        RECT 92.475 201.745 92.645 201.915 ;
        RECT 92.935 201.745 93.105 201.915 ;
        RECT 93.395 201.745 93.565 201.915 ;
        RECT 93.855 201.745 94.025 201.915 ;
        RECT 94.315 201.745 94.485 201.915 ;
        RECT 94.775 201.745 94.945 201.915 ;
        RECT 95.235 201.745 95.405 201.915 ;
        RECT 95.695 201.745 95.865 201.915 ;
        RECT 96.155 201.745 96.325 201.915 ;
        RECT 96.615 201.745 96.785 201.915 ;
        RECT 97.075 201.745 97.245 201.915 ;
        RECT 97.535 201.745 97.705 201.915 ;
        RECT 97.995 201.745 98.165 201.915 ;
        RECT 98.455 201.745 98.625 201.915 ;
        RECT 98.915 201.745 99.085 201.915 ;
        RECT 99.375 201.745 99.545 201.915 ;
        RECT 99.835 201.745 100.005 201.915 ;
        RECT 100.295 201.745 100.465 201.915 ;
        RECT 100.755 201.745 100.925 201.915 ;
        RECT 101.215 201.745 101.385 201.915 ;
        RECT 101.675 201.745 101.845 201.915 ;
        RECT 102.135 201.745 102.305 201.915 ;
        RECT 102.595 201.745 102.765 201.915 ;
        RECT 103.055 201.745 103.225 201.915 ;
        RECT 103.515 201.745 103.685 201.915 ;
        RECT 103.975 201.745 104.145 201.915 ;
        RECT 104.435 201.745 104.605 201.915 ;
        RECT 104.895 201.745 105.065 201.915 ;
        RECT 105.355 201.745 105.525 201.915 ;
        RECT 105.815 201.745 105.985 201.915 ;
        RECT 106.275 201.745 106.445 201.915 ;
        RECT 106.735 201.745 106.905 201.915 ;
        RECT 107.195 201.745 107.365 201.915 ;
        RECT 107.655 201.745 107.825 201.915 ;
        RECT 108.115 201.745 108.285 201.915 ;
        RECT 108.575 201.745 108.745 201.915 ;
        RECT 109.035 201.745 109.205 201.915 ;
        RECT 109.495 201.745 109.665 201.915 ;
        RECT 109.955 201.745 110.125 201.915 ;
        RECT 110.415 201.745 110.585 201.915 ;
        RECT 110.875 201.745 111.045 201.915 ;
        RECT 111.335 201.745 111.505 201.915 ;
        RECT 111.795 201.745 111.965 201.915 ;
        RECT 112.255 201.745 112.425 201.915 ;
        RECT 112.715 201.745 112.885 201.915 ;
        RECT 113.175 201.745 113.345 201.915 ;
        RECT 113.635 201.745 113.805 201.915 ;
        RECT 114.095 201.745 114.265 201.915 ;
        RECT 114.555 201.745 114.725 201.915 ;
        RECT 115.015 201.745 115.185 201.915 ;
        RECT 115.475 201.745 115.645 201.915 ;
        RECT 115.935 201.745 116.105 201.915 ;
        RECT 116.395 201.745 116.565 201.915 ;
        RECT 116.855 201.745 117.025 201.915 ;
        RECT 117.315 201.745 117.485 201.915 ;
        RECT 117.775 201.745 117.945 201.915 ;
        RECT 118.235 201.745 118.405 201.915 ;
        RECT 118.695 201.745 118.865 201.915 ;
        RECT 119.155 201.745 119.325 201.915 ;
        RECT 119.615 201.745 119.785 201.915 ;
        RECT 120.075 201.745 120.245 201.915 ;
        RECT 120.535 201.745 120.705 201.915 ;
        RECT 120.995 201.745 121.165 201.915 ;
        RECT 121.455 201.745 121.625 201.915 ;
        RECT 121.915 201.745 122.085 201.915 ;
        RECT 122.375 201.745 122.545 201.915 ;
        RECT 122.835 201.745 123.005 201.915 ;
        RECT 123.295 201.745 123.465 201.915 ;
        RECT 123.755 201.745 123.925 201.915 ;
        RECT 124.215 201.745 124.385 201.915 ;
        RECT 124.675 201.745 124.845 201.915 ;
        RECT 125.135 201.745 125.305 201.915 ;
        RECT 125.595 201.745 125.765 201.915 ;
        RECT 126.055 201.745 126.225 201.915 ;
        RECT 126.515 201.745 126.685 201.915 ;
        RECT 126.975 201.745 127.145 201.915 ;
        RECT 127.435 201.745 127.605 201.915 ;
        RECT 127.895 201.745 128.065 201.915 ;
        RECT 128.355 201.745 128.525 201.915 ;
        RECT 128.815 201.745 128.985 201.915 ;
        RECT 129.275 201.745 129.445 201.915 ;
        RECT 129.735 201.745 129.905 201.915 ;
        RECT 130.195 201.745 130.365 201.915 ;
        RECT 130.655 201.745 130.825 201.915 ;
        RECT 131.115 201.745 131.285 201.915 ;
        RECT 131.575 201.745 131.745 201.915 ;
        RECT 132.035 201.745 132.205 201.915 ;
        RECT 132.495 201.745 132.665 201.915 ;
        RECT 132.955 201.745 133.125 201.915 ;
        RECT 133.415 201.745 133.585 201.915 ;
        RECT 133.875 201.745 134.045 201.915 ;
        RECT 134.335 201.745 134.505 201.915 ;
        RECT 134.795 201.745 134.965 201.915 ;
        RECT 135.255 201.745 135.425 201.915 ;
        RECT 135.715 201.745 135.885 201.915 ;
        RECT 136.175 201.745 136.345 201.915 ;
        RECT 136.635 201.745 136.805 201.915 ;
        RECT 137.095 201.745 137.265 201.915 ;
        RECT 137.555 201.745 137.725 201.915 ;
        RECT 138.015 201.745 138.185 201.915 ;
        RECT 138.475 201.745 138.645 201.915 ;
        RECT 138.935 201.745 139.105 201.915 ;
        RECT 139.395 201.745 139.565 201.915 ;
        RECT 139.855 201.745 140.025 201.915 ;
        RECT 140.315 201.745 140.485 201.915 ;
        RECT 140.775 201.745 140.945 201.915 ;
        RECT 141.235 201.745 141.405 201.915 ;
        RECT 141.695 201.745 141.865 201.915 ;
        RECT 142.155 201.745 142.325 201.915 ;
        RECT 142.615 201.745 142.785 201.915 ;
        RECT 143.075 201.745 143.245 201.915 ;
        RECT 143.535 201.745 143.705 201.915 ;
        RECT 143.995 201.745 144.165 201.915 ;
        RECT 144.455 201.745 144.625 201.915 ;
        RECT 144.915 201.745 145.085 201.915 ;
        RECT 145.375 201.745 145.545 201.915 ;
        RECT 145.835 201.745 146.005 201.915 ;
        RECT 146.295 201.745 146.465 201.915 ;
        RECT 146.755 201.745 146.925 201.915 ;
        RECT 147.215 201.745 147.385 201.915 ;
        RECT 147.675 201.745 147.845 201.915 ;
        RECT 148.135 201.745 148.305 201.915 ;
        RECT 148.595 201.745 148.765 201.915 ;
        RECT 149.055 201.745 149.225 201.915 ;
        RECT 149.515 201.745 149.685 201.915 ;
        RECT 149.975 201.745 150.145 201.915 ;
        RECT 150.435 201.745 150.605 201.915 ;
        RECT 150.895 201.745 151.065 201.915 ;
        RECT 151.355 201.745 151.525 201.915 ;
        RECT 151.815 201.745 151.985 201.915 ;
        RECT 152.275 201.745 152.445 201.915 ;
        RECT 152.735 201.745 152.905 201.915 ;
        RECT 153.195 201.745 153.365 201.915 ;
        RECT 153.655 201.745 153.825 201.915 ;
        RECT 154.115 201.745 154.285 201.915 ;
        RECT 154.575 201.745 154.745 201.915 ;
        RECT 155.035 201.745 155.205 201.915 ;
        RECT 155.495 201.745 155.665 201.915 ;
        RECT 155.955 201.745 156.125 201.915 ;
        RECT 74.560 200.895 74.730 201.065 ;
        RECT 74.075 200.215 74.245 200.385 ;
        RECT 74.955 200.555 75.125 200.725 ;
        RECT 75.410 199.875 75.580 200.045 ;
        RECT 76.660 200.895 76.830 201.065 ;
        RECT 76.145 200.555 76.315 200.725 ;
        RECT 78.230 200.895 78.400 201.065 ;
        RECT 78.665 200.555 78.835 200.725 ;
        RECT 83.275 200.895 83.445 201.065 ;
        RECT 82.355 200.215 82.525 200.385 ;
        RECT 80.975 199.535 81.145 199.705 ;
        RECT 84.195 199.535 84.365 199.705 ;
        RECT 86.505 200.555 86.675 200.725 ;
        RECT 86.940 200.895 87.110 201.065 ;
        RECT 88.510 200.895 88.680 201.065 ;
        RECT 89.025 200.555 89.195 200.725 ;
        RECT 89.870 199.875 90.040 200.045 ;
        RECT 90.215 200.555 90.385 200.725 ;
        RECT 90.610 200.895 90.780 201.065 ;
        RECT 92.500 200.895 92.670 201.065 ;
        RECT 91.095 200.555 91.265 200.725 ;
        RECT 92.015 200.215 92.185 200.385 ;
        RECT 92.895 200.555 93.065 200.725 ;
        RECT 93.350 200.215 93.520 200.385 ;
        RECT 94.600 200.895 94.770 201.065 ;
        RECT 94.085 200.555 94.255 200.725 ;
        RECT 96.170 200.895 96.340 201.065 ;
        RECT 96.605 200.555 96.775 200.725 ;
        RECT 100.295 200.555 100.465 200.725 ;
        RECT 100.755 200.215 100.925 200.385 ;
        RECT 98.915 199.535 99.085 199.705 ;
        RECT 101.215 199.875 101.385 200.045 ;
        RECT 103.055 201.235 103.225 201.405 ;
        RECT 104.435 201.235 104.605 201.405 ;
        RECT 107.655 200.895 107.825 201.065 ;
        RECT 105.355 200.215 105.525 200.385 ;
        RECT 106.275 200.215 106.445 200.385 ;
        RECT 106.735 200.215 106.905 200.385 ;
        RECT 107.655 200.215 107.825 200.385 ;
        RECT 108.115 200.215 108.285 200.385 ;
        RECT 108.575 199.535 108.745 199.705 ;
        RECT 115.040 200.895 115.210 201.065 ;
        RECT 111.795 200.215 111.965 200.385 ;
        RECT 112.715 200.215 112.885 200.385 ;
        RECT 113.175 200.215 113.345 200.385 ;
        RECT 114.555 200.555 114.725 200.725 ;
        RECT 110.875 199.535 111.045 199.705 ;
        RECT 115.435 200.555 115.605 200.725 ;
        RECT 115.890 199.875 116.060 200.045 ;
        RECT 117.140 200.895 117.310 201.065 ;
        RECT 116.625 200.555 116.795 200.725 ;
        RECT 118.710 200.895 118.880 201.065 ;
        RECT 119.145 200.555 119.315 200.725 ;
        RECT 121.455 201.235 121.625 201.405 ;
        RECT 123.755 200.895 123.925 201.065 ;
        RECT 124.215 200.555 124.385 200.725 ;
        RECT 122.835 200.215 123.005 200.385 ;
        RECT 126.055 200.555 126.225 200.725 ;
        RECT 121.915 199.535 122.085 199.705 ;
        RECT 126.515 199.875 126.685 200.045 ;
        RECT 126.975 199.875 127.145 200.045 ;
        RECT 128.815 199.535 128.985 199.705 ;
        RECT 129.275 200.555 129.445 200.725 ;
        RECT 131.115 200.895 131.285 201.065 ;
        RECT 130.195 200.215 130.365 200.385 ;
        RECT 131.575 200.215 131.745 200.385 ;
        RECT 135.715 201.235 135.885 201.405 ;
        RECT 133.415 200.215 133.585 200.385 ;
        RECT 134.335 200.215 134.505 200.385 ;
        RECT 134.795 200.215 134.965 200.385 ;
        RECT 132.495 199.535 132.665 199.705 ;
        RECT 138.015 200.555 138.185 200.725 ;
        RECT 138.935 200.555 139.105 200.725 ;
        RECT 139.855 200.895 140.025 201.065 ;
        RECT 140.775 199.875 140.945 200.045 ;
        RECT 143.075 200.555 143.245 200.725 ;
        RECT 143.535 199.535 143.705 199.705 ;
        RECT 143.995 199.875 144.165 200.045 ;
        RECT 146.780 200.895 146.950 201.065 ;
        RECT 146.295 200.555 146.465 200.725 ;
        RECT 145.835 199.535 146.005 199.705 ;
        RECT 147.175 200.555 147.345 200.725 ;
        RECT 147.520 199.875 147.690 200.045 ;
        RECT 148.880 200.895 149.050 201.065 ;
        RECT 148.365 200.555 148.535 200.725 ;
        RECT 150.450 200.895 150.620 201.065 ;
        RECT 150.885 200.555 151.055 200.725 ;
        RECT 153.195 199.535 153.365 199.705 ;
        RECT 70.855 199.025 71.025 199.195 ;
        RECT 71.315 199.025 71.485 199.195 ;
        RECT 71.775 199.025 71.945 199.195 ;
        RECT 72.235 199.025 72.405 199.195 ;
        RECT 72.695 199.025 72.865 199.195 ;
        RECT 73.155 199.025 73.325 199.195 ;
        RECT 73.615 199.025 73.785 199.195 ;
        RECT 74.075 199.025 74.245 199.195 ;
        RECT 74.535 199.025 74.705 199.195 ;
        RECT 74.995 199.025 75.165 199.195 ;
        RECT 75.455 199.025 75.625 199.195 ;
        RECT 75.915 199.025 76.085 199.195 ;
        RECT 76.375 199.025 76.545 199.195 ;
        RECT 76.835 199.025 77.005 199.195 ;
        RECT 77.295 199.025 77.465 199.195 ;
        RECT 77.755 199.025 77.925 199.195 ;
        RECT 78.215 199.025 78.385 199.195 ;
        RECT 78.675 199.025 78.845 199.195 ;
        RECT 79.135 199.025 79.305 199.195 ;
        RECT 79.595 199.025 79.765 199.195 ;
        RECT 80.055 199.025 80.225 199.195 ;
        RECT 80.515 199.025 80.685 199.195 ;
        RECT 80.975 199.025 81.145 199.195 ;
        RECT 81.435 199.025 81.605 199.195 ;
        RECT 81.895 199.025 82.065 199.195 ;
        RECT 82.355 199.025 82.525 199.195 ;
        RECT 82.815 199.025 82.985 199.195 ;
        RECT 83.275 199.025 83.445 199.195 ;
        RECT 83.735 199.025 83.905 199.195 ;
        RECT 84.195 199.025 84.365 199.195 ;
        RECT 84.655 199.025 84.825 199.195 ;
        RECT 85.115 199.025 85.285 199.195 ;
        RECT 85.575 199.025 85.745 199.195 ;
        RECT 86.035 199.025 86.205 199.195 ;
        RECT 86.495 199.025 86.665 199.195 ;
        RECT 86.955 199.025 87.125 199.195 ;
        RECT 87.415 199.025 87.585 199.195 ;
        RECT 87.875 199.025 88.045 199.195 ;
        RECT 88.335 199.025 88.505 199.195 ;
        RECT 88.795 199.025 88.965 199.195 ;
        RECT 89.255 199.025 89.425 199.195 ;
        RECT 89.715 199.025 89.885 199.195 ;
        RECT 90.175 199.025 90.345 199.195 ;
        RECT 90.635 199.025 90.805 199.195 ;
        RECT 91.095 199.025 91.265 199.195 ;
        RECT 91.555 199.025 91.725 199.195 ;
        RECT 92.015 199.025 92.185 199.195 ;
        RECT 92.475 199.025 92.645 199.195 ;
        RECT 92.935 199.025 93.105 199.195 ;
        RECT 93.395 199.025 93.565 199.195 ;
        RECT 93.855 199.025 94.025 199.195 ;
        RECT 94.315 199.025 94.485 199.195 ;
        RECT 94.775 199.025 94.945 199.195 ;
        RECT 95.235 199.025 95.405 199.195 ;
        RECT 95.695 199.025 95.865 199.195 ;
        RECT 96.155 199.025 96.325 199.195 ;
        RECT 96.615 199.025 96.785 199.195 ;
        RECT 97.075 199.025 97.245 199.195 ;
        RECT 97.535 199.025 97.705 199.195 ;
        RECT 97.995 199.025 98.165 199.195 ;
        RECT 98.455 199.025 98.625 199.195 ;
        RECT 98.915 199.025 99.085 199.195 ;
        RECT 99.375 199.025 99.545 199.195 ;
        RECT 99.835 199.025 100.005 199.195 ;
        RECT 100.295 199.025 100.465 199.195 ;
        RECT 100.755 199.025 100.925 199.195 ;
        RECT 101.215 199.025 101.385 199.195 ;
        RECT 101.675 199.025 101.845 199.195 ;
        RECT 102.135 199.025 102.305 199.195 ;
        RECT 102.595 199.025 102.765 199.195 ;
        RECT 103.055 199.025 103.225 199.195 ;
        RECT 103.515 199.025 103.685 199.195 ;
        RECT 103.975 199.025 104.145 199.195 ;
        RECT 104.435 199.025 104.605 199.195 ;
        RECT 104.895 199.025 105.065 199.195 ;
        RECT 105.355 199.025 105.525 199.195 ;
        RECT 105.815 199.025 105.985 199.195 ;
        RECT 106.275 199.025 106.445 199.195 ;
        RECT 106.735 199.025 106.905 199.195 ;
        RECT 107.195 199.025 107.365 199.195 ;
        RECT 107.655 199.025 107.825 199.195 ;
        RECT 108.115 199.025 108.285 199.195 ;
        RECT 108.575 199.025 108.745 199.195 ;
        RECT 109.035 199.025 109.205 199.195 ;
        RECT 109.495 199.025 109.665 199.195 ;
        RECT 109.955 199.025 110.125 199.195 ;
        RECT 110.415 199.025 110.585 199.195 ;
        RECT 110.875 199.025 111.045 199.195 ;
        RECT 111.335 199.025 111.505 199.195 ;
        RECT 111.795 199.025 111.965 199.195 ;
        RECT 112.255 199.025 112.425 199.195 ;
        RECT 112.715 199.025 112.885 199.195 ;
        RECT 113.175 199.025 113.345 199.195 ;
        RECT 113.635 199.025 113.805 199.195 ;
        RECT 114.095 199.025 114.265 199.195 ;
        RECT 114.555 199.025 114.725 199.195 ;
        RECT 115.015 199.025 115.185 199.195 ;
        RECT 115.475 199.025 115.645 199.195 ;
        RECT 115.935 199.025 116.105 199.195 ;
        RECT 116.395 199.025 116.565 199.195 ;
        RECT 116.855 199.025 117.025 199.195 ;
        RECT 117.315 199.025 117.485 199.195 ;
        RECT 117.775 199.025 117.945 199.195 ;
        RECT 118.235 199.025 118.405 199.195 ;
        RECT 118.695 199.025 118.865 199.195 ;
        RECT 119.155 199.025 119.325 199.195 ;
        RECT 119.615 199.025 119.785 199.195 ;
        RECT 120.075 199.025 120.245 199.195 ;
        RECT 120.535 199.025 120.705 199.195 ;
        RECT 120.995 199.025 121.165 199.195 ;
        RECT 121.455 199.025 121.625 199.195 ;
        RECT 121.915 199.025 122.085 199.195 ;
        RECT 122.375 199.025 122.545 199.195 ;
        RECT 122.835 199.025 123.005 199.195 ;
        RECT 123.295 199.025 123.465 199.195 ;
        RECT 123.755 199.025 123.925 199.195 ;
        RECT 124.215 199.025 124.385 199.195 ;
        RECT 124.675 199.025 124.845 199.195 ;
        RECT 125.135 199.025 125.305 199.195 ;
        RECT 125.595 199.025 125.765 199.195 ;
        RECT 126.055 199.025 126.225 199.195 ;
        RECT 126.515 199.025 126.685 199.195 ;
        RECT 126.975 199.025 127.145 199.195 ;
        RECT 127.435 199.025 127.605 199.195 ;
        RECT 127.895 199.025 128.065 199.195 ;
        RECT 128.355 199.025 128.525 199.195 ;
        RECT 128.815 199.025 128.985 199.195 ;
        RECT 129.275 199.025 129.445 199.195 ;
        RECT 129.735 199.025 129.905 199.195 ;
        RECT 130.195 199.025 130.365 199.195 ;
        RECT 130.655 199.025 130.825 199.195 ;
        RECT 131.115 199.025 131.285 199.195 ;
        RECT 131.575 199.025 131.745 199.195 ;
        RECT 132.035 199.025 132.205 199.195 ;
        RECT 132.495 199.025 132.665 199.195 ;
        RECT 132.955 199.025 133.125 199.195 ;
        RECT 133.415 199.025 133.585 199.195 ;
        RECT 133.875 199.025 134.045 199.195 ;
        RECT 134.335 199.025 134.505 199.195 ;
        RECT 134.795 199.025 134.965 199.195 ;
        RECT 135.255 199.025 135.425 199.195 ;
        RECT 135.715 199.025 135.885 199.195 ;
        RECT 136.175 199.025 136.345 199.195 ;
        RECT 136.635 199.025 136.805 199.195 ;
        RECT 137.095 199.025 137.265 199.195 ;
        RECT 137.555 199.025 137.725 199.195 ;
        RECT 138.015 199.025 138.185 199.195 ;
        RECT 138.475 199.025 138.645 199.195 ;
        RECT 138.935 199.025 139.105 199.195 ;
        RECT 139.395 199.025 139.565 199.195 ;
        RECT 139.855 199.025 140.025 199.195 ;
        RECT 140.315 199.025 140.485 199.195 ;
        RECT 140.775 199.025 140.945 199.195 ;
        RECT 141.235 199.025 141.405 199.195 ;
        RECT 141.695 199.025 141.865 199.195 ;
        RECT 142.155 199.025 142.325 199.195 ;
        RECT 142.615 199.025 142.785 199.195 ;
        RECT 143.075 199.025 143.245 199.195 ;
        RECT 143.535 199.025 143.705 199.195 ;
        RECT 143.995 199.025 144.165 199.195 ;
        RECT 144.455 199.025 144.625 199.195 ;
        RECT 144.915 199.025 145.085 199.195 ;
        RECT 145.375 199.025 145.545 199.195 ;
        RECT 145.835 199.025 146.005 199.195 ;
        RECT 146.295 199.025 146.465 199.195 ;
        RECT 146.755 199.025 146.925 199.195 ;
        RECT 147.215 199.025 147.385 199.195 ;
        RECT 147.675 199.025 147.845 199.195 ;
        RECT 148.135 199.025 148.305 199.195 ;
        RECT 148.595 199.025 148.765 199.195 ;
        RECT 149.055 199.025 149.225 199.195 ;
        RECT 149.515 199.025 149.685 199.195 ;
        RECT 149.975 199.025 150.145 199.195 ;
        RECT 150.435 199.025 150.605 199.195 ;
        RECT 150.895 199.025 151.065 199.195 ;
        RECT 151.355 199.025 151.525 199.195 ;
        RECT 151.815 199.025 151.985 199.195 ;
        RECT 152.275 199.025 152.445 199.195 ;
        RECT 152.735 199.025 152.905 199.195 ;
        RECT 153.195 199.025 153.365 199.195 ;
        RECT 153.655 199.025 153.825 199.195 ;
        RECT 154.115 199.025 154.285 199.195 ;
        RECT 154.575 199.025 154.745 199.195 ;
        RECT 155.035 199.025 155.205 199.195 ;
        RECT 155.495 199.025 155.665 199.195 ;
        RECT 155.955 199.025 156.125 199.195 ;
        RECT 74.995 198.515 75.165 198.685 ;
        RECT 78.215 198.515 78.385 198.685 ;
        RECT 78.675 198.515 78.845 198.685 ;
        RECT 75.915 197.835 76.085 198.005 ;
        RECT 77.755 197.835 77.925 198.005 ;
        RECT 76.835 197.155 77.005 197.325 ;
        RECT 80.055 197.835 80.225 198.005 ;
        RECT 80.515 197.155 80.685 197.325 ;
        RECT 82.355 198.175 82.525 198.345 ;
        RECT 84.655 198.515 84.825 198.685 ;
        RECT 83.735 197.835 83.905 198.005 ;
        RECT 83.275 197.155 83.445 197.325 ;
        RECT 82.355 196.815 82.525 196.985 ;
        RECT 86.955 197.835 87.125 198.005 ;
        RECT 86.035 197.155 86.205 197.325 ;
        RECT 88.335 197.835 88.505 198.005 ;
        RECT 87.415 196.815 87.585 196.985 ;
        RECT 89.715 197.835 89.885 198.005 ;
        RECT 88.795 196.815 88.965 196.985 ;
        RECT 91.095 198.175 91.265 198.345 ;
        RECT 90.635 196.815 90.805 196.985 ;
        RECT 92.015 196.815 92.185 196.985 ;
        RECT 92.935 197.495 93.105 197.665 ;
        RECT 93.395 197.835 93.565 198.005 ;
        RECT 93.855 197.835 94.025 198.005 ;
        RECT 94.315 197.495 94.485 197.665 ;
        RECT 95.235 197.835 95.405 198.005 ;
        RECT 97.995 198.515 98.165 198.685 ;
        RECT 97.075 197.835 97.245 198.005 ;
        RECT 96.155 196.815 96.325 196.985 ;
        RECT 98.455 197.835 98.625 198.005 ;
        RECT 99.375 197.835 99.545 198.005 ;
        RECT 98.915 196.815 99.085 196.985 ;
        RECT 103.515 197.835 103.685 198.005 ;
        RECT 102.135 197.495 102.305 197.665 ;
        RECT 104.435 198.175 104.605 198.345 ;
        RECT 102.595 196.815 102.765 196.985 ;
        RECT 104.895 197.835 105.065 198.005 ;
        RECT 108.115 198.515 108.285 198.685 ;
        RECT 105.815 197.835 105.985 198.005 ;
        RECT 106.275 197.835 106.445 198.005 ;
        RECT 106.735 197.835 106.905 198.005 ;
        RECT 115.935 198.515 116.105 198.685 ;
        RECT 114.095 197.835 114.265 198.005 ;
        RECT 115.015 197.835 115.185 198.005 ;
        RECT 113.175 196.815 113.345 196.985 ;
        RECT 116.395 197.495 116.565 197.665 ;
        RECT 117.315 197.835 117.485 198.005 ;
        RECT 118.695 197.835 118.865 198.005 ;
        RECT 118.235 197.155 118.405 197.325 ;
        RECT 126.975 198.175 127.145 198.345 ;
        RECT 134.335 198.515 134.505 198.685 ;
        RECT 123.755 197.835 123.925 198.005 ;
        RECT 122.835 196.815 123.005 196.985 ;
        RECT 124.675 197.495 124.845 197.665 ;
        RECT 126.515 197.835 126.685 198.005 ;
        RECT 127.435 197.835 127.605 198.005 ;
        RECT 130.655 197.495 130.825 197.665 ;
        RECT 132.035 197.835 132.205 198.005 ;
        RECT 132.495 197.835 132.665 198.005 ;
        RECT 132.955 197.495 133.125 197.665 ;
        RECT 132.495 196.815 132.665 196.985 ;
        RECT 135.715 197.835 135.885 198.005 ;
        RECT 134.795 197.155 134.965 197.325 ;
        RECT 143.075 198.515 143.245 198.685 ;
        RECT 137.555 197.835 137.725 198.005 ;
        RECT 138.935 197.835 139.105 198.005 ;
        RECT 136.635 196.815 136.805 196.985 ;
        RECT 138.475 197.155 138.645 197.325 ;
        RECT 140.315 197.835 140.485 198.005 ;
        RECT 139.395 196.815 139.565 196.985 ;
        RECT 142.155 197.835 142.325 198.005 ;
        RECT 141.235 197.155 141.405 197.325 ;
        RECT 146.295 198.515 146.465 198.685 ;
        RECT 145.375 197.835 145.545 198.005 ;
        RECT 147.675 197.835 147.845 198.005 ;
        RECT 146.755 196.815 146.925 196.985 ;
        RECT 152.735 197.835 152.905 198.005 ;
        RECT 152.275 196.815 152.445 196.985 ;
        RECT 154.115 197.835 154.285 198.005 ;
        RECT 153.195 197.155 153.365 197.325 ;
        RECT 70.855 196.305 71.025 196.475 ;
        RECT 71.315 196.305 71.485 196.475 ;
        RECT 71.775 196.305 71.945 196.475 ;
        RECT 72.235 196.305 72.405 196.475 ;
        RECT 72.695 196.305 72.865 196.475 ;
        RECT 73.155 196.305 73.325 196.475 ;
        RECT 73.615 196.305 73.785 196.475 ;
        RECT 74.075 196.305 74.245 196.475 ;
        RECT 74.535 196.305 74.705 196.475 ;
        RECT 74.995 196.305 75.165 196.475 ;
        RECT 75.455 196.305 75.625 196.475 ;
        RECT 75.915 196.305 76.085 196.475 ;
        RECT 76.375 196.305 76.545 196.475 ;
        RECT 76.835 196.305 77.005 196.475 ;
        RECT 77.295 196.305 77.465 196.475 ;
        RECT 77.755 196.305 77.925 196.475 ;
        RECT 78.215 196.305 78.385 196.475 ;
        RECT 78.675 196.305 78.845 196.475 ;
        RECT 79.135 196.305 79.305 196.475 ;
        RECT 79.595 196.305 79.765 196.475 ;
        RECT 80.055 196.305 80.225 196.475 ;
        RECT 80.515 196.305 80.685 196.475 ;
        RECT 80.975 196.305 81.145 196.475 ;
        RECT 81.435 196.305 81.605 196.475 ;
        RECT 81.895 196.305 82.065 196.475 ;
        RECT 82.355 196.305 82.525 196.475 ;
        RECT 82.815 196.305 82.985 196.475 ;
        RECT 83.275 196.305 83.445 196.475 ;
        RECT 83.735 196.305 83.905 196.475 ;
        RECT 84.195 196.305 84.365 196.475 ;
        RECT 84.655 196.305 84.825 196.475 ;
        RECT 85.115 196.305 85.285 196.475 ;
        RECT 85.575 196.305 85.745 196.475 ;
        RECT 86.035 196.305 86.205 196.475 ;
        RECT 86.495 196.305 86.665 196.475 ;
        RECT 86.955 196.305 87.125 196.475 ;
        RECT 87.415 196.305 87.585 196.475 ;
        RECT 87.875 196.305 88.045 196.475 ;
        RECT 88.335 196.305 88.505 196.475 ;
        RECT 88.795 196.305 88.965 196.475 ;
        RECT 89.255 196.305 89.425 196.475 ;
        RECT 89.715 196.305 89.885 196.475 ;
        RECT 90.175 196.305 90.345 196.475 ;
        RECT 90.635 196.305 90.805 196.475 ;
        RECT 91.095 196.305 91.265 196.475 ;
        RECT 91.555 196.305 91.725 196.475 ;
        RECT 92.015 196.305 92.185 196.475 ;
        RECT 92.475 196.305 92.645 196.475 ;
        RECT 92.935 196.305 93.105 196.475 ;
        RECT 93.395 196.305 93.565 196.475 ;
        RECT 93.855 196.305 94.025 196.475 ;
        RECT 94.315 196.305 94.485 196.475 ;
        RECT 94.775 196.305 94.945 196.475 ;
        RECT 95.235 196.305 95.405 196.475 ;
        RECT 95.695 196.305 95.865 196.475 ;
        RECT 96.155 196.305 96.325 196.475 ;
        RECT 96.615 196.305 96.785 196.475 ;
        RECT 97.075 196.305 97.245 196.475 ;
        RECT 97.535 196.305 97.705 196.475 ;
        RECT 97.995 196.305 98.165 196.475 ;
        RECT 98.455 196.305 98.625 196.475 ;
        RECT 98.915 196.305 99.085 196.475 ;
        RECT 99.375 196.305 99.545 196.475 ;
        RECT 99.835 196.305 100.005 196.475 ;
        RECT 100.295 196.305 100.465 196.475 ;
        RECT 100.755 196.305 100.925 196.475 ;
        RECT 101.215 196.305 101.385 196.475 ;
        RECT 101.675 196.305 101.845 196.475 ;
        RECT 102.135 196.305 102.305 196.475 ;
        RECT 102.595 196.305 102.765 196.475 ;
        RECT 103.055 196.305 103.225 196.475 ;
        RECT 103.515 196.305 103.685 196.475 ;
        RECT 103.975 196.305 104.145 196.475 ;
        RECT 104.435 196.305 104.605 196.475 ;
        RECT 104.895 196.305 105.065 196.475 ;
        RECT 105.355 196.305 105.525 196.475 ;
        RECT 105.815 196.305 105.985 196.475 ;
        RECT 106.275 196.305 106.445 196.475 ;
        RECT 106.735 196.305 106.905 196.475 ;
        RECT 107.195 196.305 107.365 196.475 ;
        RECT 107.655 196.305 107.825 196.475 ;
        RECT 108.115 196.305 108.285 196.475 ;
        RECT 108.575 196.305 108.745 196.475 ;
        RECT 109.035 196.305 109.205 196.475 ;
        RECT 109.495 196.305 109.665 196.475 ;
        RECT 109.955 196.305 110.125 196.475 ;
        RECT 110.415 196.305 110.585 196.475 ;
        RECT 110.875 196.305 111.045 196.475 ;
        RECT 111.335 196.305 111.505 196.475 ;
        RECT 111.795 196.305 111.965 196.475 ;
        RECT 112.255 196.305 112.425 196.475 ;
        RECT 112.715 196.305 112.885 196.475 ;
        RECT 113.175 196.305 113.345 196.475 ;
        RECT 113.635 196.305 113.805 196.475 ;
        RECT 114.095 196.305 114.265 196.475 ;
        RECT 114.555 196.305 114.725 196.475 ;
        RECT 115.015 196.305 115.185 196.475 ;
        RECT 115.475 196.305 115.645 196.475 ;
        RECT 115.935 196.305 116.105 196.475 ;
        RECT 116.395 196.305 116.565 196.475 ;
        RECT 116.855 196.305 117.025 196.475 ;
        RECT 117.315 196.305 117.485 196.475 ;
        RECT 117.775 196.305 117.945 196.475 ;
        RECT 118.235 196.305 118.405 196.475 ;
        RECT 118.695 196.305 118.865 196.475 ;
        RECT 119.155 196.305 119.325 196.475 ;
        RECT 119.615 196.305 119.785 196.475 ;
        RECT 120.075 196.305 120.245 196.475 ;
        RECT 120.535 196.305 120.705 196.475 ;
        RECT 120.995 196.305 121.165 196.475 ;
        RECT 121.455 196.305 121.625 196.475 ;
        RECT 121.915 196.305 122.085 196.475 ;
        RECT 122.375 196.305 122.545 196.475 ;
        RECT 122.835 196.305 123.005 196.475 ;
        RECT 123.295 196.305 123.465 196.475 ;
        RECT 123.755 196.305 123.925 196.475 ;
        RECT 124.215 196.305 124.385 196.475 ;
        RECT 124.675 196.305 124.845 196.475 ;
        RECT 125.135 196.305 125.305 196.475 ;
        RECT 125.595 196.305 125.765 196.475 ;
        RECT 126.055 196.305 126.225 196.475 ;
        RECT 126.515 196.305 126.685 196.475 ;
        RECT 126.975 196.305 127.145 196.475 ;
        RECT 127.435 196.305 127.605 196.475 ;
        RECT 127.895 196.305 128.065 196.475 ;
        RECT 128.355 196.305 128.525 196.475 ;
        RECT 128.815 196.305 128.985 196.475 ;
        RECT 129.275 196.305 129.445 196.475 ;
        RECT 129.735 196.305 129.905 196.475 ;
        RECT 130.195 196.305 130.365 196.475 ;
        RECT 130.655 196.305 130.825 196.475 ;
        RECT 131.115 196.305 131.285 196.475 ;
        RECT 131.575 196.305 131.745 196.475 ;
        RECT 132.035 196.305 132.205 196.475 ;
        RECT 132.495 196.305 132.665 196.475 ;
        RECT 132.955 196.305 133.125 196.475 ;
        RECT 133.415 196.305 133.585 196.475 ;
        RECT 133.875 196.305 134.045 196.475 ;
        RECT 134.335 196.305 134.505 196.475 ;
        RECT 134.795 196.305 134.965 196.475 ;
        RECT 135.255 196.305 135.425 196.475 ;
        RECT 135.715 196.305 135.885 196.475 ;
        RECT 136.175 196.305 136.345 196.475 ;
        RECT 136.635 196.305 136.805 196.475 ;
        RECT 137.095 196.305 137.265 196.475 ;
        RECT 137.555 196.305 137.725 196.475 ;
        RECT 138.015 196.305 138.185 196.475 ;
        RECT 138.475 196.305 138.645 196.475 ;
        RECT 138.935 196.305 139.105 196.475 ;
        RECT 139.395 196.305 139.565 196.475 ;
        RECT 139.855 196.305 140.025 196.475 ;
        RECT 140.315 196.305 140.485 196.475 ;
        RECT 140.775 196.305 140.945 196.475 ;
        RECT 141.235 196.305 141.405 196.475 ;
        RECT 141.695 196.305 141.865 196.475 ;
        RECT 142.155 196.305 142.325 196.475 ;
        RECT 142.615 196.305 142.785 196.475 ;
        RECT 143.075 196.305 143.245 196.475 ;
        RECT 143.535 196.305 143.705 196.475 ;
        RECT 143.995 196.305 144.165 196.475 ;
        RECT 144.455 196.305 144.625 196.475 ;
        RECT 144.915 196.305 145.085 196.475 ;
        RECT 145.375 196.305 145.545 196.475 ;
        RECT 145.835 196.305 146.005 196.475 ;
        RECT 146.295 196.305 146.465 196.475 ;
        RECT 146.755 196.305 146.925 196.475 ;
        RECT 147.215 196.305 147.385 196.475 ;
        RECT 147.675 196.305 147.845 196.475 ;
        RECT 148.135 196.305 148.305 196.475 ;
        RECT 148.595 196.305 148.765 196.475 ;
        RECT 149.055 196.305 149.225 196.475 ;
        RECT 149.515 196.305 149.685 196.475 ;
        RECT 149.975 196.305 150.145 196.475 ;
        RECT 150.435 196.305 150.605 196.475 ;
        RECT 150.895 196.305 151.065 196.475 ;
        RECT 151.355 196.305 151.525 196.475 ;
        RECT 151.815 196.305 151.985 196.475 ;
        RECT 152.275 196.305 152.445 196.475 ;
        RECT 152.735 196.305 152.905 196.475 ;
        RECT 153.195 196.305 153.365 196.475 ;
        RECT 153.655 196.305 153.825 196.475 ;
        RECT 154.115 196.305 154.285 196.475 ;
        RECT 154.575 196.305 154.745 196.475 ;
        RECT 155.035 196.305 155.205 196.475 ;
        RECT 155.495 196.305 155.665 196.475 ;
        RECT 155.955 196.305 156.125 196.475 ;
        RECT 72.720 195.455 72.890 195.625 ;
        RECT 72.235 194.775 72.405 194.945 ;
        RECT 73.115 195.115 73.285 195.285 ;
        RECT 73.570 194.435 73.740 194.605 ;
        RECT 74.820 195.455 74.990 195.625 ;
        RECT 74.305 195.115 74.475 195.285 ;
        RECT 76.390 195.455 76.560 195.625 ;
        RECT 76.825 195.115 76.995 195.285 ;
        RECT 79.135 195.455 79.305 195.625 ;
        RECT 81.435 195.795 81.605 195.965 ;
        RECT 82.355 195.795 82.525 195.965 ;
        RECT 84.195 195.455 84.365 195.625 ;
        RECT 82.225 194.095 82.395 194.265 ;
        RECT 83.275 194.435 83.445 194.605 ;
        RECT 85.115 194.775 85.285 194.945 ;
        RECT 85.575 195.115 85.745 195.285 ;
        RECT 86.035 194.775 86.205 194.945 ;
        RECT 86.495 194.775 86.665 194.945 ;
        RECT 87.415 194.775 87.585 194.945 ;
        RECT 88.795 195.455 88.965 195.625 ;
        RECT 88.335 194.775 88.505 194.945 ;
        RECT 89.255 194.775 89.425 194.945 ;
        RECT 89.715 194.775 89.885 194.945 ;
        RECT 91.095 194.775 91.265 194.945 ;
        RECT 92.475 195.115 92.645 195.285 ;
        RECT 93.520 195.115 93.690 195.285 ;
        RECT 94.315 194.095 94.485 194.265 ;
        RECT 95.570 194.435 95.740 194.605 ;
        RECT 96.155 195.115 96.325 195.285 ;
        RECT 94.775 194.095 94.945 194.265 ;
        RECT 96.615 194.095 96.785 194.265 ;
        RECT 97.995 194.775 98.165 194.945 ;
        RECT 98.915 195.115 99.085 195.285 ;
        RECT 105.815 195.795 105.985 195.965 ;
        RECT 103.055 194.775 103.225 194.945 ;
        RECT 102.135 194.095 102.305 194.265 ;
        RECT 103.975 194.095 104.145 194.265 ;
        RECT 104.435 194.435 104.605 194.605 ;
        RECT 104.895 194.095 105.065 194.265 ;
        RECT 107.195 195.795 107.365 195.965 ;
        RECT 109.035 195.795 109.205 195.965 ;
        RECT 106.275 194.775 106.445 194.945 ;
        RECT 107.655 194.775 107.825 194.945 ;
        RECT 110.875 195.795 111.045 195.965 ;
        RECT 111.795 195.795 111.965 195.965 ;
        RECT 109.955 194.775 110.125 194.945 ;
        RECT 110.875 194.775 111.045 194.945 ;
        RECT 124.675 194.775 124.845 194.945 ;
        RECT 124.215 194.095 124.385 194.265 ;
        RECT 125.595 194.095 125.765 194.265 ;
        RECT 127.905 195.115 128.075 195.285 ;
        RECT 128.340 195.455 128.510 195.625 ;
        RECT 129.910 195.455 130.080 195.625 ;
        RECT 130.425 195.115 130.595 195.285 ;
        RECT 131.160 194.435 131.330 194.605 ;
        RECT 131.615 195.115 131.785 195.285 ;
        RECT 132.010 195.455 132.180 195.625 ;
        RECT 132.495 194.775 132.665 194.945 ;
        RECT 136.635 195.795 136.805 195.965 ;
        RECT 133.875 194.775 134.045 194.945 ;
        RECT 135.715 194.775 135.885 194.945 ;
        RECT 132.955 194.095 133.125 194.265 ;
        RECT 138.015 195.455 138.185 195.625 ;
        RECT 137.095 194.775 137.265 194.945 ;
        RECT 139.395 194.775 139.565 194.945 ;
        RECT 141.235 195.795 141.405 195.965 ;
        RECT 141.235 194.095 141.405 194.265 ;
        RECT 142.155 194.095 142.325 194.265 ;
        RECT 147.700 195.455 147.870 195.625 ;
        RECT 145.375 194.775 145.545 194.945 ;
        RECT 147.215 195.115 147.385 195.285 ;
        RECT 146.295 194.095 146.465 194.265 ;
        RECT 148.095 195.115 148.265 195.285 ;
        RECT 148.440 194.435 148.610 194.605 ;
        RECT 149.800 195.455 149.970 195.625 ;
        RECT 149.285 195.115 149.455 195.285 ;
        RECT 151.370 195.455 151.540 195.625 ;
        RECT 151.805 195.115 151.975 195.285 ;
        RECT 154.115 194.095 154.285 194.265 ;
        RECT 70.855 193.585 71.025 193.755 ;
        RECT 71.315 193.585 71.485 193.755 ;
        RECT 71.775 193.585 71.945 193.755 ;
        RECT 72.235 193.585 72.405 193.755 ;
        RECT 72.695 193.585 72.865 193.755 ;
        RECT 73.155 193.585 73.325 193.755 ;
        RECT 73.615 193.585 73.785 193.755 ;
        RECT 74.075 193.585 74.245 193.755 ;
        RECT 74.535 193.585 74.705 193.755 ;
        RECT 74.995 193.585 75.165 193.755 ;
        RECT 75.455 193.585 75.625 193.755 ;
        RECT 75.915 193.585 76.085 193.755 ;
        RECT 76.375 193.585 76.545 193.755 ;
        RECT 76.835 193.585 77.005 193.755 ;
        RECT 77.295 193.585 77.465 193.755 ;
        RECT 77.755 193.585 77.925 193.755 ;
        RECT 78.215 193.585 78.385 193.755 ;
        RECT 78.675 193.585 78.845 193.755 ;
        RECT 79.135 193.585 79.305 193.755 ;
        RECT 79.595 193.585 79.765 193.755 ;
        RECT 80.055 193.585 80.225 193.755 ;
        RECT 80.515 193.585 80.685 193.755 ;
        RECT 80.975 193.585 81.145 193.755 ;
        RECT 81.435 193.585 81.605 193.755 ;
        RECT 81.895 193.585 82.065 193.755 ;
        RECT 82.355 193.585 82.525 193.755 ;
        RECT 82.815 193.585 82.985 193.755 ;
        RECT 83.275 193.585 83.445 193.755 ;
        RECT 83.735 193.585 83.905 193.755 ;
        RECT 84.195 193.585 84.365 193.755 ;
        RECT 84.655 193.585 84.825 193.755 ;
        RECT 85.115 193.585 85.285 193.755 ;
        RECT 85.575 193.585 85.745 193.755 ;
        RECT 86.035 193.585 86.205 193.755 ;
        RECT 86.495 193.585 86.665 193.755 ;
        RECT 86.955 193.585 87.125 193.755 ;
        RECT 87.415 193.585 87.585 193.755 ;
        RECT 87.875 193.585 88.045 193.755 ;
        RECT 88.335 193.585 88.505 193.755 ;
        RECT 88.795 193.585 88.965 193.755 ;
        RECT 89.255 193.585 89.425 193.755 ;
        RECT 89.715 193.585 89.885 193.755 ;
        RECT 90.175 193.585 90.345 193.755 ;
        RECT 90.635 193.585 90.805 193.755 ;
        RECT 91.095 193.585 91.265 193.755 ;
        RECT 91.555 193.585 91.725 193.755 ;
        RECT 92.015 193.585 92.185 193.755 ;
        RECT 92.475 193.585 92.645 193.755 ;
        RECT 92.935 193.585 93.105 193.755 ;
        RECT 93.395 193.585 93.565 193.755 ;
        RECT 93.855 193.585 94.025 193.755 ;
        RECT 94.315 193.585 94.485 193.755 ;
        RECT 94.775 193.585 94.945 193.755 ;
        RECT 95.235 193.585 95.405 193.755 ;
        RECT 95.695 193.585 95.865 193.755 ;
        RECT 96.155 193.585 96.325 193.755 ;
        RECT 96.615 193.585 96.785 193.755 ;
        RECT 97.075 193.585 97.245 193.755 ;
        RECT 97.535 193.585 97.705 193.755 ;
        RECT 97.995 193.585 98.165 193.755 ;
        RECT 98.455 193.585 98.625 193.755 ;
        RECT 98.915 193.585 99.085 193.755 ;
        RECT 99.375 193.585 99.545 193.755 ;
        RECT 99.835 193.585 100.005 193.755 ;
        RECT 100.295 193.585 100.465 193.755 ;
        RECT 100.755 193.585 100.925 193.755 ;
        RECT 101.215 193.585 101.385 193.755 ;
        RECT 101.675 193.585 101.845 193.755 ;
        RECT 102.135 193.585 102.305 193.755 ;
        RECT 102.595 193.585 102.765 193.755 ;
        RECT 103.055 193.585 103.225 193.755 ;
        RECT 103.515 193.585 103.685 193.755 ;
        RECT 103.975 193.585 104.145 193.755 ;
        RECT 104.435 193.585 104.605 193.755 ;
        RECT 104.895 193.585 105.065 193.755 ;
        RECT 105.355 193.585 105.525 193.755 ;
        RECT 105.815 193.585 105.985 193.755 ;
        RECT 106.275 193.585 106.445 193.755 ;
        RECT 106.735 193.585 106.905 193.755 ;
        RECT 107.195 193.585 107.365 193.755 ;
        RECT 107.655 193.585 107.825 193.755 ;
        RECT 108.115 193.585 108.285 193.755 ;
        RECT 108.575 193.585 108.745 193.755 ;
        RECT 109.035 193.585 109.205 193.755 ;
        RECT 109.495 193.585 109.665 193.755 ;
        RECT 109.955 193.585 110.125 193.755 ;
        RECT 110.415 193.585 110.585 193.755 ;
        RECT 110.875 193.585 111.045 193.755 ;
        RECT 111.335 193.585 111.505 193.755 ;
        RECT 111.795 193.585 111.965 193.755 ;
        RECT 112.255 193.585 112.425 193.755 ;
        RECT 112.715 193.585 112.885 193.755 ;
        RECT 113.175 193.585 113.345 193.755 ;
        RECT 113.635 193.585 113.805 193.755 ;
        RECT 114.095 193.585 114.265 193.755 ;
        RECT 114.555 193.585 114.725 193.755 ;
        RECT 115.015 193.585 115.185 193.755 ;
        RECT 115.475 193.585 115.645 193.755 ;
        RECT 115.935 193.585 116.105 193.755 ;
        RECT 116.395 193.585 116.565 193.755 ;
        RECT 116.855 193.585 117.025 193.755 ;
        RECT 117.315 193.585 117.485 193.755 ;
        RECT 117.775 193.585 117.945 193.755 ;
        RECT 118.235 193.585 118.405 193.755 ;
        RECT 118.695 193.585 118.865 193.755 ;
        RECT 119.155 193.585 119.325 193.755 ;
        RECT 119.615 193.585 119.785 193.755 ;
        RECT 120.075 193.585 120.245 193.755 ;
        RECT 120.535 193.585 120.705 193.755 ;
        RECT 120.995 193.585 121.165 193.755 ;
        RECT 121.455 193.585 121.625 193.755 ;
        RECT 121.915 193.585 122.085 193.755 ;
        RECT 122.375 193.585 122.545 193.755 ;
        RECT 122.835 193.585 123.005 193.755 ;
        RECT 123.295 193.585 123.465 193.755 ;
        RECT 123.755 193.585 123.925 193.755 ;
        RECT 124.215 193.585 124.385 193.755 ;
        RECT 124.675 193.585 124.845 193.755 ;
        RECT 125.135 193.585 125.305 193.755 ;
        RECT 125.595 193.585 125.765 193.755 ;
        RECT 126.055 193.585 126.225 193.755 ;
        RECT 126.515 193.585 126.685 193.755 ;
        RECT 126.975 193.585 127.145 193.755 ;
        RECT 127.435 193.585 127.605 193.755 ;
        RECT 127.895 193.585 128.065 193.755 ;
        RECT 128.355 193.585 128.525 193.755 ;
        RECT 128.815 193.585 128.985 193.755 ;
        RECT 129.275 193.585 129.445 193.755 ;
        RECT 129.735 193.585 129.905 193.755 ;
        RECT 130.195 193.585 130.365 193.755 ;
        RECT 130.655 193.585 130.825 193.755 ;
        RECT 131.115 193.585 131.285 193.755 ;
        RECT 131.575 193.585 131.745 193.755 ;
        RECT 132.035 193.585 132.205 193.755 ;
        RECT 132.495 193.585 132.665 193.755 ;
        RECT 132.955 193.585 133.125 193.755 ;
        RECT 133.415 193.585 133.585 193.755 ;
        RECT 133.875 193.585 134.045 193.755 ;
        RECT 134.335 193.585 134.505 193.755 ;
        RECT 134.795 193.585 134.965 193.755 ;
        RECT 135.255 193.585 135.425 193.755 ;
        RECT 135.715 193.585 135.885 193.755 ;
        RECT 136.175 193.585 136.345 193.755 ;
        RECT 136.635 193.585 136.805 193.755 ;
        RECT 137.095 193.585 137.265 193.755 ;
        RECT 137.555 193.585 137.725 193.755 ;
        RECT 138.015 193.585 138.185 193.755 ;
        RECT 138.475 193.585 138.645 193.755 ;
        RECT 138.935 193.585 139.105 193.755 ;
        RECT 139.395 193.585 139.565 193.755 ;
        RECT 139.855 193.585 140.025 193.755 ;
        RECT 140.315 193.585 140.485 193.755 ;
        RECT 140.775 193.585 140.945 193.755 ;
        RECT 141.235 193.585 141.405 193.755 ;
        RECT 141.695 193.585 141.865 193.755 ;
        RECT 142.155 193.585 142.325 193.755 ;
        RECT 142.615 193.585 142.785 193.755 ;
        RECT 143.075 193.585 143.245 193.755 ;
        RECT 143.535 193.585 143.705 193.755 ;
        RECT 143.995 193.585 144.165 193.755 ;
        RECT 144.455 193.585 144.625 193.755 ;
        RECT 144.915 193.585 145.085 193.755 ;
        RECT 145.375 193.585 145.545 193.755 ;
        RECT 145.835 193.585 146.005 193.755 ;
        RECT 146.295 193.585 146.465 193.755 ;
        RECT 146.755 193.585 146.925 193.755 ;
        RECT 147.215 193.585 147.385 193.755 ;
        RECT 147.675 193.585 147.845 193.755 ;
        RECT 148.135 193.585 148.305 193.755 ;
        RECT 148.595 193.585 148.765 193.755 ;
        RECT 149.055 193.585 149.225 193.755 ;
        RECT 149.515 193.585 149.685 193.755 ;
        RECT 149.975 193.585 150.145 193.755 ;
        RECT 150.435 193.585 150.605 193.755 ;
        RECT 150.895 193.585 151.065 193.755 ;
        RECT 151.355 193.585 151.525 193.755 ;
        RECT 151.815 193.585 151.985 193.755 ;
        RECT 152.275 193.585 152.445 193.755 ;
        RECT 152.735 193.585 152.905 193.755 ;
        RECT 153.195 193.585 153.365 193.755 ;
        RECT 153.655 193.585 153.825 193.755 ;
        RECT 154.115 193.585 154.285 193.755 ;
        RECT 154.575 193.585 154.745 193.755 ;
        RECT 155.035 193.585 155.205 193.755 ;
        RECT 155.495 193.585 155.665 193.755 ;
        RECT 155.955 193.585 156.125 193.755 ;
        RECT 77.325 193.075 77.495 193.245 ;
        RECT 76.375 192.735 76.545 192.905 ;
        RECT 76.835 192.735 77.005 192.905 ;
        RECT 75.455 191.375 75.625 191.545 ;
        RECT 76.375 192.055 76.545 192.225 ;
        RECT 77.755 192.735 77.925 192.905 ;
        RECT 80.055 193.075 80.225 193.245 ;
        RECT 78.215 192.395 78.385 192.565 ;
        RECT 80.975 192.055 81.145 192.225 ;
        RECT 81.435 192.395 81.605 192.565 ;
        RECT 81.895 192.395 82.065 192.565 ;
        RECT 82.355 192.055 82.525 192.225 ;
        RECT 89.255 193.075 89.425 193.245 ;
        RECT 86.035 192.055 86.205 192.225 ;
        RECT 87.415 192.395 87.585 192.565 ;
        RECT 88.335 192.055 88.505 192.225 ;
        RECT 89.255 192.055 89.425 192.225 ;
        RECT 90.635 192.735 90.805 192.905 ;
        RECT 91.095 192.395 91.265 192.565 ;
        RECT 89.715 191.715 89.885 191.885 ;
        RECT 90.175 191.375 90.345 191.545 ;
        RECT 91.555 191.375 91.725 191.545 ;
        RECT 92.935 192.735 93.105 192.905 ;
        RECT 92.475 191.375 92.645 191.545 ;
        RECT 94.775 192.735 94.945 192.905 ;
        RECT 94.315 192.055 94.485 192.225 ;
        RECT 93.855 191.715 94.025 191.885 ;
        RECT 94.775 191.375 94.945 191.545 ;
        RECT 95.695 191.375 95.865 191.545 ;
        RECT 98.455 192.735 98.625 192.905 ;
        RECT 97.995 192.055 98.165 192.225 ;
        RECT 100.755 192.735 100.925 192.905 ;
        RECT 97.075 191.375 97.245 191.545 ;
        RECT 105.815 193.075 105.985 193.245 ;
        RECT 102.595 192.395 102.765 192.565 ;
        RECT 103.055 192.395 103.225 192.565 ;
        RECT 104.895 192.395 105.065 192.565 ;
        RECT 104.895 191.375 105.065 191.545 ;
        RECT 106.275 192.055 106.445 192.225 ;
        RECT 107.195 192.735 107.365 192.905 ;
        RECT 107.195 192.055 107.365 192.225 ;
        RECT 108.575 192.735 108.745 192.905 ;
        RECT 109.035 192.735 109.205 192.905 ;
        RECT 107.655 191.715 107.825 191.885 ;
        RECT 108.115 191.375 108.285 191.545 ;
        RECT 109.495 191.375 109.665 191.545 ;
        RECT 110.875 192.395 111.045 192.565 ;
        RECT 110.415 191.375 110.585 191.545 ;
        RECT 113.635 193.075 113.805 193.245 ;
        RECT 112.835 192.395 113.005 192.565 ;
        RECT 112.255 192.055 112.425 192.225 ;
        RECT 115.475 192.395 115.645 192.565 ;
        RECT 111.795 191.715 111.965 191.885 ;
        RECT 112.715 191.375 112.885 191.545 ;
        RECT 116.395 191.715 116.565 191.885 ;
        RECT 119.615 192.395 119.785 192.565 ;
        RECT 120.995 192.395 121.165 192.565 ;
        RECT 122.835 192.395 123.005 192.565 ;
        RECT 120.535 192.055 120.705 192.225 ;
        RECT 118.695 191.715 118.865 191.885 ;
        RECT 120.995 191.375 121.165 191.545 ;
        RECT 123.755 191.375 123.925 191.545 ;
        RECT 127.435 192.345 127.605 192.515 ;
        RECT 128.355 192.395 128.525 192.565 ;
        RECT 126.515 191.375 126.685 191.545 ;
        RECT 128.815 191.715 128.985 191.885 ;
        RECT 130.655 193.075 130.825 193.245 ;
        RECT 132.035 192.395 132.205 192.565 ;
        RECT 130.655 191.375 130.825 191.545 ;
        RECT 131.575 191.375 131.745 191.545 ;
        RECT 137.125 193.075 137.295 193.245 ;
        RECT 136.635 192.395 136.805 192.565 ;
        RECT 137.555 192.395 137.725 192.565 ;
        RECT 138.015 192.395 138.185 192.565 ;
        RECT 139.395 192.395 139.565 192.565 ;
        RECT 132.955 191.715 133.125 191.885 ;
        RECT 139.880 191.715 140.050 191.885 ;
        RECT 140.275 192.055 140.445 192.225 ;
        RECT 140.620 192.735 140.790 192.905 ;
        RECT 141.465 192.055 141.635 192.225 ;
        RECT 141.980 191.715 142.150 191.885 ;
        RECT 143.550 191.715 143.720 191.885 ;
        RECT 143.985 192.055 144.155 192.225 ;
        RECT 147.675 192.395 147.845 192.565 ;
        RECT 146.295 191.715 146.465 191.885 ;
        RECT 146.755 191.715 146.925 191.885 ;
        RECT 70.855 190.865 71.025 191.035 ;
        RECT 71.315 190.865 71.485 191.035 ;
        RECT 71.775 190.865 71.945 191.035 ;
        RECT 72.235 190.865 72.405 191.035 ;
        RECT 72.695 190.865 72.865 191.035 ;
        RECT 73.155 190.865 73.325 191.035 ;
        RECT 73.615 190.865 73.785 191.035 ;
        RECT 74.075 190.865 74.245 191.035 ;
        RECT 74.535 190.865 74.705 191.035 ;
        RECT 74.995 190.865 75.165 191.035 ;
        RECT 75.455 190.865 75.625 191.035 ;
        RECT 75.915 190.865 76.085 191.035 ;
        RECT 76.375 190.865 76.545 191.035 ;
        RECT 76.835 190.865 77.005 191.035 ;
        RECT 77.295 190.865 77.465 191.035 ;
        RECT 77.755 190.865 77.925 191.035 ;
        RECT 78.215 190.865 78.385 191.035 ;
        RECT 78.675 190.865 78.845 191.035 ;
        RECT 79.135 190.865 79.305 191.035 ;
        RECT 79.595 190.865 79.765 191.035 ;
        RECT 80.055 190.865 80.225 191.035 ;
        RECT 80.515 190.865 80.685 191.035 ;
        RECT 80.975 190.865 81.145 191.035 ;
        RECT 81.435 190.865 81.605 191.035 ;
        RECT 81.895 190.865 82.065 191.035 ;
        RECT 82.355 190.865 82.525 191.035 ;
        RECT 82.815 190.865 82.985 191.035 ;
        RECT 83.275 190.865 83.445 191.035 ;
        RECT 83.735 190.865 83.905 191.035 ;
        RECT 84.195 190.865 84.365 191.035 ;
        RECT 84.655 190.865 84.825 191.035 ;
        RECT 85.115 190.865 85.285 191.035 ;
        RECT 85.575 190.865 85.745 191.035 ;
        RECT 86.035 190.865 86.205 191.035 ;
        RECT 86.495 190.865 86.665 191.035 ;
        RECT 86.955 190.865 87.125 191.035 ;
        RECT 87.415 190.865 87.585 191.035 ;
        RECT 87.875 190.865 88.045 191.035 ;
        RECT 88.335 190.865 88.505 191.035 ;
        RECT 88.795 190.865 88.965 191.035 ;
        RECT 89.255 190.865 89.425 191.035 ;
        RECT 89.715 190.865 89.885 191.035 ;
        RECT 90.175 190.865 90.345 191.035 ;
        RECT 90.635 190.865 90.805 191.035 ;
        RECT 91.095 190.865 91.265 191.035 ;
        RECT 91.555 190.865 91.725 191.035 ;
        RECT 92.015 190.865 92.185 191.035 ;
        RECT 92.475 190.865 92.645 191.035 ;
        RECT 92.935 190.865 93.105 191.035 ;
        RECT 93.395 190.865 93.565 191.035 ;
        RECT 93.855 190.865 94.025 191.035 ;
        RECT 94.315 190.865 94.485 191.035 ;
        RECT 94.775 190.865 94.945 191.035 ;
        RECT 95.235 190.865 95.405 191.035 ;
        RECT 95.695 190.865 95.865 191.035 ;
        RECT 96.155 190.865 96.325 191.035 ;
        RECT 96.615 190.865 96.785 191.035 ;
        RECT 97.075 190.865 97.245 191.035 ;
        RECT 97.535 190.865 97.705 191.035 ;
        RECT 97.995 190.865 98.165 191.035 ;
        RECT 98.455 190.865 98.625 191.035 ;
        RECT 98.915 190.865 99.085 191.035 ;
        RECT 99.375 190.865 99.545 191.035 ;
        RECT 99.835 190.865 100.005 191.035 ;
        RECT 100.295 190.865 100.465 191.035 ;
        RECT 100.755 190.865 100.925 191.035 ;
        RECT 101.215 190.865 101.385 191.035 ;
        RECT 101.675 190.865 101.845 191.035 ;
        RECT 102.135 190.865 102.305 191.035 ;
        RECT 102.595 190.865 102.765 191.035 ;
        RECT 103.055 190.865 103.225 191.035 ;
        RECT 103.515 190.865 103.685 191.035 ;
        RECT 103.975 190.865 104.145 191.035 ;
        RECT 104.435 190.865 104.605 191.035 ;
        RECT 104.895 190.865 105.065 191.035 ;
        RECT 105.355 190.865 105.525 191.035 ;
        RECT 105.815 190.865 105.985 191.035 ;
        RECT 106.275 190.865 106.445 191.035 ;
        RECT 106.735 190.865 106.905 191.035 ;
        RECT 107.195 190.865 107.365 191.035 ;
        RECT 107.655 190.865 107.825 191.035 ;
        RECT 108.115 190.865 108.285 191.035 ;
        RECT 108.575 190.865 108.745 191.035 ;
        RECT 109.035 190.865 109.205 191.035 ;
        RECT 109.495 190.865 109.665 191.035 ;
        RECT 109.955 190.865 110.125 191.035 ;
        RECT 110.415 190.865 110.585 191.035 ;
        RECT 110.875 190.865 111.045 191.035 ;
        RECT 111.335 190.865 111.505 191.035 ;
        RECT 111.795 190.865 111.965 191.035 ;
        RECT 112.255 190.865 112.425 191.035 ;
        RECT 112.715 190.865 112.885 191.035 ;
        RECT 113.175 190.865 113.345 191.035 ;
        RECT 113.635 190.865 113.805 191.035 ;
        RECT 114.095 190.865 114.265 191.035 ;
        RECT 114.555 190.865 114.725 191.035 ;
        RECT 115.015 190.865 115.185 191.035 ;
        RECT 115.475 190.865 115.645 191.035 ;
        RECT 115.935 190.865 116.105 191.035 ;
        RECT 116.395 190.865 116.565 191.035 ;
        RECT 116.855 190.865 117.025 191.035 ;
        RECT 117.315 190.865 117.485 191.035 ;
        RECT 117.775 190.865 117.945 191.035 ;
        RECT 118.235 190.865 118.405 191.035 ;
        RECT 118.695 190.865 118.865 191.035 ;
        RECT 119.155 190.865 119.325 191.035 ;
        RECT 119.615 190.865 119.785 191.035 ;
        RECT 120.075 190.865 120.245 191.035 ;
        RECT 120.535 190.865 120.705 191.035 ;
        RECT 120.995 190.865 121.165 191.035 ;
        RECT 121.455 190.865 121.625 191.035 ;
        RECT 121.915 190.865 122.085 191.035 ;
        RECT 122.375 190.865 122.545 191.035 ;
        RECT 122.835 190.865 123.005 191.035 ;
        RECT 123.295 190.865 123.465 191.035 ;
        RECT 123.755 190.865 123.925 191.035 ;
        RECT 124.215 190.865 124.385 191.035 ;
        RECT 124.675 190.865 124.845 191.035 ;
        RECT 125.135 190.865 125.305 191.035 ;
        RECT 125.595 190.865 125.765 191.035 ;
        RECT 126.055 190.865 126.225 191.035 ;
        RECT 126.515 190.865 126.685 191.035 ;
        RECT 126.975 190.865 127.145 191.035 ;
        RECT 127.435 190.865 127.605 191.035 ;
        RECT 127.895 190.865 128.065 191.035 ;
        RECT 128.355 190.865 128.525 191.035 ;
        RECT 128.815 190.865 128.985 191.035 ;
        RECT 129.275 190.865 129.445 191.035 ;
        RECT 129.735 190.865 129.905 191.035 ;
        RECT 130.195 190.865 130.365 191.035 ;
        RECT 130.655 190.865 130.825 191.035 ;
        RECT 131.115 190.865 131.285 191.035 ;
        RECT 131.575 190.865 131.745 191.035 ;
        RECT 132.035 190.865 132.205 191.035 ;
        RECT 132.495 190.865 132.665 191.035 ;
        RECT 132.955 190.865 133.125 191.035 ;
        RECT 133.415 190.865 133.585 191.035 ;
        RECT 133.875 190.865 134.045 191.035 ;
        RECT 134.335 190.865 134.505 191.035 ;
        RECT 134.795 190.865 134.965 191.035 ;
        RECT 135.255 190.865 135.425 191.035 ;
        RECT 135.715 190.865 135.885 191.035 ;
        RECT 136.175 190.865 136.345 191.035 ;
        RECT 136.635 190.865 136.805 191.035 ;
        RECT 137.095 190.865 137.265 191.035 ;
        RECT 137.555 190.865 137.725 191.035 ;
        RECT 138.015 190.865 138.185 191.035 ;
        RECT 138.475 190.865 138.645 191.035 ;
        RECT 138.935 190.865 139.105 191.035 ;
        RECT 139.395 190.865 139.565 191.035 ;
        RECT 139.855 190.865 140.025 191.035 ;
        RECT 140.315 190.865 140.485 191.035 ;
        RECT 140.775 190.865 140.945 191.035 ;
        RECT 141.235 190.865 141.405 191.035 ;
        RECT 141.695 190.865 141.865 191.035 ;
        RECT 142.155 190.865 142.325 191.035 ;
        RECT 142.615 190.865 142.785 191.035 ;
        RECT 143.075 190.865 143.245 191.035 ;
        RECT 143.535 190.865 143.705 191.035 ;
        RECT 143.995 190.865 144.165 191.035 ;
        RECT 144.455 190.865 144.625 191.035 ;
        RECT 144.915 190.865 145.085 191.035 ;
        RECT 145.375 190.865 145.545 191.035 ;
        RECT 145.835 190.865 146.005 191.035 ;
        RECT 146.295 190.865 146.465 191.035 ;
        RECT 146.755 190.865 146.925 191.035 ;
        RECT 147.215 190.865 147.385 191.035 ;
        RECT 147.675 190.865 147.845 191.035 ;
        RECT 148.135 190.865 148.305 191.035 ;
        RECT 148.595 190.865 148.765 191.035 ;
        RECT 149.055 190.865 149.225 191.035 ;
        RECT 149.515 190.865 149.685 191.035 ;
        RECT 149.975 190.865 150.145 191.035 ;
        RECT 150.435 190.865 150.605 191.035 ;
        RECT 150.895 190.865 151.065 191.035 ;
        RECT 151.355 190.865 151.525 191.035 ;
        RECT 151.815 190.865 151.985 191.035 ;
        RECT 152.275 190.865 152.445 191.035 ;
        RECT 152.735 190.865 152.905 191.035 ;
        RECT 153.195 190.865 153.365 191.035 ;
        RECT 153.655 190.865 153.825 191.035 ;
        RECT 154.115 190.865 154.285 191.035 ;
        RECT 154.575 190.865 154.745 191.035 ;
        RECT 155.035 190.865 155.205 191.035 ;
        RECT 155.495 190.865 155.665 191.035 ;
        RECT 155.955 190.865 156.125 191.035 ;
        RECT 80.975 190.015 81.145 190.185 ;
        RECT 82.815 189.675 82.985 189.845 ;
        RECT 81.895 189.335 82.065 189.505 ;
        RECT 84.195 189.335 84.365 189.505 ;
        RECT 86.955 190.355 87.125 190.525 ;
        RECT 85.575 189.335 85.745 189.505 ;
        RECT 86.495 189.335 86.665 189.505 ;
        RECT 85.115 188.655 85.285 188.825 ;
        RECT 86.035 188.995 86.205 189.165 ;
        RECT 87.875 189.335 88.045 189.505 ;
        RECT 88.335 189.335 88.505 189.505 ;
        RECT 88.795 189.675 88.965 189.845 ;
        RECT 89.260 189.335 89.430 189.505 ;
        RECT 90.175 189.335 90.345 189.505 ;
        RECT 92.015 190.355 92.185 190.525 ;
        RECT 91.555 189.335 91.725 189.505 ;
        RECT 92.935 189.335 93.105 189.505 ;
        RECT 94.315 189.335 94.485 189.505 ;
        RECT 95.695 189.335 95.865 189.505 ;
        RECT 96.155 189.335 96.325 189.505 ;
        RECT 91.095 188.655 91.265 188.825 ;
        RECT 98.915 189.675 99.085 189.845 ;
        RECT 99.375 189.335 99.545 189.505 ;
        RECT 101.215 190.355 101.385 190.525 ;
        RECT 101.215 189.335 101.385 189.505 ;
        RECT 102.595 189.335 102.765 189.505 ;
        RECT 102.135 188.655 102.305 188.825 ;
        RECT 103.515 188.655 103.685 188.825 ;
        RECT 103.975 190.355 104.145 190.525 ;
        RECT 104.895 190.355 105.065 190.525 ;
        RECT 104.895 189.335 105.065 189.505 ;
        RECT 106.735 189.335 106.905 189.505 ;
        RECT 107.195 189.335 107.365 189.505 ;
        RECT 109.955 190.015 110.125 190.185 ;
        RECT 115.935 190.355 116.105 190.525 ;
        RECT 115.475 190.015 115.645 190.185 ;
        RECT 110.875 189.335 111.045 189.505 ;
        RECT 112.255 189.335 112.425 189.505 ;
        RECT 114.095 189.675 114.265 189.845 ;
        RECT 115.015 189.675 115.185 189.845 ;
        RECT 113.175 188.655 113.345 188.825 ;
        RECT 117.315 190.355 117.485 190.525 ;
        RECT 115.015 188.655 115.185 188.825 ;
        RECT 116.395 188.995 116.565 189.165 ;
        RECT 116.855 189.335 117.025 189.505 ;
        RECT 118.235 190.355 118.405 190.525 ;
        RECT 120.535 190.355 120.705 190.525 ;
        RECT 118.695 188.995 118.865 189.165 ;
        RECT 119.615 190.015 119.785 190.185 ;
        RECT 121.455 190.015 121.625 190.185 ;
        RECT 120.075 189.675 120.245 189.845 ;
        RECT 123.295 190.355 123.465 190.525 ;
        RECT 120.535 188.655 120.705 188.825 ;
        RECT 123.215 188.995 123.385 189.165 ;
        RECT 122.375 188.655 122.545 188.825 ;
        RECT 124.215 188.995 124.385 189.165 ;
        RECT 126.055 189.675 126.225 189.845 ;
        RECT 125.135 188.995 125.305 189.165 ;
        RECT 127.895 190.355 128.065 190.525 ;
        RECT 127.435 189.335 127.605 189.505 ;
        RECT 126.515 188.655 126.685 188.825 ;
        RECT 128.815 189.335 128.985 189.505 ;
        RECT 129.275 189.335 129.445 189.505 ;
        RECT 130.195 188.655 130.365 188.825 ;
        RECT 132.495 189.675 132.665 189.845 ;
        RECT 130.655 189.335 130.825 189.505 ;
        RECT 131.575 189.335 131.745 189.505 ;
        RECT 136.175 190.355 136.345 190.525 ;
        RECT 135.715 189.675 135.885 189.845 ;
        RECT 133.875 189.335 134.045 189.505 ;
        RECT 136.635 189.675 136.805 189.845 ;
        RECT 137.555 190.355 137.725 190.525 ;
        RECT 137.095 189.335 137.265 189.505 ;
        RECT 132.955 188.655 133.125 188.825 ;
        RECT 140.340 190.015 140.510 190.185 ;
        RECT 138.475 188.995 138.645 189.165 ;
        RECT 139.855 189.335 140.025 189.505 ;
        RECT 139.395 188.995 139.565 189.165 ;
        RECT 140.735 189.675 140.905 189.845 ;
        RECT 141.190 189.335 141.360 189.505 ;
        RECT 142.440 190.015 142.610 190.185 ;
        RECT 141.925 189.675 142.095 189.845 ;
        RECT 144.010 190.015 144.180 190.185 ;
        RECT 144.445 189.675 144.615 189.845 ;
        RECT 146.755 190.015 146.925 190.185 ;
        RECT 148.595 189.675 148.765 189.845 ;
        RECT 148.135 189.335 148.305 189.505 ;
        RECT 149.975 189.675 150.145 189.845 ;
        RECT 151.355 190.015 151.525 190.185 ;
        RECT 152.275 189.335 152.445 189.505 ;
        RECT 153.655 189.335 153.825 189.505 ;
        RECT 152.735 188.655 152.905 188.825 ;
        RECT 70.855 188.145 71.025 188.315 ;
        RECT 71.315 188.145 71.485 188.315 ;
        RECT 71.775 188.145 71.945 188.315 ;
        RECT 72.235 188.145 72.405 188.315 ;
        RECT 72.695 188.145 72.865 188.315 ;
        RECT 73.155 188.145 73.325 188.315 ;
        RECT 73.615 188.145 73.785 188.315 ;
        RECT 74.075 188.145 74.245 188.315 ;
        RECT 74.535 188.145 74.705 188.315 ;
        RECT 74.995 188.145 75.165 188.315 ;
        RECT 75.455 188.145 75.625 188.315 ;
        RECT 75.915 188.145 76.085 188.315 ;
        RECT 76.375 188.145 76.545 188.315 ;
        RECT 76.835 188.145 77.005 188.315 ;
        RECT 77.295 188.145 77.465 188.315 ;
        RECT 77.755 188.145 77.925 188.315 ;
        RECT 78.215 188.145 78.385 188.315 ;
        RECT 78.675 188.145 78.845 188.315 ;
        RECT 79.135 188.145 79.305 188.315 ;
        RECT 79.595 188.145 79.765 188.315 ;
        RECT 80.055 188.145 80.225 188.315 ;
        RECT 80.515 188.145 80.685 188.315 ;
        RECT 80.975 188.145 81.145 188.315 ;
        RECT 81.435 188.145 81.605 188.315 ;
        RECT 81.895 188.145 82.065 188.315 ;
        RECT 82.355 188.145 82.525 188.315 ;
        RECT 82.815 188.145 82.985 188.315 ;
        RECT 83.275 188.145 83.445 188.315 ;
        RECT 83.735 188.145 83.905 188.315 ;
        RECT 84.195 188.145 84.365 188.315 ;
        RECT 84.655 188.145 84.825 188.315 ;
        RECT 85.115 188.145 85.285 188.315 ;
        RECT 85.575 188.145 85.745 188.315 ;
        RECT 86.035 188.145 86.205 188.315 ;
        RECT 86.495 188.145 86.665 188.315 ;
        RECT 86.955 188.145 87.125 188.315 ;
        RECT 87.415 188.145 87.585 188.315 ;
        RECT 87.875 188.145 88.045 188.315 ;
        RECT 88.335 188.145 88.505 188.315 ;
        RECT 88.795 188.145 88.965 188.315 ;
        RECT 89.255 188.145 89.425 188.315 ;
        RECT 89.715 188.145 89.885 188.315 ;
        RECT 90.175 188.145 90.345 188.315 ;
        RECT 90.635 188.145 90.805 188.315 ;
        RECT 91.095 188.145 91.265 188.315 ;
        RECT 91.555 188.145 91.725 188.315 ;
        RECT 92.015 188.145 92.185 188.315 ;
        RECT 92.475 188.145 92.645 188.315 ;
        RECT 92.935 188.145 93.105 188.315 ;
        RECT 93.395 188.145 93.565 188.315 ;
        RECT 93.855 188.145 94.025 188.315 ;
        RECT 94.315 188.145 94.485 188.315 ;
        RECT 94.775 188.145 94.945 188.315 ;
        RECT 95.235 188.145 95.405 188.315 ;
        RECT 95.695 188.145 95.865 188.315 ;
        RECT 96.155 188.145 96.325 188.315 ;
        RECT 96.615 188.145 96.785 188.315 ;
        RECT 97.075 188.145 97.245 188.315 ;
        RECT 97.535 188.145 97.705 188.315 ;
        RECT 97.995 188.145 98.165 188.315 ;
        RECT 98.455 188.145 98.625 188.315 ;
        RECT 98.915 188.145 99.085 188.315 ;
        RECT 99.375 188.145 99.545 188.315 ;
        RECT 99.835 188.145 100.005 188.315 ;
        RECT 100.295 188.145 100.465 188.315 ;
        RECT 100.755 188.145 100.925 188.315 ;
        RECT 101.215 188.145 101.385 188.315 ;
        RECT 101.675 188.145 101.845 188.315 ;
        RECT 102.135 188.145 102.305 188.315 ;
        RECT 102.595 188.145 102.765 188.315 ;
        RECT 103.055 188.145 103.225 188.315 ;
        RECT 103.515 188.145 103.685 188.315 ;
        RECT 103.975 188.145 104.145 188.315 ;
        RECT 104.435 188.145 104.605 188.315 ;
        RECT 104.895 188.145 105.065 188.315 ;
        RECT 105.355 188.145 105.525 188.315 ;
        RECT 105.815 188.145 105.985 188.315 ;
        RECT 106.275 188.145 106.445 188.315 ;
        RECT 106.735 188.145 106.905 188.315 ;
        RECT 107.195 188.145 107.365 188.315 ;
        RECT 107.655 188.145 107.825 188.315 ;
        RECT 108.115 188.145 108.285 188.315 ;
        RECT 108.575 188.145 108.745 188.315 ;
        RECT 109.035 188.145 109.205 188.315 ;
        RECT 109.495 188.145 109.665 188.315 ;
        RECT 109.955 188.145 110.125 188.315 ;
        RECT 110.415 188.145 110.585 188.315 ;
        RECT 110.875 188.145 111.045 188.315 ;
        RECT 111.335 188.145 111.505 188.315 ;
        RECT 111.795 188.145 111.965 188.315 ;
        RECT 112.255 188.145 112.425 188.315 ;
        RECT 112.715 188.145 112.885 188.315 ;
        RECT 113.175 188.145 113.345 188.315 ;
        RECT 113.635 188.145 113.805 188.315 ;
        RECT 114.095 188.145 114.265 188.315 ;
        RECT 114.555 188.145 114.725 188.315 ;
        RECT 115.015 188.145 115.185 188.315 ;
        RECT 115.475 188.145 115.645 188.315 ;
        RECT 115.935 188.145 116.105 188.315 ;
        RECT 116.395 188.145 116.565 188.315 ;
        RECT 116.855 188.145 117.025 188.315 ;
        RECT 117.315 188.145 117.485 188.315 ;
        RECT 117.775 188.145 117.945 188.315 ;
        RECT 118.235 188.145 118.405 188.315 ;
        RECT 118.695 188.145 118.865 188.315 ;
        RECT 119.155 188.145 119.325 188.315 ;
        RECT 119.615 188.145 119.785 188.315 ;
        RECT 120.075 188.145 120.245 188.315 ;
        RECT 120.535 188.145 120.705 188.315 ;
        RECT 120.995 188.145 121.165 188.315 ;
        RECT 121.455 188.145 121.625 188.315 ;
        RECT 121.915 188.145 122.085 188.315 ;
        RECT 122.375 188.145 122.545 188.315 ;
        RECT 122.835 188.145 123.005 188.315 ;
        RECT 123.295 188.145 123.465 188.315 ;
        RECT 123.755 188.145 123.925 188.315 ;
        RECT 124.215 188.145 124.385 188.315 ;
        RECT 124.675 188.145 124.845 188.315 ;
        RECT 125.135 188.145 125.305 188.315 ;
        RECT 125.595 188.145 125.765 188.315 ;
        RECT 126.055 188.145 126.225 188.315 ;
        RECT 126.515 188.145 126.685 188.315 ;
        RECT 126.975 188.145 127.145 188.315 ;
        RECT 127.435 188.145 127.605 188.315 ;
        RECT 127.895 188.145 128.065 188.315 ;
        RECT 128.355 188.145 128.525 188.315 ;
        RECT 128.815 188.145 128.985 188.315 ;
        RECT 129.275 188.145 129.445 188.315 ;
        RECT 129.735 188.145 129.905 188.315 ;
        RECT 130.195 188.145 130.365 188.315 ;
        RECT 130.655 188.145 130.825 188.315 ;
        RECT 131.115 188.145 131.285 188.315 ;
        RECT 131.575 188.145 131.745 188.315 ;
        RECT 132.035 188.145 132.205 188.315 ;
        RECT 132.495 188.145 132.665 188.315 ;
        RECT 132.955 188.145 133.125 188.315 ;
        RECT 133.415 188.145 133.585 188.315 ;
        RECT 133.875 188.145 134.045 188.315 ;
        RECT 134.335 188.145 134.505 188.315 ;
        RECT 134.795 188.145 134.965 188.315 ;
        RECT 135.255 188.145 135.425 188.315 ;
        RECT 135.715 188.145 135.885 188.315 ;
        RECT 136.175 188.145 136.345 188.315 ;
        RECT 136.635 188.145 136.805 188.315 ;
        RECT 137.095 188.145 137.265 188.315 ;
        RECT 137.555 188.145 137.725 188.315 ;
        RECT 138.015 188.145 138.185 188.315 ;
        RECT 138.475 188.145 138.645 188.315 ;
        RECT 138.935 188.145 139.105 188.315 ;
        RECT 139.395 188.145 139.565 188.315 ;
        RECT 139.855 188.145 140.025 188.315 ;
        RECT 140.315 188.145 140.485 188.315 ;
        RECT 140.775 188.145 140.945 188.315 ;
        RECT 141.235 188.145 141.405 188.315 ;
        RECT 141.695 188.145 141.865 188.315 ;
        RECT 142.155 188.145 142.325 188.315 ;
        RECT 142.615 188.145 142.785 188.315 ;
        RECT 143.075 188.145 143.245 188.315 ;
        RECT 143.535 188.145 143.705 188.315 ;
        RECT 143.995 188.145 144.165 188.315 ;
        RECT 144.455 188.145 144.625 188.315 ;
        RECT 144.915 188.145 145.085 188.315 ;
        RECT 145.375 188.145 145.545 188.315 ;
        RECT 145.835 188.145 146.005 188.315 ;
        RECT 146.295 188.145 146.465 188.315 ;
        RECT 146.755 188.145 146.925 188.315 ;
        RECT 147.215 188.145 147.385 188.315 ;
        RECT 147.675 188.145 147.845 188.315 ;
        RECT 148.135 188.145 148.305 188.315 ;
        RECT 148.595 188.145 148.765 188.315 ;
        RECT 149.055 188.145 149.225 188.315 ;
        RECT 149.515 188.145 149.685 188.315 ;
        RECT 149.975 188.145 150.145 188.315 ;
        RECT 150.435 188.145 150.605 188.315 ;
        RECT 150.895 188.145 151.065 188.315 ;
        RECT 151.355 188.145 151.525 188.315 ;
        RECT 151.815 188.145 151.985 188.315 ;
        RECT 152.275 188.145 152.445 188.315 ;
        RECT 152.735 188.145 152.905 188.315 ;
        RECT 153.195 188.145 153.365 188.315 ;
        RECT 153.655 188.145 153.825 188.315 ;
        RECT 154.115 188.145 154.285 188.315 ;
        RECT 154.575 188.145 154.745 188.315 ;
        RECT 155.035 188.145 155.205 188.315 ;
        RECT 155.495 188.145 155.665 188.315 ;
        RECT 155.955 188.145 156.125 188.315 ;
        RECT 72.695 186.615 72.865 186.785 ;
        RECT 73.180 186.275 73.350 186.445 ;
        RECT 73.575 186.615 73.745 186.785 ;
        RECT 74.030 186.955 74.200 187.125 ;
        RECT 74.765 186.615 74.935 186.785 ;
        RECT 75.280 186.275 75.450 186.445 ;
        RECT 76.850 186.275 77.020 186.445 ;
        RECT 77.285 186.615 77.455 186.785 ;
        RECT 80.975 186.875 81.145 187.045 ;
        RECT 79.595 185.935 79.765 186.105 ;
        RECT 80.055 185.935 80.225 186.105 ;
        RECT 82.275 187.295 82.445 187.465 ;
        RECT 84.655 187.635 84.825 187.805 ;
        RECT 83.275 187.295 83.445 187.465 ;
        RECT 83.735 186.955 83.905 187.125 ;
        RECT 86.035 187.635 86.205 187.805 ;
        RECT 85.115 186.955 85.285 187.125 ;
        RECT 81.435 185.935 81.605 186.105 ;
        RECT 82.355 185.935 82.525 186.105 ;
        RECT 87.415 187.635 87.585 187.805 ;
        RECT 88.335 186.955 88.505 187.125 ;
        RECT 89.255 187.295 89.425 187.465 ;
        RECT 90.635 186.955 90.805 187.125 ;
        RECT 91.555 185.935 91.725 186.105 ;
        RECT 97.075 187.635 97.245 187.805 ;
        RECT 94.775 186.615 94.945 186.785 ;
        RECT 96.155 186.955 96.325 187.125 ;
        RECT 97.995 186.955 98.165 187.125 ;
        RECT 99.835 186.615 100.005 186.785 ;
        RECT 100.755 187.295 100.925 187.465 ;
        RECT 100.755 186.615 100.925 186.785 ;
        RECT 102.135 187.295 102.305 187.465 ;
        RECT 102.595 186.955 102.765 187.125 ;
        RECT 101.215 186.275 101.385 186.445 ;
        RECT 101.675 185.935 101.845 186.105 ;
        RECT 103.055 185.935 103.225 186.105 ;
        RECT 104.435 187.295 104.605 187.465 ;
        RECT 106.275 187.635 106.445 187.805 ;
        RECT 103.975 185.935 104.145 186.105 ;
        RECT 105.815 186.615 105.985 186.785 ;
        RECT 105.355 186.275 105.525 186.445 ;
        RECT 106.275 185.935 106.445 186.105 ;
        RECT 107.195 185.935 107.365 186.105 ;
        RECT 108.115 186.615 108.285 186.785 ;
        RECT 109.035 187.295 109.205 187.465 ;
        RECT 109.035 186.615 109.205 186.785 ;
        RECT 110.415 186.955 110.585 187.125 ;
        RECT 110.875 186.955 111.045 187.125 ;
        RECT 109.495 186.275 109.665 186.445 ;
        RECT 109.955 185.935 110.125 186.105 ;
        RECT 111.335 185.935 111.505 186.105 ;
        RECT 112.715 186.955 112.885 187.125 ;
        RECT 112.255 185.935 112.425 186.105 ;
        RECT 114.555 187.295 114.725 187.465 ;
        RECT 115.475 187.635 115.645 187.805 ;
        RECT 114.095 186.615 114.265 186.785 ;
        RECT 116.395 187.635 116.565 187.805 ;
        RECT 113.635 186.275 113.805 186.445 ;
        RECT 114.555 185.935 114.725 186.105 ;
        RECT 121.455 187.635 121.625 187.805 ;
        RECT 117.315 186.955 117.485 187.125 ;
        RECT 118.695 186.955 118.865 187.125 ;
        RECT 118.235 186.615 118.405 186.785 ;
        RECT 120.535 186.955 120.705 187.125 ;
        RECT 123.755 186.955 123.925 187.125 ;
        RECT 124.675 186.955 124.845 187.125 ;
        RECT 132.035 187.635 132.205 187.805 ;
        RECT 122.835 186.275 123.005 186.445 ;
        RECT 133.875 186.615 134.045 186.785 ;
        RECT 134.795 187.295 134.965 187.465 ;
        RECT 134.795 186.615 134.965 186.785 ;
        RECT 136.175 186.955 136.345 187.125 ;
        RECT 136.635 187.295 136.805 187.465 ;
        RECT 135.255 186.275 135.425 186.445 ;
        RECT 135.715 185.935 135.885 186.105 ;
        RECT 137.095 185.935 137.265 186.105 ;
        RECT 138.475 186.955 138.645 187.125 ;
        RECT 138.015 185.935 138.185 186.105 ;
        RECT 140.315 187.295 140.485 187.465 ;
        RECT 139.855 186.615 140.025 186.785 ;
        RECT 139.395 186.275 139.565 186.445 ;
        RECT 140.315 185.935 140.485 186.105 ;
        RECT 141.235 185.935 141.405 186.105 ;
        RECT 142.155 186.615 142.325 186.785 ;
        RECT 143.535 186.615 143.705 186.785 ;
        RECT 146.755 187.635 146.925 187.805 ;
        RECT 147.675 186.955 147.845 187.125 ;
        RECT 149.515 186.955 149.685 187.125 ;
        RECT 150.435 186.615 150.605 186.785 ;
        RECT 152.275 187.635 152.445 187.805 ;
        RECT 151.815 186.955 151.985 187.125 ;
        RECT 148.595 185.935 148.765 186.105 ;
        RECT 150.895 186.275 151.065 186.445 ;
        RECT 153.195 186.955 153.365 187.125 ;
        RECT 154.575 186.955 154.745 187.125 ;
        RECT 153.655 185.935 153.825 186.105 ;
        RECT 70.855 185.425 71.025 185.595 ;
        RECT 71.315 185.425 71.485 185.595 ;
        RECT 71.775 185.425 71.945 185.595 ;
        RECT 72.235 185.425 72.405 185.595 ;
        RECT 72.695 185.425 72.865 185.595 ;
        RECT 73.155 185.425 73.325 185.595 ;
        RECT 73.615 185.425 73.785 185.595 ;
        RECT 74.075 185.425 74.245 185.595 ;
        RECT 74.535 185.425 74.705 185.595 ;
        RECT 74.995 185.425 75.165 185.595 ;
        RECT 75.455 185.425 75.625 185.595 ;
        RECT 75.915 185.425 76.085 185.595 ;
        RECT 76.375 185.425 76.545 185.595 ;
        RECT 76.835 185.425 77.005 185.595 ;
        RECT 77.295 185.425 77.465 185.595 ;
        RECT 77.755 185.425 77.925 185.595 ;
        RECT 78.215 185.425 78.385 185.595 ;
        RECT 78.675 185.425 78.845 185.595 ;
        RECT 79.135 185.425 79.305 185.595 ;
        RECT 79.595 185.425 79.765 185.595 ;
        RECT 80.055 185.425 80.225 185.595 ;
        RECT 80.515 185.425 80.685 185.595 ;
        RECT 80.975 185.425 81.145 185.595 ;
        RECT 81.435 185.425 81.605 185.595 ;
        RECT 81.895 185.425 82.065 185.595 ;
        RECT 82.355 185.425 82.525 185.595 ;
        RECT 82.815 185.425 82.985 185.595 ;
        RECT 83.275 185.425 83.445 185.595 ;
        RECT 83.735 185.425 83.905 185.595 ;
        RECT 84.195 185.425 84.365 185.595 ;
        RECT 84.655 185.425 84.825 185.595 ;
        RECT 85.115 185.425 85.285 185.595 ;
        RECT 85.575 185.425 85.745 185.595 ;
        RECT 86.035 185.425 86.205 185.595 ;
        RECT 86.495 185.425 86.665 185.595 ;
        RECT 86.955 185.425 87.125 185.595 ;
        RECT 87.415 185.425 87.585 185.595 ;
        RECT 87.875 185.425 88.045 185.595 ;
        RECT 88.335 185.425 88.505 185.595 ;
        RECT 88.795 185.425 88.965 185.595 ;
        RECT 89.255 185.425 89.425 185.595 ;
        RECT 89.715 185.425 89.885 185.595 ;
        RECT 90.175 185.425 90.345 185.595 ;
        RECT 90.635 185.425 90.805 185.595 ;
        RECT 91.095 185.425 91.265 185.595 ;
        RECT 91.555 185.425 91.725 185.595 ;
        RECT 92.015 185.425 92.185 185.595 ;
        RECT 92.475 185.425 92.645 185.595 ;
        RECT 92.935 185.425 93.105 185.595 ;
        RECT 93.395 185.425 93.565 185.595 ;
        RECT 93.855 185.425 94.025 185.595 ;
        RECT 94.315 185.425 94.485 185.595 ;
        RECT 94.775 185.425 94.945 185.595 ;
        RECT 95.235 185.425 95.405 185.595 ;
        RECT 95.695 185.425 95.865 185.595 ;
        RECT 96.155 185.425 96.325 185.595 ;
        RECT 96.615 185.425 96.785 185.595 ;
        RECT 97.075 185.425 97.245 185.595 ;
        RECT 97.535 185.425 97.705 185.595 ;
        RECT 97.995 185.425 98.165 185.595 ;
        RECT 98.455 185.425 98.625 185.595 ;
        RECT 98.915 185.425 99.085 185.595 ;
        RECT 99.375 185.425 99.545 185.595 ;
        RECT 99.835 185.425 100.005 185.595 ;
        RECT 100.295 185.425 100.465 185.595 ;
        RECT 100.755 185.425 100.925 185.595 ;
        RECT 101.215 185.425 101.385 185.595 ;
        RECT 101.675 185.425 101.845 185.595 ;
        RECT 102.135 185.425 102.305 185.595 ;
        RECT 102.595 185.425 102.765 185.595 ;
        RECT 103.055 185.425 103.225 185.595 ;
        RECT 103.515 185.425 103.685 185.595 ;
        RECT 103.975 185.425 104.145 185.595 ;
        RECT 104.435 185.425 104.605 185.595 ;
        RECT 104.895 185.425 105.065 185.595 ;
        RECT 105.355 185.425 105.525 185.595 ;
        RECT 105.815 185.425 105.985 185.595 ;
        RECT 106.275 185.425 106.445 185.595 ;
        RECT 106.735 185.425 106.905 185.595 ;
        RECT 107.195 185.425 107.365 185.595 ;
        RECT 107.655 185.425 107.825 185.595 ;
        RECT 108.115 185.425 108.285 185.595 ;
        RECT 108.575 185.425 108.745 185.595 ;
        RECT 109.035 185.425 109.205 185.595 ;
        RECT 109.495 185.425 109.665 185.595 ;
        RECT 109.955 185.425 110.125 185.595 ;
        RECT 110.415 185.425 110.585 185.595 ;
        RECT 110.875 185.425 111.045 185.595 ;
        RECT 111.335 185.425 111.505 185.595 ;
        RECT 111.795 185.425 111.965 185.595 ;
        RECT 112.255 185.425 112.425 185.595 ;
        RECT 112.715 185.425 112.885 185.595 ;
        RECT 113.175 185.425 113.345 185.595 ;
        RECT 113.635 185.425 113.805 185.595 ;
        RECT 114.095 185.425 114.265 185.595 ;
        RECT 114.555 185.425 114.725 185.595 ;
        RECT 115.015 185.425 115.185 185.595 ;
        RECT 115.475 185.425 115.645 185.595 ;
        RECT 115.935 185.425 116.105 185.595 ;
        RECT 116.395 185.425 116.565 185.595 ;
        RECT 116.855 185.425 117.025 185.595 ;
        RECT 117.315 185.425 117.485 185.595 ;
        RECT 117.775 185.425 117.945 185.595 ;
        RECT 118.235 185.425 118.405 185.595 ;
        RECT 118.695 185.425 118.865 185.595 ;
        RECT 119.155 185.425 119.325 185.595 ;
        RECT 119.615 185.425 119.785 185.595 ;
        RECT 120.075 185.425 120.245 185.595 ;
        RECT 120.535 185.425 120.705 185.595 ;
        RECT 120.995 185.425 121.165 185.595 ;
        RECT 121.455 185.425 121.625 185.595 ;
        RECT 121.915 185.425 122.085 185.595 ;
        RECT 122.375 185.425 122.545 185.595 ;
        RECT 122.835 185.425 123.005 185.595 ;
        RECT 123.295 185.425 123.465 185.595 ;
        RECT 123.755 185.425 123.925 185.595 ;
        RECT 124.215 185.425 124.385 185.595 ;
        RECT 124.675 185.425 124.845 185.595 ;
        RECT 125.135 185.425 125.305 185.595 ;
        RECT 125.595 185.425 125.765 185.595 ;
        RECT 126.055 185.425 126.225 185.595 ;
        RECT 126.515 185.425 126.685 185.595 ;
        RECT 126.975 185.425 127.145 185.595 ;
        RECT 127.435 185.425 127.605 185.595 ;
        RECT 127.895 185.425 128.065 185.595 ;
        RECT 128.355 185.425 128.525 185.595 ;
        RECT 128.815 185.425 128.985 185.595 ;
        RECT 129.275 185.425 129.445 185.595 ;
        RECT 129.735 185.425 129.905 185.595 ;
        RECT 130.195 185.425 130.365 185.595 ;
        RECT 130.655 185.425 130.825 185.595 ;
        RECT 131.115 185.425 131.285 185.595 ;
        RECT 131.575 185.425 131.745 185.595 ;
        RECT 132.035 185.425 132.205 185.595 ;
        RECT 132.495 185.425 132.665 185.595 ;
        RECT 132.955 185.425 133.125 185.595 ;
        RECT 133.415 185.425 133.585 185.595 ;
        RECT 133.875 185.425 134.045 185.595 ;
        RECT 134.335 185.425 134.505 185.595 ;
        RECT 134.795 185.425 134.965 185.595 ;
        RECT 135.255 185.425 135.425 185.595 ;
        RECT 135.715 185.425 135.885 185.595 ;
        RECT 136.175 185.425 136.345 185.595 ;
        RECT 136.635 185.425 136.805 185.595 ;
        RECT 137.095 185.425 137.265 185.595 ;
        RECT 137.555 185.425 137.725 185.595 ;
        RECT 138.015 185.425 138.185 185.595 ;
        RECT 138.475 185.425 138.645 185.595 ;
        RECT 138.935 185.425 139.105 185.595 ;
        RECT 139.395 185.425 139.565 185.595 ;
        RECT 139.855 185.425 140.025 185.595 ;
        RECT 140.315 185.425 140.485 185.595 ;
        RECT 140.775 185.425 140.945 185.595 ;
        RECT 141.235 185.425 141.405 185.595 ;
        RECT 141.695 185.425 141.865 185.595 ;
        RECT 142.155 185.425 142.325 185.595 ;
        RECT 142.615 185.425 142.785 185.595 ;
        RECT 143.075 185.425 143.245 185.595 ;
        RECT 143.535 185.425 143.705 185.595 ;
        RECT 143.995 185.425 144.165 185.595 ;
        RECT 144.455 185.425 144.625 185.595 ;
        RECT 144.915 185.425 145.085 185.595 ;
        RECT 145.375 185.425 145.545 185.595 ;
        RECT 145.835 185.425 146.005 185.595 ;
        RECT 146.295 185.425 146.465 185.595 ;
        RECT 146.755 185.425 146.925 185.595 ;
        RECT 147.215 185.425 147.385 185.595 ;
        RECT 147.675 185.425 147.845 185.595 ;
        RECT 148.135 185.425 148.305 185.595 ;
        RECT 148.595 185.425 148.765 185.595 ;
        RECT 149.055 185.425 149.225 185.595 ;
        RECT 149.515 185.425 149.685 185.595 ;
        RECT 149.975 185.425 150.145 185.595 ;
        RECT 150.435 185.425 150.605 185.595 ;
        RECT 150.895 185.425 151.065 185.595 ;
        RECT 151.355 185.425 151.525 185.595 ;
        RECT 151.815 185.425 151.985 185.595 ;
        RECT 152.275 185.425 152.445 185.595 ;
        RECT 152.735 185.425 152.905 185.595 ;
        RECT 153.195 185.425 153.365 185.595 ;
        RECT 153.655 185.425 153.825 185.595 ;
        RECT 154.115 185.425 154.285 185.595 ;
        RECT 154.575 185.425 154.745 185.595 ;
        RECT 155.035 185.425 155.205 185.595 ;
        RECT 155.495 185.425 155.665 185.595 ;
        RECT 155.955 185.425 156.125 185.595 ;
        RECT 74.535 184.915 74.705 185.085 ;
        RECT 74.535 183.895 74.705 184.065 ;
        RECT 75.915 184.235 76.085 184.405 ;
        RECT 75.455 183.895 75.625 184.065 ;
        RECT 76.835 183.895 77.005 184.065 ;
        RECT 77.295 183.895 77.465 184.065 ;
        RECT 80.515 183.895 80.685 184.065 ;
        RECT 82.355 184.915 82.525 185.085 ;
        RECT 84.680 184.575 84.850 184.745 ;
        RECT 84.195 183.895 84.365 184.065 ;
        RECT 82.355 183.215 82.525 183.385 ;
        RECT 83.275 183.215 83.445 183.385 ;
        RECT 85.075 184.235 85.245 184.405 ;
        RECT 85.530 183.555 85.700 183.725 ;
        RECT 86.780 184.575 86.950 184.745 ;
        RECT 86.265 184.235 86.435 184.405 ;
        RECT 88.350 184.575 88.520 184.745 ;
        RECT 88.785 184.235 88.955 184.405 ;
        RECT 91.095 184.575 91.265 184.745 ;
        RECT 93.855 184.235 94.025 184.405 ;
        RECT 93.395 183.895 93.565 184.065 ;
        RECT 95.235 183.895 95.405 184.065 ;
        RECT 92.475 183.215 92.645 183.385 ;
        RECT 98.455 184.915 98.625 185.085 ;
        RECT 100.755 184.235 100.925 184.405 ;
        RECT 101.215 184.235 101.385 184.405 ;
        RECT 103.515 184.915 103.685 185.085 ;
        RECT 102.595 183.895 102.765 184.065 ;
        RECT 110.875 183.555 111.045 183.725 ;
        RECT 110.415 183.215 110.585 183.385 ;
        RECT 118.695 184.915 118.865 185.085 ;
        RECT 118.235 184.575 118.405 184.745 ;
        RECT 116.855 184.235 117.025 184.405 ;
        RECT 116.395 183.895 116.565 184.065 ;
        RECT 117.775 184.235 117.945 184.405 ;
        RECT 115.475 183.215 115.645 183.385 ;
        RECT 120.075 184.915 120.245 185.085 ;
        RECT 117.775 183.555 117.945 183.725 ;
        RECT 119.155 183.555 119.325 183.725 ;
        RECT 119.615 183.555 119.785 183.725 ;
        RECT 120.995 184.915 121.165 185.085 ;
        RECT 123.295 184.915 123.465 185.085 ;
        RECT 121.455 183.895 121.625 184.065 ;
        RECT 122.375 184.575 122.545 184.745 ;
        RECT 122.835 184.235 123.005 184.405 ;
        RECT 123.415 183.895 123.585 184.065 ;
        RECT 124.215 183.215 124.385 183.385 ;
        RECT 127.435 184.575 127.605 184.745 ;
        RECT 126.515 183.895 126.685 184.065 ;
        RECT 127.895 184.915 128.065 185.085 ;
        RECT 130.195 184.235 130.365 184.405 ;
        RECT 128.815 183.775 128.985 183.945 ;
        RECT 131.115 183.895 131.285 184.065 ;
        RECT 131.575 183.895 131.745 184.065 ;
        RECT 132.035 184.235 132.205 184.405 ;
        RECT 132.495 184.235 132.665 184.405 ;
        RECT 136.635 183.895 136.805 184.065 ;
        RECT 137.095 183.895 137.265 184.065 ;
        RECT 138.475 183.895 138.645 184.065 ;
        RECT 142.155 183.895 142.325 184.065 ;
        RECT 143.535 184.235 143.705 184.405 ;
        RECT 147.700 184.575 147.870 184.745 ;
        RECT 147.215 183.895 147.385 184.065 ;
        RECT 135.715 183.215 135.885 183.385 ;
        RECT 148.095 184.235 148.265 184.405 ;
        RECT 148.550 183.895 148.720 184.065 ;
        RECT 149.800 184.575 149.970 184.745 ;
        RECT 149.285 184.235 149.455 184.405 ;
        RECT 151.370 184.575 151.540 184.745 ;
        RECT 151.805 184.235 151.975 184.405 ;
        RECT 154.115 184.915 154.285 185.085 ;
        RECT 70.855 182.705 71.025 182.875 ;
        RECT 71.315 182.705 71.485 182.875 ;
        RECT 71.775 182.705 71.945 182.875 ;
        RECT 72.235 182.705 72.405 182.875 ;
        RECT 72.695 182.705 72.865 182.875 ;
        RECT 73.155 182.705 73.325 182.875 ;
        RECT 73.615 182.705 73.785 182.875 ;
        RECT 74.075 182.705 74.245 182.875 ;
        RECT 74.535 182.705 74.705 182.875 ;
        RECT 74.995 182.705 75.165 182.875 ;
        RECT 75.455 182.705 75.625 182.875 ;
        RECT 75.915 182.705 76.085 182.875 ;
        RECT 76.375 182.705 76.545 182.875 ;
        RECT 76.835 182.705 77.005 182.875 ;
        RECT 77.295 182.705 77.465 182.875 ;
        RECT 77.755 182.705 77.925 182.875 ;
        RECT 78.215 182.705 78.385 182.875 ;
        RECT 78.675 182.705 78.845 182.875 ;
        RECT 79.135 182.705 79.305 182.875 ;
        RECT 79.595 182.705 79.765 182.875 ;
        RECT 80.055 182.705 80.225 182.875 ;
        RECT 80.515 182.705 80.685 182.875 ;
        RECT 80.975 182.705 81.145 182.875 ;
        RECT 81.435 182.705 81.605 182.875 ;
        RECT 81.895 182.705 82.065 182.875 ;
        RECT 82.355 182.705 82.525 182.875 ;
        RECT 82.815 182.705 82.985 182.875 ;
        RECT 83.275 182.705 83.445 182.875 ;
        RECT 83.735 182.705 83.905 182.875 ;
        RECT 84.195 182.705 84.365 182.875 ;
        RECT 84.655 182.705 84.825 182.875 ;
        RECT 85.115 182.705 85.285 182.875 ;
        RECT 85.575 182.705 85.745 182.875 ;
        RECT 86.035 182.705 86.205 182.875 ;
        RECT 86.495 182.705 86.665 182.875 ;
        RECT 86.955 182.705 87.125 182.875 ;
        RECT 87.415 182.705 87.585 182.875 ;
        RECT 87.875 182.705 88.045 182.875 ;
        RECT 88.335 182.705 88.505 182.875 ;
        RECT 88.795 182.705 88.965 182.875 ;
        RECT 89.255 182.705 89.425 182.875 ;
        RECT 89.715 182.705 89.885 182.875 ;
        RECT 90.175 182.705 90.345 182.875 ;
        RECT 90.635 182.705 90.805 182.875 ;
        RECT 91.095 182.705 91.265 182.875 ;
        RECT 91.555 182.705 91.725 182.875 ;
        RECT 92.015 182.705 92.185 182.875 ;
        RECT 92.475 182.705 92.645 182.875 ;
        RECT 92.935 182.705 93.105 182.875 ;
        RECT 93.395 182.705 93.565 182.875 ;
        RECT 93.855 182.705 94.025 182.875 ;
        RECT 94.315 182.705 94.485 182.875 ;
        RECT 94.775 182.705 94.945 182.875 ;
        RECT 95.235 182.705 95.405 182.875 ;
        RECT 95.695 182.705 95.865 182.875 ;
        RECT 96.155 182.705 96.325 182.875 ;
        RECT 96.615 182.705 96.785 182.875 ;
        RECT 97.075 182.705 97.245 182.875 ;
        RECT 97.535 182.705 97.705 182.875 ;
        RECT 97.995 182.705 98.165 182.875 ;
        RECT 98.455 182.705 98.625 182.875 ;
        RECT 98.915 182.705 99.085 182.875 ;
        RECT 99.375 182.705 99.545 182.875 ;
        RECT 99.835 182.705 100.005 182.875 ;
        RECT 100.295 182.705 100.465 182.875 ;
        RECT 100.755 182.705 100.925 182.875 ;
        RECT 101.215 182.705 101.385 182.875 ;
        RECT 101.675 182.705 101.845 182.875 ;
        RECT 102.135 182.705 102.305 182.875 ;
        RECT 102.595 182.705 102.765 182.875 ;
        RECT 103.055 182.705 103.225 182.875 ;
        RECT 103.515 182.705 103.685 182.875 ;
        RECT 103.975 182.705 104.145 182.875 ;
        RECT 104.435 182.705 104.605 182.875 ;
        RECT 104.895 182.705 105.065 182.875 ;
        RECT 105.355 182.705 105.525 182.875 ;
        RECT 105.815 182.705 105.985 182.875 ;
        RECT 106.275 182.705 106.445 182.875 ;
        RECT 106.735 182.705 106.905 182.875 ;
        RECT 107.195 182.705 107.365 182.875 ;
        RECT 107.655 182.705 107.825 182.875 ;
        RECT 108.115 182.705 108.285 182.875 ;
        RECT 108.575 182.705 108.745 182.875 ;
        RECT 109.035 182.705 109.205 182.875 ;
        RECT 109.495 182.705 109.665 182.875 ;
        RECT 109.955 182.705 110.125 182.875 ;
        RECT 110.415 182.705 110.585 182.875 ;
        RECT 110.875 182.705 111.045 182.875 ;
        RECT 111.335 182.705 111.505 182.875 ;
        RECT 111.795 182.705 111.965 182.875 ;
        RECT 112.255 182.705 112.425 182.875 ;
        RECT 112.715 182.705 112.885 182.875 ;
        RECT 113.175 182.705 113.345 182.875 ;
        RECT 113.635 182.705 113.805 182.875 ;
        RECT 114.095 182.705 114.265 182.875 ;
        RECT 114.555 182.705 114.725 182.875 ;
        RECT 115.015 182.705 115.185 182.875 ;
        RECT 115.475 182.705 115.645 182.875 ;
        RECT 115.935 182.705 116.105 182.875 ;
        RECT 116.395 182.705 116.565 182.875 ;
        RECT 116.855 182.705 117.025 182.875 ;
        RECT 117.315 182.705 117.485 182.875 ;
        RECT 117.775 182.705 117.945 182.875 ;
        RECT 118.235 182.705 118.405 182.875 ;
        RECT 118.695 182.705 118.865 182.875 ;
        RECT 119.155 182.705 119.325 182.875 ;
        RECT 119.615 182.705 119.785 182.875 ;
        RECT 120.075 182.705 120.245 182.875 ;
        RECT 120.535 182.705 120.705 182.875 ;
        RECT 120.995 182.705 121.165 182.875 ;
        RECT 121.455 182.705 121.625 182.875 ;
        RECT 121.915 182.705 122.085 182.875 ;
        RECT 122.375 182.705 122.545 182.875 ;
        RECT 122.835 182.705 123.005 182.875 ;
        RECT 123.295 182.705 123.465 182.875 ;
        RECT 123.755 182.705 123.925 182.875 ;
        RECT 124.215 182.705 124.385 182.875 ;
        RECT 124.675 182.705 124.845 182.875 ;
        RECT 125.135 182.705 125.305 182.875 ;
        RECT 125.595 182.705 125.765 182.875 ;
        RECT 126.055 182.705 126.225 182.875 ;
        RECT 126.515 182.705 126.685 182.875 ;
        RECT 126.975 182.705 127.145 182.875 ;
        RECT 127.435 182.705 127.605 182.875 ;
        RECT 127.895 182.705 128.065 182.875 ;
        RECT 128.355 182.705 128.525 182.875 ;
        RECT 128.815 182.705 128.985 182.875 ;
        RECT 129.275 182.705 129.445 182.875 ;
        RECT 129.735 182.705 129.905 182.875 ;
        RECT 130.195 182.705 130.365 182.875 ;
        RECT 130.655 182.705 130.825 182.875 ;
        RECT 131.115 182.705 131.285 182.875 ;
        RECT 131.575 182.705 131.745 182.875 ;
        RECT 132.035 182.705 132.205 182.875 ;
        RECT 132.495 182.705 132.665 182.875 ;
        RECT 132.955 182.705 133.125 182.875 ;
        RECT 133.415 182.705 133.585 182.875 ;
        RECT 133.875 182.705 134.045 182.875 ;
        RECT 134.335 182.705 134.505 182.875 ;
        RECT 134.795 182.705 134.965 182.875 ;
        RECT 135.255 182.705 135.425 182.875 ;
        RECT 135.715 182.705 135.885 182.875 ;
        RECT 136.175 182.705 136.345 182.875 ;
        RECT 136.635 182.705 136.805 182.875 ;
        RECT 137.095 182.705 137.265 182.875 ;
        RECT 137.555 182.705 137.725 182.875 ;
        RECT 138.015 182.705 138.185 182.875 ;
        RECT 138.475 182.705 138.645 182.875 ;
        RECT 138.935 182.705 139.105 182.875 ;
        RECT 139.395 182.705 139.565 182.875 ;
        RECT 139.855 182.705 140.025 182.875 ;
        RECT 140.315 182.705 140.485 182.875 ;
        RECT 140.775 182.705 140.945 182.875 ;
        RECT 141.235 182.705 141.405 182.875 ;
        RECT 141.695 182.705 141.865 182.875 ;
        RECT 142.155 182.705 142.325 182.875 ;
        RECT 142.615 182.705 142.785 182.875 ;
        RECT 143.075 182.705 143.245 182.875 ;
        RECT 143.535 182.705 143.705 182.875 ;
        RECT 143.995 182.705 144.165 182.875 ;
        RECT 144.455 182.705 144.625 182.875 ;
        RECT 144.915 182.705 145.085 182.875 ;
        RECT 145.375 182.705 145.545 182.875 ;
        RECT 145.835 182.705 146.005 182.875 ;
        RECT 146.295 182.705 146.465 182.875 ;
        RECT 146.755 182.705 146.925 182.875 ;
        RECT 147.215 182.705 147.385 182.875 ;
        RECT 147.675 182.705 147.845 182.875 ;
        RECT 148.135 182.705 148.305 182.875 ;
        RECT 148.595 182.705 148.765 182.875 ;
        RECT 149.055 182.705 149.225 182.875 ;
        RECT 149.515 182.705 149.685 182.875 ;
        RECT 149.975 182.705 150.145 182.875 ;
        RECT 150.435 182.705 150.605 182.875 ;
        RECT 150.895 182.705 151.065 182.875 ;
        RECT 151.355 182.705 151.525 182.875 ;
        RECT 151.815 182.705 151.985 182.875 ;
        RECT 152.275 182.705 152.445 182.875 ;
        RECT 152.735 182.705 152.905 182.875 ;
        RECT 153.195 182.705 153.365 182.875 ;
        RECT 153.655 182.705 153.825 182.875 ;
        RECT 154.115 182.705 154.285 182.875 ;
        RECT 154.575 182.705 154.745 182.875 ;
        RECT 155.035 182.705 155.205 182.875 ;
        RECT 155.495 182.705 155.665 182.875 ;
        RECT 155.955 182.705 156.125 182.875 ;
        RECT 72.235 181.175 72.405 181.345 ;
        RECT 72.720 180.835 72.890 181.005 ;
        RECT 73.115 181.175 73.285 181.345 ;
        RECT 73.570 181.515 73.740 181.685 ;
        RECT 74.305 181.175 74.475 181.345 ;
        RECT 74.820 180.835 74.990 181.005 ;
        RECT 76.390 180.835 76.560 181.005 ;
        RECT 76.825 181.175 76.995 181.345 ;
        RECT 83.735 182.195 83.905 182.365 ;
        RECT 82.815 181.515 82.985 181.685 ;
        RECT 79.135 180.495 79.305 180.665 ;
        RECT 86.035 182.195 86.205 182.365 ;
        RECT 85.575 181.515 85.745 181.685 ;
        RECT 85.115 180.495 85.285 180.665 ;
        RECT 90.405 182.195 90.575 182.365 ;
        RECT 86.955 181.515 87.125 181.685 ;
        RECT 91.555 181.175 91.725 181.345 ;
        RECT 92.015 181.515 92.185 181.685 ;
        RECT 93.395 181.175 93.565 181.345 ;
        RECT 97.995 181.515 98.165 181.685 ;
        RECT 98.915 181.515 99.085 181.685 ;
        RECT 99.375 181.515 99.545 181.685 ;
        RECT 97.075 180.835 97.245 181.005 ;
        RECT 100.755 181.175 100.925 181.345 ;
        RECT 103.975 181.515 104.145 181.685 ;
        RECT 106.505 181.855 106.675 182.025 ;
        RECT 107.655 182.195 107.825 182.365 ;
        RECT 107.195 181.175 107.365 181.345 ;
        RECT 109.955 182.195 110.125 182.365 ;
        RECT 108.575 181.515 108.745 181.685 ;
        RECT 109.495 181.175 109.665 181.345 ;
        RECT 110.875 181.515 111.045 181.685 ;
        RECT 125.135 181.515 125.305 181.685 ;
        RECT 125.620 180.835 125.790 181.005 ;
        RECT 126.015 181.175 126.185 181.345 ;
        RECT 126.470 181.515 126.640 181.685 ;
        RECT 127.205 181.175 127.375 181.345 ;
        RECT 127.720 180.835 127.890 181.005 ;
        RECT 129.290 180.835 129.460 181.005 ;
        RECT 129.725 181.175 129.895 181.345 ;
        RECT 137.095 182.195 137.265 182.365 ;
        RECT 136.635 181.515 136.805 181.685 ;
        RECT 138.015 181.855 138.185 182.025 ;
        RECT 137.555 181.515 137.725 181.685 ;
        RECT 132.035 180.495 132.205 180.665 ;
        RECT 140.315 181.175 140.485 181.345 ;
        RECT 139.395 180.835 139.565 181.005 ;
        RECT 140.775 181.175 140.945 181.345 ;
        RECT 141.260 180.835 141.430 181.005 ;
        RECT 141.655 181.175 141.825 181.345 ;
        RECT 142.000 181.855 142.170 182.025 ;
        RECT 142.845 181.175 143.015 181.345 ;
        RECT 143.360 180.835 143.530 181.005 ;
        RECT 144.930 180.835 145.100 181.005 ;
        RECT 145.365 181.175 145.535 181.345 ;
        RECT 147.675 180.495 147.845 180.665 ;
        RECT 151.355 181.515 151.525 181.685 ;
        RECT 151.815 181.175 151.985 181.345 ;
        RECT 149.515 180.495 149.685 180.665 ;
        RECT 153.655 181.515 153.825 181.685 ;
        RECT 154.115 181.515 154.285 181.685 ;
        RECT 152.735 180.495 152.905 180.665 ;
        RECT 70.855 179.985 71.025 180.155 ;
        RECT 71.315 179.985 71.485 180.155 ;
        RECT 71.775 179.985 71.945 180.155 ;
        RECT 72.235 179.985 72.405 180.155 ;
        RECT 72.695 179.985 72.865 180.155 ;
        RECT 73.155 179.985 73.325 180.155 ;
        RECT 73.615 179.985 73.785 180.155 ;
        RECT 74.075 179.985 74.245 180.155 ;
        RECT 74.535 179.985 74.705 180.155 ;
        RECT 74.995 179.985 75.165 180.155 ;
        RECT 75.455 179.985 75.625 180.155 ;
        RECT 75.915 179.985 76.085 180.155 ;
        RECT 76.375 179.985 76.545 180.155 ;
        RECT 76.835 179.985 77.005 180.155 ;
        RECT 77.295 179.985 77.465 180.155 ;
        RECT 77.755 179.985 77.925 180.155 ;
        RECT 78.215 179.985 78.385 180.155 ;
        RECT 78.675 179.985 78.845 180.155 ;
        RECT 79.135 179.985 79.305 180.155 ;
        RECT 79.595 179.985 79.765 180.155 ;
        RECT 80.055 179.985 80.225 180.155 ;
        RECT 80.515 179.985 80.685 180.155 ;
        RECT 80.975 179.985 81.145 180.155 ;
        RECT 81.435 179.985 81.605 180.155 ;
        RECT 81.895 179.985 82.065 180.155 ;
        RECT 82.355 179.985 82.525 180.155 ;
        RECT 82.815 179.985 82.985 180.155 ;
        RECT 83.275 179.985 83.445 180.155 ;
        RECT 83.735 179.985 83.905 180.155 ;
        RECT 84.195 179.985 84.365 180.155 ;
        RECT 84.655 179.985 84.825 180.155 ;
        RECT 85.115 179.985 85.285 180.155 ;
        RECT 85.575 179.985 85.745 180.155 ;
        RECT 86.035 179.985 86.205 180.155 ;
        RECT 86.495 179.985 86.665 180.155 ;
        RECT 86.955 179.985 87.125 180.155 ;
        RECT 87.415 179.985 87.585 180.155 ;
        RECT 87.875 179.985 88.045 180.155 ;
        RECT 88.335 179.985 88.505 180.155 ;
        RECT 88.795 179.985 88.965 180.155 ;
        RECT 89.255 179.985 89.425 180.155 ;
        RECT 89.715 179.985 89.885 180.155 ;
        RECT 90.175 179.985 90.345 180.155 ;
        RECT 90.635 179.985 90.805 180.155 ;
        RECT 91.095 179.985 91.265 180.155 ;
        RECT 91.555 179.985 91.725 180.155 ;
        RECT 92.015 179.985 92.185 180.155 ;
        RECT 92.475 179.985 92.645 180.155 ;
        RECT 92.935 179.985 93.105 180.155 ;
        RECT 93.395 179.985 93.565 180.155 ;
        RECT 93.855 179.985 94.025 180.155 ;
        RECT 94.315 179.985 94.485 180.155 ;
        RECT 94.775 179.985 94.945 180.155 ;
        RECT 95.235 179.985 95.405 180.155 ;
        RECT 95.695 179.985 95.865 180.155 ;
        RECT 96.155 179.985 96.325 180.155 ;
        RECT 96.615 179.985 96.785 180.155 ;
        RECT 97.075 179.985 97.245 180.155 ;
        RECT 97.535 179.985 97.705 180.155 ;
        RECT 97.995 179.985 98.165 180.155 ;
        RECT 98.455 179.985 98.625 180.155 ;
        RECT 98.915 179.985 99.085 180.155 ;
        RECT 99.375 179.985 99.545 180.155 ;
        RECT 99.835 179.985 100.005 180.155 ;
        RECT 100.295 179.985 100.465 180.155 ;
        RECT 100.755 179.985 100.925 180.155 ;
        RECT 101.215 179.985 101.385 180.155 ;
        RECT 101.675 179.985 101.845 180.155 ;
        RECT 102.135 179.985 102.305 180.155 ;
        RECT 102.595 179.985 102.765 180.155 ;
        RECT 103.055 179.985 103.225 180.155 ;
        RECT 103.515 179.985 103.685 180.155 ;
        RECT 103.975 179.985 104.145 180.155 ;
        RECT 104.435 179.985 104.605 180.155 ;
        RECT 104.895 179.985 105.065 180.155 ;
        RECT 105.355 179.985 105.525 180.155 ;
        RECT 105.815 179.985 105.985 180.155 ;
        RECT 106.275 179.985 106.445 180.155 ;
        RECT 106.735 179.985 106.905 180.155 ;
        RECT 107.195 179.985 107.365 180.155 ;
        RECT 107.655 179.985 107.825 180.155 ;
        RECT 108.115 179.985 108.285 180.155 ;
        RECT 108.575 179.985 108.745 180.155 ;
        RECT 109.035 179.985 109.205 180.155 ;
        RECT 109.495 179.985 109.665 180.155 ;
        RECT 109.955 179.985 110.125 180.155 ;
        RECT 110.415 179.985 110.585 180.155 ;
        RECT 110.875 179.985 111.045 180.155 ;
        RECT 111.335 179.985 111.505 180.155 ;
        RECT 111.795 179.985 111.965 180.155 ;
        RECT 112.255 179.985 112.425 180.155 ;
        RECT 112.715 179.985 112.885 180.155 ;
        RECT 113.175 179.985 113.345 180.155 ;
        RECT 113.635 179.985 113.805 180.155 ;
        RECT 114.095 179.985 114.265 180.155 ;
        RECT 114.555 179.985 114.725 180.155 ;
        RECT 115.015 179.985 115.185 180.155 ;
        RECT 115.475 179.985 115.645 180.155 ;
        RECT 115.935 179.985 116.105 180.155 ;
        RECT 116.395 179.985 116.565 180.155 ;
        RECT 116.855 179.985 117.025 180.155 ;
        RECT 117.315 179.985 117.485 180.155 ;
        RECT 117.775 179.985 117.945 180.155 ;
        RECT 118.235 179.985 118.405 180.155 ;
        RECT 118.695 179.985 118.865 180.155 ;
        RECT 119.155 179.985 119.325 180.155 ;
        RECT 119.615 179.985 119.785 180.155 ;
        RECT 120.075 179.985 120.245 180.155 ;
        RECT 120.535 179.985 120.705 180.155 ;
        RECT 120.995 179.985 121.165 180.155 ;
        RECT 121.455 179.985 121.625 180.155 ;
        RECT 121.915 179.985 122.085 180.155 ;
        RECT 122.375 179.985 122.545 180.155 ;
        RECT 122.835 179.985 123.005 180.155 ;
        RECT 123.295 179.985 123.465 180.155 ;
        RECT 123.755 179.985 123.925 180.155 ;
        RECT 124.215 179.985 124.385 180.155 ;
        RECT 124.675 179.985 124.845 180.155 ;
        RECT 125.135 179.985 125.305 180.155 ;
        RECT 125.595 179.985 125.765 180.155 ;
        RECT 126.055 179.985 126.225 180.155 ;
        RECT 126.515 179.985 126.685 180.155 ;
        RECT 126.975 179.985 127.145 180.155 ;
        RECT 127.435 179.985 127.605 180.155 ;
        RECT 127.895 179.985 128.065 180.155 ;
        RECT 128.355 179.985 128.525 180.155 ;
        RECT 128.815 179.985 128.985 180.155 ;
        RECT 129.275 179.985 129.445 180.155 ;
        RECT 129.735 179.985 129.905 180.155 ;
        RECT 130.195 179.985 130.365 180.155 ;
        RECT 130.655 179.985 130.825 180.155 ;
        RECT 131.115 179.985 131.285 180.155 ;
        RECT 131.575 179.985 131.745 180.155 ;
        RECT 132.035 179.985 132.205 180.155 ;
        RECT 132.495 179.985 132.665 180.155 ;
        RECT 132.955 179.985 133.125 180.155 ;
        RECT 133.415 179.985 133.585 180.155 ;
        RECT 133.875 179.985 134.045 180.155 ;
        RECT 134.335 179.985 134.505 180.155 ;
        RECT 134.795 179.985 134.965 180.155 ;
        RECT 135.255 179.985 135.425 180.155 ;
        RECT 135.715 179.985 135.885 180.155 ;
        RECT 136.175 179.985 136.345 180.155 ;
        RECT 136.635 179.985 136.805 180.155 ;
        RECT 137.095 179.985 137.265 180.155 ;
        RECT 137.555 179.985 137.725 180.155 ;
        RECT 138.015 179.985 138.185 180.155 ;
        RECT 138.475 179.985 138.645 180.155 ;
        RECT 138.935 179.985 139.105 180.155 ;
        RECT 139.395 179.985 139.565 180.155 ;
        RECT 139.855 179.985 140.025 180.155 ;
        RECT 140.315 179.985 140.485 180.155 ;
        RECT 140.775 179.985 140.945 180.155 ;
        RECT 141.235 179.985 141.405 180.155 ;
        RECT 141.695 179.985 141.865 180.155 ;
        RECT 142.155 179.985 142.325 180.155 ;
        RECT 142.615 179.985 142.785 180.155 ;
        RECT 143.075 179.985 143.245 180.155 ;
        RECT 143.535 179.985 143.705 180.155 ;
        RECT 143.995 179.985 144.165 180.155 ;
        RECT 144.455 179.985 144.625 180.155 ;
        RECT 144.915 179.985 145.085 180.155 ;
        RECT 145.375 179.985 145.545 180.155 ;
        RECT 145.835 179.985 146.005 180.155 ;
        RECT 146.295 179.985 146.465 180.155 ;
        RECT 146.755 179.985 146.925 180.155 ;
        RECT 147.215 179.985 147.385 180.155 ;
        RECT 147.675 179.985 147.845 180.155 ;
        RECT 148.135 179.985 148.305 180.155 ;
        RECT 148.595 179.985 148.765 180.155 ;
        RECT 149.055 179.985 149.225 180.155 ;
        RECT 149.515 179.985 149.685 180.155 ;
        RECT 149.975 179.985 150.145 180.155 ;
        RECT 150.435 179.985 150.605 180.155 ;
        RECT 150.895 179.985 151.065 180.155 ;
        RECT 151.355 179.985 151.525 180.155 ;
        RECT 151.815 179.985 151.985 180.155 ;
        RECT 152.275 179.985 152.445 180.155 ;
        RECT 152.735 179.985 152.905 180.155 ;
        RECT 153.195 179.985 153.365 180.155 ;
        RECT 153.655 179.985 153.825 180.155 ;
        RECT 154.115 179.985 154.285 180.155 ;
        RECT 154.575 179.985 154.745 180.155 ;
        RECT 155.035 179.985 155.205 180.155 ;
        RECT 155.495 179.985 155.665 180.155 ;
        RECT 155.955 179.985 156.125 180.155 ;
        RECT 74.995 179.475 75.165 179.645 ;
        RECT 76.835 179.475 77.005 179.645 ;
        RECT 77.755 179.475 77.925 179.645 ;
        RECT 74.995 178.455 75.165 178.625 ;
        RECT 75.915 178.455 76.085 178.625 ;
        RECT 79.135 178.795 79.305 178.965 ;
        RECT 77.675 177.775 77.845 177.945 ;
        RECT 78.675 178.115 78.845 178.285 ;
        RECT 80.055 178.455 80.225 178.625 ;
        RECT 80.515 178.455 80.685 178.625 ;
        RECT 87.875 179.475 88.045 179.645 ;
        RECT 87.415 178.455 87.585 178.625 ;
        RECT 86.495 177.775 86.665 177.945 ;
        RECT 88.795 178.455 88.965 178.625 ;
        RECT 89.255 178.115 89.425 178.285 ;
        RECT 89.715 178.455 89.885 178.625 ;
        RECT 90.635 178.455 90.805 178.625 ;
        RECT 99.835 178.115 100.005 178.285 ;
        RECT 104.895 178.455 105.065 178.625 ;
        RECT 105.815 178.455 105.985 178.625 ;
        RECT 106.275 178.455 106.445 178.625 ;
        RECT 108.115 179.475 108.285 179.645 ;
        RECT 106.735 178.455 106.905 178.625 ;
        RECT 107.195 178.455 107.365 178.625 ;
        RECT 110.875 179.475 111.045 179.645 ;
        RECT 113.175 179.475 113.345 179.645 ;
        RECT 112.715 178.795 112.885 178.965 ;
        RECT 113.635 179.135 113.805 179.305 ;
        RECT 115.015 179.475 115.185 179.645 ;
        RECT 111.795 178.455 111.965 178.625 ;
        RECT 113.175 178.455 113.345 178.625 ;
        RECT 114.555 178.455 114.725 178.625 ;
        RECT 115.015 178.455 115.185 178.625 ;
        RECT 115.935 178.115 116.105 178.285 ;
        RECT 117.315 178.455 117.485 178.625 ;
        RECT 118.235 178.455 118.405 178.625 ;
        RECT 116.395 177.775 116.565 177.945 ;
        RECT 118.695 178.455 118.865 178.625 ;
        RECT 120.995 178.455 121.165 178.625 ;
        RECT 123.755 178.455 123.925 178.625 ;
        RECT 124.215 178.455 124.385 178.625 ;
        RECT 120.535 178.115 120.705 178.285 ;
        RECT 127.435 179.475 127.605 179.645 ;
        RECT 126.055 178.455 126.225 178.625 ;
        RECT 126.515 178.455 126.685 178.625 ;
        RECT 127.895 178.795 128.065 178.965 ;
        RECT 128.815 179.135 128.985 179.305 ;
        RECT 127.435 178.455 127.605 178.625 ;
        RECT 129.275 178.455 129.445 178.625 ;
        RECT 125.135 177.775 125.305 177.945 ;
        RECT 132.955 179.475 133.125 179.645 ;
        RECT 131.575 178.455 131.745 178.625 ;
        RECT 130.655 177.775 130.825 177.945 ;
        RECT 135.715 179.135 135.885 179.305 ;
        RECT 132.035 177.775 132.205 177.945 ;
        RECT 132.875 177.775 133.045 177.945 ;
        RECT 137.555 179.475 137.725 179.645 ;
        RECT 138.475 179.475 138.645 179.645 ;
        RECT 133.875 178.115 134.045 178.285 ;
        RECT 137.555 178.115 137.725 178.285 ;
        RECT 139.855 179.475 140.025 179.645 ;
        RECT 138.935 177.775 139.105 177.945 ;
        RECT 139.750 177.775 139.920 177.945 ;
        RECT 141.235 178.455 141.405 178.625 ;
        RECT 140.775 178.115 140.945 178.285 ;
        RECT 142.155 178.455 142.325 178.625 ;
        RECT 144.940 179.135 145.110 179.305 ;
        RECT 144.455 178.455 144.625 178.625 ;
        RECT 143.075 177.775 143.245 177.945 ;
        RECT 145.335 178.795 145.505 178.965 ;
        RECT 145.790 178.115 145.960 178.285 ;
        RECT 147.040 179.135 147.210 179.305 ;
        RECT 146.525 178.795 146.695 178.965 ;
        RECT 148.610 179.135 148.780 179.305 ;
        RECT 149.045 178.795 149.215 178.965 ;
        RECT 151.355 179.475 151.525 179.645 ;
        RECT 70.855 177.265 71.025 177.435 ;
        RECT 71.315 177.265 71.485 177.435 ;
        RECT 71.775 177.265 71.945 177.435 ;
        RECT 72.235 177.265 72.405 177.435 ;
        RECT 72.695 177.265 72.865 177.435 ;
        RECT 73.155 177.265 73.325 177.435 ;
        RECT 73.615 177.265 73.785 177.435 ;
        RECT 74.075 177.265 74.245 177.435 ;
        RECT 74.535 177.265 74.705 177.435 ;
        RECT 74.995 177.265 75.165 177.435 ;
        RECT 75.455 177.265 75.625 177.435 ;
        RECT 75.915 177.265 76.085 177.435 ;
        RECT 76.375 177.265 76.545 177.435 ;
        RECT 76.835 177.265 77.005 177.435 ;
        RECT 77.295 177.265 77.465 177.435 ;
        RECT 77.755 177.265 77.925 177.435 ;
        RECT 78.215 177.265 78.385 177.435 ;
        RECT 78.675 177.265 78.845 177.435 ;
        RECT 79.135 177.265 79.305 177.435 ;
        RECT 79.595 177.265 79.765 177.435 ;
        RECT 80.055 177.265 80.225 177.435 ;
        RECT 80.515 177.265 80.685 177.435 ;
        RECT 80.975 177.265 81.145 177.435 ;
        RECT 81.435 177.265 81.605 177.435 ;
        RECT 81.895 177.265 82.065 177.435 ;
        RECT 82.355 177.265 82.525 177.435 ;
        RECT 82.815 177.265 82.985 177.435 ;
        RECT 83.275 177.265 83.445 177.435 ;
        RECT 83.735 177.265 83.905 177.435 ;
        RECT 84.195 177.265 84.365 177.435 ;
        RECT 84.655 177.265 84.825 177.435 ;
        RECT 85.115 177.265 85.285 177.435 ;
        RECT 85.575 177.265 85.745 177.435 ;
        RECT 86.035 177.265 86.205 177.435 ;
        RECT 86.495 177.265 86.665 177.435 ;
        RECT 86.955 177.265 87.125 177.435 ;
        RECT 87.415 177.265 87.585 177.435 ;
        RECT 87.875 177.265 88.045 177.435 ;
        RECT 88.335 177.265 88.505 177.435 ;
        RECT 88.795 177.265 88.965 177.435 ;
        RECT 89.255 177.265 89.425 177.435 ;
        RECT 89.715 177.265 89.885 177.435 ;
        RECT 90.175 177.265 90.345 177.435 ;
        RECT 90.635 177.265 90.805 177.435 ;
        RECT 91.095 177.265 91.265 177.435 ;
        RECT 91.555 177.265 91.725 177.435 ;
        RECT 92.015 177.265 92.185 177.435 ;
        RECT 92.475 177.265 92.645 177.435 ;
        RECT 92.935 177.265 93.105 177.435 ;
        RECT 93.395 177.265 93.565 177.435 ;
        RECT 93.855 177.265 94.025 177.435 ;
        RECT 94.315 177.265 94.485 177.435 ;
        RECT 94.775 177.265 94.945 177.435 ;
        RECT 95.235 177.265 95.405 177.435 ;
        RECT 95.695 177.265 95.865 177.435 ;
        RECT 96.155 177.265 96.325 177.435 ;
        RECT 96.615 177.265 96.785 177.435 ;
        RECT 97.075 177.265 97.245 177.435 ;
        RECT 97.535 177.265 97.705 177.435 ;
        RECT 97.995 177.265 98.165 177.435 ;
        RECT 98.455 177.265 98.625 177.435 ;
        RECT 98.915 177.265 99.085 177.435 ;
        RECT 99.375 177.265 99.545 177.435 ;
        RECT 99.835 177.265 100.005 177.435 ;
        RECT 100.295 177.265 100.465 177.435 ;
        RECT 100.755 177.265 100.925 177.435 ;
        RECT 101.215 177.265 101.385 177.435 ;
        RECT 101.675 177.265 101.845 177.435 ;
        RECT 102.135 177.265 102.305 177.435 ;
        RECT 102.595 177.265 102.765 177.435 ;
        RECT 103.055 177.265 103.225 177.435 ;
        RECT 103.515 177.265 103.685 177.435 ;
        RECT 103.975 177.265 104.145 177.435 ;
        RECT 104.435 177.265 104.605 177.435 ;
        RECT 104.895 177.265 105.065 177.435 ;
        RECT 105.355 177.265 105.525 177.435 ;
        RECT 105.815 177.265 105.985 177.435 ;
        RECT 106.275 177.265 106.445 177.435 ;
        RECT 106.735 177.265 106.905 177.435 ;
        RECT 107.195 177.265 107.365 177.435 ;
        RECT 107.655 177.265 107.825 177.435 ;
        RECT 108.115 177.265 108.285 177.435 ;
        RECT 108.575 177.265 108.745 177.435 ;
        RECT 109.035 177.265 109.205 177.435 ;
        RECT 109.495 177.265 109.665 177.435 ;
        RECT 109.955 177.265 110.125 177.435 ;
        RECT 110.415 177.265 110.585 177.435 ;
        RECT 110.875 177.265 111.045 177.435 ;
        RECT 111.335 177.265 111.505 177.435 ;
        RECT 111.795 177.265 111.965 177.435 ;
        RECT 112.255 177.265 112.425 177.435 ;
        RECT 112.715 177.265 112.885 177.435 ;
        RECT 113.175 177.265 113.345 177.435 ;
        RECT 113.635 177.265 113.805 177.435 ;
        RECT 114.095 177.265 114.265 177.435 ;
        RECT 114.555 177.265 114.725 177.435 ;
        RECT 115.015 177.265 115.185 177.435 ;
        RECT 115.475 177.265 115.645 177.435 ;
        RECT 115.935 177.265 116.105 177.435 ;
        RECT 116.395 177.265 116.565 177.435 ;
        RECT 116.855 177.265 117.025 177.435 ;
        RECT 117.315 177.265 117.485 177.435 ;
        RECT 117.775 177.265 117.945 177.435 ;
        RECT 118.235 177.265 118.405 177.435 ;
        RECT 118.695 177.265 118.865 177.435 ;
        RECT 119.155 177.265 119.325 177.435 ;
        RECT 119.615 177.265 119.785 177.435 ;
        RECT 120.075 177.265 120.245 177.435 ;
        RECT 120.535 177.265 120.705 177.435 ;
        RECT 120.995 177.265 121.165 177.435 ;
        RECT 121.455 177.265 121.625 177.435 ;
        RECT 121.915 177.265 122.085 177.435 ;
        RECT 122.375 177.265 122.545 177.435 ;
        RECT 122.835 177.265 123.005 177.435 ;
        RECT 123.295 177.265 123.465 177.435 ;
        RECT 123.755 177.265 123.925 177.435 ;
        RECT 124.215 177.265 124.385 177.435 ;
        RECT 124.675 177.265 124.845 177.435 ;
        RECT 125.135 177.265 125.305 177.435 ;
        RECT 125.595 177.265 125.765 177.435 ;
        RECT 126.055 177.265 126.225 177.435 ;
        RECT 126.515 177.265 126.685 177.435 ;
        RECT 126.975 177.265 127.145 177.435 ;
        RECT 127.435 177.265 127.605 177.435 ;
        RECT 127.895 177.265 128.065 177.435 ;
        RECT 128.355 177.265 128.525 177.435 ;
        RECT 128.815 177.265 128.985 177.435 ;
        RECT 129.275 177.265 129.445 177.435 ;
        RECT 129.735 177.265 129.905 177.435 ;
        RECT 130.195 177.265 130.365 177.435 ;
        RECT 130.655 177.265 130.825 177.435 ;
        RECT 131.115 177.265 131.285 177.435 ;
        RECT 131.575 177.265 131.745 177.435 ;
        RECT 132.035 177.265 132.205 177.435 ;
        RECT 132.495 177.265 132.665 177.435 ;
        RECT 132.955 177.265 133.125 177.435 ;
        RECT 133.415 177.265 133.585 177.435 ;
        RECT 133.875 177.265 134.045 177.435 ;
        RECT 134.335 177.265 134.505 177.435 ;
        RECT 134.795 177.265 134.965 177.435 ;
        RECT 135.255 177.265 135.425 177.435 ;
        RECT 135.715 177.265 135.885 177.435 ;
        RECT 136.175 177.265 136.345 177.435 ;
        RECT 136.635 177.265 136.805 177.435 ;
        RECT 137.095 177.265 137.265 177.435 ;
        RECT 137.555 177.265 137.725 177.435 ;
        RECT 138.015 177.265 138.185 177.435 ;
        RECT 138.475 177.265 138.645 177.435 ;
        RECT 138.935 177.265 139.105 177.435 ;
        RECT 139.395 177.265 139.565 177.435 ;
        RECT 139.855 177.265 140.025 177.435 ;
        RECT 140.315 177.265 140.485 177.435 ;
        RECT 140.775 177.265 140.945 177.435 ;
        RECT 141.235 177.265 141.405 177.435 ;
        RECT 141.695 177.265 141.865 177.435 ;
        RECT 142.155 177.265 142.325 177.435 ;
        RECT 142.615 177.265 142.785 177.435 ;
        RECT 143.075 177.265 143.245 177.435 ;
        RECT 143.535 177.265 143.705 177.435 ;
        RECT 143.995 177.265 144.165 177.435 ;
        RECT 144.455 177.265 144.625 177.435 ;
        RECT 144.915 177.265 145.085 177.435 ;
        RECT 145.375 177.265 145.545 177.435 ;
        RECT 145.835 177.265 146.005 177.435 ;
        RECT 146.295 177.265 146.465 177.435 ;
        RECT 146.755 177.265 146.925 177.435 ;
        RECT 147.215 177.265 147.385 177.435 ;
        RECT 147.675 177.265 147.845 177.435 ;
        RECT 148.135 177.265 148.305 177.435 ;
        RECT 148.595 177.265 148.765 177.435 ;
        RECT 149.055 177.265 149.225 177.435 ;
        RECT 149.515 177.265 149.685 177.435 ;
        RECT 149.975 177.265 150.145 177.435 ;
        RECT 150.435 177.265 150.605 177.435 ;
        RECT 150.895 177.265 151.065 177.435 ;
        RECT 151.355 177.265 151.525 177.435 ;
        RECT 151.815 177.265 151.985 177.435 ;
        RECT 152.275 177.265 152.445 177.435 ;
        RECT 152.735 177.265 152.905 177.435 ;
        RECT 153.195 177.265 153.365 177.435 ;
        RECT 153.655 177.265 153.825 177.435 ;
        RECT 154.115 177.265 154.285 177.435 ;
        RECT 154.575 177.265 154.745 177.435 ;
        RECT 155.035 177.265 155.205 177.435 ;
        RECT 155.495 177.265 155.665 177.435 ;
        RECT 155.955 177.265 156.125 177.435 ;
        RECT 76.375 176.755 76.545 176.925 ;
        RECT 77.295 176.075 77.465 176.245 ;
        RECT 78.215 176.075 78.385 176.245 ;
        RECT 80.975 176.075 81.145 176.245 ;
        RECT 79.135 175.395 79.305 175.565 ;
        RECT 80.055 175.735 80.225 175.905 ;
        RECT 79.595 175.055 79.765 175.225 ;
        RECT 81.460 175.395 81.630 175.565 ;
        RECT 81.855 175.735 82.025 175.905 ;
        RECT 82.310 176.415 82.480 176.585 ;
        RECT 83.045 175.735 83.215 175.905 ;
        RECT 83.560 175.395 83.730 175.565 ;
        RECT 85.130 175.395 85.300 175.565 ;
        RECT 85.565 175.735 85.735 175.905 ;
        RECT 87.875 175.395 88.045 175.565 ;
        RECT 89.255 176.755 89.425 176.925 ;
        RECT 89.715 176.075 89.885 176.245 ;
        RECT 91.095 176.755 91.265 176.925 ;
        RECT 90.175 176.075 90.345 176.245 ;
        RECT 88.335 175.395 88.505 175.565 ;
        RECT 91.555 175.055 91.725 175.225 ;
        RECT 92.935 176.075 93.105 176.245 ;
        RECT 93.855 176.075 94.025 176.245 ;
        RECT 94.315 176.075 94.485 176.245 ;
        RECT 92.935 175.055 93.105 175.225 ;
        RECT 97.075 176.075 97.245 176.245 ;
        RECT 95.235 175.055 95.405 175.225 ;
        RECT 101.675 176.075 101.845 176.245 ;
        RECT 106.735 176.755 106.905 176.925 ;
        RECT 108.115 176.755 108.285 176.925 ;
        RECT 111.335 176.755 111.505 176.925 ;
        RECT 103.055 176.075 103.225 176.245 ;
        RECT 97.995 175.055 98.165 175.225 ;
        RECT 102.135 175.395 102.305 175.565 ;
        RECT 103.975 175.395 104.145 175.565 ;
        RECT 104.435 175.395 104.605 175.565 ;
        RECT 104.895 176.075 105.065 176.245 ;
        RECT 105.355 176.075 105.525 176.245 ;
        RECT 107.195 176.075 107.365 176.245 ;
        RECT 108.115 176.075 108.285 176.245 ;
        RECT 114.095 176.755 114.265 176.925 ;
        RECT 112.255 176.075 112.425 176.245 ;
        RECT 113.635 176.075 113.805 176.245 ;
        RECT 113.175 175.735 113.345 175.905 ;
        RECT 115.935 176.075 116.105 176.245 ;
        RECT 112.255 175.055 112.425 175.225 ;
        RECT 115.475 175.735 115.645 175.905 ;
        RECT 115.935 175.055 116.105 175.225 ;
        RECT 120.995 176.075 121.165 176.245 ;
        RECT 121.915 176.075 122.085 176.245 ;
        RECT 120.075 175.735 120.245 175.905 ;
        RECT 126.055 176.075 126.225 176.245 ;
        RECT 125.135 175.735 125.305 175.905 ;
        RECT 130.195 176.415 130.365 176.585 ;
        RECT 146.295 176.755 146.465 176.925 ;
        RECT 138.935 176.075 139.105 176.245 ;
        RECT 129.275 175.735 129.445 175.905 ;
        RECT 126.535 175.055 126.705 175.225 ;
        RECT 127.455 175.055 127.625 175.225 ;
        RECT 148.595 176.755 148.765 176.925 ;
        RECT 145.835 176.075 146.005 176.245 ;
        RECT 146.295 175.735 146.465 175.905 ;
        RECT 147.675 176.075 147.845 176.245 ;
        RECT 144.685 175.055 144.855 175.225 ;
        RECT 147.215 175.055 147.385 175.225 ;
        RECT 149.515 176.075 149.685 176.245 ;
        RECT 150.435 176.075 150.605 176.245 ;
        RECT 150.895 176.075 151.065 176.245 ;
        RECT 151.815 176.075 151.985 176.245 ;
        RECT 152.735 175.395 152.905 175.565 ;
        RECT 70.855 174.545 71.025 174.715 ;
        RECT 71.315 174.545 71.485 174.715 ;
        RECT 71.775 174.545 71.945 174.715 ;
        RECT 72.235 174.545 72.405 174.715 ;
        RECT 72.695 174.545 72.865 174.715 ;
        RECT 73.155 174.545 73.325 174.715 ;
        RECT 73.615 174.545 73.785 174.715 ;
        RECT 74.075 174.545 74.245 174.715 ;
        RECT 74.535 174.545 74.705 174.715 ;
        RECT 74.995 174.545 75.165 174.715 ;
        RECT 75.455 174.545 75.625 174.715 ;
        RECT 75.915 174.545 76.085 174.715 ;
        RECT 76.375 174.545 76.545 174.715 ;
        RECT 76.835 174.545 77.005 174.715 ;
        RECT 77.295 174.545 77.465 174.715 ;
        RECT 77.755 174.545 77.925 174.715 ;
        RECT 78.215 174.545 78.385 174.715 ;
        RECT 78.675 174.545 78.845 174.715 ;
        RECT 79.135 174.545 79.305 174.715 ;
        RECT 79.595 174.545 79.765 174.715 ;
        RECT 80.055 174.545 80.225 174.715 ;
        RECT 80.515 174.545 80.685 174.715 ;
        RECT 80.975 174.545 81.145 174.715 ;
        RECT 81.435 174.545 81.605 174.715 ;
        RECT 81.895 174.545 82.065 174.715 ;
        RECT 82.355 174.545 82.525 174.715 ;
        RECT 82.815 174.545 82.985 174.715 ;
        RECT 83.275 174.545 83.445 174.715 ;
        RECT 83.735 174.545 83.905 174.715 ;
        RECT 84.195 174.545 84.365 174.715 ;
        RECT 84.655 174.545 84.825 174.715 ;
        RECT 85.115 174.545 85.285 174.715 ;
        RECT 85.575 174.545 85.745 174.715 ;
        RECT 86.035 174.545 86.205 174.715 ;
        RECT 86.495 174.545 86.665 174.715 ;
        RECT 86.955 174.545 87.125 174.715 ;
        RECT 87.415 174.545 87.585 174.715 ;
        RECT 87.875 174.545 88.045 174.715 ;
        RECT 88.335 174.545 88.505 174.715 ;
        RECT 88.795 174.545 88.965 174.715 ;
        RECT 89.255 174.545 89.425 174.715 ;
        RECT 89.715 174.545 89.885 174.715 ;
        RECT 90.175 174.545 90.345 174.715 ;
        RECT 90.635 174.545 90.805 174.715 ;
        RECT 91.095 174.545 91.265 174.715 ;
        RECT 91.555 174.545 91.725 174.715 ;
        RECT 92.015 174.545 92.185 174.715 ;
        RECT 92.475 174.545 92.645 174.715 ;
        RECT 92.935 174.545 93.105 174.715 ;
        RECT 93.395 174.545 93.565 174.715 ;
        RECT 93.855 174.545 94.025 174.715 ;
        RECT 94.315 174.545 94.485 174.715 ;
        RECT 94.775 174.545 94.945 174.715 ;
        RECT 95.235 174.545 95.405 174.715 ;
        RECT 95.695 174.545 95.865 174.715 ;
        RECT 96.155 174.545 96.325 174.715 ;
        RECT 96.615 174.545 96.785 174.715 ;
        RECT 97.075 174.545 97.245 174.715 ;
        RECT 97.535 174.545 97.705 174.715 ;
        RECT 97.995 174.545 98.165 174.715 ;
        RECT 98.455 174.545 98.625 174.715 ;
        RECT 98.915 174.545 99.085 174.715 ;
        RECT 99.375 174.545 99.545 174.715 ;
        RECT 99.835 174.545 100.005 174.715 ;
        RECT 100.295 174.545 100.465 174.715 ;
        RECT 100.755 174.545 100.925 174.715 ;
        RECT 101.215 174.545 101.385 174.715 ;
        RECT 101.675 174.545 101.845 174.715 ;
        RECT 102.135 174.545 102.305 174.715 ;
        RECT 102.595 174.545 102.765 174.715 ;
        RECT 103.055 174.545 103.225 174.715 ;
        RECT 103.515 174.545 103.685 174.715 ;
        RECT 103.975 174.545 104.145 174.715 ;
        RECT 104.435 174.545 104.605 174.715 ;
        RECT 104.895 174.545 105.065 174.715 ;
        RECT 105.355 174.545 105.525 174.715 ;
        RECT 105.815 174.545 105.985 174.715 ;
        RECT 106.275 174.545 106.445 174.715 ;
        RECT 106.735 174.545 106.905 174.715 ;
        RECT 107.195 174.545 107.365 174.715 ;
        RECT 107.655 174.545 107.825 174.715 ;
        RECT 108.115 174.545 108.285 174.715 ;
        RECT 108.575 174.545 108.745 174.715 ;
        RECT 109.035 174.545 109.205 174.715 ;
        RECT 109.495 174.545 109.665 174.715 ;
        RECT 109.955 174.545 110.125 174.715 ;
        RECT 110.415 174.545 110.585 174.715 ;
        RECT 110.875 174.545 111.045 174.715 ;
        RECT 111.335 174.545 111.505 174.715 ;
        RECT 111.795 174.545 111.965 174.715 ;
        RECT 112.255 174.545 112.425 174.715 ;
        RECT 112.715 174.545 112.885 174.715 ;
        RECT 113.175 174.545 113.345 174.715 ;
        RECT 113.635 174.545 113.805 174.715 ;
        RECT 114.095 174.545 114.265 174.715 ;
        RECT 114.555 174.545 114.725 174.715 ;
        RECT 115.015 174.545 115.185 174.715 ;
        RECT 115.475 174.545 115.645 174.715 ;
        RECT 115.935 174.545 116.105 174.715 ;
        RECT 116.395 174.545 116.565 174.715 ;
        RECT 116.855 174.545 117.025 174.715 ;
        RECT 117.315 174.545 117.485 174.715 ;
        RECT 117.775 174.545 117.945 174.715 ;
        RECT 118.235 174.545 118.405 174.715 ;
        RECT 118.695 174.545 118.865 174.715 ;
        RECT 119.155 174.545 119.325 174.715 ;
        RECT 119.615 174.545 119.785 174.715 ;
        RECT 120.075 174.545 120.245 174.715 ;
        RECT 120.535 174.545 120.705 174.715 ;
        RECT 120.995 174.545 121.165 174.715 ;
        RECT 121.455 174.545 121.625 174.715 ;
        RECT 121.915 174.545 122.085 174.715 ;
        RECT 122.375 174.545 122.545 174.715 ;
        RECT 122.835 174.545 123.005 174.715 ;
        RECT 123.295 174.545 123.465 174.715 ;
        RECT 123.755 174.545 123.925 174.715 ;
        RECT 124.215 174.545 124.385 174.715 ;
        RECT 124.675 174.545 124.845 174.715 ;
        RECT 125.135 174.545 125.305 174.715 ;
        RECT 125.595 174.545 125.765 174.715 ;
        RECT 126.055 174.545 126.225 174.715 ;
        RECT 126.515 174.545 126.685 174.715 ;
        RECT 126.975 174.545 127.145 174.715 ;
        RECT 127.435 174.545 127.605 174.715 ;
        RECT 127.895 174.545 128.065 174.715 ;
        RECT 128.355 174.545 128.525 174.715 ;
        RECT 128.815 174.545 128.985 174.715 ;
        RECT 129.275 174.545 129.445 174.715 ;
        RECT 129.735 174.545 129.905 174.715 ;
        RECT 130.195 174.545 130.365 174.715 ;
        RECT 130.655 174.545 130.825 174.715 ;
        RECT 131.115 174.545 131.285 174.715 ;
        RECT 131.575 174.545 131.745 174.715 ;
        RECT 132.035 174.545 132.205 174.715 ;
        RECT 132.495 174.545 132.665 174.715 ;
        RECT 132.955 174.545 133.125 174.715 ;
        RECT 133.415 174.545 133.585 174.715 ;
        RECT 133.875 174.545 134.045 174.715 ;
        RECT 134.335 174.545 134.505 174.715 ;
        RECT 134.795 174.545 134.965 174.715 ;
        RECT 135.255 174.545 135.425 174.715 ;
        RECT 135.715 174.545 135.885 174.715 ;
        RECT 136.175 174.545 136.345 174.715 ;
        RECT 136.635 174.545 136.805 174.715 ;
        RECT 137.095 174.545 137.265 174.715 ;
        RECT 137.555 174.545 137.725 174.715 ;
        RECT 138.015 174.545 138.185 174.715 ;
        RECT 138.475 174.545 138.645 174.715 ;
        RECT 138.935 174.545 139.105 174.715 ;
        RECT 139.395 174.545 139.565 174.715 ;
        RECT 139.855 174.545 140.025 174.715 ;
        RECT 140.315 174.545 140.485 174.715 ;
        RECT 140.775 174.545 140.945 174.715 ;
        RECT 141.235 174.545 141.405 174.715 ;
        RECT 141.695 174.545 141.865 174.715 ;
        RECT 142.155 174.545 142.325 174.715 ;
        RECT 142.615 174.545 142.785 174.715 ;
        RECT 143.075 174.545 143.245 174.715 ;
        RECT 143.535 174.545 143.705 174.715 ;
        RECT 143.995 174.545 144.165 174.715 ;
        RECT 144.455 174.545 144.625 174.715 ;
        RECT 144.915 174.545 145.085 174.715 ;
        RECT 145.375 174.545 145.545 174.715 ;
        RECT 145.835 174.545 146.005 174.715 ;
        RECT 146.295 174.545 146.465 174.715 ;
        RECT 146.755 174.545 146.925 174.715 ;
        RECT 147.215 174.545 147.385 174.715 ;
        RECT 147.675 174.545 147.845 174.715 ;
        RECT 148.135 174.545 148.305 174.715 ;
        RECT 148.595 174.545 148.765 174.715 ;
        RECT 149.055 174.545 149.225 174.715 ;
        RECT 149.515 174.545 149.685 174.715 ;
        RECT 149.975 174.545 150.145 174.715 ;
        RECT 150.435 174.545 150.605 174.715 ;
        RECT 150.895 174.545 151.065 174.715 ;
        RECT 151.355 174.545 151.525 174.715 ;
        RECT 151.815 174.545 151.985 174.715 ;
        RECT 152.275 174.545 152.445 174.715 ;
        RECT 152.735 174.545 152.905 174.715 ;
        RECT 153.195 174.545 153.365 174.715 ;
        RECT 153.655 174.545 153.825 174.715 ;
        RECT 154.115 174.545 154.285 174.715 ;
        RECT 154.575 174.545 154.745 174.715 ;
        RECT 155.035 174.545 155.205 174.715 ;
        RECT 155.495 174.545 155.665 174.715 ;
        RECT 155.955 174.545 156.125 174.715 ;
        RECT 75.455 173.015 75.625 173.185 ;
        RECT 76.375 173.015 76.545 173.185 ;
        RECT 75.915 172.335 76.085 172.505 ;
        RECT 88.335 173.355 88.505 173.525 ;
        RECT 90.635 174.035 90.805 174.205 ;
        RECT 89.715 173.015 89.885 173.185 ;
        RECT 93.395 174.035 93.565 174.205 ;
        RECT 92.475 173.355 92.645 173.525 ;
        RECT 91.555 173.015 91.725 173.185 ;
        RECT 95.235 173.695 95.405 173.865 ;
        RECT 93.855 172.675 94.025 172.845 ;
        RECT 97.995 173.355 98.165 173.525 ;
        RECT 96.155 173.015 96.325 173.185 ;
        RECT 96.615 172.335 96.785 172.505 ;
        RECT 97.075 172.675 97.245 172.845 ;
        RECT 103.055 174.035 103.225 174.205 ;
        RECT 101.675 173.355 101.845 173.525 ;
        RECT 98.455 173.015 98.625 173.185 ;
        RECT 99.375 173.015 99.545 173.185 ;
        RECT 100.985 172.675 101.155 172.845 ;
        RECT 107.195 174.035 107.365 174.205 ;
        RECT 103.975 173.015 104.145 173.185 ;
        RECT 104.435 172.675 104.605 172.845 ;
        RECT 105.815 173.015 105.985 173.185 ;
        RECT 106.275 173.015 106.445 173.185 ;
        RECT 104.895 172.675 105.065 172.845 ;
        RECT 111.335 172.675 111.505 172.845 ;
        RECT 119.155 173.015 119.325 173.185 ;
        RECT 132.955 173.355 133.125 173.525 ;
        RECT 132.035 173.015 132.205 173.185 ;
        RECT 133.415 173.015 133.585 173.185 ;
        RECT 135.715 174.035 135.885 174.205 ;
        RECT 134.335 173.015 134.505 173.185 ;
        RECT 131.115 172.335 131.285 172.505 ;
        RECT 133.875 172.675 134.045 172.845 ;
        RECT 136.635 173.015 136.805 173.185 ;
        RECT 137.555 173.015 137.725 173.185 ;
        RECT 139.855 173.695 140.025 173.865 ;
        RECT 141.695 174.035 141.865 174.205 ;
        RECT 142.615 174.035 142.785 174.205 ;
        RECT 141.695 172.675 141.865 172.845 ;
        RECT 144.915 173.015 145.085 173.185 ;
        RECT 143.995 172.675 144.165 172.845 ;
        RECT 146.295 173.015 146.465 173.185 ;
        RECT 145.375 172.335 145.545 172.505 ;
        RECT 149.975 173.355 150.145 173.525 ;
        RECT 150.435 173.015 150.605 173.185 ;
        RECT 152.275 172.335 152.445 172.505 ;
        RECT 70.855 171.825 71.025 171.995 ;
        RECT 71.315 171.825 71.485 171.995 ;
        RECT 71.775 171.825 71.945 171.995 ;
        RECT 72.235 171.825 72.405 171.995 ;
        RECT 72.695 171.825 72.865 171.995 ;
        RECT 73.155 171.825 73.325 171.995 ;
        RECT 73.615 171.825 73.785 171.995 ;
        RECT 74.075 171.825 74.245 171.995 ;
        RECT 74.535 171.825 74.705 171.995 ;
        RECT 74.995 171.825 75.165 171.995 ;
        RECT 75.455 171.825 75.625 171.995 ;
        RECT 75.915 171.825 76.085 171.995 ;
        RECT 76.375 171.825 76.545 171.995 ;
        RECT 76.835 171.825 77.005 171.995 ;
        RECT 77.295 171.825 77.465 171.995 ;
        RECT 77.755 171.825 77.925 171.995 ;
        RECT 78.215 171.825 78.385 171.995 ;
        RECT 78.675 171.825 78.845 171.995 ;
        RECT 79.135 171.825 79.305 171.995 ;
        RECT 79.595 171.825 79.765 171.995 ;
        RECT 80.055 171.825 80.225 171.995 ;
        RECT 80.515 171.825 80.685 171.995 ;
        RECT 80.975 171.825 81.145 171.995 ;
        RECT 81.435 171.825 81.605 171.995 ;
        RECT 81.895 171.825 82.065 171.995 ;
        RECT 82.355 171.825 82.525 171.995 ;
        RECT 82.815 171.825 82.985 171.995 ;
        RECT 83.275 171.825 83.445 171.995 ;
        RECT 83.735 171.825 83.905 171.995 ;
        RECT 84.195 171.825 84.365 171.995 ;
        RECT 84.655 171.825 84.825 171.995 ;
        RECT 85.115 171.825 85.285 171.995 ;
        RECT 85.575 171.825 85.745 171.995 ;
        RECT 86.035 171.825 86.205 171.995 ;
        RECT 86.495 171.825 86.665 171.995 ;
        RECT 86.955 171.825 87.125 171.995 ;
        RECT 87.415 171.825 87.585 171.995 ;
        RECT 87.875 171.825 88.045 171.995 ;
        RECT 88.335 171.825 88.505 171.995 ;
        RECT 88.795 171.825 88.965 171.995 ;
        RECT 89.255 171.825 89.425 171.995 ;
        RECT 89.715 171.825 89.885 171.995 ;
        RECT 90.175 171.825 90.345 171.995 ;
        RECT 90.635 171.825 90.805 171.995 ;
        RECT 91.095 171.825 91.265 171.995 ;
        RECT 91.555 171.825 91.725 171.995 ;
        RECT 92.015 171.825 92.185 171.995 ;
        RECT 92.475 171.825 92.645 171.995 ;
        RECT 92.935 171.825 93.105 171.995 ;
        RECT 93.395 171.825 93.565 171.995 ;
        RECT 93.855 171.825 94.025 171.995 ;
        RECT 94.315 171.825 94.485 171.995 ;
        RECT 94.775 171.825 94.945 171.995 ;
        RECT 95.235 171.825 95.405 171.995 ;
        RECT 95.695 171.825 95.865 171.995 ;
        RECT 96.155 171.825 96.325 171.995 ;
        RECT 96.615 171.825 96.785 171.995 ;
        RECT 97.075 171.825 97.245 171.995 ;
        RECT 97.535 171.825 97.705 171.995 ;
        RECT 97.995 171.825 98.165 171.995 ;
        RECT 98.455 171.825 98.625 171.995 ;
        RECT 98.915 171.825 99.085 171.995 ;
        RECT 99.375 171.825 99.545 171.995 ;
        RECT 99.835 171.825 100.005 171.995 ;
        RECT 100.295 171.825 100.465 171.995 ;
        RECT 100.755 171.825 100.925 171.995 ;
        RECT 101.215 171.825 101.385 171.995 ;
        RECT 101.675 171.825 101.845 171.995 ;
        RECT 102.135 171.825 102.305 171.995 ;
        RECT 102.595 171.825 102.765 171.995 ;
        RECT 103.055 171.825 103.225 171.995 ;
        RECT 103.515 171.825 103.685 171.995 ;
        RECT 103.975 171.825 104.145 171.995 ;
        RECT 104.435 171.825 104.605 171.995 ;
        RECT 104.895 171.825 105.065 171.995 ;
        RECT 105.355 171.825 105.525 171.995 ;
        RECT 105.815 171.825 105.985 171.995 ;
        RECT 106.275 171.825 106.445 171.995 ;
        RECT 106.735 171.825 106.905 171.995 ;
        RECT 107.195 171.825 107.365 171.995 ;
        RECT 107.655 171.825 107.825 171.995 ;
        RECT 108.115 171.825 108.285 171.995 ;
        RECT 108.575 171.825 108.745 171.995 ;
        RECT 109.035 171.825 109.205 171.995 ;
        RECT 109.495 171.825 109.665 171.995 ;
        RECT 109.955 171.825 110.125 171.995 ;
        RECT 110.415 171.825 110.585 171.995 ;
        RECT 110.875 171.825 111.045 171.995 ;
        RECT 111.335 171.825 111.505 171.995 ;
        RECT 111.795 171.825 111.965 171.995 ;
        RECT 112.255 171.825 112.425 171.995 ;
        RECT 112.715 171.825 112.885 171.995 ;
        RECT 113.175 171.825 113.345 171.995 ;
        RECT 113.635 171.825 113.805 171.995 ;
        RECT 114.095 171.825 114.265 171.995 ;
        RECT 114.555 171.825 114.725 171.995 ;
        RECT 115.015 171.825 115.185 171.995 ;
        RECT 115.475 171.825 115.645 171.995 ;
        RECT 115.935 171.825 116.105 171.995 ;
        RECT 116.395 171.825 116.565 171.995 ;
        RECT 116.855 171.825 117.025 171.995 ;
        RECT 117.315 171.825 117.485 171.995 ;
        RECT 117.775 171.825 117.945 171.995 ;
        RECT 118.235 171.825 118.405 171.995 ;
        RECT 118.695 171.825 118.865 171.995 ;
        RECT 119.155 171.825 119.325 171.995 ;
        RECT 119.615 171.825 119.785 171.995 ;
        RECT 120.075 171.825 120.245 171.995 ;
        RECT 120.535 171.825 120.705 171.995 ;
        RECT 120.995 171.825 121.165 171.995 ;
        RECT 121.455 171.825 121.625 171.995 ;
        RECT 121.915 171.825 122.085 171.995 ;
        RECT 122.375 171.825 122.545 171.995 ;
        RECT 122.835 171.825 123.005 171.995 ;
        RECT 123.295 171.825 123.465 171.995 ;
        RECT 123.755 171.825 123.925 171.995 ;
        RECT 124.215 171.825 124.385 171.995 ;
        RECT 124.675 171.825 124.845 171.995 ;
        RECT 125.135 171.825 125.305 171.995 ;
        RECT 125.595 171.825 125.765 171.995 ;
        RECT 126.055 171.825 126.225 171.995 ;
        RECT 126.515 171.825 126.685 171.995 ;
        RECT 126.975 171.825 127.145 171.995 ;
        RECT 127.435 171.825 127.605 171.995 ;
        RECT 127.895 171.825 128.065 171.995 ;
        RECT 128.355 171.825 128.525 171.995 ;
        RECT 128.815 171.825 128.985 171.995 ;
        RECT 129.275 171.825 129.445 171.995 ;
        RECT 129.735 171.825 129.905 171.995 ;
        RECT 130.195 171.825 130.365 171.995 ;
        RECT 130.655 171.825 130.825 171.995 ;
        RECT 131.115 171.825 131.285 171.995 ;
        RECT 131.575 171.825 131.745 171.995 ;
        RECT 132.035 171.825 132.205 171.995 ;
        RECT 132.495 171.825 132.665 171.995 ;
        RECT 132.955 171.825 133.125 171.995 ;
        RECT 133.415 171.825 133.585 171.995 ;
        RECT 133.875 171.825 134.045 171.995 ;
        RECT 134.335 171.825 134.505 171.995 ;
        RECT 134.795 171.825 134.965 171.995 ;
        RECT 135.255 171.825 135.425 171.995 ;
        RECT 135.715 171.825 135.885 171.995 ;
        RECT 136.175 171.825 136.345 171.995 ;
        RECT 136.635 171.825 136.805 171.995 ;
        RECT 137.095 171.825 137.265 171.995 ;
        RECT 137.555 171.825 137.725 171.995 ;
        RECT 138.015 171.825 138.185 171.995 ;
        RECT 138.475 171.825 138.645 171.995 ;
        RECT 138.935 171.825 139.105 171.995 ;
        RECT 139.395 171.825 139.565 171.995 ;
        RECT 139.855 171.825 140.025 171.995 ;
        RECT 140.315 171.825 140.485 171.995 ;
        RECT 140.775 171.825 140.945 171.995 ;
        RECT 141.235 171.825 141.405 171.995 ;
        RECT 141.695 171.825 141.865 171.995 ;
        RECT 142.155 171.825 142.325 171.995 ;
        RECT 142.615 171.825 142.785 171.995 ;
        RECT 143.075 171.825 143.245 171.995 ;
        RECT 143.535 171.825 143.705 171.995 ;
        RECT 143.995 171.825 144.165 171.995 ;
        RECT 144.455 171.825 144.625 171.995 ;
        RECT 144.915 171.825 145.085 171.995 ;
        RECT 145.375 171.825 145.545 171.995 ;
        RECT 145.835 171.825 146.005 171.995 ;
        RECT 146.295 171.825 146.465 171.995 ;
        RECT 146.755 171.825 146.925 171.995 ;
        RECT 147.215 171.825 147.385 171.995 ;
        RECT 147.675 171.825 147.845 171.995 ;
        RECT 148.135 171.825 148.305 171.995 ;
        RECT 148.595 171.825 148.765 171.995 ;
        RECT 149.055 171.825 149.225 171.995 ;
        RECT 149.515 171.825 149.685 171.995 ;
        RECT 149.975 171.825 150.145 171.995 ;
        RECT 150.435 171.825 150.605 171.995 ;
        RECT 150.895 171.825 151.065 171.995 ;
        RECT 151.355 171.825 151.525 171.995 ;
        RECT 151.815 171.825 151.985 171.995 ;
        RECT 152.275 171.825 152.445 171.995 ;
        RECT 152.735 171.825 152.905 171.995 ;
        RECT 153.195 171.825 153.365 171.995 ;
        RECT 153.655 171.825 153.825 171.995 ;
        RECT 154.115 171.825 154.285 171.995 ;
        RECT 154.575 171.825 154.745 171.995 ;
        RECT 155.035 171.825 155.205 171.995 ;
        RECT 155.495 171.825 155.665 171.995 ;
        RECT 155.955 171.825 156.125 171.995 ;
        RECT 72.235 170.295 72.405 170.465 ;
        RECT 72.720 169.955 72.890 170.125 ;
        RECT 73.115 170.295 73.285 170.465 ;
        RECT 73.570 170.635 73.740 170.805 ;
        RECT 74.305 170.295 74.475 170.465 ;
        RECT 74.820 169.955 74.990 170.125 ;
        RECT 76.390 169.955 76.560 170.125 ;
        RECT 76.825 170.295 76.995 170.465 ;
        RECT 79.595 170.635 79.765 170.805 ;
        RECT 79.135 169.615 79.305 169.785 ;
        RECT 80.080 169.955 80.250 170.125 ;
        RECT 80.475 170.295 80.645 170.465 ;
        RECT 80.930 170.975 81.100 171.145 ;
        RECT 81.665 170.295 81.835 170.465 ;
        RECT 82.180 169.955 82.350 170.125 ;
        RECT 83.750 169.955 83.920 170.125 ;
        RECT 84.185 170.295 84.355 170.465 ;
        RECT 86.955 171.315 87.125 171.485 ;
        RECT 86.495 169.955 86.665 170.125 ;
        RECT 88.795 171.315 88.965 171.485 ;
        RECT 89.715 171.315 89.885 171.485 ;
        RECT 87.875 170.635 88.045 170.805 ;
        RECT 92.475 171.315 92.645 171.485 ;
        RECT 90.635 170.635 90.805 170.805 ;
        RECT 90.175 170.295 90.345 170.465 ;
        RECT 91.095 170.295 91.265 170.465 ;
        RECT 90.635 169.615 90.805 169.785 ;
        RECT 93.395 170.635 93.565 170.805 ;
        RECT 94.315 170.635 94.485 170.805 ;
        RECT 94.775 170.635 94.945 170.805 ;
        RECT 95.235 171.315 95.405 171.485 ;
        RECT 97.075 170.975 97.245 171.145 ;
        RECT 96.155 170.295 96.325 170.465 ;
        RECT 98.075 171.315 98.245 171.485 ;
        RECT 98.915 169.955 99.085 170.125 ;
        RECT 100.295 170.635 100.465 170.805 ;
        RECT 100.755 170.295 100.925 170.465 ;
        RECT 102.595 171.315 102.765 171.485 ;
        RECT 103.515 170.975 103.685 171.145 ;
        RECT 107.655 171.315 107.825 171.485 ;
        RECT 104.435 170.635 104.605 170.805 ;
        RECT 104.895 170.635 105.065 170.805 ;
        RECT 105.815 170.635 105.985 170.805 ;
        RECT 97.995 169.615 98.165 169.785 ;
        RECT 101.675 169.615 101.845 169.785 ;
        RECT 105.355 170.295 105.525 170.465 ;
        RECT 108.575 170.295 108.745 170.465 ;
        RECT 110.415 170.295 110.585 170.465 ;
        RECT 110.875 170.295 111.045 170.465 ;
        RECT 114.555 171.315 114.725 171.485 ;
        RECT 112.715 170.635 112.885 170.805 ;
        RECT 114.095 170.635 114.265 170.805 ;
        RECT 113.635 170.295 113.805 170.465 ;
        RECT 111.795 169.615 111.965 169.785 ;
        RECT 115.475 170.635 115.645 170.805 ;
        RECT 116.395 170.635 116.565 170.805 ;
        RECT 116.855 170.635 117.025 170.805 ;
        RECT 118.235 170.635 118.405 170.805 ;
        RECT 119.155 171.315 119.325 171.485 ;
        RECT 112.715 169.615 112.885 169.785 ;
        RECT 120.995 170.975 121.165 171.145 ;
        RECT 119.615 170.635 119.785 170.805 ;
        RECT 120.535 170.635 120.705 170.805 ;
        RECT 121.455 170.635 121.625 170.805 ;
        RECT 122.835 170.635 123.005 170.805 ;
        RECT 118.235 169.615 118.405 169.785 ;
        RECT 123.320 169.955 123.490 170.125 ;
        RECT 123.715 170.295 123.885 170.465 ;
        RECT 124.060 170.975 124.230 171.145 ;
        RECT 124.905 170.295 125.075 170.465 ;
        RECT 125.420 169.955 125.590 170.125 ;
        RECT 126.990 169.955 127.160 170.125 ;
        RECT 127.425 170.295 127.595 170.465 ;
        RECT 129.735 171.315 129.905 171.485 ;
        RECT 131.575 171.315 131.745 171.485 ;
        RECT 131.115 170.635 131.285 170.805 ;
        RECT 130.195 169.615 130.365 169.785 ;
        RECT 136.175 171.315 136.345 171.485 ;
        RECT 132.495 170.635 132.665 170.805 ;
        RECT 135.255 170.635 135.425 170.805 ;
        RECT 139.855 171.315 140.025 171.485 ;
        RECT 138.935 170.635 139.105 170.805 ;
        RECT 138.015 170.295 138.185 170.465 ;
        RECT 144.915 170.635 145.085 170.805 ;
        RECT 144.455 169.955 144.625 170.125 ;
        RECT 146.295 170.635 146.465 170.805 ;
        RECT 147.215 170.635 147.385 170.805 ;
        RECT 147.675 170.635 147.845 170.805 ;
        RECT 145.375 169.615 145.545 169.785 ;
        RECT 151.355 171.315 151.525 171.485 ;
        RECT 149.515 170.635 149.685 170.805 ;
        RECT 149.055 170.295 149.225 170.465 ;
        RECT 152.275 170.975 152.445 171.145 ;
        RECT 151.815 170.635 151.985 170.805 ;
        RECT 152.735 170.635 152.905 170.805 ;
        RECT 153.195 170.635 153.365 170.805 ;
        RECT 153.655 169.615 153.825 169.785 ;
        RECT 70.855 169.105 71.025 169.275 ;
        RECT 71.315 169.105 71.485 169.275 ;
        RECT 71.775 169.105 71.945 169.275 ;
        RECT 72.235 169.105 72.405 169.275 ;
        RECT 72.695 169.105 72.865 169.275 ;
        RECT 73.155 169.105 73.325 169.275 ;
        RECT 73.615 169.105 73.785 169.275 ;
        RECT 74.075 169.105 74.245 169.275 ;
        RECT 74.535 169.105 74.705 169.275 ;
        RECT 74.995 169.105 75.165 169.275 ;
        RECT 75.455 169.105 75.625 169.275 ;
        RECT 75.915 169.105 76.085 169.275 ;
        RECT 76.375 169.105 76.545 169.275 ;
        RECT 76.835 169.105 77.005 169.275 ;
        RECT 77.295 169.105 77.465 169.275 ;
        RECT 77.755 169.105 77.925 169.275 ;
        RECT 78.215 169.105 78.385 169.275 ;
        RECT 78.675 169.105 78.845 169.275 ;
        RECT 79.135 169.105 79.305 169.275 ;
        RECT 79.595 169.105 79.765 169.275 ;
        RECT 80.055 169.105 80.225 169.275 ;
        RECT 80.515 169.105 80.685 169.275 ;
        RECT 80.975 169.105 81.145 169.275 ;
        RECT 81.435 169.105 81.605 169.275 ;
        RECT 81.895 169.105 82.065 169.275 ;
        RECT 82.355 169.105 82.525 169.275 ;
        RECT 82.815 169.105 82.985 169.275 ;
        RECT 83.275 169.105 83.445 169.275 ;
        RECT 83.735 169.105 83.905 169.275 ;
        RECT 84.195 169.105 84.365 169.275 ;
        RECT 84.655 169.105 84.825 169.275 ;
        RECT 85.115 169.105 85.285 169.275 ;
        RECT 85.575 169.105 85.745 169.275 ;
        RECT 86.035 169.105 86.205 169.275 ;
        RECT 86.495 169.105 86.665 169.275 ;
        RECT 86.955 169.105 87.125 169.275 ;
        RECT 87.415 169.105 87.585 169.275 ;
        RECT 87.875 169.105 88.045 169.275 ;
        RECT 88.335 169.105 88.505 169.275 ;
        RECT 88.795 169.105 88.965 169.275 ;
        RECT 89.255 169.105 89.425 169.275 ;
        RECT 89.715 169.105 89.885 169.275 ;
        RECT 90.175 169.105 90.345 169.275 ;
        RECT 90.635 169.105 90.805 169.275 ;
        RECT 91.095 169.105 91.265 169.275 ;
        RECT 91.555 169.105 91.725 169.275 ;
        RECT 92.015 169.105 92.185 169.275 ;
        RECT 92.475 169.105 92.645 169.275 ;
        RECT 92.935 169.105 93.105 169.275 ;
        RECT 93.395 169.105 93.565 169.275 ;
        RECT 93.855 169.105 94.025 169.275 ;
        RECT 94.315 169.105 94.485 169.275 ;
        RECT 94.775 169.105 94.945 169.275 ;
        RECT 95.235 169.105 95.405 169.275 ;
        RECT 95.695 169.105 95.865 169.275 ;
        RECT 96.155 169.105 96.325 169.275 ;
        RECT 96.615 169.105 96.785 169.275 ;
        RECT 97.075 169.105 97.245 169.275 ;
        RECT 97.535 169.105 97.705 169.275 ;
        RECT 97.995 169.105 98.165 169.275 ;
        RECT 98.455 169.105 98.625 169.275 ;
        RECT 98.915 169.105 99.085 169.275 ;
        RECT 99.375 169.105 99.545 169.275 ;
        RECT 99.835 169.105 100.005 169.275 ;
        RECT 100.295 169.105 100.465 169.275 ;
        RECT 100.755 169.105 100.925 169.275 ;
        RECT 101.215 169.105 101.385 169.275 ;
        RECT 101.675 169.105 101.845 169.275 ;
        RECT 102.135 169.105 102.305 169.275 ;
        RECT 102.595 169.105 102.765 169.275 ;
        RECT 103.055 169.105 103.225 169.275 ;
        RECT 103.515 169.105 103.685 169.275 ;
        RECT 103.975 169.105 104.145 169.275 ;
        RECT 104.435 169.105 104.605 169.275 ;
        RECT 104.895 169.105 105.065 169.275 ;
        RECT 105.355 169.105 105.525 169.275 ;
        RECT 105.815 169.105 105.985 169.275 ;
        RECT 106.275 169.105 106.445 169.275 ;
        RECT 106.735 169.105 106.905 169.275 ;
        RECT 107.195 169.105 107.365 169.275 ;
        RECT 107.655 169.105 107.825 169.275 ;
        RECT 108.115 169.105 108.285 169.275 ;
        RECT 108.575 169.105 108.745 169.275 ;
        RECT 109.035 169.105 109.205 169.275 ;
        RECT 109.495 169.105 109.665 169.275 ;
        RECT 109.955 169.105 110.125 169.275 ;
        RECT 110.415 169.105 110.585 169.275 ;
        RECT 110.875 169.105 111.045 169.275 ;
        RECT 111.335 169.105 111.505 169.275 ;
        RECT 111.795 169.105 111.965 169.275 ;
        RECT 112.255 169.105 112.425 169.275 ;
        RECT 112.715 169.105 112.885 169.275 ;
        RECT 113.175 169.105 113.345 169.275 ;
        RECT 113.635 169.105 113.805 169.275 ;
        RECT 114.095 169.105 114.265 169.275 ;
        RECT 114.555 169.105 114.725 169.275 ;
        RECT 115.015 169.105 115.185 169.275 ;
        RECT 115.475 169.105 115.645 169.275 ;
        RECT 115.935 169.105 116.105 169.275 ;
        RECT 116.395 169.105 116.565 169.275 ;
        RECT 116.855 169.105 117.025 169.275 ;
        RECT 117.315 169.105 117.485 169.275 ;
        RECT 117.775 169.105 117.945 169.275 ;
        RECT 118.235 169.105 118.405 169.275 ;
        RECT 118.695 169.105 118.865 169.275 ;
        RECT 119.155 169.105 119.325 169.275 ;
        RECT 119.615 169.105 119.785 169.275 ;
        RECT 120.075 169.105 120.245 169.275 ;
        RECT 120.535 169.105 120.705 169.275 ;
        RECT 120.995 169.105 121.165 169.275 ;
        RECT 121.455 169.105 121.625 169.275 ;
        RECT 121.915 169.105 122.085 169.275 ;
        RECT 122.375 169.105 122.545 169.275 ;
        RECT 122.835 169.105 123.005 169.275 ;
        RECT 123.295 169.105 123.465 169.275 ;
        RECT 123.755 169.105 123.925 169.275 ;
        RECT 124.215 169.105 124.385 169.275 ;
        RECT 124.675 169.105 124.845 169.275 ;
        RECT 125.135 169.105 125.305 169.275 ;
        RECT 125.595 169.105 125.765 169.275 ;
        RECT 126.055 169.105 126.225 169.275 ;
        RECT 126.515 169.105 126.685 169.275 ;
        RECT 126.975 169.105 127.145 169.275 ;
        RECT 127.435 169.105 127.605 169.275 ;
        RECT 127.895 169.105 128.065 169.275 ;
        RECT 128.355 169.105 128.525 169.275 ;
        RECT 128.815 169.105 128.985 169.275 ;
        RECT 129.275 169.105 129.445 169.275 ;
        RECT 129.735 169.105 129.905 169.275 ;
        RECT 130.195 169.105 130.365 169.275 ;
        RECT 130.655 169.105 130.825 169.275 ;
        RECT 131.115 169.105 131.285 169.275 ;
        RECT 131.575 169.105 131.745 169.275 ;
        RECT 132.035 169.105 132.205 169.275 ;
        RECT 132.495 169.105 132.665 169.275 ;
        RECT 132.955 169.105 133.125 169.275 ;
        RECT 133.415 169.105 133.585 169.275 ;
        RECT 133.875 169.105 134.045 169.275 ;
        RECT 134.335 169.105 134.505 169.275 ;
        RECT 134.795 169.105 134.965 169.275 ;
        RECT 135.255 169.105 135.425 169.275 ;
        RECT 135.715 169.105 135.885 169.275 ;
        RECT 136.175 169.105 136.345 169.275 ;
        RECT 136.635 169.105 136.805 169.275 ;
        RECT 137.095 169.105 137.265 169.275 ;
        RECT 137.555 169.105 137.725 169.275 ;
        RECT 138.015 169.105 138.185 169.275 ;
        RECT 138.475 169.105 138.645 169.275 ;
        RECT 138.935 169.105 139.105 169.275 ;
        RECT 139.395 169.105 139.565 169.275 ;
        RECT 139.855 169.105 140.025 169.275 ;
        RECT 140.315 169.105 140.485 169.275 ;
        RECT 140.775 169.105 140.945 169.275 ;
        RECT 141.235 169.105 141.405 169.275 ;
        RECT 141.695 169.105 141.865 169.275 ;
        RECT 142.155 169.105 142.325 169.275 ;
        RECT 142.615 169.105 142.785 169.275 ;
        RECT 143.075 169.105 143.245 169.275 ;
        RECT 143.535 169.105 143.705 169.275 ;
        RECT 143.995 169.105 144.165 169.275 ;
        RECT 144.455 169.105 144.625 169.275 ;
        RECT 144.915 169.105 145.085 169.275 ;
        RECT 145.375 169.105 145.545 169.275 ;
        RECT 145.835 169.105 146.005 169.275 ;
        RECT 146.295 169.105 146.465 169.275 ;
        RECT 146.755 169.105 146.925 169.275 ;
        RECT 147.215 169.105 147.385 169.275 ;
        RECT 147.675 169.105 147.845 169.275 ;
        RECT 148.135 169.105 148.305 169.275 ;
        RECT 148.595 169.105 148.765 169.275 ;
        RECT 149.055 169.105 149.225 169.275 ;
        RECT 149.515 169.105 149.685 169.275 ;
        RECT 149.975 169.105 150.145 169.275 ;
        RECT 150.435 169.105 150.605 169.275 ;
        RECT 150.895 169.105 151.065 169.275 ;
        RECT 151.355 169.105 151.525 169.275 ;
        RECT 151.815 169.105 151.985 169.275 ;
        RECT 152.275 169.105 152.445 169.275 ;
        RECT 152.735 169.105 152.905 169.275 ;
        RECT 153.195 169.105 153.365 169.275 ;
        RECT 153.655 169.105 153.825 169.275 ;
        RECT 154.115 169.105 154.285 169.275 ;
        RECT 154.575 169.105 154.745 169.275 ;
        RECT 155.035 169.105 155.205 169.275 ;
        RECT 155.495 169.105 155.665 169.275 ;
        RECT 155.955 169.105 156.125 169.275 ;
        RECT 72.720 168.255 72.890 168.425 ;
        RECT 72.235 167.575 72.405 167.745 ;
        RECT 73.115 167.915 73.285 168.085 ;
        RECT 73.570 167.235 73.740 167.405 ;
        RECT 74.820 168.255 74.990 168.425 ;
        RECT 74.305 167.915 74.475 168.085 ;
        RECT 76.390 168.255 76.560 168.425 ;
        RECT 76.825 167.915 76.995 168.085 ;
        RECT 80.515 168.255 80.685 168.425 ;
        RECT 79.595 167.575 79.765 167.745 ;
        RECT 79.135 166.895 79.305 167.065 ;
        RECT 81.435 167.915 81.605 168.085 ;
        RECT 80.975 167.575 81.145 167.745 ;
        RECT 87.875 168.255 88.045 168.425 ;
        RECT 86.955 167.575 87.125 167.745 ;
        RECT 89.255 168.595 89.425 168.765 ;
        RECT 88.335 167.575 88.505 167.745 ;
        RECT 89.255 167.575 89.425 167.745 ;
        RECT 92.475 166.895 92.645 167.065 ;
        RECT 98.915 167.575 99.085 167.745 ;
        RECT 102.595 167.915 102.765 168.085 ;
        RECT 100.295 167.575 100.465 167.745 ;
        RECT 101.215 167.575 101.385 167.745 ;
        RECT 101.805 167.235 101.975 167.405 ;
        RECT 99.375 166.895 99.545 167.065 ;
        RECT 113.635 167.575 113.805 167.745 ;
        RECT 120.075 168.255 120.245 168.425 ;
        RECT 114.555 166.895 114.725 167.065 ;
        RECT 117.645 167.235 117.815 167.405 ;
        RECT 118.235 167.575 118.405 167.745 ;
        RECT 118.695 167.575 118.865 167.745 ;
        RECT 119.155 167.575 119.325 167.745 ;
        RECT 121.020 168.255 121.190 168.425 ;
        RECT 120.535 167.575 120.705 167.745 ;
        RECT 121.415 167.915 121.585 168.085 ;
        RECT 121.815 167.235 121.985 167.405 ;
        RECT 123.120 168.255 123.290 168.425 ;
        RECT 122.605 167.915 122.775 168.085 ;
        RECT 124.690 168.255 124.860 168.425 ;
        RECT 125.125 167.915 125.295 168.085 ;
        RECT 127.435 168.595 127.605 168.765 ;
        RECT 130.195 168.595 130.365 168.765 ;
        RECT 129.275 167.575 129.445 167.745 ;
        RECT 129.735 167.575 129.905 167.745 ;
        RECT 131.115 167.455 131.285 167.625 ;
        RECT 130.655 167.235 130.825 167.405 ;
        RECT 128.355 166.895 128.525 167.065 ;
        RECT 132.035 166.895 132.205 167.065 ;
        RECT 133.875 168.595 134.045 168.765 ;
        RECT 134.795 167.575 134.965 167.745 ;
        RECT 135.715 167.575 135.885 167.745 ;
        RECT 136.635 167.235 136.805 167.405 ;
        RECT 142.640 168.255 142.810 168.425 ;
        RECT 138.475 167.575 138.645 167.745 ;
        RECT 139.395 167.575 139.565 167.745 ;
        RECT 139.855 167.575 140.025 167.745 ;
        RECT 140.315 167.575 140.485 167.745 ;
        RECT 142.155 167.575 142.325 167.745 ;
        RECT 137.555 166.895 137.725 167.065 ;
        RECT 141.695 167.235 141.865 167.405 ;
        RECT 143.035 167.915 143.205 168.085 ;
        RECT 143.380 167.235 143.550 167.405 ;
        RECT 144.740 168.255 144.910 168.425 ;
        RECT 144.225 167.915 144.395 168.085 ;
        RECT 146.310 168.255 146.480 168.425 ;
        RECT 146.745 167.915 146.915 168.085 ;
        RECT 149.055 168.255 149.225 168.425 ;
        RECT 150.435 167.575 150.605 167.745 ;
        RECT 151.815 167.915 151.985 168.085 ;
        RECT 70.855 166.385 71.025 166.555 ;
        RECT 71.315 166.385 71.485 166.555 ;
        RECT 71.775 166.385 71.945 166.555 ;
        RECT 72.235 166.385 72.405 166.555 ;
        RECT 72.695 166.385 72.865 166.555 ;
        RECT 73.155 166.385 73.325 166.555 ;
        RECT 73.615 166.385 73.785 166.555 ;
        RECT 74.075 166.385 74.245 166.555 ;
        RECT 74.535 166.385 74.705 166.555 ;
        RECT 74.995 166.385 75.165 166.555 ;
        RECT 75.455 166.385 75.625 166.555 ;
        RECT 75.915 166.385 76.085 166.555 ;
        RECT 76.375 166.385 76.545 166.555 ;
        RECT 76.835 166.385 77.005 166.555 ;
        RECT 77.295 166.385 77.465 166.555 ;
        RECT 77.755 166.385 77.925 166.555 ;
        RECT 78.215 166.385 78.385 166.555 ;
        RECT 78.675 166.385 78.845 166.555 ;
        RECT 79.135 166.385 79.305 166.555 ;
        RECT 79.595 166.385 79.765 166.555 ;
        RECT 80.055 166.385 80.225 166.555 ;
        RECT 80.515 166.385 80.685 166.555 ;
        RECT 80.975 166.385 81.145 166.555 ;
        RECT 81.435 166.385 81.605 166.555 ;
        RECT 81.895 166.385 82.065 166.555 ;
        RECT 82.355 166.385 82.525 166.555 ;
        RECT 82.815 166.385 82.985 166.555 ;
        RECT 83.275 166.385 83.445 166.555 ;
        RECT 83.735 166.385 83.905 166.555 ;
        RECT 84.195 166.385 84.365 166.555 ;
        RECT 84.655 166.385 84.825 166.555 ;
        RECT 85.115 166.385 85.285 166.555 ;
        RECT 85.575 166.385 85.745 166.555 ;
        RECT 86.035 166.385 86.205 166.555 ;
        RECT 86.495 166.385 86.665 166.555 ;
        RECT 86.955 166.385 87.125 166.555 ;
        RECT 87.415 166.385 87.585 166.555 ;
        RECT 87.875 166.385 88.045 166.555 ;
        RECT 88.335 166.385 88.505 166.555 ;
        RECT 88.795 166.385 88.965 166.555 ;
        RECT 89.255 166.385 89.425 166.555 ;
        RECT 89.715 166.385 89.885 166.555 ;
        RECT 90.175 166.385 90.345 166.555 ;
        RECT 90.635 166.385 90.805 166.555 ;
        RECT 91.095 166.385 91.265 166.555 ;
        RECT 91.555 166.385 91.725 166.555 ;
        RECT 92.015 166.385 92.185 166.555 ;
        RECT 92.475 166.385 92.645 166.555 ;
        RECT 92.935 166.385 93.105 166.555 ;
        RECT 93.395 166.385 93.565 166.555 ;
        RECT 93.855 166.385 94.025 166.555 ;
        RECT 94.315 166.385 94.485 166.555 ;
        RECT 94.775 166.385 94.945 166.555 ;
        RECT 95.235 166.385 95.405 166.555 ;
        RECT 95.695 166.385 95.865 166.555 ;
        RECT 96.155 166.385 96.325 166.555 ;
        RECT 96.615 166.385 96.785 166.555 ;
        RECT 97.075 166.385 97.245 166.555 ;
        RECT 97.535 166.385 97.705 166.555 ;
        RECT 97.995 166.385 98.165 166.555 ;
        RECT 98.455 166.385 98.625 166.555 ;
        RECT 98.915 166.385 99.085 166.555 ;
        RECT 99.375 166.385 99.545 166.555 ;
        RECT 99.835 166.385 100.005 166.555 ;
        RECT 100.295 166.385 100.465 166.555 ;
        RECT 100.755 166.385 100.925 166.555 ;
        RECT 101.215 166.385 101.385 166.555 ;
        RECT 101.675 166.385 101.845 166.555 ;
        RECT 102.135 166.385 102.305 166.555 ;
        RECT 102.595 166.385 102.765 166.555 ;
        RECT 103.055 166.385 103.225 166.555 ;
        RECT 103.515 166.385 103.685 166.555 ;
        RECT 103.975 166.385 104.145 166.555 ;
        RECT 104.435 166.385 104.605 166.555 ;
        RECT 104.895 166.385 105.065 166.555 ;
        RECT 105.355 166.385 105.525 166.555 ;
        RECT 105.815 166.385 105.985 166.555 ;
        RECT 106.275 166.385 106.445 166.555 ;
        RECT 106.735 166.385 106.905 166.555 ;
        RECT 107.195 166.385 107.365 166.555 ;
        RECT 107.655 166.385 107.825 166.555 ;
        RECT 108.115 166.385 108.285 166.555 ;
        RECT 108.575 166.385 108.745 166.555 ;
        RECT 109.035 166.385 109.205 166.555 ;
        RECT 109.495 166.385 109.665 166.555 ;
        RECT 109.955 166.385 110.125 166.555 ;
        RECT 110.415 166.385 110.585 166.555 ;
        RECT 110.875 166.385 111.045 166.555 ;
        RECT 111.335 166.385 111.505 166.555 ;
        RECT 111.795 166.385 111.965 166.555 ;
        RECT 112.255 166.385 112.425 166.555 ;
        RECT 112.715 166.385 112.885 166.555 ;
        RECT 113.175 166.385 113.345 166.555 ;
        RECT 113.635 166.385 113.805 166.555 ;
        RECT 114.095 166.385 114.265 166.555 ;
        RECT 114.555 166.385 114.725 166.555 ;
        RECT 115.015 166.385 115.185 166.555 ;
        RECT 115.475 166.385 115.645 166.555 ;
        RECT 115.935 166.385 116.105 166.555 ;
        RECT 116.395 166.385 116.565 166.555 ;
        RECT 116.855 166.385 117.025 166.555 ;
        RECT 117.315 166.385 117.485 166.555 ;
        RECT 117.775 166.385 117.945 166.555 ;
        RECT 118.235 166.385 118.405 166.555 ;
        RECT 118.695 166.385 118.865 166.555 ;
        RECT 119.155 166.385 119.325 166.555 ;
        RECT 119.615 166.385 119.785 166.555 ;
        RECT 120.075 166.385 120.245 166.555 ;
        RECT 120.535 166.385 120.705 166.555 ;
        RECT 120.995 166.385 121.165 166.555 ;
        RECT 121.455 166.385 121.625 166.555 ;
        RECT 121.915 166.385 122.085 166.555 ;
        RECT 122.375 166.385 122.545 166.555 ;
        RECT 122.835 166.385 123.005 166.555 ;
        RECT 123.295 166.385 123.465 166.555 ;
        RECT 123.755 166.385 123.925 166.555 ;
        RECT 124.215 166.385 124.385 166.555 ;
        RECT 124.675 166.385 124.845 166.555 ;
        RECT 125.135 166.385 125.305 166.555 ;
        RECT 125.595 166.385 125.765 166.555 ;
        RECT 126.055 166.385 126.225 166.555 ;
        RECT 126.515 166.385 126.685 166.555 ;
        RECT 126.975 166.385 127.145 166.555 ;
        RECT 127.435 166.385 127.605 166.555 ;
        RECT 127.895 166.385 128.065 166.555 ;
        RECT 128.355 166.385 128.525 166.555 ;
        RECT 128.815 166.385 128.985 166.555 ;
        RECT 129.275 166.385 129.445 166.555 ;
        RECT 129.735 166.385 129.905 166.555 ;
        RECT 130.195 166.385 130.365 166.555 ;
        RECT 130.655 166.385 130.825 166.555 ;
        RECT 131.115 166.385 131.285 166.555 ;
        RECT 131.575 166.385 131.745 166.555 ;
        RECT 132.035 166.385 132.205 166.555 ;
        RECT 132.495 166.385 132.665 166.555 ;
        RECT 132.955 166.385 133.125 166.555 ;
        RECT 133.415 166.385 133.585 166.555 ;
        RECT 133.875 166.385 134.045 166.555 ;
        RECT 134.335 166.385 134.505 166.555 ;
        RECT 134.795 166.385 134.965 166.555 ;
        RECT 135.255 166.385 135.425 166.555 ;
        RECT 135.715 166.385 135.885 166.555 ;
        RECT 136.175 166.385 136.345 166.555 ;
        RECT 136.635 166.385 136.805 166.555 ;
        RECT 137.095 166.385 137.265 166.555 ;
        RECT 137.555 166.385 137.725 166.555 ;
        RECT 138.015 166.385 138.185 166.555 ;
        RECT 138.475 166.385 138.645 166.555 ;
        RECT 138.935 166.385 139.105 166.555 ;
        RECT 139.395 166.385 139.565 166.555 ;
        RECT 139.855 166.385 140.025 166.555 ;
        RECT 140.315 166.385 140.485 166.555 ;
        RECT 140.775 166.385 140.945 166.555 ;
        RECT 141.235 166.385 141.405 166.555 ;
        RECT 141.695 166.385 141.865 166.555 ;
        RECT 142.155 166.385 142.325 166.555 ;
        RECT 142.615 166.385 142.785 166.555 ;
        RECT 143.075 166.385 143.245 166.555 ;
        RECT 143.535 166.385 143.705 166.555 ;
        RECT 143.995 166.385 144.165 166.555 ;
        RECT 144.455 166.385 144.625 166.555 ;
        RECT 144.915 166.385 145.085 166.555 ;
        RECT 145.375 166.385 145.545 166.555 ;
        RECT 145.835 166.385 146.005 166.555 ;
        RECT 146.295 166.385 146.465 166.555 ;
        RECT 146.755 166.385 146.925 166.555 ;
        RECT 147.215 166.385 147.385 166.555 ;
        RECT 147.675 166.385 147.845 166.555 ;
        RECT 148.135 166.385 148.305 166.555 ;
        RECT 148.595 166.385 148.765 166.555 ;
        RECT 149.055 166.385 149.225 166.555 ;
        RECT 149.515 166.385 149.685 166.555 ;
        RECT 149.975 166.385 150.145 166.555 ;
        RECT 150.435 166.385 150.605 166.555 ;
        RECT 150.895 166.385 151.065 166.555 ;
        RECT 151.355 166.385 151.525 166.555 ;
        RECT 151.815 166.385 151.985 166.555 ;
        RECT 152.275 166.385 152.445 166.555 ;
        RECT 152.735 166.385 152.905 166.555 ;
        RECT 153.195 166.385 153.365 166.555 ;
        RECT 153.655 166.385 153.825 166.555 ;
        RECT 154.115 166.385 154.285 166.555 ;
        RECT 154.575 166.385 154.745 166.555 ;
        RECT 155.035 166.385 155.205 166.555 ;
        RECT 155.495 166.385 155.665 166.555 ;
        RECT 155.955 166.385 156.125 166.555 ;
        RECT 76.835 165.195 77.005 165.365 ;
        RECT 77.320 164.515 77.490 164.685 ;
        RECT 77.715 164.855 77.885 165.025 ;
        RECT 78.170 165.195 78.340 165.365 ;
        RECT 78.905 164.855 79.075 165.025 ;
        RECT 79.420 164.515 79.590 164.685 ;
        RECT 80.990 164.515 81.160 164.685 ;
        RECT 81.425 164.855 81.595 165.025 ;
        RECT 83.735 165.875 83.905 166.045 ;
        RECT 84.195 164.515 84.365 164.685 ;
        RECT 86.505 164.855 86.675 165.025 ;
        RECT 86.940 164.515 87.110 164.685 ;
        RECT 89.025 164.855 89.195 165.025 ;
        RECT 88.510 164.515 88.680 164.685 ;
        RECT 89.815 165.195 89.985 165.365 ;
        RECT 90.215 164.855 90.385 165.025 ;
        RECT 91.095 165.195 91.265 165.365 ;
        RECT 91.555 164.855 91.725 165.025 ;
        RECT 90.610 164.515 90.780 164.685 ;
        RECT 92.935 164.855 93.105 165.025 ;
        RECT 98.915 165.875 99.085 166.045 ;
        RECT 97.535 165.195 97.705 165.365 ;
        RECT 98.455 165.195 98.625 165.365 ;
        RECT 98.455 164.175 98.625 164.345 ;
        RECT 99.835 165.195 100.005 165.365 ;
        RECT 100.755 165.195 100.925 165.365 ;
        RECT 105.355 165.875 105.525 166.045 ;
        RECT 103.645 165.195 103.815 165.365 ;
        RECT 104.895 165.195 105.065 165.365 ;
        RECT 104.435 164.855 104.605 165.025 ;
        RECT 101.215 164.175 101.385 164.345 ;
        RECT 108.115 165.195 108.285 165.365 ;
        RECT 109.495 164.855 109.665 165.025 ;
        RECT 112.715 165.535 112.885 165.705 ;
        RECT 114.095 165.195 114.265 165.365 ;
        RECT 114.555 165.195 114.725 165.365 ;
        RECT 115.015 165.195 115.185 165.365 ;
        RECT 115.935 165.195 116.105 165.365 ;
        RECT 118.795 165.195 118.965 165.365 ;
        RECT 119.615 165.195 119.785 165.365 ;
        RECT 120.075 165.195 120.245 165.365 ;
        RECT 120.535 165.195 120.705 165.365 ;
        RECT 122.835 165.535 123.005 165.705 ;
        RECT 123.810 165.535 123.980 165.705 ;
        RECT 124.675 165.535 124.845 165.705 ;
        RECT 125.895 165.535 126.065 165.705 ;
        RECT 126.975 165.535 127.145 165.705 ;
        RECT 129.735 165.195 129.905 165.365 ;
        RECT 130.655 165.195 130.825 165.365 ;
        RECT 125.135 164.175 125.305 164.345 ;
        RECT 126.055 164.175 126.225 164.345 ;
        RECT 130.655 164.515 130.825 164.685 ;
        RECT 132.495 165.195 132.665 165.365 ;
        RECT 133.875 164.855 134.045 165.025 ;
        RECT 137.095 165.195 137.265 165.365 ;
        RECT 138.475 165.195 138.645 165.365 ;
        RECT 141.695 165.195 141.865 165.365 ;
        RECT 143.535 165.875 143.705 166.045 ;
        RECT 143.955 165.195 144.125 165.365 ;
        RECT 147.215 165.875 147.385 166.045 ;
        RECT 142.615 164.515 142.785 164.685 ;
        RECT 147.675 165.195 147.845 165.365 ;
        RECT 151.355 164.855 151.525 165.025 ;
        RECT 153.195 165.195 153.365 165.365 ;
        RECT 152.735 164.855 152.905 165.025 ;
        RECT 154.115 164.175 154.285 164.345 ;
        RECT 70.855 163.665 71.025 163.835 ;
        RECT 71.315 163.665 71.485 163.835 ;
        RECT 71.775 163.665 71.945 163.835 ;
        RECT 72.235 163.665 72.405 163.835 ;
        RECT 72.695 163.665 72.865 163.835 ;
        RECT 73.155 163.665 73.325 163.835 ;
        RECT 73.615 163.665 73.785 163.835 ;
        RECT 74.075 163.665 74.245 163.835 ;
        RECT 74.535 163.665 74.705 163.835 ;
        RECT 74.995 163.665 75.165 163.835 ;
        RECT 75.455 163.665 75.625 163.835 ;
        RECT 75.915 163.665 76.085 163.835 ;
        RECT 76.375 163.665 76.545 163.835 ;
        RECT 76.835 163.665 77.005 163.835 ;
        RECT 77.295 163.665 77.465 163.835 ;
        RECT 77.755 163.665 77.925 163.835 ;
        RECT 78.215 163.665 78.385 163.835 ;
        RECT 78.675 163.665 78.845 163.835 ;
        RECT 79.135 163.665 79.305 163.835 ;
        RECT 79.595 163.665 79.765 163.835 ;
        RECT 80.055 163.665 80.225 163.835 ;
        RECT 80.515 163.665 80.685 163.835 ;
        RECT 80.975 163.665 81.145 163.835 ;
        RECT 81.435 163.665 81.605 163.835 ;
        RECT 81.895 163.665 82.065 163.835 ;
        RECT 82.355 163.665 82.525 163.835 ;
        RECT 82.815 163.665 82.985 163.835 ;
        RECT 83.275 163.665 83.445 163.835 ;
        RECT 83.735 163.665 83.905 163.835 ;
        RECT 84.195 163.665 84.365 163.835 ;
        RECT 84.655 163.665 84.825 163.835 ;
        RECT 85.115 163.665 85.285 163.835 ;
        RECT 85.575 163.665 85.745 163.835 ;
        RECT 86.035 163.665 86.205 163.835 ;
        RECT 86.495 163.665 86.665 163.835 ;
        RECT 86.955 163.665 87.125 163.835 ;
        RECT 87.415 163.665 87.585 163.835 ;
        RECT 87.875 163.665 88.045 163.835 ;
        RECT 88.335 163.665 88.505 163.835 ;
        RECT 88.795 163.665 88.965 163.835 ;
        RECT 89.255 163.665 89.425 163.835 ;
        RECT 89.715 163.665 89.885 163.835 ;
        RECT 90.175 163.665 90.345 163.835 ;
        RECT 90.635 163.665 90.805 163.835 ;
        RECT 91.095 163.665 91.265 163.835 ;
        RECT 91.555 163.665 91.725 163.835 ;
        RECT 92.015 163.665 92.185 163.835 ;
        RECT 92.475 163.665 92.645 163.835 ;
        RECT 92.935 163.665 93.105 163.835 ;
        RECT 93.395 163.665 93.565 163.835 ;
        RECT 93.855 163.665 94.025 163.835 ;
        RECT 94.315 163.665 94.485 163.835 ;
        RECT 94.775 163.665 94.945 163.835 ;
        RECT 95.235 163.665 95.405 163.835 ;
        RECT 95.695 163.665 95.865 163.835 ;
        RECT 96.155 163.665 96.325 163.835 ;
        RECT 96.615 163.665 96.785 163.835 ;
        RECT 97.075 163.665 97.245 163.835 ;
        RECT 97.535 163.665 97.705 163.835 ;
        RECT 97.995 163.665 98.165 163.835 ;
        RECT 98.455 163.665 98.625 163.835 ;
        RECT 98.915 163.665 99.085 163.835 ;
        RECT 99.375 163.665 99.545 163.835 ;
        RECT 99.835 163.665 100.005 163.835 ;
        RECT 100.295 163.665 100.465 163.835 ;
        RECT 100.755 163.665 100.925 163.835 ;
        RECT 101.215 163.665 101.385 163.835 ;
        RECT 101.675 163.665 101.845 163.835 ;
        RECT 102.135 163.665 102.305 163.835 ;
        RECT 102.595 163.665 102.765 163.835 ;
        RECT 103.055 163.665 103.225 163.835 ;
        RECT 103.515 163.665 103.685 163.835 ;
        RECT 103.975 163.665 104.145 163.835 ;
        RECT 104.435 163.665 104.605 163.835 ;
        RECT 104.895 163.665 105.065 163.835 ;
        RECT 105.355 163.665 105.525 163.835 ;
        RECT 105.815 163.665 105.985 163.835 ;
        RECT 106.275 163.665 106.445 163.835 ;
        RECT 106.735 163.665 106.905 163.835 ;
        RECT 107.195 163.665 107.365 163.835 ;
        RECT 107.655 163.665 107.825 163.835 ;
        RECT 108.115 163.665 108.285 163.835 ;
        RECT 108.575 163.665 108.745 163.835 ;
        RECT 109.035 163.665 109.205 163.835 ;
        RECT 109.495 163.665 109.665 163.835 ;
        RECT 109.955 163.665 110.125 163.835 ;
        RECT 110.415 163.665 110.585 163.835 ;
        RECT 110.875 163.665 111.045 163.835 ;
        RECT 111.335 163.665 111.505 163.835 ;
        RECT 111.795 163.665 111.965 163.835 ;
        RECT 112.255 163.665 112.425 163.835 ;
        RECT 112.715 163.665 112.885 163.835 ;
        RECT 113.175 163.665 113.345 163.835 ;
        RECT 113.635 163.665 113.805 163.835 ;
        RECT 114.095 163.665 114.265 163.835 ;
        RECT 114.555 163.665 114.725 163.835 ;
        RECT 115.015 163.665 115.185 163.835 ;
        RECT 115.475 163.665 115.645 163.835 ;
        RECT 115.935 163.665 116.105 163.835 ;
        RECT 116.395 163.665 116.565 163.835 ;
        RECT 116.855 163.665 117.025 163.835 ;
        RECT 117.315 163.665 117.485 163.835 ;
        RECT 117.775 163.665 117.945 163.835 ;
        RECT 118.235 163.665 118.405 163.835 ;
        RECT 118.695 163.665 118.865 163.835 ;
        RECT 119.155 163.665 119.325 163.835 ;
        RECT 119.615 163.665 119.785 163.835 ;
        RECT 120.075 163.665 120.245 163.835 ;
        RECT 120.535 163.665 120.705 163.835 ;
        RECT 120.995 163.665 121.165 163.835 ;
        RECT 121.455 163.665 121.625 163.835 ;
        RECT 121.915 163.665 122.085 163.835 ;
        RECT 122.375 163.665 122.545 163.835 ;
        RECT 122.835 163.665 123.005 163.835 ;
        RECT 123.295 163.665 123.465 163.835 ;
        RECT 123.755 163.665 123.925 163.835 ;
        RECT 124.215 163.665 124.385 163.835 ;
        RECT 124.675 163.665 124.845 163.835 ;
        RECT 125.135 163.665 125.305 163.835 ;
        RECT 125.595 163.665 125.765 163.835 ;
        RECT 126.055 163.665 126.225 163.835 ;
        RECT 126.515 163.665 126.685 163.835 ;
        RECT 126.975 163.665 127.145 163.835 ;
        RECT 127.435 163.665 127.605 163.835 ;
        RECT 127.895 163.665 128.065 163.835 ;
        RECT 128.355 163.665 128.525 163.835 ;
        RECT 128.815 163.665 128.985 163.835 ;
        RECT 129.275 163.665 129.445 163.835 ;
        RECT 129.735 163.665 129.905 163.835 ;
        RECT 130.195 163.665 130.365 163.835 ;
        RECT 130.655 163.665 130.825 163.835 ;
        RECT 131.115 163.665 131.285 163.835 ;
        RECT 131.575 163.665 131.745 163.835 ;
        RECT 132.035 163.665 132.205 163.835 ;
        RECT 132.495 163.665 132.665 163.835 ;
        RECT 132.955 163.665 133.125 163.835 ;
        RECT 133.415 163.665 133.585 163.835 ;
        RECT 133.875 163.665 134.045 163.835 ;
        RECT 134.335 163.665 134.505 163.835 ;
        RECT 134.795 163.665 134.965 163.835 ;
        RECT 135.255 163.665 135.425 163.835 ;
        RECT 135.715 163.665 135.885 163.835 ;
        RECT 136.175 163.665 136.345 163.835 ;
        RECT 136.635 163.665 136.805 163.835 ;
        RECT 137.095 163.665 137.265 163.835 ;
        RECT 137.555 163.665 137.725 163.835 ;
        RECT 138.015 163.665 138.185 163.835 ;
        RECT 138.475 163.665 138.645 163.835 ;
        RECT 138.935 163.665 139.105 163.835 ;
        RECT 139.395 163.665 139.565 163.835 ;
        RECT 139.855 163.665 140.025 163.835 ;
        RECT 140.315 163.665 140.485 163.835 ;
        RECT 140.775 163.665 140.945 163.835 ;
        RECT 141.235 163.665 141.405 163.835 ;
        RECT 141.695 163.665 141.865 163.835 ;
        RECT 142.155 163.665 142.325 163.835 ;
        RECT 142.615 163.665 142.785 163.835 ;
        RECT 143.075 163.665 143.245 163.835 ;
        RECT 143.535 163.665 143.705 163.835 ;
        RECT 143.995 163.665 144.165 163.835 ;
        RECT 144.455 163.665 144.625 163.835 ;
        RECT 144.915 163.665 145.085 163.835 ;
        RECT 145.375 163.665 145.545 163.835 ;
        RECT 145.835 163.665 146.005 163.835 ;
        RECT 146.295 163.665 146.465 163.835 ;
        RECT 146.755 163.665 146.925 163.835 ;
        RECT 147.215 163.665 147.385 163.835 ;
        RECT 147.675 163.665 147.845 163.835 ;
        RECT 148.135 163.665 148.305 163.835 ;
        RECT 148.595 163.665 148.765 163.835 ;
        RECT 149.055 163.665 149.225 163.835 ;
        RECT 149.515 163.665 149.685 163.835 ;
        RECT 149.975 163.665 150.145 163.835 ;
        RECT 150.435 163.665 150.605 163.835 ;
        RECT 150.895 163.665 151.065 163.835 ;
        RECT 151.355 163.665 151.525 163.835 ;
        RECT 151.815 163.665 151.985 163.835 ;
        RECT 152.275 163.665 152.445 163.835 ;
        RECT 152.735 163.665 152.905 163.835 ;
        RECT 153.195 163.665 153.365 163.835 ;
        RECT 153.655 163.665 153.825 163.835 ;
        RECT 154.115 163.665 154.285 163.835 ;
        RECT 154.575 163.665 154.745 163.835 ;
        RECT 155.035 163.665 155.205 163.835 ;
        RECT 155.495 163.665 155.665 163.835 ;
        RECT 155.955 163.665 156.125 163.835 ;
        RECT 72.235 163.155 72.405 163.325 ;
        RECT 74.545 162.475 74.715 162.645 ;
        RECT 74.980 162.815 75.150 162.985 ;
        RECT 76.550 162.815 76.720 162.985 ;
        RECT 77.065 162.475 77.235 162.645 ;
        RECT 77.910 161.795 78.080 161.965 ;
        RECT 78.255 162.475 78.425 162.645 ;
        RECT 78.650 162.815 78.820 162.985 ;
        RECT 79.135 162.135 79.305 162.305 ;
        RECT 88.795 162.135 88.965 162.305 ;
        RECT 91.555 162.135 91.725 162.305 ;
        RECT 92.015 162.135 92.185 162.305 ;
        RECT 86.955 161.795 87.125 161.965 ;
        RECT 93.395 162.475 93.565 162.645 ;
        RECT 93.855 162.135 94.025 162.305 ;
        RECT 95.695 163.155 95.865 163.325 ;
        RECT 96.615 163.155 96.785 163.325 ;
        RECT 95.695 162.135 95.865 162.305 ;
        RECT 99.375 163.155 99.545 163.325 ;
        RECT 97.075 162.475 97.245 162.645 ;
        RECT 101.215 162.815 101.385 162.985 ;
        RECT 100.295 162.475 100.465 162.645 ;
        RECT 97.995 162.135 98.165 162.305 ;
        RECT 99.835 162.135 100.005 162.305 ;
        RECT 102.595 162.475 102.765 162.645 ;
        RECT 103.515 162.815 103.685 162.985 ;
        RECT 103.055 162.135 103.225 162.305 ;
        RECT 104.895 162.475 105.065 162.645 ;
        RECT 106.275 163.155 106.445 163.325 ;
        RECT 104.435 162.135 104.605 162.305 ;
        RECT 105.355 162.135 105.525 162.305 ;
        RECT 110.415 162.475 110.585 162.645 ;
        RECT 107.195 162.135 107.365 162.305 ;
        RECT 108.575 162.135 108.745 162.305 ;
        RECT 111.795 162.135 111.965 162.305 ;
        RECT 115.475 163.155 115.645 163.325 ;
        RECT 108.115 161.795 108.285 161.965 ;
        RECT 116.855 163.155 117.025 163.325 ;
        RECT 115.015 162.135 115.185 162.305 ;
        RECT 115.935 162.135 116.105 162.305 ;
        RECT 117.775 162.135 117.945 162.305 ;
        RECT 120.075 162.135 120.245 162.305 ;
        RECT 118.695 161.455 118.865 161.625 ;
        RECT 119.615 161.455 119.785 161.625 ;
        RECT 124.215 161.795 124.385 161.965 ;
        RECT 125.135 161.795 125.305 161.965 ;
        RECT 126.515 162.135 126.685 162.305 ;
        RECT 123.295 161.455 123.465 161.625 ;
        RECT 125.595 161.455 125.765 161.625 ;
        RECT 135.715 162.135 135.885 162.305 ;
        RECT 137.095 162.475 137.265 162.645 ;
        RECT 136.635 162.135 136.805 162.305 ;
        RECT 138.475 162.135 138.645 162.305 ;
        RECT 148.160 162.815 148.330 162.985 ;
        RECT 147.675 162.475 147.845 162.645 ;
        RECT 139.395 161.455 139.565 161.625 ;
        RECT 148.555 162.475 148.725 162.645 ;
        RECT 149.010 161.795 149.180 161.965 ;
        RECT 150.260 162.815 150.430 162.985 ;
        RECT 149.745 162.475 149.915 162.645 ;
        RECT 151.830 162.815 152.000 162.985 ;
        RECT 152.265 162.475 152.435 162.645 ;
        RECT 154.575 163.155 154.745 163.325 ;
        RECT 70.855 160.945 71.025 161.115 ;
        RECT 71.315 160.945 71.485 161.115 ;
        RECT 71.775 160.945 71.945 161.115 ;
        RECT 72.235 160.945 72.405 161.115 ;
        RECT 72.695 160.945 72.865 161.115 ;
        RECT 73.155 160.945 73.325 161.115 ;
        RECT 73.615 160.945 73.785 161.115 ;
        RECT 74.075 160.945 74.245 161.115 ;
        RECT 74.535 160.945 74.705 161.115 ;
        RECT 74.995 160.945 75.165 161.115 ;
        RECT 75.455 160.945 75.625 161.115 ;
        RECT 75.915 160.945 76.085 161.115 ;
        RECT 76.375 160.945 76.545 161.115 ;
        RECT 76.835 160.945 77.005 161.115 ;
        RECT 77.295 160.945 77.465 161.115 ;
        RECT 77.755 160.945 77.925 161.115 ;
        RECT 78.215 160.945 78.385 161.115 ;
        RECT 78.675 160.945 78.845 161.115 ;
        RECT 79.135 160.945 79.305 161.115 ;
        RECT 79.595 160.945 79.765 161.115 ;
        RECT 80.055 160.945 80.225 161.115 ;
        RECT 80.515 160.945 80.685 161.115 ;
        RECT 80.975 160.945 81.145 161.115 ;
        RECT 81.435 160.945 81.605 161.115 ;
        RECT 81.895 160.945 82.065 161.115 ;
        RECT 82.355 160.945 82.525 161.115 ;
        RECT 82.815 160.945 82.985 161.115 ;
        RECT 83.275 160.945 83.445 161.115 ;
        RECT 83.735 160.945 83.905 161.115 ;
        RECT 84.195 160.945 84.365 161.115 ;
        RECT 84.655 160.945 84.825 161.115 ;
        RECT 85.115 160.945 85.285 161.115 ;
        RECT 85.575 160.945 85.745 161.115 ;
        RECT 86.035 160.945 86.205 161.115 ;
        RECT 86.495 160.945 86.665 161.115 ;
        RECT 86.955 160.945 87.125 161.115 ;
        RECT 87.415 160.945 87.585 161.115 ;
        RECT 87.875 160.945 88.045 161.115 ;
        RECT 88.335 160.945 88.505 161.115 ;
        RECT 88.795 160.945 88.965 161.115 ;
        RECT 89.255 160.945 89.425 161.115 ;
        RECT 89.715 160.945 89.885 161.115 ;
        RECT 90.175 160.945 90.345 161.115 ;
        RECT 90.635 160.945 90.805 161.115 ;
        RECT 91.095 160.945 91.265 161.115 ;
        RECT 91.555 160.945 91.725 161.115 ;
        RECT 92.015 160.945 92.185 161.115 ;
        RECT 92.475 160.945 92.645 161.115 ;
        RECT 92.935 160.945 93.105 161.115 ;
        RECT 93.395 160.945 93.565 161.115 ;
        RECT 93.855 160.945 94.025 161.115 ;
        RECT 94.315 160.945 94.485 161.115 ;
        RECT 94.775 160.945 94.945 161.115 ;
        RECT 95.235 160.945 95.405 161.115 ;
        RECT 95.695 160.945 95.865 161.115 ;
        RECT 96.155 160.945 96.325 161.115 ;
        RECT 96.615 160.945 96.785 161.115 ;
        RECT 97.075 160.945 97.245 161.115 ;
        RECT 97.535 160.945 97.705 161.115 ;
        RECT 97.995 160.945 98.165 161.115 ;
        RECT 98.455 160.945 98.625 161.115 ;
        RECT 98.915 160.945 99.085 161.115 ;
        RECT 99.375 160.945 99.545 161.115 ;
        RECT 99.835 160.945 100.005 161.115 ;
        RECT 100.295 160.945 100.465 161.115 ;
        RECT 100.755 160.945 100.925 161.115 ;
        RECT 101.215 160.945 101.385 161.115 ;
        RECT 101.675 160.945 101.845 161.115 ;
        RECT 102.135 160.945 102.305 161.115 ;
        RECT 102.595 160.945 102.765 161.115 ;
        RECT 103.055 160.945 103.225 161.115 ;
        RECT 103.515 160.945 103.685 161.115 ;
        RECT 103.975 160.945 104.145 161.115 ;
        RECT 104.435 160.945 104.605 161.115 ;
        RECT 104.895 160.945 105.065 161.115 ;
        RECT 105.355 160.945 105.525 161.115 ;
        RECT 105.815 160.945 105.985 161.115 ;
        RECT 106.275 160.945 106.445 161.115 ;
        RECT 106.735 160.945 106.905 161.115 ;
        RECT 107.195 160.945 107.365 161.115 ;
        RECT 107.655 160.945 107.825 161.115 ;
        RECT 108.115 160.945 108.285 161.115 ;
        RECT 108.575 160.945 108.745 161.115 ;
        RECT 109.035 160.945 109.205 161.115 ;
        RECT 109.495 160.945 109.665 161.115 ;
        RECT 109.955 160.945 110.125 161.115 ;
        RECT 110.415 160.945 110.585 161.115 ;
        RECT 110.875 160.945 111.045 161.115 ;
        RECT 111.335 160.945 111.505 161.115 ;
        RECT 111.795 160.945 111.965 161.115 ;
        RECT 112.255 160.945 112.425 161.115 ;
        RECT 112.715 160.945 112.885 161.115 ;
        RECT 113.175 160.945 113.345 161.115 ;
        RECT 113.635 160.945 113.805 161.115 ;
        RECT 114.095 160.945 114.265 161.115 ;
        RECT 114.555 160.945 114.725 161.115 ;
        RECT 115.015 160.945 115.185 161.115 ;
        RECT 115.475 160.945 115.645 161.115 ;
        RECT 115.935 160.945 116.105 161.115 ;
        RECT 116.395 160.945 116.565 161.115 ;
        RECT 116.855 160.945 117.025 161.115 ;
        RECT 117.315 160.945 117.485 161.115 ;
        RECT 117.775 160.945 117.945 161.115 ;
        RECT 118.235 160.945 118.405 161.115 ;
        RECT 118.695 160.945 118.865 161.115 ;
        RECT 119.155 160.945 119.325 161.115 ;
        RECT 119.615 160.945 119.785 161.115 ;
        RECT 120.075 160.945 120.245 161.115 ;
        RECT 120.535 160.945 120.705 161.115 ;
        RECT 120.995 160.945 121.165 161.115 ;
        RECT 121.455 160.945 121.625 161.115 ;
        RECT 121.915 160.945 122.085 161.115 ;
        RECT 122.375 160.945 122.545 161.115 ;
        RECT 122.835 160.945 123.005 161.115 ;
        RECT 123.295 160.945 123.465 161.115 ;
        RECT 123.755 160.945 123.925 161.115 ;
        RECT 124.215 160.945 124.385 161.115 ;
        RECT 124.675 160.945 124.845 161.115 ;
        RECT 125.135 160.945 125.305 161.115 ;
        RECT 125.595 160.945 125.765 161.115 ;
        RECT 126.055 160.945 126.225 161.115 ;
        RECT 126.515 160.945 126.685 161.115 ;
        RECT 126.975 160.945 127.145 161.115 ;
        RECT 127.435 160.945 127.605 161.115 ;
        RECT 127.895 160.945 128.065 161.115 ;
        RECT 128.355 160.945 128.525 161.115 ;
        RECT 128.815 160.945 128.985 161.115 ;
        RECT 129.275 160.945 129.445 161.115 ;
        RECT 129.735 160.945 129.905 161.115 ;
        RECT 130.195 160.945 130.365 161.115 ;
        RECT 130.655 160.945 130.825 161.115 ;
        RECT 131.115 160.945 131.285 161.115 ;
        RECT 131.575 160.945 131.745 161.115 ;
        RECT 132.035 160.945 132.205 161.115 ;
        RECT 132.495 160.945 132.665 161.115 ;
        RECT 132.955 160.945 133.125 161.115 ;
        RECT 133.415 160.945 133.585 161.115 ;
        RECT 133.875 160.945 134.045 161.115 ;
        RECT 134.335 160.945 134.505 161.115 ;
        RECT 134.795 160.945 134.965 161.115 ;
        RECT 135.255 160.945 135.425 161.115 ;
        RECT 135.715 160.945 135.885 161.115 ;
        RECT 136.175 160.945 136.345 161.115 ;
        RECT 136.635 160.945 136.805 161.115 ;
        RECT 137.095 160.945 137.265 161.115 ;
        RECT 137.555 160.945 137.725 161.115 ;
        RECT 138.015 160.945 138.185 161.115 ;
        RECT 138.475 160.945 138.645 161.115 ;
        RECT 138.935 160.945 139.105 161.115 ;
        RECT 139.395 160.945 139.565 161.115 ;
        RECT 139.855 160.945 140.025 161.115 ;
        RECT 140.315 160.945 140.485 161.115 ;
        RECT 140.775 160.945 140.945 161.115 ;
        RECT 141.235 160.945 141.405 161.115 ;
        RECT 141.695 160.945 141.865 161.115 ;
        RECT 142.155 160.945 142.325 161.115 ;
        RECT 142.615 160.945 142.785 161.115 ;
        RECT 143.075 160.945 143.245 161.115 ;
        RECT 143.535 160.945 143.705 161.115 ;
        RECT 143.995 160.945 144.165 161.115 ;
        RECT 144.455 160.945 144.625 161.115 ;
        RECT 144.915 160.945 145.085 161.115 ;
        RECT 145.375 160.945 145.545 161.115 ;
        RECT 145.835 160.945 146.005 161.115 ;
        RECT 146.295 160.945 146.465 161.115 ;
        RECT 146.755 160.945 146.925 161.115 ;
        RECT 147.215 160.945 147.385 161.115 ;
        RECT 147.675 160.945 147.845 161.115 ;
        RECT 148.135 160.945 148.305 161.115 ;
        RECT 148.595 160.945 148.765 161.115 ;
        RECT 149.055 160.945 149.225 161.115 ;
        RECT 149.515 160.945 149.685 161.115 ;
        RECT 149.975 160.945 150.145 161.115 ;
        RECT 150.435 160.945 150.605 161.115 ;
        RECT 150.895 160.945 151.065 161.115 ;
        RECT 151.355 160.945 151.525 161.115 ;
        RECT 151.815 160.945 151.985 161.115 ;
        RECT 152.275 160.945 152.445 161.115 ;
        RECT 152.735 160.945 152.905 161.115 ;
        RECT 153.195 160.945 153.365 161.115 ;
        RECT 153.655 160.945 153.825 161.115 ;
        RECT 154.115 160.945 154.285 161.115 ;
        RECT 154.575 160.945 154.745 161.115 ;
        RECT 155.035 160.945 155.205 161.115 ;
        RECT 155.495 160.945 155.665 161.115 ;
        RECT 155.955 160.945 156.125 161.115 ;
        RECT 76.375 159.075 76.545 159.245 ;
        RECT 77.295 159.415 77.465 159.585 ;
        RECT 78.675 159.755 78.845 159.925 ;
        RECT 78.215 159.415 78.385 159.585 ;
        RECT 76.835 158.735 77.005 158.905 ;
        RECT 80.515 159.075 80.685 159.245 ;
        RECT 81.895 159.755 82.065 159.925 ;
        RECT 84.195 160.435 84.365 160.605 ;
        RECT 82.815 159.755 82.985 159.925 ;
        RECT 83.275 159.755 83.445 159.925 ;
        RECT 80.975 158.735 81.145 158.905 ;
        RECT 88.335 159.755 88.505 159.925 ;
        RECT 89.715 159.755 89.885 159.925 ;
        RECT 89.255 158.735 89.425 158.905 ;
        RECT 91.095 160.095 91.265 160.265 ;
        RECT 90.635 159.075 90.805 159.245 ;
        RECT 93.395 159.755 93.565 159.925 ;
        RECT 92.935 159.415 93.105 159.585 ;
        RECT 94.775 159.755 94.945 159.925 ;
        RECT 93.395 158.735 93.565 158.905 ;
        RECT 94.315 158.735 94.485 158.905 ;
        RECT 97.535 160.095 97.705 160.265 ;
        RECT 98.585 160.435 98.755 160.605 ;
        RECT 95.695 159.075 95.865 159.245 ;
        RECT 99.835 160.095 100.005 160.265 ;
        RECT 99.375 159.075 99.545 159.245 ;
        RECT 101.675 160.435 101.845 160.605 ;
        RECT 100.915 160.095 101.085 160.265 ;
        RECT 98.455 158.735 98.625 158.905 ;
        RECT 100.755 158.735 100.925 158.905 ;
        RECT 108.575 159.415 108.745 159.585 ;
        RECT 109.955 159.415 110.125 159.585 ;
        RECT 119.615 159.755 119.785 159.925 ;
        RECT 120.535 159.755 120.705 159.925 ;
        RECT 120.075 158.735 120.245 158.905 ;
        RECT 121.915 159.755 122.085 159.925 ;
        RECT 123.755 159.755 123.925 159.925 ;
        RECT 125.135 159.755 125.305 159.925 ;
        RECT 120.995 159.075 121.165 159.245 ;
        RECT 124.215 158.735 124.385 158.905 ;
        RECT 126.055 158.735 126.225 158.905 ;
        RECT 126.515 159.755 126.685 159.925 ;
        RECT 127.435 159.755 127.605 159.925 ;
        RECT 128.815 159.755 128.985 159.925 ;
        RECT 129.275 159.755 129.445 159.925 ;
        RECT 128.355 159.415 128.525 159.585 ;
        RECT 130.195 159.755 130.365 159.925 ;
        RECT 130.655 159.755 130.825 159.925 ;
        RECT 135.255 159.755 135.425 159.925 ;
        RECT 136.195 159.755 136.365 159.925 ;
        RECT 131.575 159.075 131.745 159.245 ;
        RECT 136.635 159.415 136.805 159.585 ;
        RECT 138.015 159.755 138.185 159.925 ;
        RECT 139.395 159.755 139.565 159.925 ;
        RECT 144.455 160.435 144.625 160.605 ;
        RECT 140.315 159.755 140.485 159.925 ;
        RECT 140.775 159.755 140.945 159.925 ;
        RECT 138.935 158.735 139.105 158.905 ;
        RECT 142.155 159.755 142.325 159.925 ;
        RECT 143.995 159.755 144.165 159.925 ;
        RECT 145.375 160.095 145.545 160.265 ;
        RECT 144.915 159.755 145.085 159.925 ;
        RECT 143.075 158.735 143.245 158.905 ;
        RECT 146.295 159.755 146.465 159.925 ;
        RECT 148.595 160.095 148.765 160.265 ;
        RECT 149.595 160.435 149.765 160.605 ;
        RECT 147.215 158.735 147.385 158.905 ;
        RECT 150.435 159.075 150.605 159.245 ;
        RECT 149.515 158.735 149.685 158.905 ;
        RECT 150.895 160.435 151.065 160.605 ;
        RECT 151.815 159.755 151.985 159.925 ;
        RECT 70.855 158.225 71.025 158.395 ;
        RECT 71.315 158.225 71.485 158.395 ;
        RECT 71.775 158.225 71.945 158.395 ;
        RECT 72.235 158.225 72.405 158.395 ;
        RECT 72.695 158.225 72.865 158.395 ;
        RECT 73.155 158.225 73.325 158.395 ;
        RECT 73.615 158.225 73.785 158.395 ;
        RECT 74.075 158.225 74.245 158.395 ;
        RECT 74.535 158.225 74.705 158.395 ;
        RECT 74.995 158.225 75.165 158.395 ;
        RECT 75.455 158.225 75.625 158.395 ;
        RECT 75.915 158.225 76.085 158.395 ;
        RECT 76.375 158.225 76.545 158.395 ;
        RECT 76.835 158.225 77.005 158.395 ;
        RECT 77.295 158.225 77.465 158.395 ;
        RECT 77.755 158.225 77.925 158.395 ;
        RECT 78.215 158.225 78.385 158.395 ;
        RECT 78.675 158.225 78.845 158.395 ;
        RECT 79.135 158.225 79.305 158.395 ;
        RECT 79.595 158.225 79.765 158.395 ;
        RECT 80.055 158.225 80.225 158.395 ;
        RECT 80.515 158.225 80.685 158.395 ;
        RECT 80.975 158.225 81.145 158.395 ;
        RECT 81.435 158.225 81.605 158.395 ;
        RECT 81.895 158.225 82.065 158.395 ;
        RECT 82.355 158.225 82.525 158.395 ;
        RECT 82.815 158.225 82.985 158.395 ;
        RECT 83.275 158.225 83.445 158.395 ;
        RECT 83.735 158.225 83.905 158.395 ;
        RECT 84.195 158.225 84.365 158.395 ;
        RECT 84.655 158.225 84.825 158.395 ;
        RECT 85.115 158.225 85.285 158.395 ;
        RECT 85.575 158.225 85.745 158.395 ;
        RECT 86.035 158.225 86.205 158.395 ;
        RECT 86.495 158.225 86.665 158.395 ;
        RECT 86.955 158.225 87.125 158.395 ;
        RECT 87.415 158.225 87.585 158.395 ;
        RECT 87.875 158.225 88.045 158.395 ;
        RECT 88.335 158.225 88.505 158.395 ;
        RECT 88.795 158.225 88.965 158.395 ;
        RECT 89.255 158.225 89.425 158.395 ;
        RECT 89.715 158.225 89.885 158.395 ;
        RECT 90.175 158.225 90.345 158.395 ;
        RECT 90.635 158.225 90.805 158.395 ;
        RECT 91.095 158.225 91.265 158.395 ;
        RECT 91.555 158.225 91.725 158.395 ;
        RECT 92.015 158.225 92.185 158.395 ;
        RECT 92.475 158.225 92.645 158.395 ;
        RECT 92.935 158.225 93.105 158.395 ;
        RECT 93.395 158.225 93.565 158.395 ;
        RECT 93.855 158.225 94.025 158.395 ;
        RECT 94.315 158.225 94.485 158.395 ;
        RECT 94.775 158.225 94.945 158.395 ;
        RECT 95.235 158.225 95.405 158.395 ;
        RECT 95.695 158.225 95.865 158.395 ;
        RECT 96.155 158.225 96.325 158.395 ;
        RECT 96.615 158.225 96.785 158.395 ;
        RECT 97.075 158.225 97.245 158.395 ;
        RECT 97.535 158.225 97.705 158.395 ;
        RECT 97.995 158.225 98.165 158.395 ;
        RECT 98.455 158.225 98.625 158.395 ;
        RECT 98.915 158.225 99.085 158.395 ;
        RECT 99.375 158.225 99.545 158.395 ;
        RECT 99.835 158.225 100.005 158.395 ;
        RECT 100.295 158.225 100.465 158.395 ;
        RECT 100.755 158.225 100.925 158.395 ;
        RECT 101.215 158.225 101.385 158.395 ;
        RECT 101.675 158.225 101.845 158.395 ;
        RECT 102.135 158.225 102.305 158.395 ;
        RECT 102.595 158.225 102.765 158.395 ;
        RECT 103.055 158.225 103.225 158.395 ;
        RECT 103.515 158.225 103.685 158.395 ;
        RECT 103.975 158.225 104.145 158.395 ;
        RECT 104.435 158.225 104.605 158.395 ;
        RECT 104.895 158.225 105.065 158.395 ;
        RECT 105.355 158.225 105.525 158.395 ;
        RECT 105.815 158.225 105.985 158.395 ;
        RECT 106.275 158.225 106.445 158.395 ;
        RECT 106.735 158.225 106.905 158.395 ;
        RECT 107.195 158.225 107.365 158.395 ;
        RECT 107.655 158.225 107.825 158.395 ;
        RECT 108.115 158.225 108.285 158.395 ;
        RECT 108.575 158.225 108.745 158.395 ;
        RECT 109.035 158.225 109.205 158.395 ;
        RECT 109.495 158.225 109.665 158.395 ;
        RECT 109.955 158.225 110.125 158.395 ;
        RECT 110.415 158.225 110.585 158.395 ;
        RECT 110.875 158.225 111.045 158.395 ;
        RECT 111.335 158.225 111.505 158.395 ;
        RECT 111.795 158.225 111.965 158.395 ;
        RECT 112.255 158.225 112.425 158.395 ;
        RECT 112.715 158.225 112.885 158.395 ;
        RECT 113.175 158.225 113.345 158.395 ;
        RECT 113.635 158.225 113.805 158.395 ;
        RECT 114.095 158.225 114.265 158.395 ;
        RECT 114.555 158.225 114.725 158.395 ;
        RECT 115.015 158.225 115.185 158.395 ;
        RECT 115.475 158.225 115.645 158.395 ;
        RECT 115.935 158.225 116.105 158.395 ;
        RECT 116.395 158.225 116.565 158.395 ;
        RECT 116.855 158.225 117.025 158.395 ;
        RECT 117.315 158.225 117.485 158.395 ;
        RECT 117.775 158.225 117.945 158.395 ;
        RECT 118.235 158.225 118.405 158.395 ;
        RECT 118.695 158.225 118.865 158.395 ;
        RECT 119.155 158.225 119.325 158.395 ;
        RECT 119.615 158.225 119.785 158.395 ;
        RECT 120.075 158.225 120.245 158.395 ;
        RECT 120.535 158.225 120.705 158.395 ;
        RECT 120.995 158.225 121.165 158.395 ;
        RECT 121.455 158.225 121.625 158.395 ;
        RECT 121.915 158.225 122.085 158.395 ;
        RECT 122.375 158.225 122.545 158.395 ;
        RECT 122.835 158.225 123.005 158.395 ;
        RECT 123.295 158.225 123.465 158.395 ;
        RECT 123.755 158.225 123.925 158.395 ;
        RECT 124.215 158.225 124.385 158.395 ;
        RECT 124.675 158.225 124.845 158.395 ;
        RECT 125.135 158.225 125.305 158.395 ;
        RECT 125.595 158.225 125.765 158.395 ;
        RECT 126.055 158.225 126.225 158.395 ;
        RECT 126.515 158.225 126.685 158.395 ;
        RECT 126.975 158.225 127.145 158.395 ;
        RECT 127.435 158.225 127.605 158.395 ;
        RECT 127.895 158.225 128.065 158.395 ;
        RECT 128.355 158.225 128.525 158.395 ;
        RECT 128.815 158.225 128.985 158.395 ;
        RECT 129.275 158.225 129.445 158.395 ;
        RECT 129.735 158.225 129.905 158.395 ;
        RECT 130.195 158.225 130.365 158.395 ;
        RECT 130.655 158.225 130.825 158.395 ;
        RECT 131.115 158.225 131.285 158.395 ;
        RECT 131.575 158.225 131.745 158.395 ;
        RECT 132.035 158.225 132.205 158.395 ;
        RECT 132.495 158.225 132.665 158.395 ;
        RECT 132.955 158.225 133.125 158.395 ;
        RECT 133.415 158.225 133.585 158.395 ;
        RECT 133.875 158.225 134.045 158.395 ;
        RECT 134.335 158.225 134.505 158.395 ;
        RECT 134.795 158.225 134.965 158.395 ;
        RECT 135.255 158.225 135.425 158.395 ;
        RECT 135.715 158.225 135.885 158.395 ;
        RECT 136.175 158.225 136.345 158.395 ;
        RECT 136.635 158.225 136.805 158.395 ;
        RECT 137.095 158.225 137.265 158.395 ;
        RECT 137.555 158.225 137.725 158.395 ;
        RECT 138.015 158.225 138.185 158.395 ;
        RECT 138.475 158.225 138.645 158.395 ;
        RECT 138.935 158.225 139.105 158.395 ;
        RECT 139.395 158.225 139.565 158.395 ;
        RECT 139.855 158.225 140.025 158.395 ;
        RECT 140.315 158.225 140.485 158.395 ;
        RECT 140.775 158.225 140.945 158.395 ;
        RECT 141.235 158.225 141.405 158.395 ;
        RECT 141.695 158.225 141.865 158.395 ;
        RECT 142.155 158.225 142.325 158.395 ;
        RECT 142.615 158.225 142.785 158.395 ;
        RECT 143.075 158.225 143.245 158.395 ;
        RECT 143.535 158.225 143.705 158.395 ;
        RECT 143.995 158.225 144.165 158.395 ;
        RECT 144.455 158.225 144.625 158.395 ;
        RECT 144.915 158.225 145.085 158.395 ;
        RECT 145.375 158.225 145.545 158.395 ;
        RECT 145.835 158.225 146.005 158.395 ;
        RECT 146.295 158.225 146.465 158.395 ;
        RECT 146.755 158.225 146.925 158.395 ;
        RECT 147.215 158.225 147.385 158.395 ;
        RECT 147.675 158.225 147.845 158.395 ;
        RECT 148.135 158.225 148.305 158.395 ;
        RECT 148.595 158.225 148.765 158.395 ;
        RECT 149.055 158.225 149.225 158.395 ;
        RECT 149.515 158.225 149.685 158.395 ;
        RECT 149.975 158.225 150.145 158.395 ;
        RECT 150.435 158.225 150.605 158.395 ;
        RECT 150.895 158.225 151.065 158.395 ;
        RECT 151.355 158.225 151.525 158.395 ;
        RECT 151.815 158.225 151.985 158.395 ;
        RECT 152.275 158.225 152.445 158.395 ;
        RECT 152.735 158.225 152.905 158.395 ;
        RECT 153.195 158.225 153.365 158.395 ;
        RECT 153.655 158.225 153.825 158.395 ;
        RECT 154.115 158.225 154.285 158.395 ;
        RECT 154.575 158.225 154.745 158.395 ;
        RECT 155.035 158.225 155.205 158.395 ;
        RECT 155.495 158.225 155.665 158.395 ;
        RECT 155.955 158.225 156.125 158.395 ;
        RECT 78.215 157.715 78.385 157.885 ;
        RECT 79.595 157.375 79.765 157.545 ;
        RECT 77.755 156.695 77.925 156.865 ;
        RECT 78.675 156.695 78.845 156.865 ;
        RECT 79.135 156.695 79.305 156.865 ;
        RECT 80.055 156.695 80.225 156.865 ;
        RECT 80.515 156.695 80.685 156.865 ;
        RECT 81.435 156.695 81.605 156.865 ;
        RECT 82.355 156.695 82.525 156.865 ;
        RECT 86.495 157.035 86.665 157.205 ;
        RECT 88.795 157.375 88.965 157.545 ;
        RECT 86.955 156.695 87.125 156.865 ;
        RECT 87.875 156.695 88.045 156.865 ;
        RECT 89.255 156.355 89.425 156.525 ;
        RECT 90.175 157.035 90.345 157.205 ;
        RECT 91.095 157.715 91.265 157.885 ;
        RECT 93.855 157.715 94.025 157.885 ;
        RECT 90.635 156.695 90.805 156.865 ;
        RECT 91.095 156.695 91.265 156.865 ;
        RECT 92.015 156.695 92.185 156.865 ;
        RECT 92.935 156.695 93.105 156.865 ;
        RECT 95.695 157.715 95.865 157.885 ;
        RECT 94.775 156.695 94.945 156.865 ;
        RECT 96.155 156.695 96.325 156.865 ;
        RECT 98.455 157.715 98.625 157.885 ;
        RECT 97.535 156.695 97.705 156.865 ;
        RECT 97.075 156.015 97.245 156.185 ;
        RECT 99.835 156.695 100.005 156.865 ;
        RECT 110.875 156.695 111.045 156.865 ;
        RECT 111.795 156.695 111.965 156.865 ;
        RECT 112.255 156.695 112.425 156.865 ;
        RECT 112.715 156.695 112.885 156.865 ;
        RECT 100.755 156.015 100.925 156.185 ;
        RECT 109.955 156.015 110.125 156.185 ;
        RECT 113.635 156.695 113.805 156.865 ;
        RECT 114.095 156.695 114.265 156.865 ;
        RECT 114.555 156.695 114.725 156.865 ;
        RECT 115.475 156.695 115.645 156.865 ;
        RECT 118.695 157.715 118.865 157.885 ;
        RECT 117.775 156.695 117.945 156.865 ;
        RECT 116.395 156.015 116.565 156.185 ;
        RECT 121.455 157.715 121.625 157.885 ;
        RECT 119.155 156.695 119.325 156.865 ;
        RECT 120.075 156.695 120.245 156.865 ;
        RECT 120.535 156.695 120.705 156.865 ;
        RECT 119.615 156.015 119.785 156.185 ;
        RECT 124.215 157.035 124.385 157.205 ;
        RECT 124.675 157.035 124.845 157.205 ;
        RECT 125.135 156.695 125.305 156.865 ;
        RECT 125.595 157.035 125.765 157.205 ;
        RECT 128.355 157.715 128.525 157.885 ;
        RECT 123.295 156.015 123.465 156.185 ;
        RECT 129.735 157.715 129.905 157.885 ;
        RECT 129.275 156.695 129.445 156.865 ;
        RECT 130.655 156.695 130.825 156.865 ;
        RECT 138.015 157.375 138.185 157.545 ;
        RECT 137.555 157.035 137.725 157.205 ;
        RECT 138.935 156.695 139.105 156.865 ;
        RECT 140.775 157.375 140.945 157.545 ;
        RECT 140.315 157.035 140.485 157.205 ;
        RECT 141.695 156.695 141.865 156.865 ;
        RECT 139.855 156.015 140.025 156.185 ;
        RECT 142.615 156.015 142.785 156.185 ;
        RECT 144.915 157.375 145.085 157.545 ;
        RECT 143.995 156.695 144.165 156.865 ;
        RECT 145.375 156.695 145.545 156.865 ;
        RECT 143.075 156.015 143.245 156.185 ;
        RECT 151.355 156.695 151.525 156.865 ;
        RECT 152.275 156.695 152.445 156.865 ;
        RECT 151.815 156.355 151.985 156.525 ;
        RECT 70.855 155.505 71.025 155.675 ;
        RECT 71.315 155.505 71.485 155.675 ;
        RECT 71.775 155.505 71.945 155.675 ;
        RECT 72.235 155.505 72.405 155.675 ;
        RECT 72.695 155.505 72.865 155.675 ;
        RECT 73.155 155.505 73.325 155.675 ;
        RECT 73.615 155.505 73.785 155.675 ;
        RECT 74.075 155.505 74.245 155.675 ;
        RECT 74.535 155.505 74.705 155.675 ;
        RECT 74.995 155.505 75.165 155.675 ;
        RECT 75.455 155.505 75.625 155.675 ;
        RECT 75.915 155.505 76.085 155.675 ;
        RECT 76.375 155.505 76.545 155.675 ;
        RECT 76.835 155.505 77.005 155.675 ;
        RECT 77.295 155.505 77.465 155.675 ;
        RECT 77.755 155.505 77.925 155.675 ;
        RECT 78.215 155.505 78.385 155.675 ;
        RECT 78.675 155.505 78.845 155.675 ;
        RECT 79.135 155.505 79.305 155.675 ;
        RECT 79.595 155.505 79.765 155.675 ;
        RECT 80.055 155.505 80.225 155.675 ;
        RECT 80.515 155.505 80.685 155.675 ;
        RECT 80.975 155.505 81.145 155.675 ;
        RECT 81.435 155.505 81.605 155.675 ;
        RECT 81.895 155.505 82.065 155.675 ;
        RECT 82.355 155.505 82.525 155.675 ;
        RECT 82.815 155.505 82.985 155.675 ;
        RECT 83.275 155.505 83.445 155.675 ;
        RECT 83.735 155.505 83.905 155.675 ;
        RECT 84.195 155.505 84.365 155.675 ;
        RECT 84.655 155.505 84.825 155.675 ;
        RECT 85.115 155.505 85.285 155.675 ;
        RECT 85.575 155.505 85.745 155.675 ;
        RECT 86.035 155.505 86.205 155.675 ;
        RECT 86.495 155.505 86.665 155.675 ;
        RECT 86.955 155.505 87.125 155.675 ;
        RECT 87.415 155.505 87.585 155.675 ;
        RECT 87.875 155.505 88.045 155.675 ;
        RECT 88.335 155.505 88.505 155.675 ;
        RECT 88.795 155.505 88.965 155.675 ;
        RECT 89.255 155.505 89.425 155.675 ;
        RECT 89.715 155.505 89.885 155.675 ;
        RECT 90.175 155.505 90.345 155.675 ;
        RECT 90.635 155.505 90.805 155.675 ;
        RECT 91.095 155.505 91.265 155.675 ;
        RECT 91.555 155.505 91.725 155.675 ;
        RECT 92.015 155.505 92.185 155.675 ;
        RECT 92.475 155.505 92.645 155.675 ;
        RECT 92.935 155.505 93.105 155.675 ;
        RECT 93.395 155.505 93.565 155.675 ;
        RECT 93.855 155.505 94.025 155.675 ;
        RECT 94.315 155.505 94.485 155.675 ;
        RECT 94.775 155.505 94.945 155.675 ;
        RECT 95.235 155.505 95.405 155.675 ;
        RECT 95.695 155.505 95.865 155.675 ;
        RECT 96.155 155.505 96.325 155.675 ;
        RECT 96.615 155.505 96.785 155.675 ;
        RECT 97.075 155.505 97.245 155.675 ;
        RECT 97.535 155.505 97.705 155.675 ;
        RECT 97.995 155.505 98.165 155.675 ;
        RECT 98.455 155.505 98.625 155.675 ;
        RECT 98.915 155.505 99.085 155.675 ;
        RECT 99.375 155.505 99.545 155.675 ;
        RECT 99.835 155.505 100.005 155.675 ;
        RECT 100.295 155.505 100.465 155.675 ;
        RECT 100.755 155.505 100.925 155.675 ;
        RECT 101.215 155.505 101.385 155.675 ;
        RECT 101.675 155.505 101.845 155.675 ;
        RECT 102.135 155.505 102.305 155.675 ;
        RECT 102.595 155.505 102.765 155.675 ;
        RECT 103.055 155.505 103.225 155.675 ;
        RECT 103.515 155.505 103.685 155.675 ;
        RECT 103.975 155.505 104.145 155.675 ;
        RECT 104.435 155.505 104.605 155.675 ;
        RECT 104.895 155.505 105.065 155.675 ;
        RECT 105.355 155.505 105.525 155.675 ;
        RECT 105.815 155.505 105.985 155.675 ;
        RECT 106.275 155.505 106.445 155.675 ;
        RECT 106.735 155.505 106.905 155.675 ;
        RECT 107.195 155.505 107.365 155.675 ;
        RECT 107.655 155.505 107.825 155.675 ;
        RECT 108.115 155.505 108.285 155.675 ;
        RECT 108.575 155.505 108.745 155.675 ;
        RECT 109.035 155.505 109.205 155.675 ;
        RECT 109.495 155.505 109.665 155.675 ;
        RECT 109.955 155.505 110.125 155.675 ;
        RECT 110.415 155.505 110.585 155.675 ;
        RECT 110.875 155.505 111.045 155.675 ;
        RECT 111.335 155.505 111.505 155.675 ;
        RECT 111.795 155.505 111.965 155.675 ;
        RECT 112.255 155.505 112.425 155.675 ;
        RECT 112.715 155.505 112.885 155.675 ;
        RECT 113.175 155.505 113.345 155.675 ;
        RECT 113.635 155.505 113.805 155.675 ;
        RECT 114.095 155.505 114.265 155.675 ;
        RECT 114.555 155.505 114.725 155.675 ;
        RECT 115.015 155.505 115.185 155.675 ;
        RECT 115.475 155.505 115.645 155.675 ;
        RECT 115.935 155.505 116.105 155.675 ;
        RECT 116.395 155.505 116.565 155.675 ;
        RECT 116.855 155.505 117.025 155.675 ;
        RECT 117.315 155.505 117.485 155.675 ;
        RECT 117.775 155.505 117.945 155.675 ;
        RECT 118.235 155.505 118.405 155.675 ;
        RECT 118.695 155.505 118.865 155.675 ;
        RECT 119.155 155.505 119.325 155.675 ;
        RECT 119.615 155.505 119.785 155.675 ;
        RECT 120.075 155.505 120.245 155.675 ;
        RECT 120.535 155.505 120.705 155.675 ;
        RECT 120.995 155.505 121.165 155.675 ;
        RECT 121.455 155.505 121.625 155.675 ;
        RECT 121.915 155.505 122.085 155.675 ;
        RECT 122.375 155.505 122.545 155.675 ;
        RECT 122.835 155.505 123.005 155.675 ;
        RECT 123.295 155.505 123.465 155.675 ;
        RECT 123.755 155.505 123.925 155.675 ;
        RECT 124.215 155.505 124.385 155.675 ;
        RECT 124.675 155.505 124.845 155.675 ;
        RECT 125.135 155.505 125.305 155.675 ;
        RECT 125.595 155.505 125.765 155.675 ;
        RECT 126.055 155.505 126.225 155.675 ;
        RECT 126.515 155.505 126.685 155.675 ;
        RECT 126.975 155.505 127.145 155.675 ;
        RECT 127.435 155.505 127.605 155.675 ;
        RECT 127.895 155.505 128.065 155.675 ;
        RECT 128.355 155.505 128.525 155.675 ;
        RECT 128.815 155.505 128.985 155.675 ;
        RECT 129.275 155.505 129.445 155.675 ;
        RECT 129.735 155.505 129.905 155.675 ;
        RECT 130.195 155.505 130.365 155.675 ;
        RECT 130.655 155.505 130.825 155.675 ;
        RECT 131.115 155.505 131.285 155.675 ;
        RECT 131.575 155.505 131.745 155.675 ;
        RECT 132.035 155.505 132.205 155.675 ;
        RECT 132.495 155.505 132.665 155.675 ;
        RECT 132.955 155.505 133.125 155.675 ;
        RECT 133.415 155.505 133.585 155.675 ;
        RECT 133.875 155.505 134.045 155.675 ;
        RECT 134.335 155.505 134.505 155.675 ;
        RECT 134.795 155.505 134.965 155.675 ;
        RECT 135.255 155.505 135.425 155.675 ;
        RECT 135.715 155.505 135.885 155.675 ;
        RECT 136.175 155.505 136.345 155.675 ;
        RECT 136.635 155.505 136.805 155.675 ;
        RECT 137.095 155.505 137.265 155.675 ;
        RECT 137.555 155.505 137.725 155.675 ;
        RECT 138.015 155.505 138.185 155.675 ;
        RECT 138.475 155.505 138.645 155.675 ;
        RECT 138.935 155.505 139.105 155.675 ;
        RECT 139.395 155.505 139.565 155.675 ;
        RECT 139.855 155.505 140.025 155.675 ;
        RECT 140.315 155.505 140.485 155.675 ;
        RECT 140.775 155.505 140.945 155.675 ;
        RECT 141.235 155.505 141.405 155.675 ;
        RECT 141.695 155.505 141.865 155.675 ;
        RECT 142.155 155.505 142.325 155.675 ;
        RECT 142.615 155.505 142.785 155.675 ;
        RECT 143.075 155.505 143.245 155.675 ;
        RECT 143.535 155.505 143.705 155.675 ;
        RECT 143.995 155.505 144.165 155.675 ;
        RECT 144.455 155.505 144.625 155.675 ;
        RECT 144.915 155.505 145.085 155.675 ;
        RECT 145.375 155.505 145.545 155.675 ;
        RECT 145.835 155.505 146.005 155.675 ;
        RECT 146.295 155.505 146.465 155.675 ;
        RECT 146.755 155.505 146.925 155.675 ;
        RECT 147.215 155.505 147.385 155.675 ;
        RECT 147.675 155.505 147.845 155.675 ;
        RECT 148.135 155.505 148.305 155.675 ;
        RECT 148.595 155.505 148.765 155.675 ;
        RECT 149.055 155.505 149.225 155.675 ;
        RECT 149.515 155.505 149.685 155.675 ;
        RECT 149.975 155.505 150.145 155.675 ;
        RECT 150.435 155.505 150.605 155.675 ;
        RECT 150.895 155.505 151.065 155.675 ;
        RECT 151.355 155.505 151.525 155.675 ;
        RECT 151.815 155.505 151.985 155.675 ;
        RECT 152.275 155.505 152.445 155.675 ;
        RECT 152.735 155.505 152.905 155.675 ;
        RECT 153.195 155.505 153.365 155.675 ;
        RECT 153.655 155.505 153.825 155.675 ;
        RECT 154.115 155.505 154.285 155.675 ;
        RECT 154.575 155.505 154.745 155.675 ;
        RECT 155.035 155.505 155.205 155.675 ;
        RECT 155.495 155.505 155.665 155.675 ;
        RECT 155.955 155.505 156.125 155.675 ;
        RECT 72.235 153.975 72.405 154.145 ;
        RECT 72.720 153.635 72.890 153.805 ;
        RECT 73.115 153.975 73.285 154.145 ;
        RECT 73.570 154.315 73.740 154.485 ;
        RECT 74.305 153.975 74.475 154.145 ;
        RECT 74.820 153.635 74.990 153.805 ;
        RECT 76.390 153.635 76.560 153.805 ;
        RECT 76.825 153.975 76.995 154.145 ;
        RECT 81.435 154.315 81.605 154.485 ;
        RECT 79.135 153.635 79.305 153.805 ;
        RECT 86.035 154.315 86.205 154.485 ;
        RECT 82.355 153.295 82.525 153.465 ;
        RECT 87.875 154.315 88.045 154.485 ;
        RECT 89.255 154.315 89.425 154.485 ;
        RECT 89.715 154.315 89.885 154.485 ;
        RECT 91.555 154.315 91.725 154.485 ;
        RECT 92.475 154.315 92.645 154.485 ;
        RECT 87.875 153.635 88.045 153.805 ;
        RECT 89.255 153.295 89.425 153.465 ;
        RECT 91.095 153.635 91.265 153.805 ;
        RECT 91.555 153.295 91.725 153.465 ;
        RECT 103.055 153.975 103.225 154.145 ;
        RECT 103.515 153.975 103.685 154.145 ;
        RECT 103.975 153.975 104.145 154.145 ;
        RECT 104.435 154.315 104.605 154.485 ;
        RECT 107.195 154.315 107.365 154.485 ;
        RECT 108.115 154.315 108.285 154.485 ;
        RECT 109.955 154.315 110.125 154.485 ;
        RECT 105.355 153.295 105.525 153.465 ;
        RECT 108.575 153.975 108.745 154.145 ;
        RECT 110.875 153.975 111.045 154.145 ;
        RECT 115.015 153.975 115.185 154.145 ;
        RECT 116.855 154.315 117.025 154.485 ;
        RECT 116.395 153.975 116.565 154.145 ;
        RECT 117.775 153.295 117.945 153.465 ;
        RECT 119.155 153.975 119.325 154.145 ;
        RECT 120.075 153.975 120.245 154.145 ;
        RECT 120.535 153.975 120.705 154.145 ;
        RECT 120.995 154.315 121.165 154.485 ;
        RECT 121.455 153.975 121.625 154.145 ;
        RECT 122.835 154.315 123.005 154.485 ;
        RECT 123.755 154.315 123.925 154.485 ;
        RECT 124.445 154.315 124.615 154.485 ;
        RECT 125.595 154.315 125.765 154.485 ;
        RECT 125.135 153.975 125.305 154.145 ;
        RECT 126.515 154.315 126.685 154.485 ;
        RECT 137.095 154.315 137.265 154.485 ;
        RECT 138.015 153.635 138.185 153.805 ;
        RECT 149.055 153.975 149.225 154.145 ;
        RECT 149.975 154.315 150.145 154.485 ;
        RECT 150.895 154.655 151.065 154.825 ;
        RECT 70.855 152.785 71.025 152.955 ;
        RECT 71.315 152.785 71.485 152.955 ;
        RECT 71.775 152.785 71.945 152.955 ;
        RECT 72.235 152.785 72.405 152.955 ;
        RECT 72.695 152.785 72.865 152.955 ;
        RECT 73.155 152.785 73.325 152.955 ;
        RECT 73.615 152.785 73.785 152.955 ;
        RECT 74.075 152.785 74.245 152.955 ;
        RECT 74.535 152.785 74.705 152.955 ;
        RECT 74.995 152.785 75.165 152.955 ;
        RECT 75.455 152.785 75.625 152.955 ;
        RECT 75.915 152.785 76.085 152.955 ;
        RECT 76.375 152.785 76.545 152.955 ;
        RECT 76.835 152.785 77.005 152.955 ;
        RECT 77.295 152.785 77.465 152.955 ;
        RECT 77.755 152.785 77.925 152.955 ;
        RECT 78.215 152.785 78.385 152.955 ;
        RECT 78.675 152.785 78.845 152.955 ;
        RECT 79.135 152.785 79.305 152.955 ;
        RECT 79.595 152.785 79.765 152.955 ;
        RECT 80.055 152.785 80.225 152.955 ;
        RECT 80.515 152.785 80.685 152.955 ;
        RECT 80.975 152.785 81.145 152.955 ;
        RECT 81.435 152.785 81.605 152.955 ;
        RECT 81.895 152.785 82.065 152.955 ;
        RECT 82.355 152.785 82.525 152.955 ;
        RECT 82.815 152.785 82.985 152.955 ;
        RECT 83.275 152.785 83.445 152.955 ;
        RECT 83.735 152.785 83.905 152.955 ;
        RECT 84.195 152.785 84.365 152.955 ;
        RECT 84.655 152.785 84.825 152.955 ;
        RECT 85.115 152.785 85.285 152.955 ;
        RECT 85.575 152.785 85.745 152.955 ;
        RECT 86.035 152.785 86.205 152.955 ;
        RECT 86.495 152.785 86.665 152.955 ;
        RECT 86.955 152.785 87.125 152.955 ;
        RECT 87.415 152.785 87.585 152.955 ;
        RECT 87.875 152.785 88.045 152.955 ;
        RECT 88.335 152.785 88.505 152.955 ;
        RECT 88.795 152.785 88.965 152.955 ;
        RECT 89.255 152.785 89.425 152.955 ;
        RECT 89.715 152.785 89.885 152.955 ;
        RECT 90.175 152.785 90.345 152.955 ;
        RECT 90.635 152.785 90.805 152.955 ;
        RECT 91.095 152.785 91.265 152.955 ;
        RECT 91.555 152.785 91.725 152.955 ;
        RECT 92.015 152.785 92.185 152.955 ;
        RECT 92.475 152.785 92.645 152.955 ;
        RECT 92.935 152.785 93.105 152.955 ;
        RECT 93.395 152.785 93.565 152.955 ;
        RECT 93.855 152.785 94.025 152.955 ;
        RECT 94.315 152.785 94.485 152.955 ;
        RECT 94.775 152.785 94.945 152.955 ;
        RECT 95.235 152.785 95.405 152.955 ;
        RECT 95.695 152.785 95.865 152.955 ;
        RECT 96.155 152.785 96.325 152.955 ;
        RECT 96.615 152.785 96.785 152.955 ;
        RECT 97.075 152.785 97.245 152.955 ;
        RECT 97.535 152.785 97.705 152.955 ;
        RECT 97.995 152.785 98.165 152.955 ;
        RECT 98.455 152.785 98.625 152.955 ;
        RECT 98.915 152.785 99.085 152.955 ;
        RECT 99.375 152.785 99.545 152.955 ;
        RECT 99.835 152.785 100.005 152.955 ;
        RECT 100.295 152.785 100.465 152.955 ;
        RECT 100.755 152.785 100.925 152.955 ;
        RECT 101.215 152.785 101.385 152.955 ;
        RECT 101.675 152.785 101.845 152.955 ;
        RECT 102.135 152.785 102.305 152.955 ;
        RECT 102.595 152.785 102.765 152.955 ;
        RECT 103.055 152.785 103.225 152.955 ;
        RECT 103.515 152.785 103.685 152.955 ;
        RECT 103.975 152.785 104.145 152.955 ;
        RECT 104.435 152.785 104.605 152.955 ;
        RECT 104.895 152.785 105.065 152.955 ;
        RECT 105.355 152.785 105.525 152.955 ;
        RECT 105.815 152.785 105.985 152.955 ;
        RECT 106.275 152.785 106.445 152.955 ;
        RECT 106.735 152.785 106.905 152.955 ;
        RECT 107.195 152.785 107.365 152.955 ;
        RECT 107.655 152.785 107.825 152.955 ;
        RECT 108.115 152.785 108.285 152.955 ;
        RECT 108.575 152.785 108.745 152.955 ;
        RECT 109.035 152.785 109.205 152.955 ;
        RECT 109.495 152.785 109.665 152.955 ;
        RECT 109.955 152.785 110.125 152.955 ;
        RECT 110.415 152.785 110.585 152.955 ;
        RECT 110.875 152.785 111.045 152.955 ;
        RECT 111.335 152.785 111.505 152.955 ;
        RECT 111.795 152.785 111.965 152.955 ;
        RECT 112.255 152.785 112.425 152.955 ;
        RECT 112.715 152.785 112.885 152.955 ;
        RECT 113.175 152.785 113.345 152.955 ;
        RECT 113.635 152.785 113.805 152.955 ;
        RECT 114.095 152.785 114.265 152.955 ;
        RECT 114.555 152.785 114.725 152.955 ;
        RECT 115.015 152.785 115.185 152.955 ;
        RECT 115.475 152.785 115.645 152.955 ;
        RECT 115.935 152.785 116.105 152.955 ;
        RECT 116.395 152.785 116.565 152.955 ;
        RECT 116.855 152.785 117.025 152.955 ;
        RECT 117.315 152.785 117.485 152.955 ;
        RECT 117.775 152.785 117.945 152.955 ;
        RECT 118.235 152.785 118.405 152.955 ;
        RECT 118.695 152.785 118.865 152.955 ;
        RECT 119.155 152.785 119.325 152.955 ;
        RECT 119.615 152.785 119.785 152.955 ;
        RECT 120.075 152.785 120.245 152.955 ;
        RECT 120.535 152.785 120.705 152.955 ;
        RECT 120.995 152.785 121.165 152.955 ;
        RECT 121.455 152.785 121.625 152.955 ;
        RECT 121.915 152.785 122.085 152.955 ;
        RECT 122.375 152.785 122.545 152.955 ;
        RECT 122.835 152.785 123.005 152.955 ;
        RECT 123.295 152.785 123.465 152.955 ;
        RECT 123.755 152.785 123.925 152.955 ;
        RECT 124.215 152.785 124.385 152.955 ;
        RECT 124.675 152.785 124.845 152.955 ;
        RECT 125.135 152.785 125.305 152.955 ;
        RECT 125.595 152.785 125.765 152.955 ;
        RECT 126.055 152.785 126.225 152.955 ;
        RECT 126.515 152.785 126.685 152.955 ;
        RECT 126.975 152.785 127.145 152.955 ;
        RECT 127.435 152.785 127.605 152.955 ;
        RECT 127.895 152.785 128.065 152.955 ;
        RECT 128.355 152.785 128.525 152.955 ;
        RECT 128.815 152.785 128.985 152.955 ;
        RECT 129.275 152.785 129.445 152.955 ;
        RECT 129.735 152.785 129.905 152.955 ;
        RECT 130.195 152.785 130.365 152.955 ;
        RECT 130.655 152.785 130.825 152.955 ;
        RECT 131.115 152.785 131.285 152.955 ;
        RECT 131.575 152.785 131.745 152.955 ;
        RECT 132.035 152.785 132.205 152.955 ;
        RECT 132.495 152.785 132.665 152.955 ;
        RECT 132.955 152.785 133.125 152.955 ;
        RECT 133.415 152.785 133.585 152.955 ;
        RECT 133.875 152.785 134.045 152.955 ;
        RECT 134.335 152.785 134.505 152.955 ;
        RECT 134.795 152.785 134.965 152.955 ;
        RECT 135.255 152.785 135.425 152.955 ;
        RECT 135.715 152.785 135.885 152.955 ;
        RECT 136.175 152.785 136.345 152.955 ;
        RECT 136.635 152.785 136.805 152.955 ;
        RECT 137.095 152.785 137.265 152.955 ;
        RECT 137.555 152.785 137.725 152.955 ;
        RECT 138.015 152.785 138.185 152.955 ;
        RECT 138.475 152.785 138.645 152.955 ;
        RECT 138.935 152.785 139.105 152.955 ;
        RECT 139.395 152.785 139.565 152.955 ;
        RECT 139.855 152.785 140.025 152.955 ;
        RECT 140.315 152.785 140.485 152.955 ;
        RECT 140.775 152.785 140.945 152.955 ;
        RECT 141.235 152.785 141.405 152.955 ;
        RECT 141.695 152.785 141.865 152.955 ;
        RECT 142.155 152.785 142.325 152.955 ;
        RECT 142.615 152.785 142.785 152.955 ;
        RECT 143.075 152.785 143.245 152.955 ;
        RECT 143.535 152.785 143.705 152.955 ;
        RECT 143.995 152.785 144.165 152.955 ;
        RECT 144.455 152.785 144.625 152.955 ;
        RECT 144.915 152.785 145.085 152.955 ;
        RECT 145.375 152.785 145.545 152.955 ;
        RECT 145.835 152.785 146.005 152.955 ;
        RECT 146.295 152.785 146.465 152.955 ;
        RECT 146.755 152.785 146.925 152.955 ;
        RECT 147.215 152.785 147.385 152.955 ;
        RECT 147.675 152.785 147.845 152.955 ;
        RECT 148.135 152.785 148.305 152.955 ;
        RECT 148.595 152.785 148.765 152.955 ;
        RECT 149.055 152.785 149.225 152.955 ;
        RECT 149.515 152.785 149.685 152.955 ;
        RECT 149.975 152.785 150.145 152.955 ;
        RECT 150.435 152.785 150.605 152.955 ;
        RECT 150.895 152.785 151.065 152.955 ;
        RECT 151.355 152.785 151.525 152.955 ;
        RECT 151.815 152.785 151.985 152.955 ;
        RECT 152.275 152.785 152.445 152.955 ;
        RECT 152.735 152.785 152.905 152.955 ;
        RECT 153.195 152.785 153.365 152.955 ;
        RECT 153.655 152.785 153.825 152.955 ;
        RECT 154.115 152.785 154.285 152.955 ;
        RECT 154.575 152.785 154.745 152.955 ;
        RECT 155.035 152.785 155.205 152.955 ;
        RECT 155.495 152.785 155.665 152.955 ;
        RECT 155.955 152.785 156.125 152.955 ;
        RECT 81.895 151.255 82.065 151.425 ;
        RECT 80.975 150.575 81.145 150.745 ;
        RECT 97.075 151.935 97.245 152.105 ;
        RECT 98.455 151.595 98.625 151.765 ;
        RECT 97.995 151.255 98.165 151.425 ;
        RECT 99.605 150.575 99.775 150.745 ;
        RECT 103.975 151.255 104.145 151.425 ;
        RECT 105.355 151.595 105.525 151.765 ;
        RECT 107.195 151.935 107.365 152.105 ;
        RECT 104.895 151.255 105.065 151.425 ;
        RECT 105.815 151.255 105.985 151.425 ;
        RECT 103.055 150.915 103.225 151.085 ;
        RECT 106.735 151.255 106.905 151.425 ;
        RECT 109.955 152.275 110.125 152.445 ;
        RECT 108.115 151.255 108.285 151.425 ;
        RECT 111.795 152.275 111.965 152.445 ;
        RECT 113.635 152.275 113.805 152.445 ;
        RECT 112.255 151.595 112.425 151.765 ;
        RECT 110.875 151.255 111.045 151.425 ;
        RECT 112.715 151.255 112.885 151.425 ;
        RECT 123.295 152.275 123.465 152.445 ;
        RECT 125.135 152.275 125.305 152.445 ;
        RECT 125.595 151.595 125.765 151.765 ;
        RECT 124.215 151.255 124.385 151.425 ;
        RECT 127.435 151.255 127.605 151.425 ;
        RECT 128.355 150.575 128.525 150.745 ;
        RECT 132.035 151.255 132.205 151.425 ;
        RECT 135.715 151.255 135.885 151.425 ;
        RECT 131.115 150.575 131.285 150.745 ;
        RECT 137.095 151.595 137.265 151.765 ;
        RECT 136.635 151.255 136.805 151.425 ;
        RECT 140.315 152.275 140.485 152.445 ;
        RECT 139.395 151.595 139.565 151.765 ;
        RECT 138.475 151.255 138.645 151.425 ;
        RECT 139.855 151.255 140.025 151.425 ;
        RECT 141.235 151.255 141.405 151.425 ;
        RECT 143.535 151.595 143.705 151.765 ;
        RECT 144.915 151.255 145.085 151.425 ;
        RECT 149.975 151.935 150.145 152.105 ;
        RECT 148.135 151.255 148.305 151.425 ;
        RECT 149.055 151.255 149.225 151.425 ;
        RECT 149.515 151.255 149.685 151.425 ;
        RECT 151.355 151.595 151.525 151.765 ;
        RECT 150.435 151.255 150.605 151.425 ;
        RECT 150.895 151.255 151.065 151.425 ;
        RECT 142.155 150.575 142.325 150.745 ;
        RECT 148.595 150.575 148.765 150.745 ;
        RECT 153.195 151.255 153.365 151.425 ;
        RECT 152.275 150.575 152.445 150.745 ;
        RECT 70.855 150.065 71.025 150.235 ;
        RECT 71.315 150.065 71.485 150.235 ;
        RECT 71.775 150.065 71.945 150.235 ;
        RECT 72.235 150.065 72.405 150.235 ;
        RECT 72.695 150.065 72.865 150.235 ;
        RECT 73.155 150.065 73.325 150.235 ;
        RECT 73.615 150.065 73.785 150.235 ;
        RECT 74.075 150.065 74.245 150.235 ;
        RECT 74.535 150.065 74.705 150.235 ;
        RECT 74.995 150.065 75.165 150.235 ;
        RECT 75.455 150.065 75.625 150.235 ;
        RECT 75.915 150.065 76.085 150.235 ;
        RECT 76.375 150.065 76.545 150.235 ;
        RECT 76.835 150.065 77.005 150.235 ;
        RECT 77.295 150.065 77.465 150.235 ;
        RECT 77.755 150.065 77.925 150.235 ;
        RECT 78.215 150.065 78.385 150.235 ;
        RECT 78.675 150.065 78.845 150.235 ;
        RECT 79.135 150.065 79.305 150.235 ;
        RECT 79.595 150.065 79.765 150.235 ;
        RECT 80.055 150.065 80.225 150.235 ;
        RECT 80.515 150.065 80.685 150.235 ;
        RECT 80.975 150.065 81.145 150.235 ;
        RECT 81.435 150.065 81.605 150.235 ;
        RECT 81.895 150.065 82.065 150.235 ;
        RECT 82.355 150.065 82.525 150.235 ;
        RECT 82.815 150.065 82.985 150.235 ;
        RECT 83.275 150.065 83.445 150.235 ;
        RECT 83.735 150.065 83.905 150.235 ;
        RECT 84.195 150.065 84.365 150.235 ;
        RECT 84.655 150.065 84.825 150.235 ;
        RECT 85.115 150.065 85.285 150.235 ;
        RECT 85.575 150.065 85.745 150.235 ;
        RECT 86.035 150.065 86.205 150.235 ;
        RECT 86.495 150.065 86.665 150.235 ;
        RECT 86.955 150.065 87.125 150.235 ;
        RECT 87.415 150.065 87.585 150.235 ;
        RECT 87.875 150.065 88.045 150.235 ;
        RECT 88.335 150.065 88.505 150.235 ;
        RECT 88.795 150.065 88.965 150.235 ;
        RECT 89.255 150.065 89.425 150.235 ;
        RECT 89.715 150.065 89.885 150.235 ;
        RECT 90.175 150.065 90.345 150.235 ;
        RECT 90.635 150.065 90.805 150.235 ;
        RECT 91.095 150.065 91.265 150.235 ;
        RECT 91.555 150.065 91.725 150.235 ;
        RECT 92.015 150.065 92.185 150.235 ;
        RECT 92.475 150.065 92.645 150.235 ;
        RECT 92.935 150.065 93.105 150.235 ;
        RECT 93.395 150.065 93.565 150.235 ;
        RECT 93.855 150.065 94.025 150.235 ;
        RECT 94.315 150.065 94.485 150.235 ;
        RECT 94.775 150.065 94.945 150.235 ;
        RECT 95.235 150.065 95.405 150.235 ;
        RECT 95.695 150.065 95.865 150.235 ;
        RECT 96.155 150.065 96.325 150.235 ;
        RECT 96.615 150.065 96.785 150.235 ;
        RECT 97.075 150.065 97.245 150.235 ;
        RECT 97.535 150.065 97.705 150.235 ;
        RECT 97.995 150.065 98.165 150.235 ;
        RECT 98.455 150.065 98.625 150.235 ;
        RECT 98.915 150.065 99.085 150.235 ;
        RECT 99.375 150.065 99.545 150.235 ;
        RECT 99.835 150.065 100.005 150.235 ;
        RECT 100.295 150.065 100.465 150.235 ;
        RECT 100.755 150.065 100.925 150.235 ;
        RECT 101.215 150.065 101.385 150.235 ;
        RECT 101.675 150.065 101.845 150.235 ;
        RECT 102.135 150.065 102.305 150.235 ;
        RECT 102.595 150.065 102.765 150.235 ;
        RECT 103.055 150.065 103.225 150.235 ;
        RECT 103.515 150.065 103.685 150.235 ;
        RECT 103.975 150.065 104.145 150.235 ;
        RECT 104.435 150.065 104.605 150.235 ;
        RECT 104.895 150.065 105.065 150.235 ;
        RECT 105.355 150.065 105.525 150.235 ;
        RECT 105.815 150.065 105.985 150.235 ;
        RECT 106.275 150.065 106.445 150.235 ;
        RECT 106.735 150.065 106.905 150.235 ;
        RECT 107.195 150.065 107.365 150.235 ;
        RECT 107.655 150.065 107.825 150.235 ;
        RECT 108.115 150.065 108.285 150.235 ;
        RECT 108.575 150.065 108.745 150.235 ;
        RECT 109.035 150.065 109.205 150.235 ;
        RECT 109.495 150.065 109.665 150.235 ;
        RECT 109.955 150.065 110.125 150.235 ;
        RECT 110.415 150.065 110.585 150.235 ;
        RECT 110.875 150.065 111.045 150.235 ;
        RECT 111.335 150.065 111.505 150.235 ;
        RECT 111.795 150.065 111.965 150.235 ;
        RECT 112.255 150.065 112.425 150.235 ;
        RECT 112.715 150.065 112.885 150.235 ;
        RECT 113.175 150.065 113.345 150.235 ;
        RECT 113.635 150.065 113.805 150.235 ;
        RECT 114.095 150.065 114.265 150.235 ;
        RECT 114.555 150.065 114.725 150.235 ;
        RECT 115.015 150.065 115.185 150.235 ;
        RECT 115.475 150.065 115.645 150.235 ;
        RECT 115.935 150.065 116.105 150.235 ;
        RECT 116.395 150.065 116.565 150.235 ;
        RECT 116.855 150.065 117.025 150.235 ;
        RECT 117.315 150.065 117.485 150.235 ;
        RECT 117.775 150.065 117.945 150.235 ;
        RECT 118.235 150.065 118.405 150.235 ;
        RECT 118.695 150.065 118.865 150.235 ;
        RECT 119.155 150.065 119.325 150.235 ;
        RECT 119.615 150.065 119.785 150.235 ;
        RECT 120.075 150.065 120.245 150.235 ;
        RECT 120.535 150.065 120.705 150.235 ;
        RECT 120.995 150.065 121.165 150.235 ;
        RECT 121.455 150.065 121.625 150.235 ;
        RECT 121.915 150.065 122.085 150.235 ;
        RECT 122.375 150.065 122.545 150.235 ;
        RECT 122.835 150.065 123.005 150.235 ;
        RECT 123.295 150.065 123.465 150.235 ;
        RECT 123.755 150.065 123.925 150.235 ;
        RECT 124.215 150.065 124.385 150.235 ;
        RECT 124.675 150.065 124.845 150.235 ;
        RECT 125.135 150.065 125.305 150.235 ;
        RECT 125.595 150.065 125.765 150.235 ;
        RECT 126.055 150.065 126.225 150.235 ;
        RECT 126.515 150.065 126.685 150.235 ;
        RECT 126.975 150.065 127.145 150.235 ;
        RECT 127.435 150.065 127.605 150.235 ;
        RECT 127.895 150.065 128.065 150.235 ;
        RECT 128.355 150.065 128.525 150.235 ;
        RECT 128.815 150.065 128.985 150.235 ;
        RECT 129.275 150.065 129.445 150.235 ;
        RECT 129.735 150.065 129.905 150.235 ;
        RECT 130.195 150.065 130.365 150.235 ;
        RECT 130.655 150.065 130.825 150.235 ;
        RECT 131.115 150.065 131.285 150.235 ;
        RECT 131.575 150.065 131.745 150.235 ;
        RECT 132.035 150.065 132.205 150.235 ;
        RECT 132.495 150.065 132.665 150.235 ;
        RECT 132.955 150.065 133.125 150.235 ;
        RECT 133.415 150.065 133.585 150.235 ;
        RECT 133.875 150.065 134.045 150.235 ;
        RECT 134.335 150.065 134.505 150.235 ;
        RECT 134.795 150.065 134.965 150.235 ;
        RECT 135.255 150.065 135.425 150.235 ;
        RECT 135.715 150.065 135.885 150.235 ;
        RECT 136.175 150.065 136.345 150.235 ;
        RECT 136.635 150.065 136.805 150.235 ;
        RECT 137.095 150.065 137.265 150.235 ;
        RECT 137.555 150.065 137.725 150.235 ;
        RECT 138.015 150.065 138.185 150.235 ;
        RECT 138.475 150.065 138.645 150.235 ;
        RECT 138.935 150.065 139.105 150.235 ;
        RECT 139.395 150.065 139.565 150.235 ;
        RECT 139.855 150.065 140.025 150.235 ;
        RECT 140.315 150.065 140.485 150.235 ;
        RECT 140.775 150.065 140.945 150.235 ;
        RECT 141.235 150.065 141.405 150.235 ;
        RECT 141.695 150.065 141.865 150.235 ;
        RECT 142.155 150.065 142.325 150.235 ;
        RECT 142.615 150.065 142.785 150.235 ;
        RECT 143.075 150.065 143.245 150.235 ;
        RECT 143.535 150.065 143.705 150.235 ;
        RECT 143.995 150.065 144.165 150.235 ;
        RECT 144.455 150.065 144.625 150.235 ;
        RECT 144.915 150.065 145.085 150.235 ;
        RECT 145.375 150.065 145.545 150.235 ;
        RECT 145.835 150.065 146.005 150.235 ;
        RECT 146.295 150.065 146.465 150.235 ;
        RECT 146.755 150.065 146.925 150.235 ;
        RECT 147.215 150.065 147.385 150.235 ;
        RECT 147.675 150.065 147.845 150.235 ;
        RECT 148.135 150.065 148.305 150.235 ;
        RECT 148.595 150.065 148.765 150.235 ;
        RECT 149.055 150.065 149.225 150.235 ;
        RECT 149.515 150.065 149.685 150.235 ;
        RECT 149.975 150.065 150.145 150.235 ;
        RECT 150.435 150.065 150.605 150.235 ;
        RECT 150.895 150.065 151.065 150.235 ;
        RECT 151.355 150.065 151.525 150.235 ;
        RECT 151.815 150.065 151.985 150.235 ;
        RECT 152.275 150.065 152.445 150.235 ;
        RECT 152.735 150.065 152.905 150.235 ;
        RECT 153.195 150.065 153.365 150.235 ;
        RECT 153.655 150.065 153.825 150.235 ;
        RECT 154.115 150.065 154.285 150.235 ;
        RECT 154.575 150.065 154.745 150.235 ;
        RECT 155.035 150.065 155.205 150.235 ;
        RECT 155.495 150.065 155.665 150.235 ;
        RECT 155.955 150.065 156.125 150.235 ;
        RECT 72.235 148.535 72.405 148.705 ;
        RECT 72.720 148.195 72.890 148.365 ;
        RECT 73.115 148.535 73.285 148.705 ;
        RECT 73.570 148.875 73.740 149.045 ;
        RECT 74.305 148.535 74.475 148.705 ;
        RECT 74.820 148.195 74.990 148.365 ;
        RECT 76.390 148.195 76.560 148.365 ;
        RECT 76.825 148.535 76.995 148.705 ;
        RECT 80.975 149.555 81.145 149.725 ;
        RECT 82.355 149.555 82.525 149.725 ;
        RECT 80.515 148.875 80.685 149.045 ;
        RECT 81.435 148.875 81.605 149.045 ;
        RECT 81.895 148.875 82.065 149.045 ;
        RECT 83.275 148.875 83.445 149.045 ;
        RECT 79.135 147.855 79.305 148.025 ;
        RECT 83.275 148.195 83.445 148.365 ;
        RECT 89.485 149.555 89.655 149.725 ;
        RECT 85.115 148.875 85.285 149.045 ;
        RECT 86.035 148.875 86.205 149.045 ;
        RECT 86.495 148.535 86.665 148.705 ;
        RECT 87.875 148.875 88.045 149.045 ;
        RECT 84.195 147.855 84.365 148.025 ;
        RECT 87.415 148.535 87.585 148.705 ;
        RECT 88.335 148.535 88.505 148.705 ;
        RECT 97.995 148.875 98.165 149.045 ;
        RECT 99.375 148.875 99.545 149.045 ;
        RECT 99.835 148.875 100.005 149.045 ;
        RECT 97.075 147.855 97.245 148.025 ;
        RECT 98.915 148.535 99.085 148.705 ;
        RECT 100.755 148.875 100.925 149.045 ;
        RECT 103.515 148.875 103.685 149.045 ;
        RECT 102.595 147.855 102.765 148.025 ;
        RECT 104.435 147.855 104.605 148.025 ;
        RECT 115.015 148.875 115.185 149.045 ;
        RECT 113.635 148.535 113.805 148.705 ;
        RECT 114.095 147.855 114.265 148.025 ;
        RECT 115.935 148.195 116.105 148.365 ;
        RECT 117.315 149.215 117.485 149.385 ;
        RECT 118.235 148.875 118.405 149.045 ;
        RECT 116.395 147.855 116.565 148.025 ;
        RECT 119.615 148.875 119.785 149.045 ;
        RECT 118.695 147.855 118.865 148.025 ;
        RECT 127.895 148.875 128.065 149.045 ;
        RECT 128.815 148.875 128.985 149.045 ;
        RECT 129.275 148.875 129.445 149.045 ;
        RECT 129.735 148.875 129.905 149.045 ;
        RECT 131.115 147.855 131.285 148.025 ;
        RECT 131.575 148.535 131.745 148.705 ;
        RECT 132.495 148.875 132.665 149.045 ;
        RECT 134.335 148.875 134.505 149.045 ;
        RECT 133.875 147.855 134.045 148.025 ;
        RECT 135.715 148.875 135.885 149.045 ;
        RECT 137.555 148.875 137.725 149.045 ;
        RECT 134.795 147.855 134.965 148.025 ;
        RECT 137.095 147.855 137.265 148.025 ;
        RECT 142.155 148.875 142.325 149.045 ;
        RECT 141.235 148.195 141.405 148.365 ;
        RECT 143.535 148.875 143.705 149.045 ;
        RECT 142.615 147.855 142.785 148.025 ;
        RECT 144.915 148.875 145.085 149.045 ;
        RECT 145.835 148.875 146.005 149.045 ;
        RECT 143.995 147.855 144.165 148.025 ;
        RECT 146.755 148.875 146.925 149.045 ;
        RECT 146.295 148.535 146.465 148.705 ;
        RECT 147.675 148.875 147.845 149.045 ;
        RECT 149.515 148.875 149.685 149.045 ;
        RECT 150.435 148.875 150.605 149.045 ;
        RECT 151.355 148.875 151.525 149.045 ;
        RECT 152.735 148.875 152.905 149.045 ;
        RECT 149.055 148.195 149.225 148.365 ;
        RECT 153.655 148.875 153.825 149.045 ;
        RECT 151.815 148.195 151.985 148.365 ;
        RECT 152.735 147.855 152.905 148.025 ;
        RECT 70.855 147.345 71.025 147.515 ;
        RECT 71.315 147.345 71.485 147.515 ;
        RECT 71.775 147.345 71.945 147.515 ;
        RECT 72.235 147.345 72.405 147.515 ;
        RECT 72.695 147.345 72.865 147.515 ;
        RECT 73.155 147.345 73.325 147.515 ;
        RECT 73.615 147.345 73.785 147.515 ;
        RECT 74.075 147.345 74.245 147.515 ;
        RECT 74.535 147.345 74.705 147.515 ;
        RECT 74.995 147.345 75.165 147.515 ;
        RECT 75.455 147.345 75.625 147.515 ;
        RECT 75.915 147.345 76.085 147.515 ;
        RECT 76.375 147.345 76.545 147.515 ;
        RECT 76.835 147.345 77.005 147.515 ;
        RECT 77.295 147.345 77.465 147.515 ;
        RECT 77.755 147.345 77.925 147.515 ;
        RECT 78.215 147.345 78.385 147.515 ;
        RECT 78.675 147.345 78.845 147.515 ;
        RECT 79.135 147.345 79.305 147.515 ;
        RECT 79.595 147.345 79.765 147.515 ;
        RECT 80.055 147.345 80.225 147.515 ;
        RECT 80.515 147.345 80.685 147.515 ;
        RECT 80.975 147.345 81.145 147.515 ;
        RECT 81.435 147.345 81.605 147.515 ;
        RECT 81.895 147.345 82.065 147.515 ;
        RECT 82.355 147.345 82.525 147.515 ;
        RECT 82.815 147.345 82.985 147.515 ;
        RECT 83.275 147.345 83.445 147.515 ;
        RECT 83.735 147.345 83.905 147.515 ;
        RECT 84.195 147.345 84.365 147.515 ;
        RECT 84.655 147.345 84.825 147.515 ;
        RECT 85.115 147.345 85.285 147.515 ;
        RECT 85.575 147.345 85.745 147.515 ;
        RECT 86.035 147.345 86.205 147.515 ;
        RECT 86.495 147.345 86.665 147.515 ;
        RECT 86.955 147.345 87.125 147.515 ;
        RECT 87.415 147.345 87.585 147.515 ;
        RECT 87.875 147.345 88.045 147.515 ;
        RECT 88.335 147.345 88.505 147.515 ;
        RECT 88.795 147.345 88.965 147.515 ;
        RECT 89.255 147.345 89.425 147.515 ;
        RECT 89.715 147.345 89.885 147.515 ;
        RECT 90.175 147.345 90.345 147.515 ;
        RECT 90.635 147.345 90.805 147.515 ;
        RECT 91.095 147.345 91.265 147.515 ;
        RECT 91.555 147.345 91.725 147.515 ;
        RECT 92.015 147.345 92.185 147.515 ;
        RECT 92.475 147.345 92.645 147.515 ;
        RECT 92.935 147.345 93.105 147.515 ;
        RECT 93.395 147.345 93.565 147.515 ;
        RECT 93.855 147.345 94.025 147.515 ;
        RECT 94.315 147.345 94.485 147.515 ;
        RECT 94.775 147.345 94.945 147.515 ;
        RECT 95.235 147.345 95.405 147.515 ;
        RECT 95.695 147.345 95.865 147.515 ;
        RECT 96.155 147.345 96.325 147.515 ;
        RECT 96.615 147.345 96.785 147.515 ;
        RECT 97.075 147.345 97.245 147.515 ;
        RECT 97.535 147.345 97.705 147.515 ;
        RECT 97.995 147.345 98.165 147.515 ;
        RECT 98.455 147.345 98.625 147.515 ;
        RECT 98.915 147.345 99.085 147.515 ;
        RECT 99.375 147.345 99.545 147.515 ;
        RECT 99.835 147.345 100.005 147.515 ;
        RECT 100.295 147.345 100.465 147.515 ;
        RECT 100.755 147.345 100.925 147.515 ;
        RECT 101.215 147.345 101.385 147.515 ;
        RECT 101.675 147.345 101.845 147.515 ;
        RECT 102.135 147.345 102.305 147.515 ;
        RECT 102.595 147.345 102.765 147.515 ;
        RECT 103.055 147.345 103.225 147.515 ;
        RECT 103.515 147.345 103.685 147.515 ;
        RECT 103.975 147.345 104.145 147.515 ;
        RECT 104.435 147.345 104.605 147.515 ;
        RECT 104.895 147.345 105.065 147.515 ;
        RECT 105.355 147.345 105.525 147.515 ;
        RECT 105.815 147.345 105.985 147.515 ;
        RECT 106.275 147.345 106.445 147.515 ;
        RECT 106.735 147.345 106.905 147.515 ;
        RECT 107.195 147.345 107.365 147.515 ;
        RECT 107.655 147.345 107.825 147.515 ;
        RECT 108.115 147.345 108.285 147.515 ;
        RECT 108.575 147.345 108.745 147.515 ;
        RECT 109.035 147.345 109.205 147.515 ;
        RECT 109.495 147.345 109.665 147.515 ;
        RECT 109.955 147.345 110.125 147.515 ;
        RECT 110.415 147.345 110.585 147.515 ;
        RECT 110.875 147.345 111.045 147.515 ;
        RECT 111.335 147.345 111.505 147.515 ;
        RECT 111.795 147.345 111.965 147.515 ;
        RECT 112.255 147.345 112.425 147.515 ;
        RECT 112.715 147.345 112.885 147.515 ;
        RECT 113.175 147.345 113.345 147.515 ;
        RECT 113.635 147.345 113.805 147.515 ;
        RECT 114.095 147.345 114.265 147.515 ;
        RECT 114.555 147.345 114.725 147.515 ;
        RECT 115.015 147.345 115.185 147.515 ;
        RECT 115.475 147.345 115.645 147.515 ;
        RECT 115.935 147.345 116.105 147.515 ;
        RECT 116.395 147.345 116.565 147.515 ;
        RECT 116.855 147.345 117.025 147.515 ;
        RECT 117.315 147.345 117.485 147.515 ;
        RECT 117.775 147.345 117.945 147.515 ;
        RECT 118.235 147.345 118.405 147.515 ;
        RECT 118.695 147.345 118.865 147.515 ;
        RECT 119.155 147.345 119.325 147.515 ;
        RECT 119.615 147.345 119.785 147.515 ;
        RECT 120.075 147.345 120.245 147.515 ;
        RECT 120.535 147.345 120.705 147.515 ;
        RECT 120.995 147.345 121.165 147.515 ;
        RECT 121.455 147.345 121.625 147.515 ;
        RECT 121.915 147.345 122.085 147.515 ;
        RECT 122.375 147.345 122.545 147.515 ;
        RECT 122.835 147.345 123.005 147.515 ;
        RECT 123.295 147.345 123.465 147.515 ;
        RECT 123.755 147.345 123.925 147.515 ;
        RECT 124.215 147.345 124.385 147.515 ;
        RECT 124.675 147.345 124.845 147.515 ;
        RECT 125.135 147.345 125.305 147.515 ;
        RECT 125.595 147.345 125.765 147.515 ;
        RECT 126.055 147.345 126.225 147.515 ;
        RECT 126.515 147.345 126.685 147.515 ;
        RECT 126.975 147.345 127.145 147.515 ;
        RECT 127.435 147.345 127.605 147.515 ;
        RECT 127.895 147.345 128.065 147.515 ;
        RECT 128.355 147.345 128.525 147.515 ;
        RECT 128.815 147.345 128.985 147.515 ;
        RECT 129.275 147.345 129.445 147.515 ;
        RECT 129.735 147.345 129.905 147.515 ;
        RECT 130.195 147.345 130.365 147.515 ;
        RECT 130.655 147.345 130.825 147.515 ;
        RECT 131.115 147.345 131.285 147.515 ;
        RECT 131.575 147.345 131.745 147.515 ;
        RECT 132.035 147.345 132.205 147.515 ;
        RECT 132.495 147.345 132.665 147.515 ;
        RECT 132.955 147.345 133.125 147.515 ;
        RECT 133.415 147.345 133.585 147.515 ;
        RECT 133.875 147.345 134.045 147.515 ;
        RECT 134.335 147.345 134.505 147.515 ;
        RECT 134.795 147.345 134.965 147.515 ;
        RECT 135.255 147.345 135.425 147.515 ;
        RECT 135.715 147.345 135.885 147.515 ;
        RECT 136.175 147.345 136.345 147.515 ;
        RECT 136.635 147.345 136.805 147.515 ;
        RECT 137.095 147.345 137.265 147.515 ;
        RECT 137.555 147.345 137.725 147.515 ;
        RECT 138.015 147.345 138.185 147.515 ;
        RECT 138.475 147.345 138.645 147.515 ;
        RECT 138.935 147.345 139.105 147.515 ;
        RECT 139.395 147.345 139.565 147.515 ;
        RECT 139.855 147.345 140.025 147.515 ;
        RECT 140.315 147.345 140.485 147.515 ;
        RECT 140.775 147.345 140.945 147.515 ;
        RECT 141.235 147.345 141.405 147.515 ;
        RECT 141.695 147.345 141.865 147.515 ;
        RECT 142.155 147.345 142.325 147.515 ;
        RECT 142.615 147.345 142.785 147.515 ;
        RECT 143.075 147.345 143.245 147.515 ;
        RECT 143.535 147.345 143.705 147.515 ;
        RECT 143.995 147.345 144.165 147.515 ;
        RECT 144.455 147.345 144.625 147.515 ;
        RECT 144.915 147.345 145.085 147.515 ;
        RECT 145.375 147.345 145.545 147.515 ;
        RECT 145.835 147.345 146.005 147.515 ;
        RECT 146.295 147.345 146.465 147.515 ;
        RECT 146.755 147.345 146.925 147.515 ;
        RECT 147.215 147.345 147.385 147.515 ;
        RECT 147.675 147.345 147.845 147.515 ;
        RECT 148.135 147.345 148.305 147.515 ;
        RECT 148.595 147.345 148.765 147.515 ;
        RECT 149.055 147.345 149.225 147.515 ;
        RECT 149.515 147.345 149.685 147.515 ;
        RECT 149.975 147.345 150.145 147.515 ;
        RECT 150.435 147.345 150.605 147.515 ;
        RECT 150.895 147.345 151.065 147.515 ;
        RECT 151.355 147.345 151.525 147.515 ;
        RECT 151.815 147.345 151.985 147.515 ;
        RECT 152.275 147.345 152.445 147.515 ;
        RECT 152.735 147.345 152.905 147.515 ;
        RECT 153.195 147.345 153.365 147.515 ;
        RECT 153.655 147.345 153.825 147.515 ;
        RECT 154.115 147.345 154.285 147.515 ;
        RECT 154.575 147.345 154.745 147.515 ;
        RECT 155.035 147.345 155.205 147.515 ;
        RECT 155.495 147.345 155.665 147.515 ;
        RECT 155.955 147.345 156.125 147.515 ;
        RECT 72.695 146.835 72.865 147.005 ;
        RECT 72.235 145.815 72.405 145.985 ;
        RECT 73.155 145.815 73.325 145.985 ;
        RECT 74.535 145.815 74.705 145.985 ;
        RECT 74.995 145.815 75.165 145.985 ;
        RECT 74.075 145.135 74.245 145.305 ;
        RECT 75.915 145.475 76.085 145.645 ;
        RECT 76.835 145.475 77.005 145.645 ;
        RECT 78.215 146.835 78.385 147.005 ;
        RECT 80.055 146.495 80.225 146.665 ;
        RECT 82.355 146.835 82.525 147.005 ;
        RECT 77.295 145.135 77.465 145.305 ;
        RECT 79.595 145.815 79.765 145.985 ;
        RECT 79.135 145.475 79.305 145.645 ;
        RECT 80.975 145.815 81.145 145.985 ;
        RECT 80.515 145.475 80.685 145.645 ;
        RECT 85.115 146.835 85.285 147.005 ;
        RECT 81.435 145.135 81.605 145.305 ;
        RECT 83.275 145.475 83.445 145.645 ;
        RECT 86.035 145.815 86.205 145.985 ;
        RECT 86.495 145.815 86.665 145.985 ;
        RECT 86.955 146.155 87.125 146.325 ;
        RECT 87.415 145.815 87.585 145.985 ;
        RECT 89.255 146.495 89.425 146.665 ;
        RECT 88.335 145.815 88.505 145.985 ;
        RECT 92.475 145.815 92.645 145.985 ;
        RECT 93.855 146.155 94.025 146.325 ;
        RECT 96.155 146.835 96.325 147.005 ;
        RECT 93.395 145.815 93.565 145.985 ;
        RECT 95.235 145.815 95.405 145.985 ;
        RECT 98.915 146.155 99.085 146.325 ;
        RECT 100.295 146.155 100.465 146.325 ;
        RECT 105.815 146.835 105.985 147.005 ;
        RECT 104.435 145.815 104.605 145.985 ;
        RECT 106.275 145.815 106.445 145.985 ;
        RECT 103.515 145.135 103.685 145.305 ;
        RECT 109.955 145.815 110.125 145.985 ;
        RECT 112.255 146.495 112.425 146.665 ;
        RECT 110.875 145.815 111.045 145.985 ;
        RECT 112.715 145.815 112.885 145.985 ;
        RECT 113.175 145.815 113.345 145.985 ;
        RECT 115.015 146.495 115.185 146.665 ;
        RECT 114.555 145.815 114.725 145.985 ;
        RECT 115.935 145.815 116.105 145.985 ;
        RECT 116.395 145.815 116.565 145.985 ;
        RECT 114.095 145.135 114.265 145.305 ;
        RECT 117.315 145.135 117.485 145.305 ;
        RECT 119.615 145.815 119.785 145.985 ;
        RECT 120.995 146.155 121.165 146.325 ;
        RECT 120.535 145.815 120.705 145.985 ;
        RECT 121.455 145.815 121.625 145.985 ;
        RECT 118.695 145.135 118.865 145.305 ;
        RECT 122.375 145.815 122.545 145.985 ;
        RECT 122.835 145.815 123.005 145.985 ;
        RECT 124.675 146.495 124.845 146.665 ;
        RECT 125.135 146.155 125.305 146.325 ;
        RECT 123.755 145.815 123.925 145.985 ;
        RECT 127.435 145.815 127.605 145.985 ;
        RECT 128.815 146.155 128.985 146.325 ;
        RECT 128.355 145.815 128.525 145.985 ;
        RECT 130.195 145.815 130.365 145.985 ;
        RECT 131.115 145.475 131.285 145.645 ;
        RECT 132.495 145.815 132.665 145.985 ;
        RECT 136.175 146.835 136.345 147.005 ;
        RECT 135.715 145.815 135.885 145.985 ;
        RECT 137.095 145.815 137.265 145.985 ;
        RECT 137.555 145.815 137.725 145.985 ;
        RECT 131.575 145.135 131.745 145.305 ;
        RECT 138.475 146.155 138.645 146.325 ;
        RECT 70.855 144.625 71.025 144.795 ;
        RECT 71.315 144.625 71.485 144.795 ;
        RECT 71.775 144.625 71.945 144.795 ;
        RECT 72.235 144.625 72.405 144.795 ;
        RECT 72.695 144.625 72.865 144.795 ;
        RECT 73.155 144.625 73.325 144.795 ;
        RECT 73.615 144.625 73.785 144.795 ;
        RECT 74.075 144.625 74.245 144.795 ;
        RECT 74.535 144.625 74.705 144.795 ;
        RECT 74.995 144.625 75.165 144.795 ;
        RECT 75.455 144.625 75.625 144.795 ;
        RECT 75.915 144.625 76.085 144.795 ;
        RECT 76.375 144.625 76.545 144.795 ;
        RECT 76.835 144.625 77.005 144.795 ;
        RECT 77.295 144.625 77.465 144.795 ;
        RECT 77.755 144.625 77.925 144.795 ;
        RECT 78.215 144.625 78.385 144.795 ;
        RECT 78.675 144.625 78.845 144.795 ;
        RECT 79.135 144.625 79.305 144.795 ;
        RECT 79.595 144.625 79.765 144.795 ;
        RECT 80.055 144.625 80.225 144.795 ;
        RECT 80.515 144.625 80.685 144.795 ;
        RECT 80.975 144.625 81.145 144.795 ;
        RECT 81.435 144.625 81.605 144.795 ;
        RECT 81.895 144.625 82.065 144.795 ;
        RECT 82.355 144.625 82.525 144.795 ;
        RECT 82.815 144.625 82.985 144.795 ;
        RECT 83.275 144.625 83.445 144.795 ;
        RECT 83.735 144.625 83.905 144.795 ;
        RECT 84.195 144.625 84.365 144.795 ;
        RECT 84.655 144.625 84.825 144.795 ;
        RECT 85.115 144.625 85.285 144.795 ;
        RECT 85.575 144.625 85.745 144.795 ;
        RECT 86.035 144.625 86.205 144.795 ;
        RECT 86.495 144.625 86.665 144.795 ;
        RECT 86.955 144.625 87.125 144.795 ;
        RECT 87.415 144.625 87.585 144.795 ;
        RECT 87.875 144.625 88.045 144.795 ;
        RECT 88.335 144.625 88.505 144.795 ;
        RECT 88.795 144.625 88.965 144.795 ;
        RECT 89.255 144.625 89.425 144.795 ;
        RECT 89.715 144.625 89.885 144.795 ;
        RECT 90.175 144.625 90.345 144.795 ;
        RECT 90.635 144.625 90.805 144.795 ;
        RECT 91.095 144.625 91.265 144.795 ;
        RECT 91.555 144.625 91.725 144.795 ;
        RECT 92.015 144.625 92.185 144.795 ;
        RECT 92.475 144.625 92.645 144.795 ;
        RECT 92.935 144.625 93.105 144.795 ;
        RECT 93.395 144.625 93.565 144.795 ;
        RECT 93.855 144.625 94.025 144.795 ;
        RECT 94.315 144.625 94.485 144.795 ;
        RECT 94.775 144.625 94.945 144.795 ;
        RECT 95.235 144.625 95.405 144.795 ;
        RECT 95.695 144.625 95.865 144.795 ;
        RECT 96.155 144.625 96.325 144.795 ;
        RECT 96.615 144.625 96.785 144.795 ;
        RECT 97.075 144.625 97.245 144.795 ;
        RECT 97.535 144.625 97.705 144.795 ;
        RECT 97.995 144.625 98.165 144.795 ;
        RECT 98.455 144.625 98.625 144.795 ;
        RECT 98.915 144.625 99.085 144.795 ;
        RECT 99.375 144.625 99.545 144.795 ;
        RECT 99.835 144.625 100.005 144.795 ;
        RECT 100.295 144.625 100.465 144.795 ;
        RECT 100.755 144.625 100.925 144.795 ;
        RECT 101.215 144.625 101.385 144.795 ;
        RECT 101.675 144.625 101.845 144.795 ;
        RECT 102.135 144.625 102.305 144.795 ;
        RECT 102.595 144.625 102.765 144.795 ;
        RECT 103.055 144.625 103.225 144.795 ;
        RECT 103.515 144.625 103.685 144.795 ;
        RECT 103.975 144.625 104.145 144.795 ;
        RECT 104.435 144.625 104.605 144.795 ;
        RECT 104.895 144.625 105.065 144.795 ;
        RECT 105.355 144.625 105.525 144.795 ;
        RECT 105.815 144.625 105.985 144.795 ;
        RECT 106.275 144.625 106.445 144.795 ;
        RECT 106.735 144.625 106.905 144.795 ;
        RECT 107.195 144.625 107.365 144.795 ;
        RECT 107.655 144.625 107.825 144.795 ;
        RECT 108.115 144.625 108.285 144.795 ;
        RECT 108.575 144.625 108.745 144.795 ;
        RECT 109.035 144.625 109.205 144.795 ;
        RECT 109.495 144.625 109.665 144.795 ;
        RECT 109.955 144.625 110.125 144.795 ;
        RECT 110.415 144.625 110.585 144.795 ;
        RECT 110.875 144.625 111.045 144.795 ;
        RECT 111.335 144.625 111.505 144.795 ;
        RECT 111.795 144.625 111.965 144.795 ;
        RECT 112.255 144.625 112.425 144.795 ;
        RECT 112.715 144.625 112.885 144.795 ;
        RECT 113.175 144.625 113.345 144.795 ;
        RECT 113.635 144.625 113.805 144.795 ;
        RECT 114.095 144.625 114.265 144.795 ;
        RECT 114.555 144.625 114.725 144.795 ;
        RECT 115.015 144.625 115.185 144.795 ;
        RECT 115.475 144.625 115.645 144.795 ;
        RECT 115.935 144.625 116.105 144.795 ;
        RECT 116.395 144.625 116.565 144.795 ;
        RECT 116.855 144.625 117.025 144.795 ;
        RECT 117.315 144.625 117.485 144.795 ;
        RECT 117.775 144.625 117.945 144.795 ;
        RECT 118.235 144.625 118.405 144.795 ;
        RECT 118.695 144.625 118.865 144.795 ;
        RECT 119.155 144.625 119.325 144.795 ;
        RECT 119.615 144.625 119.785 144.795 ;
        RECT 120.075 144.625 120.245 144.795 ;
        RECT 120.535 144.625 120.705 144.795 ;
        RECT 120.995 144.625 121.165 144.795 ;
        RECT 121.455 144.625 121.625 144.795 ;
        RECT 121.915 144.625 122.085 144.795 ;
        RECT 122.375 144.625 122.545 144.795 ;
        RECT 122.835 144.625 123.005 144.795 ;
        RECT 123.295 144.625 123.465 144.795 ;
        RECT 123.755 144.625 123.925 144.795 ;
        RECT 124.215 144.625 124.385 144.795 ;
        RECT 124.675 144.625 124.845 144.795 ;
        RECT 125.135 144.625 125.305 144.795 ;
        RECT 125.595 144.625 125.765 144.795 ;
        RECT 126.055 144.625 126.225 144.795 ;
        RECT 126.515 144.625 126.685 144.795 ;
        RECT 126.975 144.625 127.145 144.795 ;
        RECT 127.435 144.625 127.605 144.795 ;
        RECT 127.895 144.625 128.065 144.795 ;
        RECT 128.355 144.625 128.525 144.795 ;
        RECT 128.815 144.625 128.985 144.795 ;
        RECT 129.275 144.625 129.445 144.795 ;
        RECT 129.735 144.625 129.905 144.795 ;
        RECT 130.195 144.625 130.365 144.795 ;
        RECT 130.655 144.625 130.825 144.795 ;
        RECT 131.115 144.625 131.285 144.795 ;
        RECT 131.575 144.625 131.745 144.795 ;
        RECT 132.035 144.625 132.205 144.795 ;
        RECT 132.495 144.625 132.665 144.795 ;
        RECT 132.955 144.625 133.125 144.795 ;
        RECT 133.415 144.625 133.585 144.795 ;
        RECT 133.875 144.625 134.045 144.795 ;
        RECT 134.335 144.625 134.505 144.795 ;
        RECT 134.795 144.625 134.965 144.795 ;
        RECT 135.255 144.625 135.425 144.795 ;
        RECT 135.715 144.625 135.885 144.795 ;
        RECT 136.175 144.625 136.345 144.795 ;
        RECT 136.635 144.625 136.805 144.795 ;
        RECT 137.095 144.625 137.265 144.795 ;
        RECT 137.555 144.625 137.725 144.795 ;
        RECT 138.015 144.625 138.185 144.795 ;
        RECT 138.475 144.625 138.645 144.795 ;
        RECT 138.935 144.625 139.105 144.795 ;
        RECT 139.395 144.625 139.565 144.795 ;
        RECT 139.855 144.625 140.025 144.795 ;
        RECT 140.315 144.625 140.485 144.795 ;
        RECT 140.775 144.625 140.945 144.795 ;
        RECT 141.235 144.625 141.405 144.795 ;
        RECT 141.695 144.625 141.865 144.795 ;
        RECT 142.155 144.625 142.325 144.795 ;
        RECT 142.615 144.625 142.785 144.795 ;
        RECT 143.075 144.625 143.245 144.795 ;
        RECT 143.535 144.625 143.705 144.795 ;
        RECT 143.995 144.625 144.165 144.795 ;
        RECT 144.455 144.625 144.625 144.795 ;
        RECT 144.915 144.625 145.085 144.795 ;
        RECT 145.375 144.625 145.545 144.795 ;
        RECT 145.835 144.625 146.005 144.795 ;
        RECT 146.295 144.625 146.465 144.795 ;
        RECT 146.755 144.625 146.925 144.795 ;
        RECT 147.215 144.625 147.385 144.795 ;
        RECT 147.675 144.625 147.845 144.795 ;
        RECT 148.135 144.625 148.305 144.795 ;
        RECT 148.595 144.625 148.765 144.795 ;
        RECT 149.055 144.625 149.225 144.795 ;
        RECT 149.515 144.625 149.685 144.795 ;
        RECT 149.975 144.625 150.145 144.795 ;
        RECT 150.435 144.625 150.605 144.795 ;
        RECT 150.895 144.625 151.065 144.795 ;
        RECT 151.355 144.625 151.525 144.795 ;
        RECT 151.815 144.625 151.985 144.795 ;
        RECT 152.275 144.625 152.445 144.795 ;
        RECT 152.735 144.625 152.905 144.795 ;
        RECT 153.195 144.625 153.365 144.795 ;
        RECT 153.655 144.625 153.825 144.795 ;
        RECT 154.115 144.625 154.285 144.795 ;
        RECT 154.575 144.625 154.745 144.795 ;
        RECT 155.035 144.625 155.205 144.795 ;
        RECT 155.495 144.625 155.665 144.795 ;
        RECT 155.955 144.625 156.125 144.795 ;
        RECT 76.375 144.115 76.545 144.285 ;
        RECT 74.995 143.435 75.165 143.605 ;
        RECT 74.075 142.415 74.245 142.585 ;
        RECT 76.835 143.435 77.005 143.605 ;
        RECT 83.275 144.115 83.445 144.285 ;
        RECT 83.275 143.095 83.445 143.265 ;
        RECT 84.655 143.435 84.825 143.605 ;
        RECT 85.115 143.435 85.285 143.605 ;
        RECT 84.195 143.095 84.365 143.265 ;
        RECT 86.035 142.415 86.205 142.585 ;
        RECT 92.475 143.435 92.645 143.605 ;
        RECT 93.395 143.435 93.565 143.605 ;
        RECT 93.855 143.435 94.025 143.605 ;
        RECT 95.235 143.435 95.405 143.605 ;
        RECT 97.075 143.485 97.245 143.655 ;
        RECT 97.995 143.435 98.165 143.605 ;
        RECT 96.155 142.415 96.325 142.585 ;
        RECT 98.455 143.095 98.625 143.265 ;
        RECT 99.835 143.435 100.005 143.605 ;
        RECT 100.755 142.415 100.925 142.585 ;
        RECT 102.595 143.435 102.765 143.605 ;
        RECT 103.975 143.435 104.145 143.605 ;
        RECT 103.055 143.095 103.225 143.265 ;
        RECT 104.895 143.095 105.065 143.265 ;
        RECT 106.275 143.435 106.445 143.605 ;
        RECT 108.115 143.435 108.285 143.605 ;
        RECT 105.355 142.415 105.525 142.585 ;
        RECT 107.195 143.095 107.365 143.265 ;
        RECT 107.655 143.095 107.825 143.265 ;
        RECT 109.095 143.435 109.265 143.605 ;
        RECT 115.935 143.435 116.105 143.605 ;
        RECT 115.015 143.095 115.185 143.265 ;
        RECT 117.315 143.435 117.485 143.605 ;
        RECT 117.835 143.435 118.005 143.605 ;
        RECT 116.855 143.095 117.025 143.265 ;
        RECT 124.675 144.115 124.845 144.285 ;
        RECT 127.895 144.115 128.065 144.285 ;
        RECT 118.695 143.435 118.865 143.605 ;
        RECT 126.055 143.775 126.225 143.945 ;
        RECT 125.595 143.435 125.765 143.605 ;
        RECT 126.975 143.775 127.145 143.945 ;
        RECT 128.355 143.095 128.525 143.265 ;
        RECT 129.735 143.435 129.905 143.605 ;
        RECT 136.635 143.435 136.805 143.605 ;
        RECT 137.095 143.095 137.265 143.265 ;
        RECT 137.555 143.095 137.725 143.265 ;
        RECT 138.015 143.095 138.185 143.265 ;
        RECT 138.935 142.415 139.105 142.585 ;
        RECT 141.235 143.775 141.405 143.945 ;
        RECT 142.155 143.435 142.325 143.605 ;
        RECT 142.615 143.435 142.785 143.605 ;
        RECT 143.535 143.435 143.705 143.605 ;
        RECT 140.315 142.415 140.485 142.585 ;
        RECT 143.075 142.415 143.245 142.585 ;
        RECT 150.895 143.435 151.065 143.605 ;
        RECT 151.355 143.095 151.525 143.265 ;
        RECT 149.055 142.415 149.225 142.585 ;
        RECT 70.855 141.905 71.025 142.075 ;
        RECT 71.315 141.905 71.485 142.075 ;
        RECT 71.775 141.905 71.945 142.075 ;
        RECT 72.235 141.905 72.405 142.075 ;
        RECT 72.695 141.905 72.865 142.075 ;
        RECT 73.155 141.905 73.325 142.075 ;
        RECT 73.615 141.905 73.785 142.075 ;
        RECT 74.075 141.905 74.245 142.075 ;
        RECT 74.535 141.905 74.705 142.075 ;
        RECT 74.995 141.905 75.165 142.075 ;
        RECT 75.455 141.905 75.625 142.075 ;
        RECT 75.915 141.905 76.085 142.075 ;
        RECT 76.375 141.905 76.545 142.075 ;
        RECT 76.835 141.905 77.005 142.075 ;
        RECT 77.295 141.905 77.465 142.075 ;
        RECT 77.755 141.905 77.925 142.075 ;
        RECT 78.215 141.905 78.385 142.075 ;
        RECT 78.675 141.905 78.845 142.075 ;
        RECT 79.135 141.905 79.305 142.075 ;
        RECT 79.595 141.905 79.765 142.075 ;
        RECT 80.055 141.905 80.225 142.075 ;
        RECT 80.515 141.905 80.685 142.075 ;
        RECT 80.975 141.905 81.145 142.075 ;
        RECT 81.435 141.905 81.605 142.075 ;
        RECT 81.895 141.905 82.065 142.075 ;
        RECT 82.355 141.905 82.525 142.075 ;
        RECT 82.815 141.905 82.985 142.075 ;
        RECT 83.275 141.905 83.445 142.075 ;
        RECT 83.735 141.905 83.905 142.075 ;
        RECT 84.195 141.905 84.365 142.075 ;
        RECT 84.655 141.905 84.825 142.075 ;
        RECT 85.115 141.905 85.285 142.075 ;
        RECT 85.575 141.905 85.745 142.075 ;
        RECT 86.035 141.905 86.205 142.075 ;
        RECT 86.495 141.905 86.665 142.075 ;
        RECT 86.955 141.905 87.125 142.075 ;
        RECT 87.415 141.905 87.585 142.075 ;
        RECT 87.875 141.905 88.045 142.075 ;
        RECT 88.335 141.905 88.505 142.075 ;
        RECT 88.795 141.905 88.965 142.075 ;
        RECT 89.255 141.905 89.425 142.075 ;
        RECT 89.715 141.905 89.885 142.075 ;
        RECT 90.175 141.905 90.345 142.075 ;
        RECT 90.635 141.905 90.805 142.075 ;
        RECT 91.095 141.905 91.265 142.075 ;
        RECT 91.555 141.905 91.725 142.075 ;
        RECT 92.015 141.905 92.185 142.075 ;
        RECT 92.475 141.905 92.645 142.075 ;
        RECT 92.935 141.905 93.105 142.075 ;
        RECT 93.395 141.905 93.565 142.075 ;
        RECT 93.855 141.905 94.025 142.075 ;
        RECT 94.315 141.905 94.485 142.075 ;
        RECT 94.775 141.905 94.945 142.075 ;
        RECT 95.235 141.905 95.405 142.075 ;
        RECT 95.695 141.905 95.865 142.075 ;
        RECT 96.155 141.905 96.325 142.075 ;
        RECT 96.615 141.905 96.785 142.075 ;
        RECT 97.075 141.905 97.245 142.075 ;
        RECT 97.535 141.905 97.705 142.075 ;
        RECT 97.995 141.905 98.165 142.075 ;
        RECT 98.455 141.905 98.625 142.075 ;
        RECT 98.915 141.905 99.085 142.075 ;
        RECT 99.375 141.905 99.545 142.075 ;
        RECT 99.835 141.905 100.005 142.075 ;
        RECT 100.295 141.905 100.465 142.075 ;
        RECT 100.755 141.905 100.925 142.075 ;
        RECT 101.215 141.905 101.385 142.075 ;
        RECT 101.675 141.905 101.845 142.075 ;
        RECT 102.135 141.905 102.305 142.075 ;
        RECT 102.595 141.905 102.765 142.075 ;
        RECT 103.055 141.905 103.225 142.075 ;
        RECT 103.515 141.905 103.685 142.075 ;
        RECT 103.975 141.905 104.145 142.075 ;
        RECT 104.435 141.905 104.605 142.075 ;
        RECT 104.895 141.905 105.065 142.075 ;
        RECT 105.355 141.905 105.525 142.075 ;
        RECT 105.815 141.905 105.985 142.075 ;
        RECT 106.275 141.905 106.445 142.075 ;
        RECT 106.735 141.905 106.905 142.075 ;
        RECT 107.195 141.905 107.365 142.075 ;
        RECT 107.655 141.905 107.825 142.075 ;
        RECT 108.115 141.905 108.285 142.075 ;
        RECT 108.575 141.905 108.745 142.075 ;
        RECT 109.035 141.905 109.205 142.075 ;
        RECT 109.495 141.905 109.665 142.075 ;
        RECT 109.955 141.905 110.125 142.075 ;
        RECT 110.415 141.905 110.585 142.075 ;
        RECT 110.875 141.905 111.045 142.075 ;
        RECT 111.335 141.905 111.505 142.075 ;
        RECT 111.795 141.905 111.965 142.075 ;
        RECT 112.255 141.905 112.425 142.075 ;
        RECT 112.715 141.905 112.885 142.075 ;
        RECT 113.175 141.905 113.345 142.075 ;
        RECT 113.635 141.905 113.805 142.075 ;
        RECT 114.095 141.905 114.265 142.075 ;
        RECT 114.555 141.905 114.725 142.075 ;
        RECT 115.015 141.905 115.185 142.075 ;
        RECT 115.475 141.905 115.645 142.075 ;
        RECT 115.935 141.905 116.105 142.075 ;
        RECT 116.395 141.905 116.565 142.075 ;
        RECT 116.855 141.905 117.025 142.075 ;
        RECT 117.315 141.905 117.485 142.075 ;
        RECT 117.775 141.905 117.945 142.075 ;
        RECT 118.235 141.905 118.405 142.075 ;
        RECT 118.695 141.905 118.865 142.075 ;
        RECT 119.155 141.905 119.325 142.075 ;
        RECT 119.615 141.905 119.785 142.075 ;
        RECT 120.075 141.905 120.245 142.075 ;
        RECT 120.535 141.905 120.705 142.075 ;
        RECT 120.995 141.905 121.165 142.075 ;
        RECT 121.455 141.905 121.625 142.075 ;
        RECT 121.915 141.905 122.085 142.075 ;
        RECT 122.375 141.905 122.545 142.075 ;
        RECT 122.835 141.905 123.005 142.075 ;
        RECT 123.295 141.905 123.465 142.075 ;
        RECT 123.755 141.905 123.925 142.075 ;
        RECT 124.215 141.905 124.385 142.075 ;
        RECT 124.675 141.905 124.845 142.075 ;
        RECT 125.135 141.905 125.305 142.075 ;
        RECT 125.595 141.905 125.765 142.075 ;
        RECT 126.055 141.905 126.225 142.075 ;
        RECT 126.515 141.905 126.685 142.075 ;
        RECT 126.975 141.905 127.145 142.075 ;
        RECT 127.435 141.905 127.605 142.075 ;
        RECT 127.895 141.905 128.065 142.075 ;
        RECT 128.355 141.905 128.525 142.075 ;
        RECT 128.815 141.905 128.985 142.075 ;
        RECT 129.275 141.905 129.445 142.075 ;
        RECT 129.735 141.905 129.905 142.075 ;
        RECT 130.195 141.905 130.365 142.075 ;
        RECT 130.655 141.905 130.825 142.075 ;
        RECT 131.115 141.905 131.285 142.075 ;
        RECT 131.575 141.905 131.745 142.075 ;
        RECT 132.035 141.905 132.205 142.075 ;
        RECT 132.495 141.905 132.665 142.075 ;
        RECT 132.955 141.905 133.125 142.075 ;
        RECT 133.415 141.905 133.585 142.075 ;
        RECT 133.875 141.905 134.045 142.075 ;
        RECT 134.335 141.905 134.505 142.075 ;
        RECT 134.795 141.905 134.965 142.075 ;
        RECT 135.255 141.905 135.425 142.075 ;
        RECT 135.715 141.905 135.885 142.075 ;
        RECT 136.175 141.905 136.345 142.075 ;
        RECT 136.635 141.905 136.805 142.075 ;
        RECT 137.095 141.905 137.265 142.075 ;
        RECT 137.555 141.905 137.725 142.075 ;
        RECT 138.015 141.905 138.185 142.075 ;
        RECT 138.475 141.905 138.645 142.075 ;
        RECT 138.935 141.905 139.105 142.075 ;
        RECT 139.395 141.905 139.565 142.075 ;
        RECT 139.855 141.905 140.025 142.075 ;
        RECT 140.315 141.905 140.485 142.075 ;
        RECT 140.775 141.905 140.945 142.075 ;
        RECT 141.235 141.905 141.405 142.075 ;
        RECT 141.695 141.905 141.865 142.075 ;
        RECT 142.155 141.905 142.325 142.075 ;
        RECT 142.615 141.905 142.785 142.075 ;
        RECT 143.075 141.905 143.245 142.075 ;
        RECT 143.535 141.905 143.705 142.075 ;
        RECT 143.995 141.905 144.165 142.075 ;
        RECT 144.455 141.905 144.625 142.075 ;
        RECT 144.915 141.905 145.085 142.075 ;
        RECT 145.375 141.905 145.545 142.075 ;
        RECT 145.835 141.905 146.005 142.075 ;
        RECT 146.295 141.905 146.465 142.075 ;
        RECT 146.755 141.905 146.925 142.075 ;
        RECT 147.215 141.905 147.385 142.075 ;
        RECT 147.675 141.905 147.845 142.075 ;
        RECT 148.135 141.905 148.305 142.075 ;
        RECT 148.595 141.905 148.765 142.075 ;
        RECT 149.055 141.905 149.225 142.075 ;
        RECT 149.515 141.905 149.685 142.075 ;
        RECT 149.975 141.905 150.145 142.075 ;
        RECT 150.435 141.905 150.605 142.075 ;
        RECT 150.895 141.905 151.065 142.075 ;
        RECT 151.355 141.905 151.525 142.075 ;
        RECT 151.815 141.905 151.985 142.075 ;
        RECT 152.275 141.905 152.445 142.075 ;
        RECT 152.735 141.905 152.905 142.075 ;
        RECT 153.195 141.905 153.365 142.075 ;
        RECT 153.655 141.905 153.825 142.075 ;
        RECT 154.115 141.905 154.285 142.075 ;
        RECT 154.575 141.905 154.745 142.075 ;
        RECT 155.035 141.905 155.205 142.075 ;
        RECT 155.495 141.905 155.665 142.075 ;
        RECT 155.955 141.905 156.125 142.075 ;
        RECT 72.720 141.055 72.890 141.225 ;
        RECT 72.235 140.375 72.405 140.545 ;
        RECT 73.115 140.715 73.285 140.885 ;
        RECT 73.570 140.035 73.740 140.205 ;
        RECT 74.820 141.055 74.990 141.225 ;
        RECT 74.305 140.715 74.475 140.885 ;
        RECT 76.390 141.055 76.560 141.225 ;
        RECT 76.825 140.715 76.995 140.885 ;
        RECT 79.135 139.695 79.305 139.865 ;
        RECT 80.515 140.375 80.685 140.545 ;
        RECT 81.435 140.375 81.605 140.545 ;
        RECT 79.595 139.695 79.765 139.865 ;
        RECT 82.355 140.035 82.525 140.205 ;
        RECT 84.680 141.055 84.850 141.225 ;
        RECT 84.195 140.715 84.365 140.885 ;
        RECT 82.815 139.695 82.985 139.865 ;
        RECT 85.075 140.715 85.245 140.885 ;
        RECT 85.530 140.375 85.700 140.545 ;
        RECT 86.780 141.055 86.950 141.225 ;
        RECT 86.265 140.715 86.435 140.885 ;
        RECT 88.350 141.055 88.520 141.225 ;
        RECT 88.785 140.715 88.955 140.885 ;
        RECT 91.095 141.395 91.265 141.565 ;
        RECT 98.915 141.395 99.085 141.565 ;
        RECT 96.155 140.375 96.325 140.545 ;
        RECT 96.615 140.375 96.785 140.545 ;
        RECT 97.075 140.375 97.245 140.545 ;
        RECT 94.775 139.695 94.945 139.865 ;
        RECT 97.995 140.375 98.165 140.545 ;
        RECT 98.455 140.375 98.625 140.545 ;
        RECT 99.835 140.375 100.005 140.545 ;
        RECT 100.755 139.695 100.925 139.865 ;
        RECT 105.815 141.055 105.985 141.225 ;
        RECT 106.275 140.715 106.445 140.885 ;
        RECT 104.895 140.375 105.065 140.545 ;
        RECT 103.975 139.695 104.145 139.865 ;
        RECT 115.935 140.375 116.105 140.545 ;
        RECT 116.855 140.375 117.025 140.545 ;
        RECT 116.855 139.695 117.025 139.865 ;
        RECT 125.135 141.395 125.305 141.565 ;
        RECT 123.295 140.375 123.465 140.545 ;
        RECT 124.675 140.715 124.845 140.885 ;
        RECT 126.055 140.375 126.225 140.545 ;
        RECT 129.735 140.375 129.905 140.545 ;
        RECT 131.115 140.715 131.285 140.885 ;
        RECT 132.495 140.715 132.665 140.885 ;
        RECT 132.955 140.375 133.125 140.545 ;
        RECT 133.415 140.375 133.585 140.545 ;
        RECT 133.875 140.375 134.045 140.545 ;
        RECT 135.715 141.395 135.885 141.565 ;
        RECT 137.095 140.375 137.265 140.545 ;
        RECT 137.555 140.375 137.725 140.545 ;
        RECT 138.015 140.375 138.185 140.545 ;
        RECT 134.795 139.695 134.965 139.865 ;
        RECT 138.935 140.375 139.105 140.545 ;
        RECT 140.315 140.715 140.485 140.885 ;
        RECT 140.775 140.375 140.945 140.545 ;
        RECT 141.235 140.715 141.405 140.885 ;
        RECT 141.695 140.715 141.865 140.885 ;
        RECT 144.455 140.375 144.625 140.545 ;
        RECT 144.915 140.375 145.085 140.545 ;
        RECT 139.395 139.695 139.565 139.865 ;
        RECT 143.535 139.695 143.705 139.865 ;
        RECT 146.295 140.375 146.465 140.545 ;
        RECT 146.755 140.035 146.925 140.205 ;
        RECT 147.215 140.375 147.385 140.545 ;
        RECT 148.595 141.055 148.765 141.225 ;
        RECT 148.135 140.375 148.305 140.545 ;
        RECT 149.055 140.715 149.225 140.885 ;
        RECT 149.515 140.375 149.685 140.545 ;
        RECT 151.815 140.375 151.985 140.545 ;
        RECT 152.735 140.375 152.905 140.545 ;
        RECT 154.115 140.035 154.285 140.205 ;
        RECT 154.575 140.375 154.745 140.545 ;
        RECT 70.855 139.185 71.025 139.355 ;
        RECT 71.315 139.185 71.485 139.355 ;
        RECT 71.775 139.185 71.945 139.355 ;
        RECT 72.235 139.185 72.405 139.355 ;
        RECT 72.695 139.185 72.865 139.355 ;
        RECT 73.155 139.185 73.325 139.355 ;
        RECT 73.615 139.185 73.785 139.355 ;
        RECT 74.075 139.185 74.245 139.355 ;
        RECT 74.535 139.185 74.705 139.355 ;
        RECT 74.995 139.185 75.165 139.355 ;
        RECT 75.455 139.185 75.625 139.355 ;
        RECT 75.915 139.185 76.085 139.355 ;
        RECT 76.375 139.185 76.545 139.355 ;
        RECT 76.835 139.185 77.005 139.355 ;
        RECT 77.295 139.185 77.465 139.355 ;
        RECT 77.755 139.185 77.925 139.355 ;
        RECT 78.215 139.185 78.385 139.355 ;
        RECT 78.675 139.185 78.845 139.355 ;
        RECT 79.135 139.185 79.305 139.355 ;
        RECT 79.595 139.185 79.765 139.355 ;
        RECT 80.055 139.185 80.225 139.355 ;
        RECT 80.515 139.185 80.685 139.355 ;
        RECT 80.975 139.185 81.145 139.355 ;
        RECT 81.435 139.185 81.605 139.355 ;
        RECT 81.895 139.185 82.065 139.355 ;
        RECT 82.355 139.185 82.525 139.355 ;
        RECT 82.815 139.185 82.985 139.355 ;
        RECT 83.275 139.185 83.445 139.355 ;
        RECT 83.735 139.185 83.905 139.355 ;
        RECT 84.195 139.185 84.365 139.355 ;
        RECT 84.655 139.185 84.825 139.355 ;
        RECT 85.115 139.185 85.285 139.355 ;
        RECT 85.575 139.185 85.745 139.355 ;
        RECT 86.035 139.185 86.205 139.355 ;
        RECT 86.495 139.185 86.665 139.355 ;
        RECT 86.955 139.185 87.125 139.355 ;
        RECT 87.415 139.185 87.585 139.355 ;
        RECT 87.875 139.185 88.045 139.355 ;
        RECT 88.335 139.185 88.505 139.355 ;
        RECT 88.795 139.185 88.965 139.355 ;
        RECT 89.255 139.185 89.425 139.355 ;
        RECT 89.715 139.185 89.885 139.355 ;
        RECT 90.175 139.185 90.345 139.355 ;
        RECT 90.635 139.185 90.805 139.355 ;
        RECT 91.095 139.185 91.265 139.355 ;
        RECT 91.555 139.185 91.725 139.355 ;
        RECT 92.015 139.185 92.185 139.355 ;
        RECT 92.475 139.185 92.645 139.355 ;
        RECT 92.935 139.185 93.105 139.355 ;
        RECT 93.395 139.185 93.565 139.355 ;
        RECT 93.855 139.185 94.025 139.355 ;
        RECT 94.315 139.185 94.485 139.355 ;
        RECT 94.775 139.185 94.945 139.355 ;
        RECT 95.235 139.185 95.405 139.355 ;
        RECT 95.695 139.185 95.865 139.355 ;
        RECT 96.155 139.185 96.325 139.355 ;
        RECT 96.615 139.185 96.785 139.355 ;
        RECT 97.075 139.185 97.245 139.355 ;
        RECT 97.535 139.185 97.705 139.355 ;
        RECT 97.995 139.185 98.165 139.355 ;
        RECT 98.455 139.185 98.625 139.355 ;
        RECT 98.915 139.185 99.085 139.355 ;
        RECT 99.375 139.185 99.545 139.355 ;
        RECT 99.835 139.185 100.005 139.355 ;
        RECT 100.295 139.185 100.465 139.355 ;
        RECT 100.755 139.185 100.925 139.355 ;
        RECT 101.215 139.185 101.385 139.355 ;
        RECT 101.675 139.185 101.845 139.355 ;
        RECT 102.135 139.185 102.305 139.355 ;
        RECT 102.595 139.185 102.765 139.355 ;
        RECT 103.055 139.185 103.225 139.355 ;
        RECT 103.515 139.185 103.685 139.355 ;
        RECT 103.975 139.185 104.145 139.355 ;
        RECT 104.435 139.185 104.605 139.355 ;
        RECT 104.895 139.185 105.065 139.355 ;
        RECT 105.355 139.185 105.525 139.355 ;
        RECT 105.815 139.185 105.985 139.355 ;
        RECT 106.275 139.185 106.445 139.355 ;
        RECT 106.735 139.185 106.905 139.355 ;
        RECT 107.195 139.185 107.365 139.355 ;
        RECT 107.655 139.185 107.825 139.355 ;
        RECT 108.115 139.185 108.285 139.355 ;
        RECT 108.575 139.185 108.745 139.355 ;
        RECT 109.035 139.185 109.205 139.355 ;
        RECT 109.495 139.185 109.665 139.355 ;
        RECT 109.955 139.185 110.125 139.355 ;
        RECT 110.415 139.185 110.585 139.355 ;
        RECT 110.875 139.185 111.045 139.355 ;
        RECT 111.335 139.185 111.505 139.355 ;
        RECT 111.795 139.185 111.965 139.355 ;
        RECT 112.255 139.185 112.425 139.355 ;
        RECT 112.715 139.185 112.885 139.355 ;
        RECT 113.175 139.185 113.345 139.355 ;
        RECT 113.635 139.185 113.805 139.355 ;
        RECT 114.095 139.185 114.265 139.355 ;
        RECT 114.555 139.185 114.725 139.355 ;
        RECT 115.015 139.185 115.185 139.355 ;
        RECT 115.475 139.185 115.645 139.355 ;
        RECT 115.935 139.185 116.105 139.355 ;
        RECT 116.395 139.185 116.565 139.355 ;
        RECT 116.855 139.185 117.025 139.355 ;
        RECT 117.315 139.185 117.485 139.355 ;
        RECT 117.775 139.185 117.945 139.355 ;
        RECT 118.235 139.185 118.405 139.355 ;
        RECT 118.695 139.185 118.865 139.355 ;
        RECT 119.155 139.185 119.325 139.355 ;
        RECT 119.615 139.185 119.785 139.355 ;
        RECT 120.075 139.185 120.245 139.355 ;
        RECT 120.535 139.185 120.705 139.355 ;
        RECT 120.995 139.185 121.165 139.355 ;
        RECT 121.455 139.185 121.625 139.355 ;
        RECT 121.915 139.185 122.085 139.355 ;
        RECT 122.375 139.185 122.545 139.355 ;
        RECT 122.835 139.185 123.005 139.355 ;
        RECT 123.295 139.185 123.465 139.355 ;
        RECT 123.755 139.185 123.925 139.355 ;
        RECT 124.215 139.185 124.385 139.355 ;
        RECT 124.675 139.185 124.845 139.355 ;
        RECT 125.135 139.185 125.305 139.355 ;
        RECT 125.595 139.185 125.765 139.355 ;
        RECT 126.055 139.185 126.225 139.355 ;
        RECT 126.515 139.185 126.685 139.355 ;
        RECT 126.975 139.185 127.145 139.355 ;
        RECT 127.435 139.185 127.605 139.355 ;
        RECT 127.895 139.185 128.065 139.355 ;
        RECT 128.355 139.185 128.525 139.355 ;
        RECT 128.815 139.185 128.985 139.355 ;
        RECT 129.275 139.185 129.445 139.355 ;
        RECT 129.735 139.185 129.905 139.355 ;
        RECT 130.195 139.185 130.365 139.355 ;
        RECT 130.655 139.185 130.825 139.355 ;
        RECT 131.115 139.185 131.285 139.355 ;
        RECT 131.575 139.185 131.745 139.355 ;
        RECT 132.035 139.185 132.205 139.355 ;
        RECT 132.495 139.185 132.665 139.355 ;
        RECT 132.955 139.185 133.125 139.355 ;
        RECT 133.415 139.185 133.585 139.355 ;
        RECT 133.875 139.185 134.045 139.355 ;
        RECT 134.335 139.185 134.505 139.355 ;
        RECT 134.795 139.185 134.965 139.355 ;
        RECT 135.255 139.185 135.425 139.355 ;
        RECT 135.715 139.185 135.885 139.355 ;
        RECT 136.175 139.185 136.345 139.355 ;
        RECT 136.635 139.185 136.805 139.355 ;
        RECT 137.095 139.185 137.265 139.355 ;
        RECT 137.555 139.185 137.725 139.355 ;
        RECT 138.015 139.185 138.185 139.355 ;
        RECT 138.475 139.185 138.645 139.355 ;
        RECT 138.935 139.185 139.105 139.355 ;
        RECT 139.395 139.185 139.565 139.355 ;
        RECT 139.855 139.185 140.025 139.355 ;
        RECT 140.315 139.185 140.485 139.355 ;
        RECT 140.775 139.185 140.945 139.355 ;
        RECT 141.235 139.185 141.405 139.355 ;
        RECT 141.695 139.185 141.865 139.355 ;
        RECT 142.155 139.185 142.325 139.355 ;
        RECT 142.615 139.185 142.785 139.355 ;
        RECT 143.075 139.185 143.245 139.355 ;
        RECT 143.535 139.185 143.705 139.355 ;
        RECT 143.995 139.185 144.165 139.355 ;
        RECT 144.455 139.185 144.625 139.355 ;
        RECT 144.915 139.185 145.085 139.355 ;
        RECT 145.375 139.185 145.545 139.355 ;
        RECT 145.835 139.185 146.005 139.355 ;
        RECT 146.295 139.185 146.465 139.355 ;
        RECT 146.755 139.185 146.925 139.355 ;
        RECT 147.215 139.185 147.385 139.355 ;
        RECT 147.675 139.185 147.845 139.355 ;
        RECT 148.135 139.185 148.305 139.355 ;
        RECT 148.595 139.185 148.765 139.355 ;
        RECT 149.055 139.185 149.225 139.355 ;
        RECT 149.515 139.185 149.685 139.355 ;
        RECT 149.975 139.185 150.145 139.355 ;
        RECT 150.435 139.185 150.605 139.355 ;
        RECT 150.895 139.185 151.065 139.355 ;
        RECT 151.355 139.185 151.525 139.355 ;
        RECT 151.815 139.185 151.985 139.355 ;
        RECT 152.275 139.185 152.445 139.355 ;
        RECT 152.735 139.185 152.905 139.355 ;
        RECT 153.195 139.185 153.365 139.355 ;
        RECT 153.655 139.185 153.825 139.355 ;
        RECT 154.115 139.185 154.285 139.355 ;
        RECT 154.575 139.185 154.745 139.355 ;
        RECT 155.035 139.185 155.205 139.355 ;
        RECT 155.495 139.185 155.665 139.355 ;
        RECT 155.955 139.185 156.125 139.355 ;
        RECT 79.135 138.675 79.305 138.845 ;
        RECT 78.215 137.995 78.385 138.165 ;
        RECT 79.595 137.995 79.765 138.165 ;
        RECT 80.055 137.995 80.225 138.165 ;
        RECT 81.895 138.675 82.065 138.845 ;
        RECT 80.975 137.995 81.145 138.165 ;
        RECT 82.355 137.995 82.525 138.165 ;
        RECT 77.295 136.975 77.465 137.145 ;
        RECT 80.055 136.975 80.225 137.145 ;
        RECT 85.575 137.655 85.745 137.825 ;
        RECT 86.955 137.995 87.125 138.165 ;
        RECT 94.315 138.335 94.485 138.505 ;
        RECT 95.235 137.995 95.405 138.165 ;
        RECT 96.155 137.315 96.325 137.485 ;
        RECT 98.455 138.335 98.625 138.505 ;
        RECT 99.375 138.335 99.545 138.505 ;
        RECT 99.835 137.995 100.005 138.165 ;
        RECT 97.535 136.975 97.705 137.145 ;
        RECT 100.755 137.315 100.925 137.485 ;
        RECT 107.195 137.995 107.365 138.165 ;
        RECT 107.655 137.995 107.825 138.165 ;
        RECT 108.115 137.995 108.285 138.165 ;
        RECT 109.035 137.995 109.205 138.165 ;
        RECT 112.715 138.335 112.885 138.505 ;
        RECT 105.815 136.975 105.985 137.145 ;
        RECT 113.635 137.995 113.805 138.165 ;
        RECT 114.555 137.315 114.725 137.485 ;
        RECT 115.475 138.335 115.645 138.505 ;
        RECT 116.855 137.995 117.025 138.165 ;
        RECT 117.315 137.995 117.485 138.165 ;
        RECT 117.775 137.995 117.945 138.165 ;
        RECT 118.695 137.995 118.865 138.165 ;
        RECT 119.615 137.995 119.785 138.165 ;
        RECT 120.075 137.655 120.245 137.825 ;
        RECT 120.535 137.995 120.705 138.165 ;
        RECT 120.995 137.655 121.165 137.825 ;
        RECT 121.915 137.655 122.085 137.825 ;
        RECT 126.515 137.315 126.685 137.485 ;
        RECT 126.055 136.975 126.225 137.145 ;
        RECT 128.355 138.335 128.525 138.505 ;
        RECT 128.815 137.995 128.985 138.165 ;
        RECT 130.155 137.995 130.325 138.165 ;
        RECT 131.115 137.995 131.285 138.165 ;
        RECT 129.735 137.315 129.905 137.485 ;
        RECT 130.655 136.975 130.825 137.145 ;
        RECT 133.415 137.995 133.585 138.165 ;
        RECT 137.555 138.675 137.725 138.845 ;
        RECT 134.335 137.995 134.505 138.165 ;
        RECT 134.795 137.995 134.965 138.165 ;
        RECT 135.255 137.995 135.425 138.165 ;
        RECT 137.095 137.995 137.265 138.165 ;
        RECT 138.015 137.995 138.185 138.165 ;
        RECT 136.635 136.975 136.805 137.145 ;
        RECT 138.935 137.655 139.105 137.825 ;
        RECT 139.395 137.655 139.565 137.825 ;
        RECT 139.855 137.655 140.025 137.825 ;
        RECT 140.315 137.995 140.485 138.165 ;
        RECT 141.695 137.995 141.865 138.165 ;
        RECT 141.235 136.975 141.405 137.145 ;
        RECT 143.075 137.655 143.245 137.825 ;
        RECT 150.435 137.995 150.605 138.165 ;
        RECT 149.975 137.655 150.145 137.825 ;
        RECT 151.815 137.995 151.985 138.165 ;
        RECT 148.595 137.315 148.765 137.485 ;
        RECT 152.275 136.975 152.445 137.145 ;
        RECT 154.115 136.975 154.285 137.145 ;
        RECT 70.855 136.465 71.025 136.635 ;
        RECT 71.315 136.465 71.485 136.635 ;
        RECT 71.775 136.465 71.945 136.635 ;
        RECT 72.235 136.465 72.405 136.635 ;
        RECT 72.695 136.465 72.865 136.635 ;
        RECT 73.155 136.465 73.325 136.635 ;
        RECT 73.615 136.465 73.785 136.635 ;
        RECT 74.075 136.465 74.245 136.635 ;
        RECT 74.535 136.465 74.705 136.635 ;
        RECT 74.995 136.465 75.165 136.635 ;
        RECT 75.455 136.465 75.625 136.635 ;
        RECT 75.915 136.465 76.085 136.635 ;
        RECT 76.375 136.465 76.545 136.635 ;
        RECT 76.835 136.465 77.005 136.635 ;
        RECT 77.295 136.465 77.465 136.635 ;
        RECT 77.755 136.465 77.925 136.635 ;
        RECT 78.215 136.465 78.385 136.635 ;
        RECT 78.675 136.465 78.845 136.635 ;
        RECT 79.135 136.465 79.305 136.635 ;
        RECT 79.595 136.465 79.765 136.635 ;
        RECT 80.055 136.465 80.225 136.635 ;
        RECT 80.515 136.465 80.685 136.635 ;
        RECT 80.975 136.465 81.145 136.635 ;
        RECT 81.435 136.465 81.605 136.635 ;
        RECT 81.895 136.465 82.065 136.635 ;
        RECT 82.355 136.465 82.525 136.635 ;
        RECT 82.815 136.465 82.985 136.635 ;
        RECT 83.275 136.465 83.445 136.635 ;
        RECT 83.735 136.465 83.905 136.635 ;
        RECT 84.195 136.465 84.365 136.635 ;
        RECT 84.655 136.465 84.825 136.635 ;
        RECT 85.115 136.465 85.285 136.635 ;
        RECT 85.575 136.465 85.745 136.635 ;
        RECT 86.035 136.465 86.205 136.635 ;
        RECT 86.495 136.465 86.665 136.635 ;
        RECT 86.955 136.465 87.125 136.635 ;
        RECT 87.415 136.465 87.585 136.635 ;
        RECT 87.875 136.465 88.045 136.635 ;
        RECT 88.335 136.465 88.505 136.635 ;
        RECT 88.795 136.465 88.965 136.635 ;
        RECT 89.255 136.465 89.425 136.635 ;
        RECT 89.715 136.465 89.885 136.635 ;
        RECT 90.175 136.465 90.345 136.635 ;
        RECT 90.635 136.465 90.805 136.635 ;
        RECT 91.095 136.465 91.265 136.635 ;
        RECT 91.555 136.465 91.725 136.635 ;
        RECT 92.015 136.465 92.185 136.635 ;
        RECT 92.475 136.465 92.645 136.635 ;
        RECT 92.935 136.465 93.105 136.635 ;
        RECT 93.395 136.465 93.565 136.635 ;
        RECT 93.855 136.465 94.025 136.635 ;
        RECT 94.315 136.465 94.485 136.635 ;
        RECT 94.775 136.465 94.945 136.635 ;
        RECT 95.235 136.465 95.405 136.635 ;
        RECT 95.695 136.465 95.865 136.635 ;
        RECT 96.155 136.465 96.325 136.635 ;
        RECT 96.615 136.465 96.785 136.635 ;
        RECT 97.075 136.465 97.245 136.635 ;
        RECT 97.535 136.465 97.705 136.635 ;
        RECT 97.995 136.465 98.165 136.635 ;
        RECT 98.455 136.465 98.625 136.635 ;
        RECT 98.915 136.465 99.085 136.635 ;
        RECT 99.375 136.465 99.545 136.635 ;
        RECT 99.835 136.465 100.005 136.635 ;
        RECT 100.295 136.465 100.465 136.635 ;
        RECT 100.755 136.465 100.925 136.635 ;
        RECT 101.215 136.465 101.385 136.635 ;
        RECT 101.675 136.465 101.845 136.635 ;
        RECT 102.135 136.465 102.305 136.635 ;
        RECT 102.595 136.465 102.765 136.635 ;
        RECT 103.055 136.465 103.225 136.635 ;
        RECT 103.515 136.465 103.685 136.635 ;
        RECT 103.975 136.465 104.145 136.635 ;
        RECT 104.435 136.465 104.605 136.635 ;
        RECT 104.895 136.465 105.065 136.635 ;
        RECT 105.355 136.465 105.525 136.635 ;
        RECT 105.815 136.465 105.985 136.635 ;
        RECT 106.275 136.465 106.445 136.635 ;
        RECT 106.735 136.465 106.905 136.635 ;
        RECT 107.195 136.465 107.365 136.635 ;
        RECT 107.655 136.465 107.825 136.635 ;
        RECT 108.115 136.465 108.285 136.635 ;
        RECT 108.575 136.465 108.745 136.635 ;
        RECT 109.035 136.465 109.205 136.635 ;
        RECT 109.495 136.465 109.665 136.635 ;
        RECT 109.955 136.465 110.125 136.635 ;
        RECT 110.415 136.465 110.585 136.635 ;
        RECT 110.875 136.465 111.045 136.635 ;
        RECT 111.335 136.465 111.505 136.635 ;
        RECT 111.795 136.465 111.965 136.635 ;
        RECT 112.255 136.465 112.425 136.635 ;
        RECT 112.715 136.465 112.885 136.635 ;
        RECT 113.175 136.465 113.345 136.635 ;
        RECT 113.635 136.465 113.805 136.635 ;
        RECT 114.095 136.465 114.265 136.635 ;
        RECT 114.555 136.465 114.725 136.635 ;
        RECT 115.015 136.465 115.185 136.635 ;
        RECT 115.475 136.465 115.645 136.635 ;
        RECT 115.935 136.465 116.105 136.635 ;
        RECT 116.395 136.465 116.565 136.635 ;
        RECT 116.855 136.465 117.025 136.635 ;
        RECT 117.315 136.465 117.485 136.635 ;
        RECT 117.775 136.465 117.945 136.635 ;
        RECT 118.235 136.465 118.405 136.635 ;
        RECT 118.695 136.465 118.865 136.635 ;
        RECT 119.155 136.465 119.325 136.635 ;
        RECT 119.615 136.465 119.785 136.635 ;
        RECT 120.075 136.465 120.245 136.635 ;
        RECT 120.535 136.465 120.705 136.635 ;
        RECT 120.995 136.465 121.165 136.635 ;
        RECT 121.455 136.465 121.625 136.635 ;
        RECT 121.915 136.465 122.085 136.635 ;
        RECT 122.375 136.465 122.545 136.635 ;
        RECT 122.835 136.465 123.005 136.635 ;
        RECT 123.295 136.465 123.465 136.635 ;
        RECT 123.755 136.465 123.925 136.635 ;
        RECT 124.215 136.465 124.385 136.635 ;
        RECT 124.675 136.465 124.845 136.635 ;
        RECT 125.135 136.465 125.305 136.635 ;
        RECT 125.595 136.465 125.765 136.635 ;
        RECT 126.055 136.465 126.225 136.635 ;
        RECT 126.515 136.465 126.685 136.635 ;
        RECT 126.975 136.465 127.145 136.635 ;
        RECT 127.435 136.465 127.605 136.635 ;
        RECT 127.895 136.465 128.065 136.635 ;
        RECT 128.355 136.465 128.525 136.635 ;
        RECT 128.815 136.465 128.985 136.635 ;
        RECT 129.275 136.465 129.445 136.635 ;
        RECT 129.735 136.465 129.905 136.635 ;
        RECT 130.195 136.465 130.365 136.635 ;
        RECT 130.655 136.465 130.825 136.635 ;
        RECT 131.115 136.465 131.285 136.635 ;
        RECT 131.575 136.465 131.745 136.635 ;
        RECT 132.035 136.465 132.205 136.635 ;
        RECT 132.495 136.465 132.665 136.635 ;
        RECT 132.955 136.465 133.125 136.635 ;
        RECT 133.415 136.465 133.585 136.635 ;
        RECT 133.875 136.465 134.045 136.635 ;
        RECT 134.335 136.465 134.505 136.635 ;
        RECT 134.795 136.465 134.965 136.635 ;
        RECT 135.255 136.465 135.425 136.635 ;
        RECT 135.715 136.465 135.885 136.635 ;
        RECT 136.175 136.465 136.345 136.635 ;
        RECT 136.635 136.465 136.805 136.635 ;
        RECT 137.095 136.465 137.265 136.635 ;
        RECT 137.555 136.465 137.725 136.635 ;
        RECT 138.015 136.465 138.185 136.635 ;
        RECT 138.475 136.465 138.645 136.635 ;
        RECT 138.935 136.465 139.105 136.635 ;
        RECT 139.395 136.465 139.565 136.635 ;
        RECT 139.855 136.465 140.025 136.635 ;
        RECT 140.315 136.465 140.485 136.635 ;
        RECT 140.775 136.465 140.945 136.635 ;
        RECT 141.235 136.465 141.405 136.635 ;
        RECT 141.695 136.465 141.865 136.635 ;
        RECT 142.155 136.465 142.325 136.635 ;
        RECT 142.615 136.465 142.785 136.635 ;
        RECT 143.075 136.465 143.245 136.635 ;
        RECT 143.535 136.465 143.705 136.635 ;
        RECT 143.995 136.465 144.165 136.635 ;
        RECT 144.455 136.465 144.625 136.635 ;
        RECT 144.915 136.465 145.085 136.635 ;
        RECT 145.375 136.465 145.545 136.635 ;
        RECT 145.835 136.465 146.005 136.635 ;
        RECT 146.295 136.465 146.465 136.635 ;
        RECT 146.755 136.465 146.925 136.635 ;
        RECT 147.215 136.465 147.385 136.635 ;
        RECT 147.675 136.465 147.845 136.635 ;
        RECT 148.135 136.465 148.305 136.635 ;
        RECT 148.595 136.465 148.765 136.635 ;
        RECT 149.055 136.465 149.225 136.635 ;
        RECT 149.515 136.465 149.685 136.635 ;
        RECT 149.975 136.465 150.145 136.635 ;
        RECT 150.435 136.465 150.605 136.635 ;
        RECT 150.895 136.465 151.065 136.635 ;
        RECT 151.355 136.465 151.525 136.635 ;
        RECT 151.815 136.465 151.985 136.635 ;
        RECT 152.275 136.465 152.445 136.635 ;
        RECT 152.735 136.465 152.905 136.635 ;
        RECT 153.195 136.465 153.365 136.635 ;
        RECT 153.655 136.465 153.825 136.635 ;
        RECT 154.115 136.465 154.285 136.635 ;
        RECT 154.575 136.465 154.745 136.635 ;
        RECT 155.035 136.465 155.205 136.635 ;
        RECT 155.495 136.465 155.665 136.635 ;
        RECT 155.955 136.465 156.125 136.635 ;
        RECT 78.675 135.955 78.845 136.125 ;
        RECT 76.835 135.275 77.005 135.445 ;
        RECT 76.375 134.935 76.545 135.105 ;
        RECT 78.675 134.935 78.845 135.105 ;
        RECT 79.595 134.935 79.765 135.105 ;
        RECT 78.215 134.255 78.385 134.425 ;
        RECT 86.495 134.935 86.665 135.105 ;
        RECT 87.875 135.275 88.045 135.445 ;
        RECT 87.415 134.935 87.585 135.105 ;
        RECT 88.795 134.935 88.965 135.105 ;
        RECT 86.955 134.255 87.125 134.425 ;
        RECT 89.715 134.255 89.885 134.425 ;
        RECT 91.095 134.935 91.265 135.105 ;
        RECT 91.555 134.935 91.725 135.105 ;
        RECT 90.175 134.255 90.345 134.425 ;
        RECT 94.315 134.935 94.485 135.105 ;
        RECT 95.235 134.935 95.405 135.105 ;
        RECT 94.775 134.595 94.945 134.765 ;
        RECT 96.615 134.935 96.785 135.105 ;
        RECT 97.075 134.935 97.245 135.105 ;
        RECT 97.535 134.935 97.705 135.105 ;
        RECT 98.125 134.935 98.295 135.105 ;
        RECT 98.915 134.935 99.085 135.105 ;
        RECT 99.835 134.935 100.005 135.105 ;
        RECT 100.295 134.935 100.465 135.105 ;
        RECT 100.755 134.935 100.925 135.105 ;
        RECT 101.255 135.275 101.425 135.445 ;
        RECT 95.695 134.255 95.865 134.425 ;
        RECT 103.975 135.955 104.145 136.125 ;
        RECT 103.055 134.935 103.225 135.105 ;
        RECT 102.135 134.255 102.305 134.425 ;
        RECT 104.435 134.935 104.605 135.105 ;
        RECT 106.275 135.275 106.445 135.445 ;
        RECT 106.735 134.935 106.905 135.105 ;
        RECT 107.195 134.935 107.365 135.105 ;
        RECT 107.655 135.275 107.825 135.445 ;
        RECT 105.355 134.255 105.525 134.425 ;
        RECT 108.575 134.255 108.745 134.425 ;
        RECT 115.935 134.935 116.105 135.105 ;
        RECT 116.395 134.935 116.565 135.105 ;
        RECT 116.855 135.275 117.025 135.445 ;
        RECT 117.315 135.275 117.485 135.445 ;
        RECT 115.015 134.255 115.185 134.425 ;
        RECT 126.975 134.935 127.145 135.105 ;
        RECT 127.895 134.935 128.065 135.105 ;
        RECT 128.355 134.935 128.525 135.105 ;
        RECT 129.275 134.935 129.445 135.105 ;
        RECT 129.735 134.935 129.905 135.105 ;
        RECT 133.875 134.935 134.045 135.105 ;
        RECT 135.715 135.275 135.885 135.445 ;
        RECT 136.635 134.935 136.805 135.105 ;
        RECT 137.095 135.275 137.265 135.445 ;
        RECT 137.555 134.935 137.725 135.105 ;
        RECT 138.015 135.275 138.185 135.445 ;
        RECT 134.795 134.255 134.965 134.425 ;
        RECT 139.855 134.595 140.025 134.765 ;
        RECT 140.775 134.595 140.945 134.765 ;
        RECT 144.455 134.935 144.625 135.105 ;
        RECT 145.835 135.275 146.005 135.445 ;
        RECT 138.935 134.255 139.105 134.425 ;
        RECT 149.975 134.935 150.145 135.105 ;
        RECT 152.275 135.955 152.445 136.125 ;
        RECT 151.815 134.935 151.985 135.105 ;
        RECT 153.195 135.275 153.365 135.445 ;
        RECT 153.655 134.935 153.825 135.105 ;
        RECT 150.895 134.255 151.065 134.425 ;
        RECT 153.195 134.595 153.365 134.765 ;
        RECT 154.575 134.935 154.745 135.105 ;
        RECT 154.575 134.255 154.745 134.425 ;
        RECT 70.855 133.745 71.025 133.915 ;
        RECT 71.315 133.745 71.485 133.915 ;
        RECT 71.775 133.745 71.945 133.915 ;
        RECT 72.235 133.745 72.405 133.915 ;
        RECT 72.695 133.745 72.865 133.915 ;
        RECT 73.155 133.745 73.325 133.915 ;
        RECT 73.615 133.745 73.785 133.915 ;
        RECT 74.075 133.745 74.245 133.915 ;
        RECT 74.535 133.745 74.705 133.915 ;
        RECT 74.995 133.745 75.165 133.915 ;
        RECT 75.455 133.745 75.625 133.915 ;
        RECT 75.915 133.745 76.085 133.915 ;
        RECT 76.375 133.745 76.545 133.915 ;
        RECT 76.835 133.745 77.005 133.915 ;
        RECT 77.295 133.745 77.465 133.915 ;
        RECT 77.755 133.745 77.925 133.915 ;
        RECT 78.215 133.745 78.385 133.915 ;
        RECT 78.675 133.745 78.845 133.915 ;
        RECT 79.135 133.745 79.305 133.915 ;
        RECT 79.595 133.745 79.765 133.915 ;
        RECT 80.055 133.745 80.225 133.915 ;
        RECT 80.515 133.745 80.685 133.915 ;
        RECT 80.975 133.745 81.145 133.915 ;
        RECT 81.435 133.745 81.605 133.915 ;
        RECT 81.895 133.745 82.065 133.915 ;
        RECT 82.355 133.745 82.525 133.915 ;
        RECT 82.815 133.745 82.985 133.915 ;
        RECT 83.275 133.745 83.445 133.915 ;
        RECT 83.735 133.745 83.905 133.915 ;
        RECT 84.195 133.745 84.365 133.915 ;
        RECT 84.655 133.745 84.825 133.915 ;
        RECT 85.115 133.745 85.285 133.915 ;
        RECT 85.575 133.745 85.745 133.915 ;
        RECT 86.035 133.745 86.205 133.915 ;
        RECT 86.495 133.745 86.665 133.915 ;
        RECT 86.955 133.745 87.125 133.915 ;
        RECT 87.415 133.745 87.585 133.915 ;
        RECT 87.875 133.745 88.045 133.915 ;
        RECT 88.335 133.745 88.505 133.915 ;
        RECT 88.795 133.745 88.965 133.915 ;
        RECT 89.255 133.745 89.425 133.915 ;
        RECT 89.715 133.745 89.885 133.915 ;
        RECT 90.175 133.745 90.345 133.915 ;
        RECT 90.635 133.745 90.805 133.915 ;
        RECT 91.095 133.745 91.265 133.915 ;
        RECT 91.555 133.745 91.725 133.915 ;
        RECT 92.015 133.745 92.185 133.915 ;
        RECT 92.475 133.745 92.645 133.915 ;
        RECT 92.935 133.745 93.105 133.915 ;
        RECT 93.395 133.745 93.565 133.915 ;
        RECT 93.855 133.745 94.025 133.915 ;
        RECT 94.315 133.745 94.485 133.915 ;
        RECT 94.775 133.745 94.945 133.915 ;
        RECT 95.235 133.745 95.405 133.915 ;
        RECT 95.695 133.745 95.865 133.915 ;
        RECT 96.155 133.745 96.325 133.915 ;
        RECT 96.615 133.745 96.785 133.915 ;
        RECT 97.075 133.745 97.245 133.915 ;
        RECT 97.535 133.745 97.705 133.915 ;
        RECT 97.995 133.745 98.165 133.915 ;
        RECT 98.455 133.745 98.625 133.915 ;
        RECT 98.915 133.745 99.085 133.915 ;
        RECT 99.375 133.745 99.545 133.915 ;
        RECT 99.835 133.745 100.005 133.915 ;
        RECT 100.295 133.745 100.465 133.915 ;
        RECT 100.755 133.745 100.925 133.915 ;
        RECT 101.215 133.745 101.385 133.915 ;
        RECT 101.675 133.745 101.845 133.915 ;
        RECT 102.135 133.745 102.305 133.915 ;
        RECT 102.595 133.745 102.765 133.915 ;
        RECT 103.055 133.745 103.225 133.915 ;
        RECT 103.515 133.745 103.685 133.915 ;
        RECT 103.975 133.745 104.145 133.915 ;
        RECT 104.435 133.745 104.605 133.915 ;
        RECT 104.895 133.745 105.065 133.915 ;
        RECT 105.355 133.745 105.525 133.915 ;
        RECT 105.815 133.745 105.985 133.915 ;
        RECT 106.275 133.745 106.445 133.915 ;
        RECT 106.735 133.745 106.905 133.915 ;
        RECT 107.195 133.745 107.365 133.915 ;
        RECT 107.655 133.745 107.825 133.915 ;
        RECT 108.115 133.745 108.285 133.915 ;
        RECT 108.575 133.745 108.745 133.915 ;
        RECT 109.035 133.745 109.205 133.915 ;
        RECT 109.495 133.745 109.665 133.915 ;
        RECT 109.955 133.745 110.125 133.915 ;
        RECT 110.415 133.745 110.585 133.915 ;
        RECT 110.875 133.745 111.045 133.915 ;
        RECT 111.335 133.745 111.505 133.915 ;
        RECT 111.795 133.745 111.965 133.915 ;
        RECT 112.255 133.745 112.425 133.915 ;
        RECT 112.715 133.745 112.885 133.915 ;
        RECT 113.175 133.745 113.345 133.915 ;
        RECT 113.635 133.745 113.805 133.915 ;
        RECT 114.095 133.745 114.265 133.915 ;
        RECT 114.555 133.745 114.725 133.915 ;
        RECT 115.015 133.745 115.185 133.915 ;
        RECT 115.475 133.745 115.645 133.915 ;
        RECT 115.935 133.745 116.105 133.915 ;
        RECT 116.395 133.745 116.565 133.915 ;
        RECT 116.855 133.745 117.025 133.915 ;
        RECT 117.315 133.745 117.485 133.915 ;
        RECT 117.775 133.745 117.945 133.915 ;
        RECT 118.235 133.745 118.405 133.915 ;
        RECT 118.695 133.745 118.865 133.915 ;
        RECT 119.155 133.745 119.325 133.915 ;
        RECT 119.615 133.745 119.785 133.915 ;
        RECT 120.075 133.745 120.245 133.915 ;
        RECT 120.535 133.745 120.705 133.915 ;
        RECT 120.995 133.745 121.165 133.915 ;
        RECT 121.455 133.745 121.625 133.915 ;
        RECT 121.915 133.745 122.085 133.915 ;
        RECT 122.375 133.745 122.545 133.915 ;
        RECT 122.835 133.745 123.005 133.915 ;
        RECT 123.295 133.745 123.465 133.915 ;
        RECT 123.755 133.745 123.925 133.915 ;
        RECT 124.215 133.745 124.385 133.915 ;
        RECT 124.675 133.745 124.845 133.915 ;
        RECT 125.135 133.745 125.305 133.915 ;
        RECT 125.595 133.745 125.765 133.915 ;
        RECT 126.055 133.745 126.225 133.915 ;
        RECT 126.515 133.745 126.685 133.915 ;
        RECT 126.975 133.745 127.145 133.915 ;
        RECT 127.435 133.745 127.605 133.915 ;
        RECT 127.895 133.745 128.065 133.915 ;
        RECT 128.355 133.745 128.525 133.915 ;
        RECT 128.815 133.745 128.985 133.915 ;
        RECT 129.275 133.745 129.445 133.915 ;
        RECT 129.735 133.745 129.905 133.915 ;
        RECT 130.195 133.745 130.365 133.915 ;
        RECT 130.655 133.745 130.825 133.915 ;
        RECT 131.115 133.745 131.285 133.915 ;
        RECT 131.575 133.745 131.745 133.915 ;
        RECT 132.035 133.745 132.205 133.915 ;
        RECT 132.495 133.745 132.665 133.915 ;
        RECT 132.955 133.745 133.125 133.915 ;
        RECT 133.415 133.745 133.585 133.915 ;
        RECT 133.875 133.745 134.045 133.915 ;
        RECT 134.335 133.745 134.505 133.915 ;
        RECT 134.795 133.745 134.965 133.915 ;
        RECT 135.255 133.745 135.425 133.915 ;
        RECT 135.715 133.745 135.885 133.915 ;
        RECT 136.175 133.745 136.345 133.915 ;
        RECT 136.635 133.745 136.805 133.915 ;
        RECT 137.095 133.745 137.265 133.915 ;
        RECT 137.555 133.745 137.725 133.915 ;
        RECT 138.015 133.745 138.185 133.915 ;
        RECT 138.475 133.745 138.645 133.915 ;
        RECT 138.935 133.745 139.105 133.915 ;
        RECT 139.395 133.745 139.565 133.915 ;
        RECT 139.855 133.745 140.025 133.915 ;
        RECT 140.315 133.745 140.485 133.915 ;
        RECT 140.775 133.745 140.945 133.915 ;
        RECT 141.235 133.745 141.405 133.915 ;
        RECT 141.695 133.745 141.865 133.915 ;
        RECT 142.155 133.745 142.325 133.915 ;
        RECT 142.615 133.745 142.785 133.915 ;
        RECT 143.075 133.745 143.245 133.915 ;
        RECT 143.535 133.745 143.705 133.915 ;
        RECT 143.995 133.745 144.165 133.915 ;
        RECT 144.455 133.745 144.625 133.915 ;
        RECT 144.915 133.745 145.085 133.915 ;
        RECT 145.375 133.745 145.545 133.915 ;
        RECT 145.835 133.745 146.005 133.915 ;
        RECT 146.295 133.745 146.465 133.915 ;
        RECT 146.755 133.745 146.925 133.915 ;
        RECT 147.215 133.745 147.385 133.915 ;
        RECT 147.675 133.745 147.845 133.915 ;
        RECT 148.135 133.745 148.305 133.915 ;
        RECT 148.595 133.745 148.765 133.915 ;
        RECT 149.055 133.745 149.225 133.915 ;
        RECT 149.515 133.745 149.685 133.915 ;
        RECT 149.975 133.745 150.145 133.915 ;
        RECT 150.435 133.745 150.605 133.915 ;
        RECT 150.895 133.745 151.065 133.915 ;
        RECT 151.355 133.745 151.525 133.915 ;
        RECT 151.815 133.745 151.985 133.915 ;
        RECT 152.275 133.745 152.445 133.915 ;
        RECT 152.735 133.745 152.905 133.915 ;
        RECT 153.195 133.745 153.365 133.915 ;
        RECT 153.655 133.745 153.825 133.915 ;
        RECT 154.115 133.745 154.285 133.915 ;
        RECT 154.575 133.745 154.745 133.915 ;
        RECT 155.035 133.745 155.205 133.915 ;
        RECT 155.495 133.745 155.665 133.915 ;
        RECT 155.955 133.745 156.125 133.915 ;
        RECT 73.155 132.555 73.325 132.725 ;
        RECT 73.615 132.215 73.785 132.385 ;
        RECT 74.995 131.875 75.165 132.045 ;
        RECT 83.735 132.895 83.905 133.065 ;
        RECT 84.195 133.235 84.365 133.405 ;
        RECT 83.275 132.555 83.445 132.725 ;
        RECT 85.115 132.555 85.285 132.725 ;
        RECT 88.335 132.555 88.505 132.725 ;
        RECT 89.255 132.555 89.425 132.725 ;
        RECT 97.075 133.235 97.245 133.405 ;
        RECT 84.655 131.535 84.825 131.705 ;
        RECT 88.335 131.535 88.505 131.705 ;
        RECT 97.995 132.555 98.165 132.725 ;
        RECT 98.915 132.555 99.085 132.725 ;
        RECT 100.755 132.555 100.925 132.725 ;
        RECT 99.835 131.875 100.005 132.045 ;
        RECT 105.355 132.895 105.525 133.065 ;
        RECT 106.275 132.895 106.445 133.065 ;
        RECT 104.435 131.535 104.605 131.705 ;
        RECT 113.175 132.555 113.345 132.725 ;
        RECT 113.635 132.555 113.805 132.725 ;
        RECT 114.555 132.555 114.725 132.725 ;
        RECT 115.015 132.555 115.185 132.725 ;
        RECT 112.255 131.535 112.425 131.705 ;
        RECT 123.755 133.235 123.925 133.405 ;
        RECT 123.295 132.895 123.465 133.065 ;
        RECT 124.675 132.555 124.845 132.725 ;
        RECT 125.595 131.535 125.765 131.705 ;
        RECT 130.150 132.555 130.320 132.725 ;
        RECT 130.655 132.555 130.825 132.725 ;
        RECT 129.275 131.875 129.445 132.045 ;
        RECT 132.035 132.555 132.205 132.725 ;
        RECT 131.575 131.535 131.745 131.705 ;
        RECT 132.955 131.875 133.125 132.045 ;
        RECT 139.395 132.555 139.565 132.725 ;
        RECT 138.475 131.535 138.645 131.705 ;
        RECT 139.855 132.215 140.025 132.385 ;
        RECT 140.270 132.555 140.440 132.725 ;
        RECT 140.775 132.555 140.945 132.725 ;
        RECT 141.695 132.555 141.865 132.725 ;
        RECT 142.615 132.555 142.785 132.725 ;
        RECT 143.535 132.555 143.705 132.725 ;
        RECT 142.155 132.215 142.325 132.385 ;
        RECT 144.455 132.555 144.625 132.725 ;
        RECT 144.915 132.555 145.085 132.725 ;
        RECT 145.835 132.555 146.005 132.725 ;
        RECT 146.295 132.555 146.465 132.725 ;
        RECT 144.455 131.535 144.625 131.705 ;
        RECT 145.375 132.215 145.545 132.385 ;
        RECT 148.595 132.895 148.765 133.065 ;
        RECT 149.595 133.235 149.765 133.405 ;
        RECT 147.215 131.535 147.385 131.705 ;
        RECT 149.515 131.535 149.685 131.705 ;
        RECT 150.435 131.535 150.605 131.705 ;
        RECT 153.655 133.235 153.825 133.405 ;
        RECT 152.275 132.555 152.445 132.725 ;
        RECT 153.195 132.895 153.365 133.065 ;
        RECT 153.655 132.555 153.825 132.725 ;
        RECT 154.575 132.555 154.745 132.725 ;
        RECT 151.355 131.535 151.525 131.705 ;
        RECT 70.855 131.025 71.025 131.195 ;
        RECT 71.315 131.025 71.485 131.195 ;
        RECT 71.775 131.025 71.945 131.195 ;
        RECT 72.235 131.025 72.405 131.195 ;
        RECT 72.695 131.025 72.865 131.195 ;
        RECT 73.155 131.025 73.325 131.195 ;
        RECT 73.615 131.025 73.785 131.195 ;
        RECT 74.075 131.025 74.245 131.195 ;
        RECT 74.535 131.025 74.705 131.195 ;
        RECT 74.995 131.025 75.165 131.195 ;
        RECT 75.455 131.025 75.625 131.195 ;
        RECT 75.915 131.025 76.085 131.195 ;
        RECT 76.375 131.025 76.545 131.195 ;
        RECT 76.835 131.025 77.005 131.195 ;
        RECT 77.295 131.025 77.465 131.195 ;
        RECT 77.755 131.025 77.925 131.195 ;
        RECT 78.215 131.025 78.385 131.195 ;
        RECT 78.675 131.025 78.845 131.195 ;
        RECT 79.135 131.025 79.305 131.195 ;
        RECT 79.595 131.025 79.765 131.195 ;
        RECT 80.055 131.025 80.225 131.195 ;
        RECT 80.515 131.025 80.685 131.195 ;
        RECT 80.975 131.025 81.145 131.195 ;
        RECT 81.435 131.025 81.605 131.195 ;
        RECT 81.895 131.025 82.065 131.195 ;
        RECT 82.355 131.025 82.525 131.195 ;
        RECT 82.815 131.025 82.985 131.195 ;
        RECT 83.275 131.025 83.445 131.195 ;
        RECT 83.735 131.025 83.905 131.195 ;
        RECT 84.195 131.025 84.365 131.195 ;
        RECT 84.655 131.025 84.825 131.195 ;
        RECT 85.115 131.025 85.285 131.195 ;
        RECT 85.575 131.025 85.745 131.195 ;
        RECT 86.035 131.025 86.205 131.195 ;
        RECT 86.495 131.025 86.665 131.195 ;
        RECT 86.955 131.025 87.125 131.195 ;
        RECT 87.415 131.025 87.585 131.195 ;
        RECT 87.875 131.025 88.045 131.195 ;
        RECT 88.335 131.025 88.505 131.195 ;
        RECT 88.795 131.025 88.965 131.195 ;
        RECT 89.255 131.025 89.425 131.195 ;
        RECT 89.715 131.025 89.885 131.195 ;
        RECT 90.175 131.025 90.345 131.195 ;
        RECT 90.635 131.025 90.805 131.195 ;
        RECT 91.095 131.025 91.265 131.195 ;
        RECT 91.555 131.025 91.725 131.195 ;
        RECT 92.015 131.025 92.185 131.195 ;
        RECT 92.475 131.025 92.645 131.195 ;
        RECT 92.935 131.025 93.105 131.195 ;
        RECT 93.395 131.025 93.565 131.195 ;
        RECT 93.855 131.025 94.025 131.195 ;
        RECT 94.315 131.025 94.485 131.195 ;
        RECT 94.775 131.025 94.945 131.195 ;
        RECT 95.235 131.025 95.405 131.195 ;
        RECT 95.695 131.025 95.865 131.195 ;
        RECT 96.155 131.025 96.325 131.195 ;
        RECT 96.615 131.025 96.785 131.195 ;
        RECT 97.075 131.025 97.245 131.195 ;
        RECT 97.535 131.025 97.705 131.195 ;
        RECT 97.995 131.025 98.165 131.195 ;
        RECT 98.455 131.025 98.625 131.195 ;
        RECT 98.915 131.025 99.085 131.195 ;
        RECT 99.375 131.025 99.545 131.195 ;
        RECT 99.835 131.025 100.005 131.195 ;
        RECT 100.295 131.025 100.465 131.195 ;
        RECT 100.755 131.025 100.925 131.195 ;
        RECT 101.215 131.025 101.385 131.195 ;
        RECT 101.675 131.025 101.845 131.195 ;
        RECT 102.135 131.025 102.305 131.195 ;
        RECT 102.595 131.025 102.765 131.195 ;
        RECT 103.055 131.025 103.225 131.195 ;
        RECT 103.515 131.025 103.685 131.195 ;
        RECT 103.975 131.025 104.145 131.195 ;
        RECT 104.435 131.025 104.605 131.195 ;
        RECT 104.895 131.025 105.065 131.195 ;
        RECT 105.355 131.025 105.525 131.195 ;
        RECT 105.815 131.025 105.985 131.195 ;
        RECT 106.275 131.025 106.445 131.195 ;
        RECT 106.735 131.025 106.905 131.195 ;
        RECT 107.195 131.025 107.365 131.195 ;
        RECT 107.655 131.025 107.825 131.195 ;
        RECT 108.115 131.025 108.285 131.195 ;
        RECT 108.575 131.025 108.745 131.195 ;
        RECT 109.035 131.025 109.205 131.195 ;
        RECT 109.495 131.025 109.665 131.195 ;
        RECT 109.955 131.025 110.125 131.195 ;
        RECT 110.415 131.025 110.585 131.195 ;
        RECT 110.875 131.025 111.045 131.195 ;
        RECT 111.335 131.025 111.505 131.195 ;
        RECT 111.795 131.025 111.965 131.195 ;
        RECT 112.255 131.025 112.425 131.195 ;
        RECT 112.715 131.025 112.885 131.195 ;
        RECT 113.175 131.025 113.345 131.195 ;
        RECT 113.635 131.025 113.805 131.195 ;
        RECT 114.095 131.025 114.265 131.195 ;
        RECT 114.555 131.025 114.725 131.195 ;
        RECT 115.015 131.025 115.185 131.195 ;
        RECT 115.475 131.025 115.645 131.195 ;
        RECT 115.935 131.025 116.105 131.195 ;
        RECT 116.395 131.025 116.565 131.195 ;
        RECT 116.855 131.025 117.025 131.195 ;
        RECT 117.315 131.025 117.485 131.195 ;
        RECT 117.775 131.025 117.945 131.195 ;
        RECT 118.235 131.025 118.405 131.195 ;
        RECT 118.695 131.025 118.865 131.195 ;
        RECT 119.155 131.025 119.325 131.195 ;
        RECT 119.615 131.025 119.785 131.195 ;
        RECT 120.075 131.025 120.245 131.195 ;
        RECT 120.535 131.025 120.705 131.195 ;
        RECT 120.995 131.025 121.165 131.195 ;
        RECT 121.455 131.025 121.625 131.195 ;
        RECT 121.915 131.025 122.085 131.195 ;
        RECT 122.375 131.025 122.545 131.195 ;
        RECT 122.835 131.025 123.005 131.195 ;
        RECT 123.295 131.025 123.465 131.195 ;
        RECT 123.755 131.025 123.925 131.195 ;
        RECT 124.215 131.025 124.385 131.195 ;
        RECT 124.675 131.025 124.845 131.195 ;
        RECT 125.135 131.025 125.305 131.195 ;
        RECT 125.595 131.025 125.765 131.195 ;
        RECT 126.055 131.025 126.225 131.195 ;
        RECT 126.515 131.025 126.685 131.195 ;
        RECT 126.975 131.025 127.145 131.195 ;
        RECT 127.435 131.025 127.605 131.195 ;
        RECT 127.895 131.025 128.065 131.195 ;
        RECT 128.355 131.025 128.525 131.195 ;
        RECT 128.815 131.025 128.985 131.195 ;
        RECT 129.275 131.025 129.445 131.195 ;
        RECT 129.735 131.025 129.905 131.195 ;
        RECT 130.195 131.025 130.365 131.195 ;
        RECT 130.655 131.025 130.825 131.195 ;
        RECT 131.115 131.025 131.285 131.195 ;
        RECT 131.575 131.025 131.745 131.195 ;
        RECT 132.035 131.025 132.205 131.195 ;
        RECT 132.495 131.025 132.665 131.195 ;
        RECT 132.955 131.025 133.125 131.195 ;
        RECT 133.415 131.025 133.585 131.195 ;
        RECT 133.875 131.025 134.045 131.195 ;
        RECT 134.335 131.025 134.505 131.195 ;
        RECT 134.795 131.025 134.965 131.195 ;
        RECT 135.255 131.025 135.425 131.195 ;
        RECT 135.715 131.025 135.885 131.195 ;
        RECT 136.175 131.025 136.345 131.195 ;
        RECT 136.635 131.025 136.805 131.195 ;
        RECT 137.095 131.025 137.265 131.195 ;
        RECT 137.555 131.025 137.725 131.195 ;
        RECT 138.015 131.025 138.185 131.195 ;
        RECT 138.475 131.025 138.645 131.195 ;
        RECT 138.935 131.025 139.105 131.195 ;
        RECT 139.395 131.025 139.565 131.195 ;
        RECT 139.855 131.025 140.025 131.195 ;
        RECT 140.315 131.025 140.485 131.195 ;
        RECT 140.775 131.025 140.945 131.195 ;
        RECT 141.235 131.025 141.405 131.195 ;
        RECT 141.695 131.025 141.865 131.195 ;
        RECT 142.155 131.025 142.325 131.195 ;
        RECT 142.615 131.025 142.785 131.195 ;
        RECT 143.075 131.025 143.245 131.195 ;
        RECT 143.535 131.025 143.705 131.195 ;
        RECT 143.995 131.025 144.165 131.195 ;
        RECT 144.455 131.025 144.625 131.195 ;
        RECT 144.915 131.025 145.085 131.195 ;
        RECT 145.375 131.025 145.545 131.195 ;
        RECT 145.835 131.025 146.005 131.195 ;
        RECT 146.295 131.025 146.465 131.195 ;
        RECT 146.755 131.025 146.925 131.195 ;
        RECT 147.215 131.025 147.385 131.195 ;
        RECT 147.675 131.025 147.845 131.195 ;
        RECT 148.135 131.025 148.305 131.195 ;
        RECT 148.595 131.025 148.765 131.195 ;
        RECT 149.055 131.025 149.225 131.195 ;
        RECT 149.515 131.025 149.685 131.195 ;
        RECT 149.975 131.025 150.145 131.195 ;
        RECT 150.435 131.025 150.605 131.195 ;
        RECT 150.895 131.025 151.065 131.195 ;
        RECT 151.355 131.025 151.525 131.195 ;
        RECT 151.815 131.025 151.985 131.195 ;
        RECT 152.275 131.025 152.445 131.195 ;
        RECT 152.735 131.025 152.905 131.195 ;
        RECT 153.195 131.025 153.365 131.195 ;
        RECT 153.655 131.025 153.825 131.195 ;
        RECT 154.115 131.025 154.285 131.195 ;
        RECT 154.575 131.025 154.745 131.195 ;
        RECT 155.035 131.025 155.205 131.195 ;
        RECT 155.495 131.025 155.665 131.195 ;
        RECT 155.955 131.025 156.125 131.195 ;
        RECT 75.455 129.835 75.625 130.005 ;
        RECT 74.995 129.495 75.165 129.665 ;
        RECT 77.755 129.495 77.925 129.665 ;
        RECT 78.675 129.495 78.845 129.665 ;
        RECT 79.135 129.495 79.305 129.665 ;
        RECT 80.515 129.495 80.685 129.665 ;
        RECT 76.835 128.815 77.005 128.985 ;
        RECT 78.675 128.815 78.845 128.985 ;
        RECT 79.595 128.815 79.765 128.985 ;
        RECT 81.895 129.495 82.065 129.665 ;
        RECT 85.115 130.515 85.285 130.685 ;
        RECT 86.035 130.175 86.205 130.345 ;
        RECT 82.815 129.495 82.985 129.665 ;
        RECT 81.435 128.815 81.605 128.985 ;
        RECT 82.815 128.815 82.985 128.985 ;
        RECT 84.195 129.155 84.365 129.325 ;
        RECT 85.345 129.325 85.515 129.495 ;
        RECT 86.495 129.495 86.665 129.665 ;
        RECT 86.955 129.495 87.125 129.665 ;
        RECT 87.875 129.495 88.045 129.665 ;
        RECT 88.335 129.495 88.505 129.665 ;
        RECT 89.715 129.835 89.885 130.005 ;
        RECT 89.255 128.815 89.425 128.985 ;
        RECT 90.635 128.815 90.805 128.985 ;
        RECT 91.095 129.495 91.265 129.665 ;
        RECT 91.555 129.495 91.725 129.665 ;
        RECT 92.475 128.815 92.645 128.985 ;
        RECT 92.935 129.495 93.105 129.665 ;
        RECT 94.315 130.175 94.485 130.345 ;
        RECT 93.855 129.495 94.025 129.665 ;
        RECT 94.775 130.175 94.945 130.345 ;
        RECT 95.235 129.495 95.405 129.665 ;
        RECT 98.455 130.515 98.625 130.685 ;
        RECT 99.375 129.495 99.545 129.665 ;
        RECT 99.835 129.495 100.005 129.665 ;
        RECT 100.295 130.175 100.465 130.345 ;
        RECT 100.755 129.495 100.925 129.665 ;
        RECT 102.135 129.495 102.305 129.665 ;
        RECT 102.595 129.835 102.765 130.005 ;
        RECT 103.055 129.495 103.225 129.665 ;
        RECT 103.515 129.835 103.685 130.005 ;
        RECT 104.895 129.835 105.065 130.005 ;
        RECT 106.275 129.495 106.445 129.665 ;
        RECT 109.955 129.495 110.125 129.665 ;
        RECT 104.435 128.815 104.605 128.985 ;
        RECT 110.875 128.815 111.045 128.985 ;
        RECT 113.635 130.175 113.805 130.345 ;
        RECT 111.335 129.495 111.505 129.665 ;
        RECT 112.255 129.495 112.425 129.665 ;
        RECT 113.175 129.495 113.345 129.665 ;
        RECT 115.935 129.835 116.105 130.005 ;
        RECT 114.555 129.495 114.725 129.665 ;
        RECT 115.475 129.495 115.645 129.665 ;
        RECT 116.395 129.495 116.565 129.665 ;
        RECT 116.855 129.495 117.025 129.665 ;
        RECT 117.775 129.495 117.945 129.665 ;
        RECT 118.695 128.815 118.865 128.985 ;
        RECT 120.535 130.175 120.705 130.345 ;
        RECT 120.075 129.495 120.245 129.665 ;
        RECT 119.155 128.815 119.325 128.985 ;
        RECT 121.915 130.515 122.085 130.685 ;
        RECT 121.455 129.495 121.625 129.665 ;
        RECT 123.755 130.175 123.925 130.345 ;
        RECT 122.835 129.495 123.005 129.665 ;
        RECT 124.675 129.495 124.845 129.665 ;
        RECT 127.895 129.835 128.065 130.005 ;
        RECT 130.655 130.175 130.825 130.345 ;
        RECT 129.275 129.835 129.445 130.005 ;
        RECT 129.735 129.495 129.905 129.665 ;
        RECT 132.495 129.495 132.665 129.665 ;
        RECT 132.955 129.495 133.125 129.665 ;
        RECT 133.415 129.495 133.585 129.665 ;
        RECT 131.115 128.815 131.285 128.985 ;
        RECT 134.335 129.495 134.505 129.665 ;
        RECT 136.175 129.835 136.345 130.005 ;
        RECT 136.635 129.835 136.805 130.005 ;
        RECT 137.095 129.495 137.265 129.665 ;
        RECT 137.555 129.835 137.725 130.005 ;
        RECT 138.475 130.175 138.645 130.345 ;
        RECT 141.235 130.175 141.405 130.345 ;
        RECT 139.855 129.495 140.025 129.665 ;
        RECT 140.315 129.495 140.485 129.665 ;
        RECT 139.395 128.815 139.565 128.985 ;
        RECT 141.235 129.495 141.405 129.665 ;
        RECT 145.375 130.515 145.545 130.685 ;
        RECT 143.535 129.835 143.705 130.005 ;
        RECT 143.075 129.495 143.245 129.665 ;
        RECT 144.455 129.495 144.625 129.665 ;
        RECT 142.155 128.815 142.325 128.985 ;
        RECT 152.735 130.515 152.905 130.685 ;
        RECT 147.215 129.495 147.385 129.665 ;
        RECT 146.295 128.815 146.465 128.985 ;
        RECT 147.675 129.155 147.845 129.325 ;
        RECT 148.595 129.495 148.765 129.665 ;
        RECT 149.515 129.495 149.685 129.665 ;
        RECT 148.135 129.155 148.305 129.325 ;
        RECT 150.895 129.495 151.065 129.665 ;
        RECT 153.655 130.515 153.825 130.685 ;
        RECT 151.355 129.495 151.525 129.665 ;
        RECT 149.975 128.815 150.145 128.985 ;
        RECT 153.195 129.495 153.365 129.665 ;
        RECT 153.655 129.495 153.825 129.665 ;
        RECT 154.545 129.495 154.715 129.665 ;
        RECT 70.855 128.305 71.025 128.475 ;
        RECT 71.315 128.305 71.485 128.475 ;
        RECT 71.775 128.305 71.945 128.475 ;
        RECT 72.235 128.305 72.405 128.475 ;
        RECT 72.695 128.305 72.865 128.475 ;
        RECT 73.155 128.305 73.325 128.475 ;
        RECT 73.615 128.305 73.785 128.475 ;
        RECT 74.075 128.305 74.245 128.475 ;
        RECT 74.535 128.305 74.705 128.475 ;
        RECT 74.995 128.305 75.165 128.475 ;
        RECT 75.455 128.305 75.625 128.475 ;
        RECT 75.915 128.305 76.085 128.475 ;
        RECT 76.375 128.305 76.545 128.475 ;
        RECT 76.835 128.305 77.005 128.475 ;
        RECT 77.295 128.305 77.465 128.475 ;
        RECT 77.755 128.305 77.925 128.475 ;
        RECT 78.215 128.305 78.385 128.475 ;
        RECT 78.675 128.305 78.845 128.475 ;
        RECT 79.135 128.305 79.305 128.475 ;
        RECT 79.595 128.305 79.765 128.475 ;
        RECT 80.055 128.305 80.225 128.475 ;
        RECT 80.515 128.305 80.685 128.475 ;
        RECT 80.975 128.305 81.145 128.475 ;
        RECT 81.435 128.305 81.605 128.475 ;
        RECT 81.895 128.305 82.065 128.475 ;
        RECT 82.355 128.305 82.525 128.475 ;
        RECT 82.815 128.305 82.985 128.475 ;
        RECT 83.275 128.305 83.445 128.475 ;
        RECT 83.735 128.305 83.905 128.475 ;
        RECT 84.195 128.305 84.365 128.475 ;
        RECT 84.655 128.305 84.825 128.475 ;
        RECT 85.115 128.305 85.285 128.475 ;
        RECT 85.575 128.305 85.745 128.475 ;
        RECT 86.035 128.305 86.205 128.475 ;
        RECT 86.495 128.305 86.665 128.475 ;
        RECT 86.955 128.305 87.125 128.475 ;
        RECT 87.415 128.305 87.585 128.475 ;
        RECT 87.875 128.305 88.045 128.475 ;
        RECT 88.335 128.305 88.505 128.475 ;
        RECT 88.795 128.305 88.965 128.475 ;
        RECT 89.255 128.305 89.425 128.475 ;
        RECT 89.715 128.305 89.885 128.475 ;
        RECT 90.175 128.305 90.345 128.475 ;
        RECT 90.635 128.305 90.805 128.475 ;
        RECT 91.095 128.305 91.265 128.475 ;
        RECT 91.555 128.305 91.725 128.475 ;
        RECT 92.015 128.305 92.185 128.475 ;
        RECT 92.475 128.305 92.645 128.475 ;
        RECT 92.935 128.305 93.105 128.475 ;
        RECT 93.395 128.305 93.565 128.475 ;
        RECT 93.855 128.305 94.025 128.475 ;
        RECT 94.315 128.305 94.485 128.475 ;
        RECT 94.775 128.305 94.945 128.475 ;
        RECT 95.235 128.305 95.405 128.475 ;
        RECT 95.695 128.305 95.865 128.475 ;
        RECT 96.155 128.305 96.325 128.475 ;
        RECT 96.615 128.305 96.785 128.475 ;
        RECT 97.075 128.305 97.245 128.475 ;
        RECT 97.535 128.305 97.705 128.475 ;
        RECT 97.995 128.305 98.165 128.475 ;
        RECT 98.455 128.305 98.625 128.475 ;
        RECT 98.915 128.305 99.085 128.475 ;
        RECT 99.375 128.305 99.545 128.475 ;
        RECT 99.835 128.305 100.005 128.475 ;
        RECT 100.295 128.305 100.465 128.475 ;
        RECT 100.755 128.305 100.925 128.475 ;
        RECT 101.215 128.305 101.385 128.475 ;
        RECT 101.675 128.305 101.845 128.475 ;
        RECT 102.135 128.305 102.305 128.475 ;
        RECT 102.595 128.305 102.765 128.475 ;
        RECT 103.055 128.305 103.225 128.475 ;
        RECT 103.515 128.305 103.685 128.475 ;
        RECT 103.975 128.305 104.145 128.475 ;
        RECT 104.435 128.305 104.605 128.475 ;
        RECT 104.895 128.305 105.065 128.475 ;
        RECT 105.355 128.305 105.525 128.475 ;
        RECT 105.815 128.305 105.985 128.475 ;
        RECT 106.275 128.305 106.445 128.475 ;
        RECT 106.735 128.305 106.905 128.475 ;
        RECT 107.195 128.305 107.365 128.475 ;
        RECT 107.655 128.305 107.825 128.475 ;
        RECT 108.115 128.305 108.285 128.475 ;
        RECT 108.575 128.305 108.745 128.475 ;
        RECT 109.035 128.305 109.205 128.475 ;
        RECT 109.495 128.305 109.665 128.475 ;
        RECT 109.955 128.305 110.125 128.475 ;
        RECT 110.415 128.305 110.585 128.475 ;
        RECT 110.875 128.305 111.045 128.475 ;
        RECT 111.335 128.305 111.505 128.475 ;
        RECT 111.795 128.305 111.965 128.475 ;
        RECT 112.255 128.305 112.425 128.475 ;
        RECT 112.715 128.305 112.885 128.475 ;
        RECT 113.175 128.305 113.345 128.475 ;
        RECT 113.635 128.305 113.805 128.475 ;
        RECT 114.095 128.305 114.265 128.475 ;
        RECT 114.555 128.305 114.725 128.475 ;
        RECT 115.015 128.305 115.185 128.475 ;
        RECT 115.475 128.305 115.645 128.475 ;
        RECT 115.935 128.305 116.105 128.475 ;
        RECT 116.395 128.305 116.565 128.475 ;
        RECT 116.855 128.305 117.025 128.475 ;
        RECT 117.315 128.305 117.485 128.475 ;
        RECT 117.775 128.305 117.945 128.475 ;
        RECT 118.235 128.305 118.405 128.475 ;
        RECT 118.695 128.305 118.865 128.475 ;
        RECT 119.155 128.305 119.325 128.475 ;
        RECT 119.615 128.305 119.785 128.475 ;
        RECT 120.075 128.305 120.245 128.475 ;
        RECT 120.535 128.305 120.705 128.475 ;
        RECT 120.995 128.305 121.165 128.475 ;
        RECT 121.455 128.305 121.625 128.475 ;
        RECT 121.915 128.305 122.085 128.475 ;
        RECT 122.375 128.305 122.545 128.475 ;
        RECT 122.835 128.305 123.005 128.475 ;
        RECT 123.295 128.305 123.465 128.475 ;
        RECT 123.755 128.305 123.925 128.475 ;
        RECT 124.215 128.305 124.385 128.475 ;
        RECT 124.675 128.305 124.845 128.475 ;
        RECT 125.135 128.305 125.305 128.475 ;
        RECT 125.595 128.305 125.765 128.475 ;
        RECT 126.055 128.305 126.225 128.475 ;
        RECT 126.515 128.305 126.685 128.475 ;
        RECT 126.975 128.305 127.145 128.475 ;
        RECT 127.435 128.305 127.605 128.475 ;
        RECT 127.895 128.305 128.065 128.475 ;
        RECT 128.355 128.305 128.525 128.475 ;
        RECT 128.815 128.305 128.985 128.475 ;
        RECT 129.275 128.305 129.445 128.475 ;
        RECT 129.735 128.305 129.905 128.475 ;
        RECT 130.195 128.305 130.365 128.475 ;
        RECT 130.655 128.305 130.825 128.475 ;
        RECT 131.115 128.305 131.285 128.475 ;
        RECT 131.575 128.305 131.745 128.475 ;
        RECT 132.035 128.305 132.205 128.475 ;
        RECT 132.495 128.305 132.665 128.475 ;
        RECT 132.955 128.305 133.125 128.475 ;
        RECT 133.415 128.305 133.585 128.475 ;
        RECT 133.875 128.305 134.045 128.475 ;
        RECT 134.335 128.305 134.505 128.475 ;
        RECT 134.795 128.305 134.965 128.475 ;
        RECT 135.255 128.305 135.425 128.475 ;
        RECT 135.715 128.305 135.885 128.475 ;
        RECT 136.175 128.305 136.345 128.475 ;
        RECT 136.635 128.305 136.805 128.475 ;
        RECT 137.095 128.305 137.265 128.475 ;
        RECT 137.555 128.305 137.725 128.475 ;
        RECT 138.015 128.305 138.185 128.475 ;
        RECT 138.475 128.305 138.645 128.475 ;
        RECT 138.935 128.305 139.105 128.475 ;
        RECT 139.395 128.305 139.565 128.475 ;
        RECT 139.855 128.305 140.025 128.475 ;
        RECT 140.315 128.305 140.485 128.475 ;
        RECT 140.775 128.305 140.945 128.475 ;
        RECT 141.235 128.305 141.405 128.475 ;
        RECT 141.695 128.305 141.865 128.475 ;
        RECT 142.155 128.305 142.325 128.475 ;
        RECT 142.615 128.305 142.785 128.475 ;
        RECT 143.075 128.305 143.245 128.475 ;
        RECT 143.535 128.305 143.705 128.475 ;
        RECT 143.995 128.305 144.165 128.475 ;
        RECT 144.455 128.305 144.625 128.475 ;
        RECT 144.915 128.305 145.085 128.475 ;
        RECT 145.375 128.305 145.545 128.475 ;
        RECT 145.835 128.305 146.005 128.475 ;
        RECT 146.295 128.305 146.465 128.475 ;
        RECT 146.755 128.305 146.925 128.475 ;
        RECT 147.215 128.305 147.385 128.475 ;
        RECT 147.675 128.305 147.845 128.475 ;
        RECT 148.135 128.305 148.305 128.475 ;
        RECT 148.595 128.305 148.765 128.475 ;
        RECT 149.055 128.305 149.225 128.475 ;
        RECT 149.515 128.305 149.685 128.475 ;
        RECT 149.975 128.305 150.145 128.475 ;
        RECT 150.435 128.305 150.605 128.475 ;
        RECT 150.895 128.305 151.065 128.475 ;
        RECT 151.355 128.305 151.525 128.475 ;
        RECT 151.815 128.305 151.985 128.475 ;
        RECT 152.275 128.305 152.445 128.475 ;
        RECT 152.735 128.305 152.905 128.475 ;
        RECT 153.195 128.305 153.365 128.475 ;
        RECT 153.655 128.305 153.825 128.475 ;
        RECT 154.115 128.305 154.285 128.475 ;
        RECT 154.575 128.305 154.745 128.475 ;
        RECT 155.035 128.305 155.205 128.475 ;
        RECT 155.495 128.305 155.665 128.475 ;
        RECT 155.955 128.305 156.125 128.475 ;
        RECT 74.535 127.115 74.705 127.285 ;
        RECT 73.615 126.095 73.785 126.265 ;
        RECT 80.055 127.795 80.225 127.965 ;
        RECT 76.375 127.115 76.545 127.285 ;
        RECT 78.215 127.115 78.385 127.285 ;
        RECT 79.135 127.455 79.305 127.625 ;
        RECT 75.455 126.095 75.625 126.265 ;
        RECT 80.975 127.455 81.145 127.625 ;
        RECT 82.815 127.795 82.985 127.965 ;
        RECT 86.495 127.795 86.665 127.965 ;
        RECT 81.975 127.455 82.145 127.625 ;
        RECT 81.895 126.095 82.065 126.265 ;
        RECT 84.195 127.115 84.365 127.285 ;
        RECT 84.655 127.115 84.825 127.285 ;
        RECT 85.115 126.775 85.285 126.945 ;
        RECT 85.575 126.775 85.745 126.945 ;
        RECT 86.955 127.455 87.125 127.625 ;
        RECT 87.875 127.115 88.045 127.285 ;
        RECT 88.335 127.115 88.505 127.285 ;
        RECT 88.795 127.115 88.965 127.285 ;
        RECT 89.715 127.115 89.885 127.285 ;
        RECT 87.415 126.435 87.585 126.605 ;
        RECT 89.255 126.095 89.425 126.265 ;
        RECT 92.015 127.115 92.185 127.285 ;
        RECT 91.555 126.775 91.725 126.945 ;
        RECT 93.855 126.775 94.025 126.945 ;
        RECT 95.695 127.115 95.865 127.285 ;
        RECT 94.775 126.095 94.945 126.265 ;
        RECT 97.995 127.115 98.165 127.285 ;
        RECT 97.075 126.095 97.245 126.265 ;
        RECT 98.455 126.775 98.625 126.945 ;
        RECT 99.375 127.115 99.545 127.285 ;
        RECT 98.915 126.775 99.085 126.945 ;
        RECT 100.295 127.115 100.465 127.285 ;
        RECT 101.215 126.095 101.385 126.265 ;
        RECT 103.055 127.795 103.225 127.965 ;
        RECT 102.595 127.115 102.765 127.285 ;
        RECT 103.055 127.115 103.225 127.285 ;
        RECT 103.975 127.115 104.145 127.285 ;
        RECT 101.675 126.095 101.845 126.265 ;
        RECT 104.435 126.775 104.605 126.945 ;
        RECT 105.355 127.115 105.525 127.285 ;
        RECT 106.275 127.115 106.445 127.285 ;
        RECT 108.575 127.115 108.745 127.285 ;
        RECT 107.195 126.775 107.365 126.945 ;
        RECT 109.495 126.775 109.665 126.945 ;
        RECT 113.175 127.115 113.345 127.285 ;
        RECT 114.095 127.115 114.265 127.285 ;
        RECT 112.255 126.435 112.425 126.605 ;
        RECT 116.395 127.115 116.565 127.285 ;
        RECT 116.855 127.115 117.025 127.285 ;
        RECT 117.315 127.115 117.485 127.285 ;
        RECT 118.235 127.115 118.405 127.285 ;
        RECT 115.015 126.095 115.185 126.265 ;
        RECT 119.615 127.115 119.785 127.285 ;
        RECT 118.695 126.435 118.865 126.605 ;
        RECT 120.075 126.435 120.245 126.605 ;
        RECT 120.995 127.115 121.165 127.285 ;
        RECT 120.535 126.775 120.705 126.945 ;
        RECT 124.215 127.115 124.385 127.285 ;
        RECT 122.835 126.775 123.005 126.945 ;
        RECT 123.295 126.095 123.465 126.265 ;
        RECT 127.435 127.455 127.605 127.625 ;
        RECT 125.135 126.095 125.305 126.265 ;
        RECT 129.735 127.115 129.905 127.285 ;
        RECT 128.355 126.775 128.525 126.945 ;
        RECT 126.055 126.095 126.225 126.265 ;
        RECT 128.815 126.095 128.985 126.265 ;
        RECT 130.655 126.095 130.825 126.265 ;
        RECT 131.115 127.795 131.285 127.965 ;
        RECT 133.875 127.455 134.045 127.625 ;
        RECT 132.035 127.115 132.205 127.285 ;
        RECT 132.955 127.115 133.125 127.285 ;
        RECT 134.795 127.115 134.965 127.285 ;
        RECT 135.715 127.115 135.885 127.285 ;
        RECT 137.555 127.115 137.725 127.285 ;
        RECT 138.475 127.115 138.645 127.285 ;
        RECT 136.635 126.435 136.805 126.605 ;
        RECT 140.775 127.115 140.945 127.285 ;
        RECT 139.395 126.775 139.565 126.945 ;
        RECT 143.075 127.795 143.245 127.965 ;
        RECT 142.155 127.115 142.325 127.285 ;
        RECT 141.695 126.435 141.865 126.605 ;
        RECT 146.755 127.795 146.925 127.965 ;
        RECT 144.915 127.115 145.085 127.285 ;
        RECT 144.455 126.775 144.625 126.945 ;
        RECT 149.055 127.455 149.225 127.625 ;
        RECT 152.275 127.455 152.445 127.625 ;
        RECT 151.355 126.775 151.525 126.945 ;
        RECT 149.515 126.095 149.685 126.265 ;
        RECT 153.195 127.115 153.365 127.285 ;
        RECT 70.855 125.585 71.025 125.755 ;
        RECT 71.315 125.585 71.485 125.755 ;
        RECT 71.775 125.585 71.945 125.755 ;
        RECT 72.235 125.585 72.405 125.755 ;
        RECT 72.695 125.585 72.865 125.755 ;
        RECT 73.155 125.585 73.325 125.755 ;
        RECT 73.615 125.585 73.785 125.755 ;
        RECT 74.075 125.585 74.245 125.755 ;
        RECT 74.535 125.585 74.705 125.755 ;
        RECT 74.995 125.585 75.165 125.755 ;
        RECT 75.455 125.585 75.625 125.755 ;
        RECT 75.915 125.585 76.085 125.755 ;
        RECT 76.375 125.585 76.545 125.755 ;
        RECT 76.835 125.585 77.005 125.755 ;
        RECT 77.295 125.585 77.465 125.755 ;
        RECT 77.755 125.585 77.925 125.755 ;
        RECT 78.215 125.585 78.385 125.755 ;
        RECT 78.675 125.585 78.845 125.755 ;
        RECT 79.135 125.585 79.305 125.755 ;
        RECT 79.595 125.585 79.765 125.755 ;
        RECT 80.055 125.585 80.225 125.755 ;
        RECT 80.515 125.585 80.685 125.755 ;
        RECT 80.975 125.585 81.145 125.755 ;
        RECT 81.435 125.585 81.605 125.755 ;
        RECT 81.895 125.585 82.065 125.755 ;
        RECT 82.355 125.585 82.525 125.755 ;
        RECT 82.815 125.585 82.985 125.755 ;
        RECT 83.275 125.585 83.445 125.755 ;
        RECT 83.735 125.585 83.905 125.755 ;
        RECT 84.195 125.585 84.365 125.755 ;
        RECT 84.655 125.585 84.825 125.755 ;
        RECT 85.115 125.585 85.285 125.755 ;
        RECT 85.575 125.585 85.745 125.755 ;
        RECT 86.035 125.585 86.205 125.755 ;
        RECT 86.495 125.585 86.665 125.755 ;
        RECT 86.955 125.585 87.125 125.755 ;
        RECT 87.415 125.585 87.585 125.755 ;
        RECT 87.875 125.585 88.045 125.755 ;
        RECT 88.335 125.585 88.505 125.755 ;
        RECT 88.795 125.585 88.965 125.755 ;
        RECT 89.255 125.585 89.425 125.755 ;
        RECT 89.715 125.585 89.885 125.755 ;
        RECT 90.175 125.585 90.345 125.755 ;
        RECT 90.635 125.585 90.805 125.755 ;
        RECT 91.095 125.585 91.265 125.755 ;
        RECT 91.555 125.585 91.725 125.755 ;
        RECT 92.015 125.585 92.185 125.755 ;
        RECT 92.475 125.585 92.645 125.755 ;
        RECT 92.935 125.585 93.105 125.755 ;
        RECT 93.395 125.585 93.565 125.755 ;
        RECT 93.855 125.585 94.025 125.755 ;
        RECT 94.315 125.585 94.485 125.755 ;
        RECT 94.775 125.585 94.945 125.755 ;
        RECT 95.235 125.585 95.405 125.755 ;
        RECT 95.695 125.585 95.865 125.755 ;
        RECT 96.155 125.585 96.325 125.755 ;
        RECT 96.615 125.585 96.785 125.755 ;
        RECT 97.075 125.585 97.245 125.755 ;
        RECT 97.535 125.585 97.705 125.755 ;
        RECT 97.995 125.585 98.165 125.755 ;
        RECT 98.455 125.585 98.625 125.755 ;
        RECT 98.915 125.585 99.085 125.755 ;
        RECT 99.375 125.585 99.545 125.755 ;
        RECT 99.835 125.585 100.005 125.755 ;
        RECT 100.295 125.585 100.465 125.755 ;
        RECT 100.755 125.585 100.925 125.755 ;
        RECT 101.215 125.585 101.385 125.755 ;
        RECT 101.675 125.585 101.845 125.755 ;
        RECT 102.135 125.585 102.305 125.755 ;
        RECT 102.595 125.585 102.765 125.755 ;
        RECT 103.055 125.585 103.225 125.755 ;
        RECT 103.515 125.585 103.685 125.755 ;
        RECT 103.975 125.585 104.145 125.755 ;
        RECT 104.435 125.585 104.605 125.755 ;
        RECT 104.895 125.585 105.065 125.755 ;
        RECT 105.355 125.585 105.525 125.755 ;
        RECT 105.815 125.585 105.985 125.755 ;
        RECT 106.275 125.585 106.445 125.755 ;
        RECT 106.735 125.585 106.905 125.755 ;
        RECT 107.195 125.585 107.365 125.755 ;
        RECT 107.655 125.585 107.825 125.755 ;
        RECT 108.115 125.585 108.285 125.755 ;
        RECT 108.575 125.585 108.745 125.755 ;
        RECT 109.035 125.585 109.205 125.755 ;
        RECT 109.495 125.585 109.665 125.755 ;
        RECT 109.955 125.585 110.125 125.755 ;
        RECT 110.415 125.585 110.585 125.755 ;
        RECT 110.875 125.585 111.045 125.755 ;
        RECT 111.335 125.585 111.505 125.755 ;
        RECT 111.795 125.585 111.965 125.755 ;
        RECT 112.255 125.585 112.425 125.755 ;
        RECT 112.715 125.585 112.885 125.755 ;
        RECT 113.175 125.585 113.345 125.755 ;
        RECT 113.635 125.585 113.805 125.755 ;
        RECT 114.095 125.585 114.265 125.755 ;
        RECT 114.555 125.585 114.725 125.755 ;
        RECT 115.015 125.585 115.185 125.755 ;
        RECT 115.475 125.585 115.645 125.755 ;
        RECT 115.935 125.585 116.105 125.755 ;
        RECT 116.395 125.585 116.565 125.755 ;
        RECT 116.855 125.585 117.025 125.755 ;
        RECT 117.315 125.585 117.485 125.755 ;
        RECT 117.775 125.585 117.945 125.755 ;
        RECT 118.235 125.585 118.405 125.755 ;
        RECT 118.695 125.585 118.865 125.755 ;
        RECT 119.155 125.585 119.325 125.755 ;
        RECT 119.615 125.585 119.785 125.755 ;
        RECT 120.075 125.585 120.245 125.755 ;
        RECT 120.535 125.585 120.705 125.755 ;
        RECT 120.995 125.585 121.165 125.755 ;
        RECT 121.455 125.585 121.625 125.755 ;
        RECT 121.915 125.585 122.085 125.755 ;
        RECT 122.375 125.585 122.545 125.755 ;
        RECT 122.835 125.585 123.005 125.755 ;
        RECT 123.295 125.585 123.465 125.755 ;
        RECT 123.755 125.585 123.925 125.755 ;
        RECT 124.215 125.585 124.385 125.755 ;
        RECT 124.675 125.585 124.845 125.755 ;
        RECT 125.135 125.585 125.305 125.755 ;
        RECT 125.595 125.585 125.765 125.755 ;
        RECT 126.055 125.585 126.225 125.755 ;
        RECT 126.515 125.585 126.685 125.755 ;
        RECT 126.975 125.585 127.145 125.755 ;
        RECT 127.435 125.585 127.605 125.755 ;
        RECT 127.895 125.585 128.065 125.755 ;
        RECT 128.355 125.585 128.525 125.755 ;
        RECT 128.815 125.585 128.985 125.755 ;
        RECT 129.275 125.585 129.445 125.755 ;
        RECT 129.735 125.585 129.905 125.755 ;
        RECT 130.195 125.585 130.365 125.755 ;
        RECT 130.655 125.585 130.825 125.755 ;
        RECT 131.115 125.585 131.285 125.755 ;
        RECT 131.575 125.585 131.745 125.755 ;
        RECT 132.035 125.585 132.205 125.755 ;
        RECT 132.495 125.585 132.665 125.755 ;
        RECT 132.955 125.585 133.125 125.755 ;
        RECT 133.415 125.585 133.585 125.755 ;
        RECT 133.875 125.585 134.045 125.755 ;
        RECT 134.335 125.585 134.505 125.755 ;
        RECT 134.795 125.585 134.965 125.755 ;
        RECT 135.255 125.585 135.425 125.755 ;
        RECT 135.715 125.585 135.885 125.755 ;
        RECT 136.175 125.585 136.345 125.755 ;
        RECT 136.635 125.585 136.805 125.755 ;
        RECT 137.095 125.585 137.265 125.755 ;
        RECT 137.555 125.585 137.725 125.755 ;
        RECT 138.015 125.585 138.185 125.755 ;
        RECT 138.475 125.585 138.645 125.755 ;
        RECT 138.935 125.585 139.105 125.755 ;
        RECT 139.395 125.585 139.565 125.755 ;
        RECT 139.855 125.585 140.025 125.755 ;
        RECT 140.315 125.585 140.485 125.755 ;
        RECT 140.775 125.585 140.945 125.755 ;
        RECT 141.235 125.585 141.405 125.755 ;
        RECT 141.695 125.585 141.865 125.755 ;
        RECT 142.155 125.585 142.325 125.755 ;
        RECT 142.615 125.585 142.785 125.755 ;
        RECT 143.075 125.585 143.245 125.755 ;
        RECT 143.535 125.585 143.705 125.755 ;
        RECT 143.995 125.585 144.165 125.755 ;
        RECT 144.455 125.585 144.625 125.755 ;
        RECT 144.915 125.585 145.085 125.755 ;
        RECT 145.375 125.585 145.545 125.755 ;
        RECT 145.835 125.585 146.005 125.755 ;
        RECT 146.295 125.585 146.465 125.755 ;
        RECT 146.755 125.585 146.925 125.755 ;
        RECT 147.215 125.585 147.385 125.755 ;
        RECT 147.675 125.585 147.845 125.755 ;
        RECT 148.135 125.585 148.305 125.755 ;
        RECT 148.595 125.585 148.765 125.755 ;
        RECT 149.055 125.585 149.225 125.755 ;
        RECT 149.515 125.585 149.685 125.755 ;
        RECT 149.975 125.585 150.145 125.755 ;
        RECT 150.435 125.585 150.605 125.755 ;
        RECT 150.895 125.585 151.065 125.755 ;
        RECT 151.355 125.585 151.525 125.755 ;
        RECT 151.815 125.585 151.985 125.755 ;
        RECT 152.275 125.585 152.445 125.755 ;
        RECT 152.735 125.585 152.905 125.755 ;
        RECT 153.195 125.585 153.365 125.755 ;
        RECT 153.655 125.585 153.825 125.755 ;
        RECT 154.115 125.585 154.285 125.755 ;
        RECT 154.575 125.585 154.745 125.755 ;
        RECT 155.035 125.585 155.205 125.755 ;
        RECT 155.495 125.585 155.665 125.755 ;
        RECT 155.955 125.585 156.125 125.755 ;
        RECT 73.615 124.055 73.785 124.225 ;
        RECT 75.915 124.055 76.085 124.225 ;
        RECT 72.695 123.375 72.865 123.545 ;
        RECT 74.535 123.375 74.705 123.545 ;
        RECT 80.515 125.075 80.685 125.245 ;
        RECT 79.135 124.055 79.305 124.225 ;
        RECT 81.435 124.735 81.605 124.905 ;
        RECT 80.515 124.055 80.685 124.225 ;
        RECT 80.055 123.715 80.225 123.885 ;
        RECT 82.355 124.055 82.525 124.225 ;
        RECT 85.575 124.055 85.745 124.225 ;
        RECT 84.655 123.375 84.825 123.545 ;
        RECT 87.415 124.055 87.585 124.225 ;
        RECT 86.495 123.375 86.665 123.545 ;
        RECT 91.095 124.055 91.265 124.225 ;
        RECT 90.175 123.375 90.345 123.545 ;
        RECT 94.775 124.055 94.945 124.225 ;
        RECT 93.855 123.375 94.025 123.545 ;
        RECT 98.455 124.055 98.625 124.225 ;
        RECT 97.535 123.375 97.705 123.545 ;
        RECT 102.135 124.055 102.305 124.225 ;
        RECT 104.435 124.055 104.605 124.225 ;
        RECT 101.215 123.375 101.385 123.545 ;
        RECT 105.355 123.375 105.525 123.545 ;
        RECT 109.035 124.055 109.205 124.225 ;
        RECT 108.115 123.375 108.285 123.545 ;
        RECT 110.415 124.055 110.585 124.225 ;
        RECT 117.315 125.075 117.485 125.245 ;
        RECT 115.935 124.055 116.105 124.225 ;
        RECT 110.875 123.375 111.045 123.545 ;
        RECT 115.475 123.375 115.645 123.545 ;
        RECT 116.855 124.055 117.025 124.225 ;
        RECT 118.235 124.055 118.405 124.225 ;
        RECT 119.155 123.715 119.325 123.885 ;
        RECT 120.535 125.075 120.705 125.245 ;
        RECT 123.295 125.075 123.465 125.245 ;
        RECT 120.075 123.715 120.245 123.885 ;
        RECT 122.835 124.055 123.005 124.225 ;
        RECT 124.215 124.055 124.385 124.225 ;
        RECT 125.135 123.375 125.305 123.545 ;
        RECT 126.055 125.075 126.225 125.245 ;
        RECT 126.975 124.055 127.145 124.225 ;
        RECT 127.895 124.055 128.065 124.225 ;
        RECT 130.195 124.055 130.365 124.225 ;
        RECT 128.815 123.375 128.985 123.545 ;
        RECT 131.575 125.075 131.745 125.245 ;
        RECT 133.415 124.735 133.585 124.905 ;
        RECT 133.875 124.395 134.045 124.565 ;
        RECT 132.495 124.055 132.665 124.225 ;
        RECT 136.175 124.055 136.345 124.225 ;
        RECT 139.855 125.075 140.025 125.245 ;
        RECT 139.395 124.055 139.565 124.225 ;
        RECT 140.775 124.055 140.945 124.225 ;
        RECT 142.615 125.075 142.785 125.245 ;
        RECT 144.455 125.075 144.625 125.245 ;
        RECT 142.155 124.055 142.325 124.225 ;
        RECT 143.535 124.055 143.705 124.225 ;
        RECT 136.635 123.375 136.805 123.545 ;
        RECT 141.695 123.715 141.865 123.885 ;
        RECT 146.755 124.395 146.925 124.565 ;
        RECT 149.515 125.075 149.685 125.245 ;
        RECT 145.375 123.715 145.545 123.885 ;
        RECT 153.195 125.075 153.365 125.245 ;
        RECT 149.055 123.715 149.225 123.885 ;
        RECT 151.355 124.395 151.525 124.565 ;
        RECT 152.275 124.055 152.445 124.225 ;
        RECT 70.855 122.865 71.025 123.035 ;
        RECT 71.315 122.865 71.485 123.035 ;
        RECT 71.775 122.865 71.945 123.035 ;
        RECT 72.235 122.865 72.405 123.035 ;
        RECT 72.695 122.865 72.865 123.035 ;
        RECT 73.155 122.865 73.325 123.035 ;
        RECT 73.615 122.865 73.785 123.035 ;
        RECT 74.075 122.865 74.245 123.035 ;
        RECT 74.535 122.865 74.705 123.035 ;
        RECT 74.995 122.865 75.165 123.035 ;
        RECT 75.455 122.865 75.625 123.035 ;
        RECT 75.915 122.865 76.085 123.035 ;
        RECT 76.375 122.865 76.545 123.035 ;
        RECT 76.835 122.865 77.005 123.035 ;
        RECT 77.295 122.865 77.465 123.035 ;
        RECT 77.755 122.865 77.925 123.035 ;
        RECT 78.215 122.865 78.385 123.035 ;
        RECT 78.675 122.865 78.845 123.035 ;
        RECT 79.135 122.865 79.305 123.035 ;
        RECT 79.595 122.865 79.765 123.035 ;
        RECT 80.055 122.865 80.225 123.035 ;
        RECT 80.515 122.865 80.685 123.035 ;
        RECT 80.975 122.865 81.145 123.035 ;
        RECT 81.435 122.865 81.605 123.035 ;
        RECT 81.895 122.865 82.065 123.035 ;
        RECT 82.355 122.865 82.525 123.035 ;
        RECT 82.815 122.865 82.985 123.035 ;
        RECT 83.275 122.865 83.445 123.035 ;
        RECT 83.735 122.865 83.905 123.035 ;
        RECT 84.195 122.865 84.365 123.035 ;
        RECT 84.655 122.865 84.825 123.035 ;
        RECT 85.115 122.865 85.285 123.035 ;
        RECT 85.575 122.865 85.745 123.035 ;
        RECT 86.035 122.865 86.205 123.035 ;
        RECT 86.495 122.865 86.665 123.035 ;
        RECT 86.955 122.865 87.125 123.035 ;
        RECT 87.415 122.865 87.585 123.035 ;
        RECT 87.875 122.865 88.045 123.035 ;
        RECT 88.335 122.865 88.505 123.035 ;
        RECT 88.795 122.865 88.965 123.035 ;
        RECT 89.255 122.865 89.425 123.035 ;
        RECT 89.715 122.865 89.885 123.035 ;
        RECT 90.175 122.865 90.345 123.035 ;
        RECT 90.635 122.865 90.805 123.035 ;
        RECT 91.095 122.865 91.265 123.035 ;
        RECT 91.555 122.865 91.725 123.035 ;
        RECT 92.015 122.865 92.185 123.035 ;
        RECT 92.475 122.865 92.645 123.035 ;
        RECT 92.935 122.865 93.105 123.035 ;
        RECT 93.395 122.865 93.565 123.035 ;
        RECT 93.855 122.865 94.025 123.035 ;
        RECT 94.315 122.865 94.485 123.035 ;
        RECT 94.775 122.865 94.945 123.035 ;
        RECT 95.235 122.865 95.405 123.035 ;
        RECT 95.695 122.865 95.865 123.035 ;
        RECT 96.155 122.865 96.325 123.035 ;
        RECT 96.615 122.865 96.785 123.035 ;
        RECT 97.075 122.865 97.245 123.035 ;
        RECT 97.535 122.865 97.705 123.035 ;
        RECT 97.995 122.865 98.165 123.035 ;
        RECT 98.455 122.865 98.625 123.035 ;
        RECT 98.915 122.865 99.085 123.035 ;
        RECT 99.375 122.865 99.545 123.035 ;
        RECT 99.835 122.865 100.005 123.035 ;
        RECT 100.295 122.865 100.465 123.035 ;
        RECT 100.755 122.865 100.925 123.035 ;
        RECT 101.215 122.865 101.385 123.035 ;
        RECT 101.675 122.865 101.845 123.035 ;
        RECT 102.135 122.865 102.305 123.035 ;
        RECT 102.595 122.865 102.765 123.035 ;
        RECT 103.055 122.865 103.225 123.035 ;
        RECT 103.515 122.865 103.685 123.035 ;
        RECT 103.975 122.865 104.145 123.035 ;
        RECT 104.435 122.865 104.605 123.035 ;
        RECT 104.895 122.865 105.065 123.035 ;
        RECT 105.355 122.865 105.525 123.035 ;
        RECT 105.815 122.865 105.985 123.035 ;
        RECT 106.275 122.865 106.445 123.035 ;
        RECT 106.735 122.865 106.905 123.035 ;
        RECT 107.195 122.865 107.365 123.035 ;
        RECT 107.655 122.865 107.825 123.035 ;
        RECT 108.115 122.865 108.285 123.035 ;
        RECT 108.575 122.865 108.745 123.035 ;
        RECT 109.035 122.865 109.205 123.035 ;
        RECT 109.495 122.865 109.665 123.035 ;
        RECT 109.955 122.865 110.125 123.035 ;
        RECT 110.415 122.865 110.585 123.035 ;
        RECT 110.875 122.865 111.045 123.035 ;
        RECT 111.335 122.865 111.505 123.035 ;
        RECT 111.795 122.865 111.965 123.035 ;
        RECT 112.255 122.865 112.425 123.035 ;
        RECT 112.715 122.865 112.885 123.035 ;
        RECT 113.175 122.865 113.345 123.035 ;
        RECT 113.635 122.865 113.805 123.035 ;
        RECT 114.095 122.865 114.265 123.035 ;
        RECT 114.555 122.865 114.725 123.035 ;
        RECT 115.015 122.865 115.185 123.035 ;
        RECT 115.475 122.865 115.645 123.035 ;
        RECT 115.935 122.865 116.105 123.035 ;
        RECT 116.395 122.865 116.565 123.035 ;
        RECT 116.855 122.865 117.025 123.035 ;
        RECT 117.315 122.865 117.485 123.035 ;
        RECT 117.775 122.865 117.945 123.035 ;
        RECT 118.235 122.865 118.405 123.035 ;
        RECT 118.695 122.865 118.865 123.035 ;
        RECT 119.155 122.865 119.325 123.035 ;
        RECT 119.615 122.865 119.785 123.035 ;
        RECT 120.075 122.865 120.245 123.035 ;
        RECT 120.535 122.865 120.705 123.035 ;
        RECT 120.995 122.865 121.165 123.035 ;
        RECT 121.455 122.865 121.625 123.035 ;
        RECT 121.915 122.865 122.085 123.035 ;
        RECT 122.375 122.865 122.545 123.035 ;
        RECT 122.835 122.865 123.005 123.035 ;
        RECT 123.295 122.865 123.465 123.035 ;
        RECT 123.755 122.865 123.925 123.035 ;
        RECT 124.215 122.865 124.385 123.035 ;
        RECT 124.675 122.865 124.845 123.035 ;
        RECT 125.135 122.865 125.305 123.035 ;
        RECT 125.595 122.865 125.765 123.035 ;
        RECT 126.055 122.865 126.225 123.035 ;
        RECT 126.515 122.865 126.685 123.035 ;
        RECT 126.975 122.865 127.145 123.035 ;
        RECT 127.435 122.865 127.605 123.035 ;
        RECT 127.895 122.865 128.065 123.035 ;
        RECT 128.355 122.865 128.525 123.035 ;
        RECT 128.815 122.865 128.985 123.035 ;
        RECT 129.275 122.865 129.445 123.035 ;
        RECT 129.735 122.865 129.905 123.035 ;
        RECT 130.195 122.865 130.365 123.035 ;
        RECT 130.655 122.865 130.825 123.035 ;
        RECT 131.115 122.865 131.285 123.035 ;
        RECT 131.575 122.865 131.745 123.035 ;
        RECT 132.035 122.865 132.205 123.035 ;
        RECT 132.495 122.865 132.665 123.035 ;
        RECT 132.955 122.865 133.125 123.035 ;
        RECT 133.415 122.865 133.585 123.035 ;
        RECT 133.875 122.865 134.045 123.035 ;
        RECT 134.335 122.865 134.505 123.035 ;
        RECT 134.795 122.865 134.965 123.035 ;
        RECT 135.255 122.865 135.425 123.035 ;
        RECT 135.715 122.865 135.885 123.035 ;
        RECT 136.175 122.865 136.345 123.035 ;
        RECT 136.635 122.865 136.805 123.035 ;
        RECT 137.095 122.865 137.265 123.035 ;
        RECT 137.555 122.865 137.725 123.035 ;
        RECT 138.015 122.865 138.185 123.035 ;
        RECT 138.475 122.865 138.645 123.035 ;
        RECT 138.935 122.865 139.105 123.035 ;
        RECT 139.395 122.865 139.565 123.035 ;
        RECT 139.855 122.865 140.025 123.035 ;
        RECT 140.315 122.865 140.485 123.035 ;
        RECT 140.775 122.865 140.945 123.035 ;
        RECT 141.235 122.865 141.405 123.035 ;
        RECT 141.695 122.865 141.865 123.035 ;
        RECT 142.155 122.865 142.325 123.035 ;
        RECT 142.615 122.865 142.785 123.035 ;
        RECT 143.075 122.865 143.245 123.035 ;
        RECT 143.535 122.865 143.705 123.035 ;
        RECT 143.995 122.865 144.165 123.035 ;
        RECT 144.455 122.865 144.625 123.035 ;
        RECT 144.915 122.865 145.085 123.035 ;
        RECT 145.375 122.865 145.545 123.035 ;
        RECT 145.835 122.865 146.005 123.035 ;
        RECT 146.295 122.865 146.465 123.035 ;
        RECT 146.755 122.865 146.925 123.035 ;
        RECT 147.215 122.865 147.385 123.035 ;
        RECT 147.675 122.865 147.845 123.035 ;
        RECT 148.135 122.865 148.305 123.035 ;
        RECT 148.595 122.865 148.765 123.035 ;
        RECT 149.055 122.865 149.225 123.035 ;
        RECT 149.515 122.865 149.685 123.035 ;
        RECT 149.975 122.865 150.145 123.035 ;
        RECT 150.435 122.865 150.605 123.035 ;
        RECT 150.895 122.865 151.065 123.035 ;
        RECT 151.355 122.865 151.525 123.035 ;
        RECT 151.815 122.865 151.985 123.035 ;
        RECT 152.275 122.865 152.445 123.035 ;
        RECT 152.735 122.865 152.905 123.035 ;
        RECT 153.195 122.865 153.365 123.035 ;
        RECT 153.655 122.865 153.825 123.035 ;
        RECT 154.115 122.865 154.285 123.035 ;
        RECT 154.575 122.865 154.745 123.035 ;
        RECT 155.035 122.865 155.205 123.035 ;
        RECT 155.495 122.865 155.665 123.035 ;
        RECT 155.955 122.865 156.125 123.035 ;
        RECT 51.840 100.925 52.370 102.910 ;
        RECT 55.840 100.925 56.370 102.910 ;
        RECT 59.840 100.925 60.370 102.910 ;
        RECT 63.840 100.925 64.370 102.910 ;
        RECT 67.840 100.925 68.370 102.910 ;
        RECT 71.840 100.925 72.370 102.910 ;
        RECT 75.840 100.925 76.370 102.910 ;
        RECT 79.840 100.925 80.370 102.910 ;
        RECT 88.840 100.925 89.370 102.910 ;
        RECT 92.840 100.925 93.370 102.910 ;
        RECT 96.840 100.925 97.370 102.910 ;
        RECT 100.840 100.925 101.370 102.910 ;
        RECT 104.840 100.925 105.370 102.910 ;
        RECT 108.840 100.925 109.370 102.910 ;
        RECT 112.840 100.925 113.370 102.910 ;
        RECT 116.840 100.925 117.370 102.910 ;
        RECT 125.840 100.925 126.370 102.910 ;
        RECT 129.840 100.925 130.370 102.910 ;
        RECT 133.840 100.925 134.370 102.910 ;
        RECT 137.840 100.925 138.370 102.910 ;
        RECT 141.840 100.925 142.370 102.910 ;
        RECT 145.840 100.925 146.370 102.910 ;
        RECT 149.840 100.925 150.370 102.910 ;
        RECT 153.840 100.925 154.370 102.910 ;
        RECT 51.030 79.170 51.370 79.970 ;
        RECT 52.830 79.170 53.170 79.970 ;
        RECT 55.030 79.170 55.370 79.970 ;
        RECT 56.830 79.170 57.170 79.970 ;
        RECT 59.030 79.170 59.370 79.970 ;
        RECT 60.830 79.170 61.170 79.970 ;
        RECT 63.030 79.170 63.370 79.970 ;
        RECT 64.830 79.170 65.170 79.970 ;
        RECT 67.030 79.170 67.370 79.970 ;
        RECT 68.830 79.170 69.170 79.970 ;
        RECT 71.030 79.170 71.370 79.970 ;
        RECT 72.830 79.170 73.170 79.970 ;
        RECT 75.030 79.170 75.370 79.970 ;
        RECT 76.830 79.170 77.170 79.970 ;
        RECT 79.030 79.170 79.370 79.970 ;
        RECT 80.830 79.170 81.170 79.970 ;
        RECT 88.030 79.170 88.370 79.970 ;
        RECT 89.830 79.170 90.170 79.970 ;
        RECT 92.030 79.170 92.370 79.970 ;
        RECT 93.830 79.170 94.170 79.970 ;
        RECT 96.030 79.170 96.370 79.970 ;
        RECT 97.830 79.170 98.170 79.970 ;
        RECT 100.030 79.170 100.370 79.970 ;
        RECT 101.830 79.170 102.170 79.970 ;
        RECT 104.030 79.170 104.370 79.970 ;
        RECT 105.830 79.170 106.170 79.970 ;
        RECT 108.030 79.170 108.370 79.970 ;
        RECT 109.830 79.170 110.170 79.970 ;
        RECT 112.030 79.170 112.370 79.970 ;
        RECT 113.830 79.170 114.170 79.970 ;
        RECT 116.030 79.170 116.370 79.970 ;
        RECT 117.830 79.170 118.170 79.970 ;
        RECT 125.030 79.170 125.370 79.970 ;
        RECT 126.830 79.170 127.170 79.970 ;
        RECT 129.030 79.170 129.370 79.970 ;
        RECT 130.830 79.170 131.170 79.970 ;
        RECT 133.030 79.170 133.370 79.970 ;
        RECT 134.830 79.170 135.170 79.970 ;
        RECT 137.030 79.170 137.370 79.970 ;
        RECT 138.830 79.170 139.170 79.970 ;
        RECT 141.030 79.170 141.370 79.970 ;
        RECT 142.830 79.170 143.170 79.970 ;
        RECT 145.030 79.170 145.370 79.970 ;
        RECT 146.830 79.170 147.170 79.970 ;
        RECT 149.030 79.170 149.370 79.970 ;
        RECT 150.830 79.170 151.170 79.970 ;
        RECT 153.030 79.170 153.370 79.970 ;
        RECT 154.830 79.170 155.170 79.970 ;
        RECT 51.840 59.030 52.370 61.015 ;
        RECT 55.840 59.030 56.370 61.015 ;
        RECT 59.840 59.030 60.370 61.015 ;
        RECT 63.840 59.030 64.370 61.015 ;
        RECT 67.840 59.030 68.370 61.015 ;
        RECT 71.840 59.030 72.370 61.015 ;
        RECT 75.840 59.030 76.370 61.015 ;
        RECT 79.840 59.030 80.370 61.015 ;
        RECT 88.840 59.030 89.370 61.015 ;
        RECT 92.840 59.030 93.370 61.015 ;
        RECT 96.840 59.030 97.370 61.015 ;
        RECT 100.840 59.030 101.370 61.015 ;
        RECT 104.840 59.030 105.370 61.015 ;
        RECT 108.840 59.030 109.370 61.015 ;
        RECT 112.840 59.030 113.370 61.015 ;
        RECT 116.840 59.030 117.370 61.015 ;
        RECT 125.840 59.030 126.370 61.015 ;
        RECT 129.840 59.030 130.370 61.015 ;
        RECT 133.840 59.030 134.370 61.015 ;
        RECT 137.840 59.030 138.370 61.015 ;
        RECT 141.840 59.030 142.370 61.015 ;
        RECT 145.840 59.030 146.370 61.015 ;
        RECT 149.840 59.030 150.370 61.015 ;
        RECT 153.840 59.030 154.370 61.015 ;
        RECT 51.840 52.925 52.370 54.910 ;
        RECT 51.840 31.380 52.370 33.365 ;
        RECT 55.840 52.925 56.370 54.910 ;
        RECT 55.840 31.380 56.370 33.365 ;
        RECT 59.840 52.925 60.370 54.910 ;
        RECT 59.840 31.380 60.370 33.365 ;
        RECT 63.840 52.925 64.370 54.910 ;
        RECT 63.840 31.380 64.370 33.365 ;
        RECT 67.840 52.925 68.370 54.910 ;
        RECT 67.840 31.380 68.370 33.365 ;
        RECT 71.840 52.925 72.370 54.910 ;
        RECT 71.840 31.380 72.370 33.365 ;
        RECT 75.840 52.925 76.370 54.910 ;
        RECT 75.840 31.380 76.370 33.365 ;
        RECT 79.840 52.925 80.370 54.910 ;
        RECT 79.840 31.380 80.370 33.365 ;
        RECT 88.840 52.925 89.370 54.910 ;
        RECT 88.840 31.380 89.370 33.365 ;
        RECT 92.840 52.925 93.370 54.910 ;
        RECT 92.840 31.380 93.370 33.365 ;
        RECT 96.840 52.925 97.370 54.910 ;
        RECT 96.840 31.380 97.370 33.365 ;
        RECT 100.840 52.925 101.370 54.910 ;
        RECT 100.840 31.380 101.370 33.365 ;
        RECT 104.840 52.925 105.370 54.910 ;
        RECT 104.840 31.380 105.370 33.365 ;
        RECT 108.840 52.925 109.370 54.910 ;
        RECT 108.840 31.380 109.370 33.365 ;
        RECT 112.840 52.925 113.370 54.910 ;
        RECT 112.840 31.380 113.370 33.365 ;
        RECT 116.840 52.925 117.370 54.910 ;
        RECT 116.840 31.380 117.370 33.365 ;
        RECT 125.840 52.925 126.370 54.910 ;
        RECT 125.840 31.380 126.370 33.365 ;
        RECT 129.840 52.925 130.370 54.910 ;
        RECT 129.840 31.380 130.370 33.365 ;
        RECT 133.840 52.925 134.370 54.910 ;
        RECT 133.840 31.380 134.370 33.365 ;
        RECT 137.840 52.925 138.370 54.910 ;
        RECT 137.840 31.380 138.370 33.365 ;
        RECT 141.840 52.925 142.370 54.910 ;
        RECT 141.840 31.380 142.370 33.365 ;
        RECT 145.840 52.925 146.370 54.910 ;
        RECT 145.840 31.380 146.370 33.365 ;
        RECT 149.840 52.925 150.370 54.910 ;
        RECT 149.840 31.380 150.370 33.365 ;
        RECT 153.840 52.925 154.370 54.910 ;
        RECT 153.840 31.380 154.370 33.365 ;
        RECT 32.075 26.110 32.245 26.280 ;
        RECT 31.220 21.745 31.520 22.445 ;
        RECT 31.855 17.935 32.025 25.815 ;
        RECT 32.295 17.935 32.465 25.815 ;
        RECT 32.075 17.470 32.245 17.640 ;
        RECT 34.890 24.085 35.060 24.255 ;
        RECT 34.670 19.955 34.840 23.835 ;
        RECT 35.110 19.955 35.280 23.835 ;
        RECT 35.620 22.845 35.920 23.645 ;
        RECT 34.890 19.535 35.060 19.705 ;
      LAYER met1 ;
        RECT 131.960 208.530 132.280 208.590 ;
        RECT 138.400 208.530 138.720 208.590 ;
        RECT 131.960 208.390 138.720 208.530 ;
        RECT 131.960 208.330 132.280 208.390 ;
        RECT 138.400 208.330 138.720 208.390 ;
        RECT 104.360 208.190 104.680 208.250 ;
        RECT 126.900 208.190 127.220 208.250 ;
        RECT 142.080 208.190 142.400 208.250 ;
        RECT 104.360 208.050 142.400 208.190 ;
        RECT 104.360 207.990 104.680 208.050 ;
        RECT 126.900 207.990 127.220 208.050 ;
        RECT 142.080 207.990 142.400 208.050 ;
        RECT 82.740 207.850 83.060 207.910 ;
        RECT 103.900 207.850 104.220 207.910 ;
        RECT 82.740 207.710 104.220 207.850 ;
        RECT 82.740 207.650 83.060 207.710 ;
        RECT 103.900 207.650 104.220 207.710 ;
        RECT 125.060 207.850 125.380 207.910 ;
        RECT 132.880 207.850 133.200 207.910 ;
        RECT 125.060 207.710 133.200 207.850 ;
        RECT 125.060 207.650 125.380 207.710 ;
        RECT 132.880 207.650 133.200 207.710 ;
        RECT 136.100 207.850 136.420 207.910 ;
        RECT 140.700 207.850 141.020 207.910 ;
        RECT 136.100 207.710 141.020 207.850 ;
        RECT 136.100 207.650 136.420 207.710 ;
        RECT 140.700 207.650 141.020 207.710 ;
        RECT 70.710 207.030 156.270 207.510 ;
        RECT 74.000 206.630 74.320 206.890 ;
        RECT 78.140 206.630 78.460 206.890 ;
        RECT 82.280 206.630 82.600 206.890 ;
        RECT 86.420 206.830 86.740 206.890 ;
        RECT 88.275 206.830 88.565 206.875 ;
        RECT 86.420 206.690 88.565 206.830 ;
        RECT 86.420 206.630 86.740 206.690 ;
        RECT 88.275 206.645 88.565 206.690 ;
        RECT 90.560 206.830 90.880 206.890 ;
        RECT 91.495 206.830 91.785 206.875 ;
        RECT 90.560 206.690 91.785 206.830 ;
        RECT 90.560 206.630 90.880 206.690 ;
        RECT 91.495 206.645 91.785 206.690 ;
        RECT 94.700 206.830 95.020 206.890 ;
        RECT 97.475 206.830 97.765 206.875 ;
        RECT 94.700 206.690 97.765 206.830 ;
        RECT 94.700 206.630 95.020 206.690 ;
        RECT 97.475 206.645 97.765 206.690 ;
        RECT 98.840 206.830 99.160 206.890 ;
        RECT 102.980 206.830 103.300 206.890 ;
        RECT 104.375 206.830 104.665 206.875 ;
        RECT 98.840 206.690 102.750 206.830 ;
        RECT 98.840 206.630 99.160 206.690 ;
        RECT 82.370 206.490 82.510 206.630 ;
        RECT 94.255 206.490 94.545 206.535 ;
        RECT 82.370 206.350 94.545 206.490 ;
        RECT 94.255 206.305 94.545 206.350 ;
        RECT 100.695 206.490 100.985 206.535 ;
        RECT 101.600 206.490 101.920 206.550 ;
        RECT 100.695 206.350 101.920 206.490 ;
        RECT 102.610 206.490 102.750 206.690 ;
        RECT 102.980 206.690 104.665 206.830 ;
        RECT 102.980 206.630 103.300 206.690 ;
        RECT 104.375 206.645 104.665 206.690 ;
        RECT 107.120 206.830 107.440 206.890 ;
        RECT 108.515 206.830 108.805 206.875 ;
        RECT 107.120 206.690 108.805 206.830 ;
        RECT 107.120 206.630 107.440 206.690 ;
        RECT 108.515 206.645 108.805 206.690 ;
        RECT 111.260 206.830 111.580 206.890 ;
        RECT 112.195 206.830 112.485 206.875 ;
        RECT 111.260 206.690 112.485 206.830 ;
        RECT 111.260 206.630 111.580 206.690 ;
        RECT 112.195 206.645 112.485 206.690 ;
        RECT 123.680 206.830 124.000 206.890 ;
        RECT 144.380 206.830 144.700 206.890 ;
        RECT 148.980 206.830 149.300 206.890 ;
        RECT 123.680 206.690 136.330 206.830 ;
        RECT 123.680 206.630 124.000 206.690 ;
        RECT 106.215 206.490 106.505 206.535 ;
        RECT 131.515 206.490 131.805 206.535 ;
        RECT 102.610 206.350 106.505 206.490 ;
        RECT 100.695 206.305 100.985 206.350 ;
        RECT 101.600 206.290 101.920 206.350 ;
        RECT 106.215 206.305 106.505 206.350 ;
        RECT 125.610 206.350 131.805 206.490 ;
        RECT 75.470 206.010 82.510 206.150 ;
        RECT 75.470 205.855 75.610 206.010 ;
        RECT 75.395 205.625 75.685 205.855 ;
        RECT 77.235 205.625 77.525 205.855 ;
        RECT 79.075 205.810 79.365 205.855 ;
        RECT 81.820 205.810 82.140 205.870 ;
        RECT 79.075 205.670 82.140 205.810 ;
        RECT 82.370 205.810 82.510 206.010 ;
        RECT 82.740 205.950 83.060 206.210 ;
        RECT 83.200 205.950 83.520 206.210 ;
        RECT 104.360 206.150 104.680 206.210 ;
        RECT 125.610 206.195 125.750 206.350 ;
        RECT 131.515 206.305 131.805 206.350 ;
        RECT 132.880 206.490 133.200 206.550 ;
        RECT 135.655 206.490 135.945 206.535 ;
        RECT 132.880 206.350 135.945 206.490 ;
        RECT 132.880 206.290 133.200 206.350 ;
        RECT 135.655 206.305 135.945 206.350 ;
        RECT 110.355 206.150 110.645 206.195 ;
        RECT 86.510 206.010 104.680 206.150 ;
        RECT 83.290 205.810 83.430 205.950 ;
        RECT 82.370 205.670 83.430 205.810 ;
        RECT 79.075 205.625 79.365 205.670 ;
        RECT 77.310 205.470 77.450 205.625 ;
        RECT 81.820 205.610 82.140 205.670 ;
        RECT 81.375 205.470 81.665 205.515 ;
        RECT 84.135 205.470 84.425 205.515 ;
        RECT 77.310 205.330 79.750 205.470 ;
        RECT 76.300 204.930 76.620 205.190 ;
        RECT 79.610 205.175 79.750 205.330 ;
        RECT 81.375 205.330 84.425 205.470 ;
        RECT 81.375 205.285 81.665 205.330 ;
        RECT 84.135 205.285 84.425 205.330 ;
        RECT 79.535 204.945 79.825 205.175 ;
        RECT 81.835 205.130 82.125 205.175 ;
        RECT 86.510 205.130 86.650 206.010 ;
        RECT 104.360 205.950 104.680 206.010 ;
        RECT 104.910 206.010 110.645 206.150 ;
        RECT 86.895 205.625 87.185 205.855 ;
        RECT 86.970 205.470 87.110 205.625 ;
        RECT 89.180 205.610 89.500 205.870 ;
        RECT 92.400 205.610 92.720 205.870 ;
        RECT 102.060 205.610 102.380 205.870 ;
        RECT 103.440 205.610 103.760 205.870 ;
        RECT 93.335 205.470 93.625 205.515 ;
        RECT 86.970 205.330 93.625 205.470 ;
        RECT 86.970 205.190 87.110 205.330 ;
        RECT 93.335 205.285 93.625 205.330 ;
        RECT 98.855 205.470 99.145 205.515 ;
        RECT 100.220 205.470 100.540 205.530 ;
        RECT 98.855 205.330 100.540 205.470 ;
        RECT 98.855 205.285 99.145 205.330 ;
        RECT 100.220 205.270 100.540 205.330 ;
        RECT 100.680 205.270 101.000 205.530 ;
        RECT 101.615 205.470 101.905 205.515 ;
        RECT 104.910 205.470 105.050 206.010 ;
        RECT 110.355 205.965 110.645 206.010 ;
        RECT 125.535 205.965 125.825 206.195 ;
        RECT 125.980 206.150 126.300 206.210 ;
        RECT 130.135 206.150 130.425 206.195 ;
        RECT 125.980 206.010 130.425 206.150 ;
        RECT 125.980 205.950 126.300 206.010 ;
        RECT 130.135 205.965 130.425 206.010 ;
        RECT 105.295 205.625 105.585 205.855 ;
        RECT 101.615 205.330 105.050 205.470 ;
        RECT 101.615 205.285 101.905 205.330 ;
        RECT 81.835 204.990 86.650 205.130 ;
        RECT 81.835 204.945 82.125 204.990 ;
        RECT 86.880 204.930 87.200 205.190 ;
        RECT 89.180 205.130 89.500 205.190 ;
        RECT 95.160 205.130 95.480 205.190 ;
        RECT 89.180 204.990 95.480 205.130 ;
        RECT 89.180 204.930 89.500 204.990 ;
        RECT 95.160 204.930 95.480 204.990 ;
        RECT 99.760 205.130 100.080 205.190 ;
        RECT 105.370 205.130 105.510 205.625 ;
        RECT 107.580 205.610 107.900 205.870 ;
        RECT 110.815 205.625 111.105 205.855 ;
        RECT 110.890 205.190 111.030 205.625 ;
        RECT 113.100 205.610 113.420 205.870 ;
        RECT 113.575 205.625 113.865 205.855 ;
        RECT 115.400 205.810 115.720 205.870 ;
        RECT 116.795 205.810 117.085 205.855 ;
        RECT 115.400 205.670 117.085 205.810 ;
        RECT 113.650 205.470 113.790 205.625 ;
        RECT 115.400 205.610 115.720 205.670 ;
        RECT 116.795 205.625 117.085 205.670 ;
        RECT 117.255 205.810 117.545 205.855 ;
        RECT 119.540 205.810 119.860 205.870 ;
        RECT 117.255 205.670 119.860 205.810 ;
        RECT 117.255 205.625 117.545 205.670 ;
        RECT 119.540 205.610 119.860 205.670 ;
        RECT 121.840 205.610 122.160 205.870 ;
        RECT 125.060 205.610 125.380 205.870 ;
        RECT 127.820 205.810 128.140 205.870 ;
        RECT 134.735 205.810 135.025 205.855 ;
        RECT 135.180 205.810 135.500 205.870 ;
        RECT 127.820 205.670 134.030 205.810 ;
        RECT 127.820 205.610 128.140 205.670 ;
        RECT 129.215 205.470 129.505 205.515 ;
        RECT 131.500 205.470 131.820 205.530 ;
        RECT 133.890 205.470 134.030 205.670 ;
        RECT 134.735 205.670 135.500 205.810 ;
        RECT 136.190 205.810 136.330 206.690 ;
        RECT 144.380 206.690 149.300 206.830 ;
        RECT 144.380 206.630 144.700 206.690 ;
        RECT 148.980 206.630 149.300 206.690 ;
        RECT 137.020 206.290 137.340 206.550 ;
        RECT 141.200 206.490 141.490 206.535 ;
        RECT 143.300 206.490 143.590 206.535 ;
        RECT 144.870 206.490 145.160 206.535 ;
        RECT 141.200 206.350 145.160 206.490 ;
        RECT 141.200 206.305 141.490 206.350 ;
        RECT 143.300 206.305 143.590 206.350 ;
        RECT 144.870 206.305 145.160 206.350 ;
        RECT 141.595 206.150 141.885 206.195 ;
        RECT 142.785 206.150 143.075 206.195 ;
        RECT 145.305 206.150 145.595 206.195 ;
        RECT 141.595 206.010 145.595 206.150 ;
        RECT 141.595 205.965 141.885 206.010 ;
        RECT 142.785 205.965 143.075 206.010 ;
        RECT 145.305 205.965 145.595 206.010 ;
        RECT 148.520 206.150 148.840 206.210 ;
        RECT 148.995 206.150 149.285 206.195 ;
        RECT 148.520 206.010 149.285 206.150 ;
        RECT 148.520 205.950 148.840 206.010 ;
        RECT 148.995 205.965 149.285 206.010 ;
        RECT 136.575 205.810 136.865 205.855 ;
        RECT 136.190 205.670 136.865 205.810 ;
        RECT 134.735 205.625 135.025 205.670 ;
        RECT 135.180 205.610 135.500 205.670 ;
        RECT 136.575 205.625 136.865 205.670 ;
        RECT 137.955 205.625 138.245 205.855 ;
        RECT 138.400 205.810 138.720 205.870 ;
        RECT 139.335 205.810 139.625 205.855 ;
        RECT 138.400 205.670 139.625 205.810 ;
        RECT 138.030 205.470 138.170 205.625 ;
        RECT 138.400 205.610 138.720 205.670 ;
        RECT 139.335 205.625 139.625 205.670 ;
        RECT 139.780 205.810 140.100 205.870 ;
        RECT 140.715 205.810 141.005 205.855 ;
        RECT 139.780 205.670 141.005 205.810 ;
        RECT 139.780 205.610 140.100 205.670 ;
        RECT 140.715 205.625 141.005 205.670 ;
        RECT 144.840 205.810 145.160 205.870 ;
        RECT 150.375 205.810 150.665 205.855 ;
        RECT 144.840 205.670 150.665 205.810 ;
        RECT 144.840 205.610 145.160 205.670 ;
        RECT 150.375 205.625 150.665 205.670 ;
        RECT 113.650 205.330 127.590 205.470 ;
        RECT 99.760 204.990 105.510 205.130 ;
        RECT 99.760 204.930 100.080 204.990 ;
        RECT 110.800 204.930 111.120 205.190 ;
        RECT 114.480 204.930 114.800 205.190 ;
        RECT 114.940 205.130 115.260 205.190 ;
        RECT 115.875 205.130 116.165 205.175 ;
        RECT 114.940 204.990 116.165 205.130 ;
        RECT 114.940 204.930 115.260 204.990 ;
        RECT 115.875 204.945 116.165 204.990 ;
        RECT 118.160 204.930 118.480 205.190 ;
        RECT 118.620 204.930 118.940 205.190 ;
        RECT 123.220 204.930 123.540 205.190 ;
        RECT 127.450 205.175 127.590 205.330 ;
        RECT 129.215 205.330 133.570 205.470 ;
        RECT 133.890 205.330 138.170 205.470 ;
        RECT 142.050 205.470 142.340 205.515 ;
        RECT 143.460 205.470 143.780 205.530 ;
        RECT 142.050 205.330 143.780 205.470 ;
        RECT 129.215 205.285 129.505 205.330 ;
        RECT 131.500 205.270 131.820 205.330 ;
        RECT 127.375 204.945 127.665 205.175 ;
        RECT 128.280 205.130 128.600 205.190 ;
        RECT 129.675 205.130 129.965 205.175 ;
        RECT 128.280 204.990 129.965 205.130 ;
        RECT 133.430 205.130 133.570 205.330 ;
        RECT 142.050 205.285 142.340 205.330 ;
        RECT 143.460 205.270 143.780 205.330 ;
        RECT 138.415 205.130 138.705 205.175 ;
        RECT 133.430 204.990 138.705 205.130 ;
        RECT 128.280 204.930 128.600 204.990 ;
        RECT 129.675 204.945 129.965 204.990 ;
        RECT 138.415 204.945 138.705 204.990 ;
        RECT 147.140 205.130 147.460 205.190 ;
        RECT 147.615 205.130 147.905 205.175 ;
        RECT 147.140 204.990 147.905 205.130 ;
        RECT 147.140 204.930 147.460 204.990 ;
        RECT 147.615 204.945 147.905 204.990 ;
        RECT 70.710 204.310 156.270 204.790 ;
        RECT 76.300 203.910 76.620 204.170 ;
        RECT 79.995 204.110 80.285 204.155 ;
        RECT 86.880 204.110 87.200 204.170 ;
        RECT 79.995 203.970 87.200 204.110 ;
        RECT 79.995 203.925 80.285 203.970 ;
        RECT 86.880 203.910 87.200 203.970 ;
        RECT 94.255 204.110 94.545 204.155 ;
        RECT 95.620 204.110 95.940 204.170 ;
        RECT 94.255 203.970 95.940 204.110 ;
        RECT 94.255 203.925 94.545 203.970 ;
        RECT 95.620 203.910 95.940 203.970 ;
        RECT 99.760 203.910 100.080 204.170 ;
        RECT 100.680 203.910 101.000 204.170 ;
        RECT 104.835 204.110 105.125 204.155 ;
        RECT 101.230 203.970 105.125 204.110 ;
        RECT 74.430 203.770 74.720 203.815 ;
        RECT 76.390 203.770 76.530 203.910 ;
        RECT 101.230 203.770 101.370 203.970 ;
        RECT 104.835 203.925 105.125 203.970 ;
        RECT 114.480 203.910 114.800 204.170 ;
        RECT 118.620 204.110 118.940 204.170 ;
        RECT 120.015 204.110 120.305 204.155 ;
        RECT 118.620 203.970 120.305 204.110 ;
        RECT 118.620 203.910 118.940 203.970 ;
        RECT 120.015 203.925 120.305 203.970 ;
        RECT 131.960 204.110 132.280 204.170 ;
        RECT 136.560 204.110 136.880 204.170 ;
        RECT 131.960 203.970 136.880 204.110 ;
        RECT 131.960 203.910 132.280 203.970 ;
        RECT 136.560 203.910 136.880 203.970 ;
        RECT 140.240 204.110 140.560 204.170 ;
        RECT 140.240 203.970 146.910 204.110 ;
        RECT 140.240 203.910 140.560 203.970 ;
        RECT 74.430 203.630 76.530 203.770 ;
        RECT 92.030 203.630 101.370 203.770 ;
        RECT 74.430 203.585 74.720 203.630 ;
        RECT 81.820 203.430 82.140 203.490 ;
        RECT 82.295 203.430 82.585 203.475 ;
        RECT 82.740 203.430 83.060 203.490 ;
        RECT 81.820 203.290 83.060 203.430 ;
        RECT 81.820 203.230 82.140 203.290 ;
        RECT 82.295 203.245 82.585 203.290 ;
        RECT 82.740 203.230 83.060 203.290 ;
        RECT 83.200 203.230 83.520 203.490 ;
        RECT 84.120 203.430 84.440 203.490 ;
        RECT 92.030 203.475 92.170 203.630 ;
        RECT 101.615 203.585 101.905 203.815 ;
        RECT 106.675 203.770 106.965 203.815 ;
        RECT 114.020 203.770 114.340 203.830 ;
        RECT 106.675 203.630 114.340 203.770 ;
        RECT 106.675 203.585 106.965 203.630 ;
        RECT 84.955 203.430 85.245 203.475 ;
        RECT 84.120 203.290 85.245 203.430 ;
        RECT 84.120 203.230 84.440 203.290 ;
        RECT 84.955 203.245 85.245 203.290 ;
        RECT 91.955 203.245 92.245 203.475 ;
        RECT 93.335 203.245 93.625 203.475 ;
        RECT 95.635 203.430 95.925 203.475 ;
        RECT 97.460 203.430 97.780 203.490 ;
        RECT 95.635 203.290 97.780 203.430 ;
        RECT 95.635 203.245 95.925 203.290 ;
        RECT 72.160 203.090 72.480 203.150 ;
        RECT 73.095 203.090 73.385 203.135 ;
        RECT 72.160 202.950 73.385 203.090 ;
        RECT 72.160 202.890 72.480 202.950 ;
        RECT 73.095 202.905 73.385 202.950 ;
        RECT 73.975 203.090 74.265 203.135 ;
        RECT 75.165 203.090 75.455 203.135 ;
        RECT 77.685 203.090 77.975 203.135 ;
        RECT 83.675 203.090 83.965 203.135 ;
        RECT 73.975 202.950 77.975 203.090 ;
        RECT 73.975 202.905 74.265 202.950 ;
        RECT 75.165 202.905 75.455 202.950 ;
        RECT 77.685 202.905 77.975 202.950 ;
        RECT 81.910 202.950 83.965 203.090 ;
        RECT 73.580 202.750 73.870 202.795 ;
        RECT 75.680 202.750 75.970 202.795 ;
        RECT 77.250 202.750 77.540 202.795 ;
        RECT 73.580 202.610 77.540 202.750 ;
        RECT 73.580 202.565 73.870 202.610 ;
        RECT 75.680 202.565 75.970 202.610 ;
        RECT 77.250 202.565 77.540 202.610 ;
        RECT 81.910 202.470 82.050 202.950 ;
        RECT 83.675 202.905 83.965 202.950 ;
        RECT 84.555 203.090 84.845 203.135 ;
        RECT 85.745 203.090 86.035 203.135 ;
        RECT 88.265 203.090 88.555 203.135 ;
        RECT 84.555 202.950 88.555 203.090 ;
        RECT 84.555 202.905 84.845 202.950 ;
        RECT 85.745 202.905 86.035 202.950 ;
        RECT 88.265 202.905 88.555 202.950 ;
        RECT 89.180 203.090 89.500 203.150 ;
        RECT 93.410 203.090 93.550 203.245 ;
        RECT 97.460 203.230 97.780 203.290 ;
        RECT 97.920 203.230 98.240 203.490 ;
        RECT 99.300 203.430 99.620 203.490 ;
        RECT 101.690 203.430 101.830 203.585 ;
        RECT 114.020 203.570 114.340 203.630 ;
        RECT 114.570 203.475 114.710 203.910 ;
        RECT 139.780 203.770 140.100 203.830 ;
        RECT 115.950 203.630 140.100 203.770 ;
        RECT 115.950 203.490 116.090 203.630 ;
        RECT 99.300 203.290 101.830 203.430 ;
        RECT 102.610 203.290 109.190 203.430 ;
        RECT 99.300 203.230 99.620 203.290 ;
        RECT 89.180 202.950 93.550 203.090 ;
        RECT 98.395 203.090 98.685 203.135 ;
        RECT 98.840 203.090 99.160 203.150 ;
        RECT 98.395 202.950 99.160 203.090 ;
        RECT 89.180 202.890 89.500 202.950 ;
        RECT 98.395 202.905 98.685 202.950 ;
        RECT 98.840 202.890 99.160 202.950 ;
        RECT 84.160 202.750 84.450 202.795 ;
        RECT 86.260 202.750 86.550 202.795 ;
        RECT 87.830 202.750 88.120 202.795 ;
        RECT 99.760 202.750 100.080 202.810 ;
        RECT 84.160 202.610 88.120 202.750 ;
        RECT 84.160 202.565 84.450 202.610 ;
        RECT 86.260 202.565 86.550 202.610 ;
        RECT 87.830 202.565 88.120 202.610 ;
        RECT 88.810 202.610 100.080 202.750 ;
        RECT 81.820 202.210 82.140 202.470 ;
        RECT 83.215 202.410 83.505 202.455 ;
        RECT 88.810 202.410 88.950 202.610 ;
        RECT 99.760 202.550 100.080 202.610 ;
        RECT 83.215 202.270 88.950 202.410 ;
        RECT 89.180 202.410 89.500 202.470 ;
        RECT 90.575 202.410 90.865 202.455 ;
        RECT 89.180 202.270 90.865 202.410 ;
        RECT 83.215 202.225 83.505 202.270 ;
        RECT 89.180 202.210 89.500 202.270 ;
        RECT 90.575 202.225 90.865 202.270 ;
        RECT 91.020 202.210 91.340 202.470 ;
        RECT 94.700 202.210 95.020 202.470 ;
        RECT 101.615 202.410 101.905 202.455 ;
        RECT 102.610 202.410 102.750 203.290 ;
        RECT 102.980 203.090 103.300 203.150 ;
        RECT 107.135 203.090 107.425 203.135 ;
        RECT 102.980 202.950 107.425 203.090 ;
        RECT 102.980 202.890 103.300 202.950 ;
        RECT 107.135 202.905 107.425 202.950 ;
        RECT 107.595 202.905 107.885 203.135 ;
        RECT 103.455 202.750 103.745 202.795 ;
        RECT 104.820 202.750 105.140 202.810 ;
        RECT 103.455 202.610 105.140 202.750 ;
        RECT 103.455 202.565 103.745 202.610 ;
        RECT 104.820 202.550 105.140 202.610 ;
        RECT 101.615 202.270 102.750 202.410 ;
        RECT 102.980 202.410 103.300 202.470 ;
        RECT 107.670 202.410 107.810 202.905 ;
        RECT 109.050 202.455 109.190 203.290 ;
        RECT 114.540 203.245 114.830 203.475 ;
        RECT 115.860 203.230 116.180 203.490 ;
        RECT 117.255 203.430 117.545 203.475 ;
        RECT 118.160 203.430 118.480 203.490 ;
        RECT 119.555 203.430 119.845 203.475 ;
        RECT 117.255 203.290 117.930 203.430 ;
        RECT 117.255 203.245 117.545 203.290 ;
        RECT 111.285 203.090 111.575 203.135 ;
        RECT 113.805 203.090 114.095 203.135 ;
        RECT 114.995 203.090 115.285 203.135 ;
        RECT 111.285 202.950 115.285 203.090 ;
        RECT 111.285 202.905 111.575 202.950 ;
        RECT 113.805 202.905 114.095 202.950 ;
        RECT 114.995 202.905 115.285 202.950 ;
        RECT 117.790 202.795 117.930 203.290 ;
        RECT 118.160 203.290 119.845 203.430 ;
        RECT 118.160 203.230 118.480 203.290 ;
        RECT 119.555 203.245 119.845 203.290 ;
        RECT 123.220 203.430 123.540 203.490 ;
        RECT 125.610 203.475 125.750 203.630 ;
        RECT 124.155 203.430 124.445 203.475 ;
        RECT 123.220 203.290 124.445 203.430 ;
        RECT 123.220 203.230 123.540 203.290 ;
        RECT 124.155 203.245 124.445 203.290 ;
        RECT 125.535 203.245 125.825 203.475 ;
        RECT 126.815 203.430 127.105 203.475 ;
        RECT 126.070 203.290 127.105 203.430 ;
        RECT 120.935 202.905 121.225 203.135 ;
        RECT 126.070 203.090 126.210 203.290 ;
        RECT 126.815 203.245 127.105 203.290 ;
        RECT 133.800 203.430 134.120 203.490 ;
        RECT 134.275 203.430 134.565 203.475 ;
        RECT 133.800 203.290 134.565 203.430 ;
        RECT 133.800 203.230 134.120 203.290 ;
        RECT 134.275 203.245 134.565 203.290 ;
        RECT 134.720 203.430 135.040 203.490 ;
        RECT 137.110 203.475 137.250 203.630 ;
        RECT 139.780 203.570 140.100 203.630 ;
        RECT 135.655 203.430 135.945 203.475 ;
        RECT 134.720 203.290 135.945 203.430 ;
        RECT 134.720 203.230 135.040 203.290 ;
        RECT 135.655 203.245 135.945 203.290 ;
        RECT 137.035 203.245 137.325 203.475 ;
        RECT 138.315 203.430 138.605 203.475 ;
        RECT 137.570 203.290 138.605 203.430 ;
        RECT 125.150 202.950 126.210 203.090 ;
        RECT 126.415 203.090 126.705 203.135 ;
        RECT 127.605 203.090 127.895 203.135 ;
        RECT 130.125 203.090 130.415 203.135 ;
        RECT 135.180 203.090 135.500 203.150 ;
        RECT 137.570 203.090 137.710 203.290 ;
        RECT 138.315 203.245 138.605 203.290 ;
        RECT 140.700 203.430 141.020 203.490 ;
        RECT 146.770 203.475 146.910 203.970 ;
        RECT 148.980 203.910 149.300 204.170 ;
        RECT 149.070 203.770 149.210 203.910 ;
        RECT 149.070 203.630 153.810 203.770 ;
        RECT 145.315 203.430 145.605 203.475 ;
        RECT 140.700 203.290 145.605 203.430 ;
        RECT 140.700 203.230 141.020 203.290 ;
        RECT 145.315 203.245 145.605 203.290 ;
        RECT 146.695 203.245 146.985 203.475 ;
        RECT 148.060 203.430 148.380 203.490 ;
        RECT 153.670 203.475 153.810 203.630 ;
        RECT 150.375 203.430 150.665 203.475 ;
        RECT 148.060 203.290 152.890 203.430 ;
        RECT 148.060 203.230 148.380 203.290 ;
        RECT 150.375 203.245 150.665 203.290 ;
        RECT 126.415 202.950 130.415 203.090 ;
        RECT 111.720 202.750 112.010 202.795 ;
        RECT 113.290 202.750 113.580 202.795 ;
        RECT 115.390 202.750 115.680 202.795 ;
        RECT 111.720 202.610 115.680 202.750 ;
        RECT 111.720 202.565 112.010 202.610 ;
        RECT 113.290 202.565 113.580 202.610 ;
        RECT 115.390 202.565 115.680 202.610 ;
        RECT 117.715 202.565 118.005 202.795 ;
        RECT 102.980 202.270 107.810 202.410 ;
        RECT 108.975 202.410 109.265 202.455 ;
        RECT 110.800 202.410 111.120 202.470 ;
        RECT 114.020 202.410 114.340 202.470 ;
        RECT 108.975 202.270 114.340 202.410 ;
        RECT 101.615 202.225 101.905 202.270 ;
        RECT 102.980 202.210 103.300 202.270 ;
        RECT 108.975 202.225 109.265 202.270 ;
        RECT 110.800 202.210 111.120 202.270 ;
        RECT 114.020 202.210 114.340 202.270 ;
        RECT 116.320 202.210 116.640 202.470 ;
        RECT 121.010 202.410 121.150 202.905 ;
        RECT 125.150 202.795 125.290 202.950 ;
        RECT 126.415 202.905 126.705 202.950 ;
        RECT 127.605 202.905 127.895 202.950 ;
        RECT 130.125 202.905 130.415 202.950 ;
        RECT 132.510 202.950 135.500 203.090 ;
        RECT 125.075 202.565 125.365 202.795 ;
        RECT 125.520 202.550 125.840 202.810 ;
        RECT 132.510 202.795 132.650 202.950 ;
        RECT 135.180 202.890 135.500 202.950 ;
        RECT 137.110 202.950 137.710 203.090 ;
        RECT 137.915 203.090 138.205 203.135 ;
        RECT 139.105 203.090 139.395 203.135 ;
        RECT 141.625 203.090 141.915 203.135 ;
        RECT 137.915 202.950 141.915 203.090 ;
        RECT 126.020 202.750 126.310 202.795 ;
        RECT 128.120 202.750 128.410 202.795 ;
        RECT 129.690 202.750 129.980 202.795 ;
        RECT 126.020 202.610 129.980 202.750 ;
        RECT 126.020 202.565 126.310 202.610 ;
        RECT 128.120 202.565 128.410 202.610 ;
        RECT 129.690 202.565 129.980 202.610 ;
        RECT 132.435 202.565 132.725 202.795 ;
        RECT 136.575 202.750 136.865 202.795 ;
        RECT 137.110 202.750 137.250 202.950 ;
        RECT 137.915 202.905 138.205 202.950 ;
        RECT 139.105 202.905 139.395 202.950 ;
        RECT 141.625 202.905 141.915 202.950 ;
        RECT 142.080 202.890 142.400 203.150 ;
        RECT 147.140 203.090 147.460 203.150 ;
        RECT 150.835 203.090 151.125 203.135 ;
        RECT 147.140 202.950 151.125 203.090 ;
        RECT 147.140 202.890 147.460 202.950 ;
        RECT 150.835 202.905 151.125 202.950 ;
        RECT 151.295 202.905 151.585 203.135 ;
        RECT 136.575 202.610 137.250 202.750 ;
        RECT 137.520 202.750 137.810 202.795 ;
        RECT 139.620 202.750 139.910 202.795 ;
        RECT 141.190 202.750 141.480 202.795 ;
        RECT 137.520 202.610 141.480 202.750 ;
        RECT 136.575 202.565 136.865 202.610 ;
        RECT 137.520 202.565 137.810 202.610 ;
        RECT 139.620 202.565 139.910 202.610 ;
        RECT 141.190 202.565 141.480 202.610 ;
        RECT 125.610 202.410 125.750 202.550 ;
        RECT 121.010 202.270 125.750 202.410 ;
        RECT 130.580 202.410 130.900 202.470 ;
        RECT 132.510 202.410 132.650 202.565 ;
        RECT 130.580 202.270 132.650 202.410 ;
        RECT 133.340 202.410 133.660 202.470 ;
        RECT 138.860 202.410 139.180 202.470 ;
        RECT 133.340 202.270 139.180 202.410 ;
        RECT 142.170 202.410 142.310 202.890 ;
        RECT 143.000 202.750 143.320 202.810 ;
        RECT 151.370 202.750 151.510 202.905 ;
        RECT 152.750 202.795 152.890 203.290 ;
        RECT 153.595 203.245 153.885 203.475 ;
        RECT 143.000 202.610 151.510 202.750 ;
        RECT 143.000 202.550 143.320 202.610 ;
        RECT 152.675 202.565 152.965 202.795 ;
        RECT 143.935 202.410 144.225 202.455 ;
        RECT 142.170 202.270 144.225 202.410 ;
        RECT 130.580 202.210 130.900 202.270 ;
        RECT 133.340 202.210 133.660 202.270 ;
        RECT 138.860 202.210 139.180 202.270 ;
        RECT 143.935 202.225 144.225 202.270 ;
        RECT 144.380 202.210 144.700 202.470 ;
        RECT 145.760 202.210 146.080 202.470 ;
        RECT 148.520 202.210 148.840 202.470 ;
        RECT 70.710 201.590 156.270 202.070 ;
        RECT 101.600 201.190 101.920 201.450 ;
        RECT 102.060 201.390 102.380 201.450 ;
        RECT 102.995 201.390 103.285 201.435 ;
        RECT 102.060 201.250 103.285 201.390 ;
        RECT 102.060 201.190 102.380 201.250 ;
        RECT 102.995 201.205 103.285 201.250 ;
        RECT 103.900 201.190 104.220 201.450 ;
        RECT 104.360 201.190 104.680 201.450 ;
        RECT 115.860 201.390 116.180 201.450 ;
        RECT 114.570 201.250 116.180 201.390 ;
        RECT 74.500 201.050 74.790 201.095 ;
        RECT 76.600 201.050 76.890 201.095 ;
        RECT 78.170 201.050 78.460 201.095 ;
        RECT 74.500 200.910 78.460 201.050 ;
        RECT 74.500 200.865 74.790 200.910 ;
        RECT 76.600 200.865 76.890 200.910 ;
        RECT 78.170 200.865 78.460 200.910 ;
        RECT 83.215 201.050 83.505 201.095 ;
        RECT 84.120 201.050 84.440 201.110 ;
        RECT 83.215 200.910 84.440 201.050 ;
        RECT 83.215 200.865 83.505 200.910 ;
        RECT 84.120 200.850 84.440 200.910 ;
        RECT 86.880 201.050 87.170 201.095 ;
        RECT 88.450 201.050 88.740 201.095 ;
        RECT 90.550 201.050 90.840 201.095 ;
        RECT 86.880 200.910 90.840 201.050 ;
        RECT 86.880 200.865 87.170 200.910 ;
        RECT 88.450 200.865 88.740 200.910 ;
        RECT 90.550 200.865 90.840 200.910 ;
        RECT 92.440 201.050 92.730 201.095 ;
        RECT 94.540 201.050 94.830 201.095 ;
        RECT 96.110 201.050 96.400 201.095 ;
        RECT 92.440 200.910 96.400 201.050 ;
        RECT 92.440 200.865 92.730 200.910 ;
        RECT 94.540 200.865 94.830 200.910 ;
        RECT 96.110 200.865 96.400 200.910 ;
        RECT 74.895 200.710 75.185 200.755 ;
        RECT 76.085 200.710 76.375 200.755 ;
        RECT 78.605 200.710 78.895 200.755 ;
        RECT 81.820 200.710 82.140 200.770 ;
        RECT 86.445 200.710 86.735 200.755 ;
        RECT 88.965 200.710 89.255 200.755 ;
        RECT 90.155 200.710 90.445 200.755 ;
        RECT 74.895 200.570 78.895 200.710 ;
        RECT 74.895 200.525 75.185 200.570 ;
        RECT 76.085 200.525 76.375 200.570 ;
        RECT 78.605 200.525 78.895 200.570 ;
        RECT 80.945 200.570 83.890 200.710 ;
        RECT 72.160 200.370 72.480 200.430 ;
        RECT 74.015 200.370 74.305 200.415 ;
        RECT 80.945 200.370 81.085 200.570 ;
        RECT 81.820 200.510 82.140 200.570 ;
        RECT 72.160 200.230 81.085 200.370 ;
        RECT 82.295 200.370 82.585 200.415 ;
        RECT 83.200 200.370 83.520 200.430 ;
        RECT 82.295 200.230 83.520 200.370 ;
        RECT 83.750 200.370 83.890 200.570 ;
        RECT 86.445 200.570 90.445 200.710 ;
        RECT 86.445 200.525 86.735 200.570 ;
        RECT 88.965 200.525 89.255 200.570 ;
        RECT 90.155 200.525 90.445 200.570 ;
        RECT 91.035 200.525 91.325 200.755 ;
        RECT 92.835 200.710 93.125 200.755 ;
        RECT 94.025 200.710 94.315 200.755 ;
        RECT 96.545 200.710 96.835 200.755 ;
        RECT 92.835 200.570 96.835 200.710 ;
        RECT 92.835 200.525 93.125 200.570 ;
        RECT 94.025 200.525 94.315 200.570 ;
        RECT 96.545 200.525 96.835 200.570 ;
        RECT 91.110 200.370 91.250 200.525 ;
        RECT 100.220 200.510 100.540 200.770 ;
        RECT 101.690 200.710 101.830 201.190 ;
        RECT 103.990 201.050 104.130 201.190 ;
        RECT 107.595 201.050 107.885 201.095 ;
        RECT 103.990 200.910 107.885 201.050 ;
        RECT 107.595 200.865 107.885 200.910 ;
        RECT 114.570 200.755 114.710 201.250 ;
        RECT 115.860 201.190 116.180 201.250 ;
        RECT 121.395 201.390 121.685 201.435 ;
        RECT 121.840 201.390 122.160 201.450 ;
        RECT 125.520 201.390 125.840 201.450 ;
        RECT 129.660 201.390 129.980 201.450 ;
        RECT 121.395 201.250 125.840 201.390 ;
        RECT 121.395 201.205 121.685 201.250 ;
        RECT 121.840 201.190 122.160 201.250 ;
        RECT 125.520 201.190 125.840 201.250 ;
        RECT 129.290 201.250 129.980 201.390 ;
        RECT 114.980 201.050 115.270 201.095 ;
        RECT 117.080 201.050 117.370 201.095 ;
        RECT 118.650 201.050 118.940 201.095 ;
        RECT 114.980 200.910 118.940 201.050 ;
        RECT 114.980 200.865 115.270 200.910 ;
        RECT 117.080 200.865 117.370 200.910 ;
        RECT 118.650 200.865 118.940 200.910 ;
        RECT 123.680 201.050 124.000 201.110 ;
        RECT 129.290 201.050 129.430 201.250 ;
        RECT 129.660 201.190 129.980 201.250 ;
        RECT 134.260 201.390 134.580 201.450 ;
        RECT 135.655 201.390 135.945 201.435 ;
        RECT 134.260 201.250 135.945 201.390 ;
        RECT 134.260 201.190 134.580 201.250 ;
        RECT 135.655 201.205 135.945 201.250 ;
        RECT 123.680 200.910 129.430 201.050 ;
        RECT 131.040 201.050 131.360 201.110 ;
        RECT 133.340 201.050 133.660 201.110 ;
        RECT 139.795 201.050 140.085 201.095 ;
        RECT 131.040 200.910 133.660 201.050 ;
        RECT 123.680 200.850 124.000 200.910 ;
        RECT 131.040 200.850 131.360 200.910 ;
        RECT 133.340 200.850 133.660 200.910 ;
        RECT 138.030 200.910 140.085 201.050 ;
        RECT 101.690 200.570 108.270 200.710 ;
        RECT 91.955 200.370 92.245 200.415 ;
        RECT 83.750 200.230 92.245 200.370 ;
        RECT 72.160 200.170 72.480 200.230 ;
        RECT 74.015 200.185 74.305 200.230 ;
        RECT 82.295 200.185 82.585 200.230 ;
        RECT 83.200 200.170 83.520 200.230 ;
        RECT 91.955 200.185 92.245 200.230 ;
        RECT 93.290 200.370 93.580 200.415 ;
        RECT 94.700 200.370 95.020 200.430 ;
        RECT 100.695 200.370 100.985 200.415 ;
        RECT 93.290 200.230 95.020 200.370 ;
        RECT 93.290 200.185 93.580 200.230 ;
        RECT 94.700 200.170 95.020 200.230 ;
        RECT 95.710 200.230 100.985 200.370 ;
        RECT 95.710 200.090 95.850 200.230 ;
        RECT 100.695 200.185 100.985 200.230 ;
        RECT 105.295 200.185 105.585 200.415 ;
        RECT 106.215 200.185 106.505 200.415 ;
        RECT 106.675 200.370 106.965 200.415 ;
        RECT 107.120 200.370 107.440 200.430 ;
        RECT 106.675 200.230 107.440 200.370 ;
        RECT 106.675 200.185 106.965 200.230 ;
        RECT 75.380 200.075 75.700 200.090 ;
        RECT 75.350 199.845 75.700 200.075 ;
        RECT 89.810 200.030 90.100 200.075 ;
        RECT 91.020 200.030 91.340 200.090 ;
        RECT 75.380 199.830 75.700 199.845 ;
        RECT 80.990 199.890 89.410 200.030 ;
        RECT 80.990 199.750 81.130 199.890 ;
        RECT 80.900 199.490 81.220 199.750 ;
        RECT 84.120 199.490 84.440 199.750 ;
        RECT 89.270 199.690 89.410 199.890 ;
        RECT 89.810 199.890 91.340 200.030 ;
        RECT 89.810 199.845 90.100 199.890 ;
        RECT 91.020 199.830 91.340 199.890 ;
        RECT 95.620 199.830 95.940 200.090 ;
        RECT 96.080 200.030 96.400 200.090 ;
        RECT 101.155 200.030 101.445 200.075 ;
        RECT 96.080 199.890 101.445 200.030 ;
        RECT 96.080 199.830 96.400 199.890 ;
        RECT 101.155 199.845 101.445 199.890 ;
        RECT 105.370 199.750 105.510 200.185 ;
        RECT 106.290 200.030 106.430 200.185 ;
        RECT 107.120 200.170 107.440 200.230 ;
        RECT 107.580 200.170 107.900 200.430 ;
        RECT 108.130 200.415 108.270 200.570 ;
        RECT 114.495 200.525 114.785 200.755 ;
        RECT 115.375 200.710 115.665 200.755 ;
        RECT 116.565 200.710 116.855 200.755 ;
        RECT 119.085 200.710 119.375 200.755 ;
        RECT 115.375 200.570 119.375 200.710 ;
        RECT 115.375 200.525 115.665 200.570 ;
        RECT 116.565 200.525 116.855 200.570 ;
        RECT 119.085 200.525 119.375 200.570 ;
        RECT 124.155 200.710 124.445 200.755 ;
        RECT 125.060 200.710 125.380 200.770 ;
        RECT 124.155 200.570 125.380 200.710 ;
        RECT 124.155 200.525 124.445 200.570 ;
        RECT 125.060 200.510 125.380 200.570 ;
        RECT 125.980 200.510 126.300 200.770 ;
        RECT 129.200 200.510 129.520 200.770 ;
        RECT 137.020 200.710 137.340 200.770 ;
        RECT 138.030 200.755 138.170 200.910 ;
        RECT 139.795 200.865 140.085 200.910 ;
        RECT 140.240 201.050 140.560 201.110 ;
        RECT 146.720 201.050 147.010 201.095 ;
        RECT 148.820 201.050 149.110 201.095 ;
        RECT 150.390 201.050 150.680 201.095 ;
        RECT 140.240 200.910 146.450 201.050 ;
        RECT 140.240 200.850 140.560 200.910 ;
        RECT 137.955 200.710 138.245 200.755 ;
        RECT 130.210 200.570 134.030 200.710 ;
        RECT 108.055 200.185 108.345 200.415 ;
        RECT 108.960 200.170 109.280 200.430 ;
        RECT 111.735 200.185 112.025 200.415 ;
        RECT 112.655 200.185 112.945 200.415 ;
        RECT 113.115 200.370 113.405 200.415 ;
        RECT 114.940 200.370 115.260 200.430 ;
        RECT 113.115 200.230 115.260 200.370 ;
        RECT 113.115 200.185 113.405 200.230 ;
        RECT 109.050 200.030 109.190 200.170 ;
        RECT 106.290 199.890 109.190 200.030 ;
        RECT 111.810 200.030 111.950 200.185 ;
        RECT 112.180 200.030 112.500 200.090 ;
        RECT 111.810 199.890 112.500 200.030 ;
        RECT 112.730 200.030 112.870 200.185 ;
        RECT 114.940 200.170 115.260 200.230 ;
        RECT 122.760 200.370 123.080 200.430 ;
        RECT 130.210 200.415 130.350 200.570 ;
        RECT 130.135 200.370 130.425 200.415 ;
        RECT 122.760 200.230 130.635 200.370 ;
        RECT 122.760 200.170 123.080 200.230 ;
        RECT 130.135 200.185 130.425 200.230 ;
        RECT 131.500 200.170 131.820 200.430 ;
        RECT 133.355 200.185 133.645 200.415 ;
        RECT 114.480 200.030 114.800 200.090 ;
        RECT 112.730 199.890 114.800 200.030 ;
        RECT 112.180 199.830 112.500 199.890 ;
        RECT 114.480 199.830 114.800 199.890 ;
        RECT 115.830 200.030 116.120 200.075 ;
        RECT 116.320 200.030 116.640 200.090 ;
        RECT 115.830 199.890 116.640 200.030 ;
        RECT 115.830 199.845 116.120 199.890 ;
        RECT 116.320 199.830 116.640 199.890 ;
        RECT 126.440 199.830 126.760 200.090 ;
        RECT 126.915 200.030 127.205 200.075 ;
        RECT 131.960 200.030 132.280 200.090 ;
        RECT 126.915 199.890 132.280 200.030 ;
        RECT 126.915 199.845 127.205 199.890 ;
        RECT 131.960 199.830 132.280 199.890 ;
        RECT 133.430 199.750 133.570 200.185 ;
        RECT 133.890 200.030 134.030 200.570 ;
        RECT 137.020 200.570 138.245 200.710 ;
        RECT 137.020 200.510 137.340 200.570 ;
        RECT 137.955 200.525 138.245 200.570 ;
        RECT 138.875 200.710 139.165 200.755 ;
        RECT 143.000 200.710 143.320 200.770 ;
        RECT 146.310 200.755 146.450 200.910 ;
        RECT 146.720 200.910 150.680 201.050 ;
        RECT 146.720 200.865 147.010 200.910 ;
        RECT 148.820 200.865 149.110 200.910 ;
        RECT 150.390 200.865 150.680 200.910 ;
        RECT 138.875 200.570 143.320 200.710 ;
        RECT 138.875 200.525 139.165 200.570 ;
        RECT 143.000 200.510 143.320 200.570 ;
        RECT 146.235 200.525 146.525 200.755 ;
        RECT 147.115 200.710 147.405 200.755 ;
        RECT 148.305 200.710 148.595 200.755 ;
        RECT 150.825 200.710 151.115 200.755 ;
        RECT 147.115 200.570 151.115 200.710 ;
        RECT 147.115 200.525 147.405 200.570 ;
        RECT 148.305 200.525 148.595 200.570 ;
        RECT 150.825 200.525 151.115 200.570 ;
        RECT 134.260 200.170 134.580 200.430 ;
        RECT 134.735 200.370 135.025 200.415 ;
        RECT 137.495 200.370 137.785 200.415 ;
        RECT 144.380 200.370 144.700 200.430 ;
        RECT 134.735 200.230 144.700 200.370 ;
        RECT 134.735 200.185 135.025 200.230 ;
        RECT 137.495 200.185 137.785 200.230 ;
        RECT 144.380 200.170 144.700 200.230 ;
        RECT 145.760 200.170 146.080 200.430 ;
        RECT 140.715 200.030 141.005 200.075 ;
        RECT 142.080 200.030 142.400 200.090 ;
        RECT 133.890 199.890 139.550 200.030 ;
        RECT 139.410 199.750 139.550 199.890 ;
        RECT 140.715 199.890 142.400 200.030 ;
        RECT 140.715 199.845 141.005 199.890 ;
        RECT 142.080 199.830 142.400 199.890 ;
        RECT 143.920 200.030 144.240 200.090 ;
        RECT 145.850 200.030 145.990 200.170 ;
        RECT 143.920 199.890 145.990 200.030 ;
        RECT 146.680 200.030 147.000 200.090 ;
        RECT 147.460 200.030 147.750 200.075 ;
        RECT 146.680 199.890 147.750 200.030 ;
        RECT 143.920 199.830 144.240 199.890 ;
        RECT 146.680 199.830 147.000 199.890 ;
        RECT 147.460 199.845 147.750 199.890 ;
        RECT 96.540 199.690 96.860 199.750 ;
        RECT 89.270 199.550 96.860 199.690 ;
        RECT 96.540 199.490 96.860 199.550 ;
        RECT 98.840 199.490 99.160 199.750 ;
        RECT 105.280 199.490 105.600 199.750 ;
        RECT 108.515 199.690 108.805 199.735 ;
        RECT 110.340 199.690 110.660 199.750 ;
        RECT 108.515 199.550 110.660 199.690 ;
        RECT 108.515 199.505 108.805 199.550 ;
        RECT 110.340 199.490 110.660 199.550 ;
        RECT 110.815 199.690 111.105 199.735 ;
        RECT 112.640 199.690 112.960 199.750 ;
        RECT 110.815 199.550 112.960 199.690 ;
        RECT 110.815 199.505 111.105 199.550 ;
        RECT 112.640 199.490 112.960 199.550 ;
        RECT 121.840 199.490 122.160 199.750 ;
        RECT 128.740 199.490 129.060 199.750 ;
        RECT 132.420 199.490 132.740 199.750 ;
        RECT 133.340 199.690 133.660 199.750 ;
        RECT 137.480 199.690 137.800 199.750 ;
        RECT 133.340 199.550 137.800 199.690 ;
        RECT 133.340 199.490 133.660 199.550 ;
        RECT 137.480 199.490 137.800 199.550 ;
        RECT 139.320 199.490 139.640 199.750 ;
        RECT 143.475 199.690 143.765 199.735 ;
        RECT 145.300 199.690 145.620 199.750 ;
        RECT 143.475 199.550 145.620 199.690 ;
        RECT 143.475 199.505 143.765 199.550 ;
        RECT 145.300 199.490 145.620 199.550 ;
        RECT 145.760 199.490 146.080 199.750 ;
        RECT 153.120 199.490 153.440 199.750 ;
        RECT 70.710 198.870 156.270 199.350 ;
        RECT 74.935 198.670 75.225 198.715 ;
        RECT 75.380 198.670 75.700 198.730 ;
        RECT 74.935 198.530 75.700 198.670 ;
        RECT 74.935 198.485 75.225 198.530 ;
        RECT 75.380 198.470 75.700 198.530 ;
        RECT 78.140 198.470 78.460 198.730 ;
        RECT 78.615 198.485 78.905 198.715 ;
        RECT 80.900 198.670 81.220 198.730 ;
        RECT 84.120 198.670 84.440 198.730 ;
        RECT 84.595 198.670 84.885 198.715 ;
        RECT 87.800 198.670 88.120 198.730 ;
        RECT 80.900 198.530 83.890 198.670 ;
        RECT 78.690 198.330 78.830 198.485 ;
        RECT 80.900 198.470 81.220 198.530 ;
        RECT 81.820 198.330 82.140 198.390 ;
        RECT 82.295 198.330 82.585 198.375 ;
        RECT 75.930 198.190 78.830 198.330 ;
        RECT 80.070 198.190 82.585 198.330 ;
        RECT 75.930 198.035 76.070 198.190 ;
        RECT 75.855 197.805 76.145 198.035 ;
        RECT 77.695 197.990 77.985 198.035 ;
        RECT 76.850 197.850 77.985 197.990 ;
        RECT 76.850 197.355 76.990 197.850 ;
        RECT 77.695 197.805 77.985 197.850 ;
        RECT 78.140 197.790 78.460 198.050 ;
        RECT 80.070 198.035 80.210 198.190 ;
        RECT 81.820 198.130 82.140 198.190 ;
        RECT 82.295 198.145 82.585 198.190 ;
        RECT 83.200 198.130 83.520 198.390 ;
        RECT 79.995 197.805 80.285 198.035 ;
        RECT 77.235 197.650 77.525 197.695 ;
        RECT 78.230 197.650 78.370 197.790 ;
        RECT 77.235 197.510 78.370 197.650 ;
        RECT 77.235 197.465 77.525 197.510 ;
        RECT 76.775 197.310 77.065 197.355 ;
        RECT 80.455 197.310 80.745 197.355 ;
        RECT 81.360 197.310 81.680 197.370 ;
        RECT 83.290 197.355 83.430 198.130 ;
        RECT 83.750 198.035 83.890 198.530 ;
        RECT 84.120 198.530 88.120 198.670 ;
        RECT 84.120 198.470 84.440 198.530 ;
        RECT 84.595 198.485 84.885 198.530 ;
        RECT 87.800 198.470 88.120 198.530 ;
        RECT 92.400 198.670 92.720 198.730 ;
        RECT 97.000 198.670 97.320 198.730 ;
        RECT 97.935 198.670 98.225 198.715 ;
        RECT 99.300 198.670 99.620 198.730 ;
        RECT 92.400 198.530 94.930 198.670 ;
        RECT 92.400 198.470 92.720 198.530 ;
        RECT 91.020 198.330 91.340 198.390 ;
        RECT 92.860 198.330 93.180 198.390 ;
        RECT 94.240 198.330 94.560 198.390 ;
        RECT 86.970 198.190 88.950 198.330 ;
        RECT 86.970 198.035 87.110 198.190 ;
        RECT 88.810 198.050 88.950 198.190 ;
        RECT 91.020 198.190 93.180 198.330 ;
        RECT 91.020 198.130 91.340 198.190 ;
        RECT 92.860 198.130 93.180 198.190 ;
        RECT 93.415 198.190 94.560 198.330 ;
        RECT 94.790 198.330 94.930 198.530 ;
        RECT 97.000 198.530 99.620 198.670 ;
        RECT 97.000 198.470 97.320 198.530 ;
        RECT 97.935 198.485 98.225 198.530 ;
        RECT 99.300 198.470 99.620 198.530 ;
        RECT 99.760 198.670 100.080 198.730 ;
        RECT 107.580 198.670 107.900 198.730 ;
        RECT 108.055 198.670 108.345 198.715 ;
        RECT 99.760 198.530 107.350 198.670 ;
        RECT 99.760 198.470 100.080 198.530 ;
        RECT 100.220 198.330 100.540 198.390 ;
        RECT 104.375 198.330 104.665 198.375 ;
        RECT 105.280 198.330 105.600 198.390 ;
        RECT 107.210 198.330 107.350 198.530 ;
        RECT 107.580 198.530 108.345 198.670 ;
        RECT 107.580 198.470 107.900 198.530 ;
        RECT 108.055 198.485 108.345 198.530 ;
        RECT 114.480 198.470 114.800 198.730 ;
        RECT 115.875 198.670 116.165 198.715 ;
        RECT 115.875 198.530 117.470 198.670 ;
        RECT 115.875 198.485 116.165 198.530 ;
        RECT 114.570 198.330 114.710 198.470 ;
        RECT 117.330 198.330 117.470 198.530 ;
        RECT 122.760 198.470 123.080 198.730 ;
        RECT 133.340 198.670 133.660 198.730 ;
        RECT 123.770 198.530 133.660 198.670 ;
        RECT 122.850 198.330 122.990 198.470 ;
        RECT 94.790 198.190 98.610 198.330 ;
        RECT 83.675 197.805 83.965 198.035 ;
        RECT 86.895 197.805 87.185 198.035 ;
        RECT 88.260 197.790 88.580 198.050 ;
        RECT 88.720 197.790 89.040 198.050 ;
        RECT 89.180 197.990 89.500 198.050 ;
        RECT 93.415 198.035 93.555 198.190 ;
        RECT 94.240 198.130 94.560 198.190 ;
        RECT 89.655 197.990 89.945 198.035 ;
        RECT 89.180 197.850 89.945 197.990 ;
        RECT 89.180 197.790 89.500 197.850 ;
        RECT 89.655 197.805 89.945 197.850 ;
        RECT 93.335 197.805 93.625 198.035 ;
        RECT 93.795 197.805 94.085 198.035 ;
        RECT 94.700 197.990 95.020 198.050 ;
        RECT 95.175 197.990 95.465 198.035 ;
        RECT 94.700 197.850 95.465 197.990 ;
        RECT 87.340 197.650 87.660 197.710 ;
        RECT 92.875 197.650 93.165 197.695 ;
        RECT 93.870 197.650 94.010 197.805 ;
        RECT 94.700 197.790 95.020 197.850 ;
        RECT 95.175 197.805 95.465 197.850 ;
        RECT 96.540 197.990 96.860 198.050 ;
        RECT 98.470 198.035 98.610 198.190 ;
        RECT 100.220 198.190 104.130 198.330 ;
        RECT 100.220 198.130 100.540 198.190 ;
        RECT 97.015 197.990 97.305 198.035 ;
        RECT 96.540 197.850 97.305 197.990 ;
        RECT 96.540 197.790 96.860 197.850 ;
        RECT 97.015 197.805 97.305 197.850 ;
        RECT 98.395 197.805 98.685 198.035 ;
        RECT 87.340 197.510 93.165 197.650 ;
        RECT 87.340 197.450 87.660 197.510 ;
        RECT 92.875 197.465 93.165 197.510 ;
        RECT 93.535 197.510 94.010 197.650 ;
        RECT 76.775 197.170 81.680 197.310 ;
        RECT 76.775 197.125 77.065 197.170 ;
        RECT 80.455 197.125 80.745 197.170 ;
        RECT 81.360 197.110 81.680 197.170 ;
        RECT 83.215 197.125 83.505 197.355 ;
        RECT 85.975 197.310 86.265 197.355 ;
        RECT 86.880 197.310 87.200 197.370 ;
        RECT 93.535 197.310 93.675 197.510 ;
        RECT 94.255 197.465 94.545 197.695 ;
        RECT 97.090 197.650 97.230 197.805 ;
        RECT 99.300 197.790 99.620 198.050 ;
        RECT 103.455 197.805 103.745 198.035 ;
        RECT 103.990 197.990 104.130 198.190 ;
        RECT 104.375 198.190 105.970 198.330 ;
        RECT 107.210 198.190 114.250 198.330 ;
        RECT 114.570 198.190 116.320 198.330 ;
        RECT 104.375 198.145 104.665 198.190 ;
        RECT 105.280 198.130 105.600 198.190 ;
        RECT 105.830 198.035 105.970 198.190 ;
        RECT 104.835 197.990 105.125 198.035 ;
        RECT 103.990 197.850 105.125 197.990 ;
        RECT 104.835 197.805 105.125 197.850 ;
        RECT 105.755 197.805 106.045 198.035 ;
        RECT 106.215 197.805 106.505 198.035 ;
        RECT 106.675 197.990 106.965 198.035 ;
        RECT 111.720 197.990 112.040 198.050 ;
        RECT 114.110 198.035 114.250 198.190 ;
        RECT 106.675 197.850 112.040 197.990 ;
        RECT 106.675 197.805 106.965 197.850 ;
        RECT 101.140 197.650 101.460 197.710 ;
        RECT 97.090 197.510 101.460 197.650 ;
        RECT 94.330 197.310 94.470 197.465 ;
        RECT 101.140 197.450 101.460 197.510 ;
        RECT 102.075 197.465 102.365 197.695 ;
        RECT 103.530 197.650 103.670 197.805 ;
        RECT 103.900 197.650 104.220 197.710 ;
        RECT 103.530 197.510 104.220 197.650 ;
        RECT 85.975 197.170 87.200 197.310 ;
        RECT 85.975 197.125 86.265 197.170 ;
        RECT 86.880 197.110 87.200 197.170 ;
        RECT 92.950 197.170 93.675 197.310 ;
        RECT 93.870 197.170 94.470 197.310 ;
        RECT 102.150 197.310 102.290 197.465 ;
        RECT 103.900 197.450 104.220 197.510 ;
        RECT 104.360 197.650 104.680 197.710 ;
        RECT 106.290 197.650 106.430 197.805 ;
        RECT 104.360 197.510 106.430 197.650 ;
        RECT 104.360 197.450 104.680 197.510 ;
        RECT 106.750 197.310 106.890 197.805 ;
        RECT 111.720 197.790 112.040 197.850 ;
        RECT 114.035 197.990 114.325 198.035 ;
        RECT 114.955 197.990 115.245 198.035 ;
        RECT 114.035 197.850 115.245 197.990 ;
        RECT 116.180 197.990 116.320 198.190 ;
        RECT 117.330 198.190 122.990 198.330 ;
        RECT 117.330 198.035 117.470 198.190 ;
        RECT 116.180 197.850 117.010 197.990 ;
        RECT 114.035 197.805 114.325 197.850 ;
        RECT 114.955 197.805 115.245 197.850 ;
        RECT 113.560 197.650 113.880 197.710 ;
        RECT 116.335 197.650 116.625 197.695 ;
        RECT 113.560 197.510 116.625 197.650 ;
        RECT 116.870 197.650 117.010 197.850 ;
        RECT 117.255 197.805 117.545 198.035 ;
        RECT 118.160 197.990 118.480 198.050 ;
        RECT 118.635 197.990 118.925 198.035 ;
        RECT 118.160 197.850 118.925 197.990 ;
        RECT 118.160 197.790 118.480 197.850 ;
        RECT 118.635 197.805 118.925 197.850 ;
        RECT 119.080 197.990 119.400 198.050 ;
        RECT 123.770 198.035 123.910 198.530 ;
        RECT 133.340 198.470 133.660 198.530 ;
        RECT 133.800 198.670 134.120 198.730 ;
        RECT 134.275 198.670 134.565 198.715 ;
        RECT 133.800 198.530 134.565 198.670 ;
        RECT 133.800 198.470 134.120 198.530 ;
        RECT 134.275 198.485 134.565 198.530 ;
        RECT 143.000 198.470 143.320 198.730 ;
        RECT 145.760 198.470 146.080 198.730 ;
        RECT 146.235 198.670 146.525 198.715 ;
        RECT 146.680 198.670 147.000 198.730 ;
        RECT 146.235 198.530 147.000 198.670 ;
        RECT 146.235 198.485 146.525 198.530 ;
        RECT 146.680 198.470 147.000 198.530 ;
        RECT 148.520 198.470 148.840 198.730 ;
        RECT 153.120 198.470 153.440 198.730 ;
        RECT 126.915 198.330 127.205 198.375 ;
        RECT 127.820 198.330 128.140 198.390 ;
        RECT 126.915 198.190 128.140 198.330 ;
        RECT 126.915 198.145 127.205 198.190 ;
        RECT 127.820 198.130 128.140 198.190 ;
        RECT 128.740 198.330 129.060 198.390 ;
        RECT 128.740 198.190 135.870 198.330 ;
        RECT 128.740 198.130 129.060 198.190 ;
        RECT 123.695 197.990 123.985 198.035 ;
        RECT 119.080 197.850 123.985 197.990 ;
        RECT 119.080 197.790 119.400 197.850 ;
        RECT 123.695 197.805 123.985 197.850 ;
        RECT 125.520 197.990 125.840 198.050 ;
        RECT 126.455 197.990 126.745 198.035 ;
        RECT 125.520 197.850 126.745 197.990 ;
        RECT 125.520 197.790 125.840 197.850 ;
        RECT 126.455 197.805 126.745 197.850 ;
        RECT 127.375 197.990 127.665 198.035 ;
        RECT 129.660 197.990 129.980 198.050 ;
        RECT 131.500 197.990 131.820 198.050 ;
        RECT 127.375 197.850 129.980 197.990 ;
        RECT 127.375 197.805 127.665 197.850 ;
        RECT 129.660 197.790 129.980 197.850 ;
        RECT 130.210 197.850 131.820 197.990 ;
        RECT 124.600 197.650 124.920 197.710 ;
        RECT 116.870 197.510 124.920 197.650 ;
        RECT 113.560 197.450 113.880 197.510 ;
        RECT 116.335 197.465 116.625 197.510 ;
        RECT 124.600 197.450 124.920 197.510 ;
        RECT 125.075 197.650 125.365 197.695 ;
        RECT 130.210 197.650 130.350 197.850 ;
        RECT 131.500 197.790 131.820 197.850 ;
        RECT 131.975 197.805 132.265 198.035 ;
        RECT 132.435 197.990 132.725 198.035 ;
        RECT 133.340 197.990 133.660 198.050 ;
        RECT 135.730 198.035 135.870 198.190 ;
        RECT 138.950 198.190 144.150 198.330 ;
        RECT 132.435 197.850 133.660 197.990 ;
        RECT 132.435 197.805 132.725 197.850 ;
        RECT 125.075 197.510 130.350 197.650 ;
        RECT 125.075 197.465 125.365 197.510 ;
        RECT 130.595 197.465 130.885 197.695 ;
        RECT 102.150 197.170 106.890 197.310 ;
        RECT 92.950 197.030 93.090 197.170 ;
        RECT 93.870 197.030 94.010 197.170 ;
        RECT 117.700 197.110 118.020 197.370 ;
        RECT 118.175 197.310 118.465 197.355 ;
        RECT 123.680 197.310 124.000 197.370 ;
        RECT 118.175 197.170 124.000 197.310 ;
        RECT 118.175 197.125 118.465 197.170 ;
        RECT 123.680 197.110 124.000 197.170 ;
        RECT 125.980 197.310 126.300 197.370 ;
        RECT 130.670 197.310 130.810 197.465 ;
        RECT 132.050 197.370 132.190 197.805 ;
        RECT 133.340 197.790 133.660 197.850 ;
        RECT 135.655 197.805 135.945 198.035 ;
        RECT 137.480 197.790 137.800 198.050 ;
        RECT 138.950 198.035 139.090 198.190 ;
        RECT 144.010 198.050 144.150 198.190 ;
        RECT 138.875 197.805 139.165 198.035 ;
        RECT 139.320 197.990 139.640 198.050 ;
        RECT 140.255 197.990 140.545 198.035 ;
        RECT 142.095 197.990 142.385 198.035 ;
        RECT 139.320 197.850 140.545 197.990 ;
        RECT 139.320 197.790 139.640 197.850 ;
        RECT 140.255 197.805 140.545 197.850 ;
        RECT 140.790 197.850 142.385 197.990 ;
        RECT 140.790 197.710 140.930 197.850 ;
        RECT 142.095 197.805 142.385 197.850 ;
        RECT 143.920 197.790 144.240 198.050 ;
        RECT 145.315 197.990 145.605 198.035 ;
        RECT 145.850 197.990 145.990 198.470 ;
        RECT 145.315 197.850 145.990 197.990 ;
        RECT 147.615 197.990 147.905 198.035 ;
        RECT 148.610 197.990 148.750 198.470 ;
        RECT 147.615 197.850 148.750 197.990 ;
        RECT 152.675 197.990 152.965 198.035 ;
        RECT 153.210 197.990 153.350 198.470 ;
        RECT 154.055 197.990 154.345 198.035 ;
        RECT 152.675 197.850 154.345 197.990 ;
        RECT 145.315 197.805 145.605 197.850 ;
        RECT 147.615 197.805 147.905 197.850 ;
        RECT 152.675 197.805 152.965 197.850 ;
        RECT 154.055 197.805 154.345 197.850 ;
        RECT 132.880 197.450 133.200 197.710 ;
        RECT 140.700 197.450 141.020 197.710 ;
        RECT 141.635 197.650 141.925 197.695 ;
        RECT 148.060 197.650 148.380 197.710 ;
        RECT 141.635 197.510 148.380 197.650 ;
        RECT 141.635 197.465 141.925 197.510 ;
        RECT 148.060 197.450 148.380 197.510 ;
        RECT 125.980 197.170 130.810 197.310 ;
        RECT 125.980 197.110 126.300 197.170 ;
        RECT 131.960 197.110 132.280 197.370 ;
        RECT 134.260 197.310 134.580 197.370 ;
        RECT 134.735 197.310 135.025 197.355 ;
        RECT 134.260 197.170 135.025 197.310 ;
        RECT 134.260 197.110 134.580 197.170 ;
        RECT 134.735 197.125 135.025 197.170 ;
        RECT 135.180 197.310 135.500 197.370 ;
        RECT 137.480 197.310 137.800 197.370 ;
        RECT 138.415 197.310 138.705 197.355 ;
        RECT 135.180 197.170 138.705 197.310 ;
        RECT 135.180 197.110 135.500 197.170 ;
        RECT 137.480 197.110 137.800 197.170 ;
        RECT 138.415 197.125 138.705 197.170 ;
        RECT 138.860 197.310 139.180 197.370 ;
        RECT 141.175 197.310 141.465 197.355 ;
        RECT 138.860 197.170 141.465 197.310 ;
        RECT 138.860 197.110 139.180 197.170 ;
        RECT 141.175 197.125 141.465 197.170 ;
        RECT 145.300 197.310 145.620 197.370 ;
        RECT 153.135 197.310 153.425 197.355 ;
        RECT 145.300 197.170 153.425 197.310 ;
        RECT 145.300 197.110 145.620 197.170 ;
        RECT 82.280 196.770 82.600 197.030 ;
        RECT 85.500 196.970 85.820 197.030 ;
        RECT 87.355 196.970 87.645 197.015 ;
        RECT 85.500 196.830 87.645 196.970 ;
        RECT 85.500 196.770 85.820 196.830 ;
        RECT 87.355 196.785 87.645 196.830 ;
        RECT 88.720 196.770 89.040 197.030 ;
        RECT 89.180 196.970 89.500 197.030 ;
        RECT 90.575 196.970 90.865 197.015 ;
        RECT 89.180 196.830 90.865 196.970 ;
        RECT 89.180 196.770 89.500 196.830 ;
        RECT 90.575 196.785 90.865 196.830 ;
        RECT 91.940 196.770 92.260 197.030 ;
        RECT 92.860 196.770 93.180 197.030 ;
        RECT 93.780 196.770 94.100 197.030 ;
        RECT 96.080 196.770 96.400 197.030 ;
        RECT 98.855 196.970 99.145 197.015 ;
        RECT 102.535 196.970 102.825 197.015 ;
        RECT 98.855 196.830 102.825 196.970 ;
        RECT 98.855 196.785 99.145 196.830 ;
        RECT 102.535 196.785 102.825 196.830 ;
        RECT 107.580 196.970 107.900 197.030 ;
        RECT 110.800 196.970 111.120 197.030 ;
        RECT 107.580 196.830 111.120 196.970 ;
        RECT 107.580 196.770 107.900 196.830 ;
        RECT 110.800 196.770 111.120 196.830 ;
        RECT 112.180 196.970 112.500 197.030 ;
        RECT 113.115 196.970 113.405 197.015 ;
        RECT 117.790 196.970 117.930 197.110 ;
        RECT 147.690 197.030 147.830 197.170 ;
        RECT 153.135 197.125 153.425 197.170 ;
        RECT 112.180 196.830 117.930 196.970 ;
        RECT 118.620 196.970 118.940 197.030 ;
        RECT 122.775 196.970 123.065 197.015 ;
        RECT 118.620 196.830 123.065 196.970 ;
        RECT 112.180 196.770 112.500 196.830 ;
        RECT 113.115 196.785 113.405 196.830 ;
        RECT 118.620 196.770 118.940 196.830 ;
        RECT 122.775 196.785 123.065 196.830 ;
        RECT 131.500 196.970 131.820 197.030 ;
        RECT 132.435 196.970 132.725 197.015 ;
        RECT 131.500 196.830 132.725 196.970 ;
        RECT 131.500 196.770 131.820 196.830 ;
        RECT 132.435 196.785 132.725 196.830 ;
        RECT 132.880 196.970 133.200 197.030 ;
        RECT 136.575 196.970 136.865 197.015 ;
        RECT 132.880 196.830 136.865 196.970 ;
        RECT 132.880 196.770 133.200 196.830 ;
        RECT 136.575 196.785 136.865 196.830 ;
        RECT 139.320 196.770 139.640 197.030 ;
        RECT 143.460 196.970 143.780 197.030 ;
        RECT 146.695 196.970 146.985 197.015 ;
        RECT 143.460 196.830 146.985 196.970 ;
        RECT 143.460 196.770 143.780 196.830 ;
        RECT 146.695 196.785 146.985 196.830 ;
        RECT 147.600 196.770 147.920 197.030 ;
        RECT 152.200 196.770 152.520 197.030 ;
        RECT 70.710 196.150 156.270 196.630 ;
        RECT 81.360 195.750 81.680 196.010 ;
        RECT 82.295 195.950 82.585 195.995 ;
        RECT 82.740 195.950 83.060 196.010 ;
        RECT 85.500 195.950 85.820 196.010 ;
        RECT 93.780 195.950 94.100 196.010 ;
        RECT 82.295 195.810 85.820 195.950 ;
        RECT 82.295 195.765 82.585 195.810 ;
        RECT 82.740 195.750 83.060 195.810 ;
        RECT 85.500 195.750 85.820 195.810 ;
        RECT 88.350 195.810 94.100 195.950 ;
        RECT 72.660 195.610 72.950 195.655 ;
        RECT 74.760 195.610 75.050 195.655 ;
        RECT 76.330 195.610 76.620 195.655 ;
        RECT 72.660 195.470 76.620 195.610 ;
        RECT 72.660 195.425 72.950 195.470 ;
        RECT 74.760 195.425 75.050 195.470 ;
        RECT 76.330 195.425 76.620 195.470 ;
        RECT 79.075 195.610 79.365 195.655 ;
        RECT 83.660 195.610 83.980 195.670 ;
        RECT 84.135 195.610 84.425 195.655 ;
        RECT 79.075 195.470 82.970 195.610 ;
        RECT 79.075 195.425 79.365 195.470 ;
        RECT 73.055 195.270 73.345 195.315 ;
        RECT 74.245 195.270 74.535 195.315 ;
        RECT 76.765 195.270 77.055 195.315 ;
        RECT 73.055 195.130 77.055 195.270 ;
        RECT 73.055 195.085 73.345 195.130 ;
        RECT 74.245 195.085 74.535 195.130 ;
        RECT 76.765 195.085 77.055 195.130 ;
        RECT 72.160 194.730 72.480 194.990 ;
        RECT 73.510 194.590 73.800 194.635 ;
        RECT 74.920 194.590 75.240 194.650 ;
        RECT 73.510 194.450 75.240 194.590 ;
        RECT 73.510 194.405 73.800 194.450 ;
        RECT 74.920 194.390 75.240 194.450 ;
        RECT 78.140 194.250 78.460 194.310 ;
        RECT 82.165 194.250 82.455 194.295 ;
        RECT 78.140 194.110 82.455 194.250 ;
        RECT 82.830 194.250 82.970 195.470 ;
        RECT 83.660 195.470 84.425 195.610 ;
        RECT 83.660 195.410 83.980 195.470 ;
        RECT 84.135 195.425 84.425 195.470 ;
        RECT 85.500 195.070 85.820 195.330 ;
        RECT 88.350 195.270 88.490 195.810 ;
        RECT 93.780 195.750 94.100 195.810 ;
        RECT 97.920 195.950 98.240 196.010 ;
        RECT 100.680 195.950 101.000 196.010 ;
        RECT 97.920 195.810 101.000 195.950 ;
        RECT 97.920 195.750 98.240 195.810 ;
        RECT 100.680 195.750 101.000 195.810 ;
        RECT 105.755 195.950 106.045 195.995 ;
        RECT 106.200 195.950 106.520 196.010 ;
        RECT 105.755 195.810 106.520 195.950 ;
        RECT 105.755 195.765 106.045 195.810 ;
        RECT 106.200 195.750 106.520 195.810 ;
        RECT 107.135 195.765 107.425 195.995 ;
        RECT 108.975 195.950 109.265 195.995 ;
        RECT 108.975 195.810 109.650 195.950 ;
        RECT 108.975 195.765 109.265 195.810 ;
        RECT 88.735 195.610 89.025 195.655 ;
        RECT 89.180 195.610 89.500 195.670 ;
        RECT 101.140 195.610 101.460 195.670 ;
        RECT 107.210 195.610 107.350 195.765 ;
        RECT 108.040 195.610 108.360 195.670 ;
        RECT 88.735 195.470 89.500 195.610 ;
        RECT 88.735 195.425 89.025 195.470 ;
        RECT 89.180 195.410 89.500 195.470 ;
        RECT 92.030 195.470 99.530 195.610 ;
        RECT 92.030 195.270 92.170 195.470 ;
        RECT 86.050 195.130 88.490 195.270 ;
        RECT 85.040 194.730 85.360 194.990 ;
        RECT 86.050 194.975 86.190 195.130 ;
        RECT 85.975 194.745 86.265 194.975 ;
        RECT 86.435 194.930 86.725 194.975 ;
        RECT 87.355 194.930 87.645 194.975 ;
        RECT 86.435 194.790 87.645 194.930 ;
        RECT 86.435 194.745 86.725 194.790 ;
        RECT 87.355 194.745 87.645 194.790 ;
        RECT 87.800 194.730 88.120 194.990 ;
        RECT 88.350 194.975 88.490 195.130 ;
        RECT 89.270 195.130 92.170 195.270 ;
        RECT 88.275 194.745 88.565 194.975 ;
        RECT 88.720 194.930 89.040 194.990 ;
        RECT 89.270 194.975 89.410 195.130 ;
        RECT 92.400 195.070 92.720 195.330 ;
        RECT 93.460 195.270 93.750 195.315 ;
        RECT 95.620 195.270 95.940 195.330 ;
        RECT 96.095 195.270 96.385 195.315 ;
        RECT 98.380 195.270 98.700 195.330 ;
        RECT 93.460 195.130 98.700 195.270 ;
        RECT 93.460 195.085 93.750 195.130 ;
        RECT 95.620 195.070 95.940 195.130 ;
        RECT 96.095 195.085 96.385 195.130 ;
        RECT 98.380 195.070 98.700 195.130 ;
        RECT 98.840 195.070 99.160 195.330 ;
        RECT 99.390 195.270 99.530 195.470 ;
        RECT 101.140 195.470 106.430 195.610 ;
        RECT 107.210 195.470 108.360 195.610 ;
        RECT 101.140 195.410 101.460 195.470 ;
        RECT 104.820 195.270 105.140 195.330 ;
        RECT 99.390 195.130 105.140 195.270 ;
        RECT 104.820 195.070 105.140 195.130 ;
        RECT 89.195 194.930 89.485 194.975 ;
        RECT 88.720 194.790 89.485 194.930 ;
        RECT 88.720 194.730 89.040 194.790 ;
        RECT 89.195 194.745 89.485 194.790 ;
        RECT 89.655 194.745 89.945 194.975 ;
        RECT 91.035 194.930 91.325 194.975 ;
        RECT 94.240 194.930 94.560 194.990 ;
        RECT 97.000 194.930 97.320 194.990 ;
        RECT 91.035 194.790 97.320 194.930 ;
        RECT 91.035 194.745 91.325 194.790 ;
        RECT 83.215 194.590 83.505 194.635 ;
        RECT 86.880 194.590 87.200 194.650 ;
        RECT 83.215 194.450 87.200 194.590 ;
        RECT 87.890 194.590 88.030 194.730 ;
        RECT 89.730 194.590 89.870 194.745 ;
        RECT 94.240 194.730 94.560 194.790 ;
        RECT 97.000 194.730 97.320 194.790 ;
        RECT 97.935 194.930 98.225 194.975 ;
        RECT 99.300 194.930 99.620 194.990 ;
        RECT 97.935 194.790 99.620 194.930 ;
        RECT 97.935 194.745 98.225 194.790 ;
        RECT 99.300 194.730 99.620 194.790 ;
        RECT 100.680 194.930 101.000 194.990 ;
        RECT 101.600 194.930 101.920 194.990 ;
        RECT 102.520 194.930 102.840 194.990 ;
        RECT 106.290 194.975 106.430 195.470 ;
        RECT 108.040 195.410 108.360 195.470 ;
        RECT 102.995 194.930 103.285 194.975 ;
        RECT 100.680 194.790 103.285 194.930 ;
        RECT 100.680 194.730 101.000 194.790 ;
        RECT 101.600 194.730 101.920 194.790 ;
        RECT 102.520 194.730 102.840 194.790 ;
        RECT 102.995 194.745 103.285 194.790 ;
        RECT 106.215 194.745 106.505 194.975 ;
        RECT 106.660 194.940 106.980 194.990 ;
        RECT 109.510 194.980 109.650 195.810 ;
        RECT 110.800 195.750 111.120 196.010 ;
        RECT 111.720 195.750 112.040 196.010 ;
        RECT 135.180 195.950 135.500 196.010 ;
        RECT 116.180 195.810 135.500 195.950 ;
        RECT 109.880 195.410 110.200 195.670 ;
        RECT 110.890 195.610 111.030 195.750 ;
        RECT 116.180 195.610 116.320 195.810 ;
        RECT 135.180 195.750 135.500 195.810 ;
        RECT 136.575 195.950 136.865 195.995 ;
        RECT 137.480 195.950 137.800 196.010 ;
        RECT 136.575 195.810 137.800 195.950 ;
        RECT 136.575 195.765 136.865 195.810 ;
        RECT 137.480 195.750 137.800 195.810 ;
        RECT 141.175 195.950 141.465 195.995 ;
        RECT 143.000 195.950 143.320 196.010 ;
        RECT 141.175 195.810 143.320 195.950 ;
        RECT 141.175 195.765 141.465 195.810 ;
        RECT 143.000 195.750 143.320 195.810 ;
        RECT 144.840 195.750 145.160 196.010 ;
        RECT 110.890 195.470 116.320 195.610 ;
        RECT 126.900 195.410 127.220 195.670 ;
        RECT 128.280 195.610 128.570 195.655 ;
        RECT 129.850 195.610 130.140 195.655 ;
        RECT 131.950 195.610 132.240 195.655 ;
        RECT 128.280 195.470 132.240 195.610 ;
        RECT 128.280 195.425 128.570 195.470 ;
        RECT 129.850 195.425 130.140 195.470 ;
        RECT 131.950 195.425 132.240 195.470 ;
        RECT 132.420 195.610 132.740 195.670 ;
        RECT 137.955 195.610 138.245 195.655 ;
        RECT 140.700 195.610 141.020 195.670 ;
        RECT 132.420 195.470 141.020 195.610 ;
        RECT 132.420 195.410 132.740 195.470 ;
        RECT 137.955 195.425 138.245 195.470 ;
        RECT 109.970 195.270 110.110 195.410 ;
        RECT 118.160 195.270 118.480 195.330 ;
        RECT 109.970 195.130 118.480 195.270 ;
        RECT 118.160 195.070 118.480 195.130 ;
        RECT 109.510 194.975 110.110 194.980 ;
        RECT 106.660 194.930 107.350 194.940 ;
        RECT 107.595 194.930 107.885 194.975 ;
        RECT 106.660 194.800 107.885 194.930 ;
        RECT 109.510 194.840 110.185 194.975 ;
        RECT 106.660 194.730 106.980 194.800 ;
        RECT 107.210 194.790 107.885 194.800 ;
        RECT 107.595 194.745 107.885 194.790 ;
        RECT 109.895 194.745 110.185 194.840 ;
        RECT 110.800 194.730 111.120 194.990 ;
        RECT 112.180 194.930 112.500 194.990 ;
        RECT 115.860 194.930 116.180 194.990 ;
        RECT 124.615 194.930 124.905 194.975 ;
        RECT 126.990 194.930 127.130 195.410 ;
        RECT 138.950 195.330 139.090 195.470 ;
        RECT 140.700 195.410 141.020 195.470 ;
        RECT 141.620 195.610 141.940 195.670 ;
        RECT 144.930 195.610 145.070 195.750 ;
        RECT 141.620 195.470 145.070 195.610 ;
        RECT 147.640 195.610 147.930 195.655 ;
        RECT 149.740 195.610 150.030 195.655 ;
        RECT 151.310 195.610 151.600 195.655 ;
        RECT 147.640 195.470 151.600 195.610 ;
        RECT 141.620 195.410 141.940 195.470 ;
        RECT 147.640 195.425 147.930 195.470 ;
        RECT 149.740 195.425 150.030 195.470 ;
        RECT 151.310 195.425 151.600 195.470 ;
        RECT 127.845 195.270 128.135 195.315 ;
        RECT 130.365 195.270 130.655 195.315 ;
        RECT 131.555 195.270 131.845 195.315 ;
        RECT 127.845 195.130 131.845 195.270 ;
        RECT 127.845 195.085 128.135 195.130 ;
        RECT 130.365 195.085 130.655 195.130 ;
        RECT 131.555 195.085 131.845 195.130 ;
        RECT 134.260 195.070 134.580 195.330 ;
        RECT 138.860 195.070 139.180 195.330 ;
        RECT 139.780 195.270 140.100 195.330 ;
        RECT 147.155 195.270 147.445 195.315 ;
        RECT 139.780 195.130 147.445 195.270 ;
        RECT 139.780 195.070 140.100 195.130 ;
        RECT 147.155 195.085 147.445 195.130 ;
        RECT 148.035 195.270 148.325 195.315 ;
        RECT 149.225 195.270 149.515 195.315 ;
        RECT 151.745 195.270 152.035 195.315 ;
        RECT 148.035 195.130 152.035 195.270 ;
        RECT 148.035 195.085 148.325 195.130 ;
        RECT 149.225 195.085 149.515 195.130 ;
        RECT 151.745 195.085 152.035 195.130 ;
        RECT 112.180 194.790 124.370 194.930 ;
        RECT 112.180 194.730 112.500 194.790 ;
        RECT 115.860 194.730 116.180 194.790 ;
        RECT 87.890 194.450 89.870 194.590 ;
        RECT 95.510 194.590 95.800 194.635 ;
        RECT 99.760 194.590 100.080 194.650 ;
        RECT 95.510 194.450 100.080 194.590 ;
        RECT 83.215 194.405 83.505 194.450 ;
        RECT 86.880 194.390 87.200 194.450 ;
        RECT 95.510 194.405 95.800 194.450 ;
        RECT 99.760 194.390 100.080 194.450 ;
        RECT 104.375 194.590 104.665 194.635 ;
        RECT 108.960 194.590 109.280 194.650 ;
        RECT 104.375 194.450 117.470 194.590 ;
        RECT 104.375 194.405 104.665 194.450 ;
        RECT 108.960 194.390 109.280 194.450 ;
        RECT 117.330 194.310 117.470 194.450 ;
        RECT 86.420 194.250 86.740 194.310 ;
        RECT 91.020 194.250 91.340 194.310 ;
        RECT 82.830 194.110 91.340 194.250 ;
        RECT 78.140 194.050 78.460 194.110 ;
        RECT 82.165 194.065 82.455 194.110 ;
        RECT 86.420 194.050 86.740 194.110 ;
        RECT 91.020 194.050 91.340 194.110 ;
        RECT 92.860 194.050 93.180 194.310 ;
        RECT 94.240 194.050 94.560 194.310 ;
        RECT 94.700 194.050 95.020 194.310 ;
        RECT 96.555 194.250 96.845 194.295 ;
        RECT 97.920 194.250 98.240 194.310 ;
        RECT 96.555 194.110 98.240 194.250 ;
        RECT 96.555 194.065 96.845 194.110 ;
        RECT 97.920 194.050 98.240 194.110 ;
        RECT 100.680 194.250 101.000 194.310 ;
        RECT 102.075 194.250 102.365 194.295 ;
        RECT 100.680 194.110 102.365 194.250 ;
        RECT 100.680 194.050 101.000 194.110 ;
        RECT 102.075 194.065 102.365 194.110 ;
        RECT 103.440 194.250 103.760 194.310 ;
        RECT 103.915 194.250 104.205 194.295 ;
        RECT 103.440 194.110 104.205 194.250 ;
        RECT 103.440 194.050 103.760 194.110 ;
        RECT 103.915 194.065 104.205 194.110 ;
        RECT 104.820 194.050 105.140 194.310 ;
        RECT 117.240 194.050 117.560 194.310 ;
        RECT 124.230 194.295 124.370 194.790 ;
        RECT 124.615 194.790 127.130 194.930 ;
        RECT 127.360 194.930 127.680 194.990 ;
        RECT 129.200 194.930 129.520 194.990 ;
        RECT 127.360 194.790 129.520 194.930 ;
        RECT 124.615 194.745 124.905 194.790 ;
        RECT 127.360 194.730 127.680 194.790 ;
        RECT 129.200 194.730 129.520 194.790 ;
        RECT 129.980 194.790 131.730 194.930 ;
        RECT 129.980 194.650 130.120 194.790 ;
        RECT 129.660 194.590 130.120 194.650 ;
        RECT 131.040 194.635 131.360 194.650 ;
        RECT 131.040 194.590 131.390 194.635 ;
        RECT 125.610 194.450 130.120 194.590 ;
        RECT 130.890 194.450 131.390 194.590 ;
        RECT 131.590 194.590 131.730 194.790 ;
        RECT 132.420 194.730 132.740 194.990 ;
        RECT 133.815 194.745 134.105 194.975 ;
        RECT 134.350 194.930 134.490 195.070 ;
        RECT 135.655 194.930 135.945 194.975 ;
        RECT 134.350 194.790 135.945 194.930 ;
        RECT 135.655 194.745 135.945 194.790 ;
        RECT 137.035 194.745 137.325 194.975 ;
        RECT 137.940 194.930 138.260 194.990 ;
        RECT 139.335 194.930 139.625 194.975 ;
        RECT 137.940 194.790 139.625 194.930 ;
        RECT 133.890 194.590 134.030 194.745 ;
        RECT 131.590 194.450 134.030 194.590 ;
        RECT 124.155 194.250 124.445 194.295 ;
        RECT 125.060 194.250 125.380 194.310 ;
        RECT 125.610 194.295 125.750 194.450 ;
        RECT 129.660 194.390 129.980 194.450 ;
        RECT 131.040 194.405 131.390 194.450 ;
        RECT 131.040 194.390 131.360 194.405 ;
        RECT 135.180 194.390 135.500 194.650 ;
        RECT 137.110 194.590 137.250 194.745 ;
        RECT 137.940 194.730 138.260 194.790 ;
        RECT 139.335 194.745 139.625 194.790 ;
        RECT 140.700 194.730 141.020 194.990 ;
        RECT 145.315 194.930 145.605 194.975 ;
        RECT 142.170 194.790 145.605 194.930 ;
        RECT 137.480 194.590 137.800 194.650 ;
        RECT 140.790 194.590 140.930 194.730 ;
        RECT 137.110 194.450 140.930 194.590 ;
        RECT 137.480 194.390 137.800 194.450 ;
        RECT 124.155 194.110 125.380 194.250 ;
        RECT 124.155 194.065 124.445 194.110 ;
        RECT 125.060 194.050 125.380 194.110 ;
        RECT 125.535 194.065 125.825 194.295 ;
        RECT 126.440 194.250 126.760 194.310 ;
        RECT 132.895 194.250 133.185 194.295 ;
        RECT 133.340 194.250 133.660 194.310 ;
        RECT 126.440 194.110 133.660 194.250 ;
        RECT 135.270 194.250 135.410 194.390 ;
        RECT 138.400 194.250 138.720 194.310 ;
        RECT 142.170 194.295 142.310 194.790 ;
        RECT 145.315 194.745 145.605 194.790 ;
        RECT 148.380 194.590 148.670 194.635 ;
        RECT 146.310 194.450 148.670 194.590 ;
        RECT 146.310 194.295 146.450 194.450 ;
        RECT 148.380 194.405 148.670 194.450 ;
        RECT 141.175 194.250 141.465 194.295 ;
        RECT 135.270 194.110 141.465 194.250 ;
        RECT 126.440 194.050 126.760 194.110 ;
        RECT 132.895 194.065 133.185 194.110 ;
        RECT 133.340 194.050 133.660 194.110 ;
        RECT 138.400 194.050 138.720 194.110 ;
        RECT 141.175 194.065 141.465 194.110 ;
        RECT 142.095 194.065 142.385 194.295 ;
        RECT 146.235 194.065 146.525 194.295 ;
        RECT 153.120 194.250 153.440 194.310 ;
        RECT 154.055 194.250 154.345 194.295 ;
        RECT 153.120 194.110 154.345 194.250 ;
        RECT 153.120 194.050 153.440 194.110 ;
        RECT 154.055 194.065 154.345 194.110 ;
        RECT 70.710 193.430 156.270 193.910 ;
        RECT 74.920 193.230 75.240 193.290 ;
        RECT 77.265 193.230 77.555 193.275 ;
        RECT 74.920 193.090 77.555 193.230 ;
        RECT 74.920 193.030 75.240 193.090 ;
        RECT 77.265 193.045 77.555 193.090 ;
        RECT 79.995 193.230 80.285 193.275 ;
        RECT 82.280 193.230 82.600 193.290 ;
        RECT 79.995 193.090 82.600 193.230 ;
        RECT 79.995 193.045 80.285 193.090 ;
        RECT 82.280 193.030 82.600 193.090 ;
        RECT 85.500 193.230 85.820 193.290 ;
        RECT 89.195 193.230 89.485 193.275 ;
        RECT 93.320 193.230 93.640 193.290 ;
        RECT 85.500 193.090 89.485 193.230 ;
        RECT 85.500 193.030 85.820 193.090 ;
        RECT 89.195 193.045 89.485 193.090 ;
        RECT 89.885 193.090 93.640 193.230 ;
        RECT 76.315 192.890 76.605 192.935 ;
        RECT 76.775 192.890 77.065 192.935 ;
        RECT 76.315 192.750 77.065 192.890 ;
        RECT 76.315 192.705 76.605 192.750 ;
        RECT 76.775 192.705 77.065 192.750 ;
        RECT 77.695 192.890 77.985 192.935 ;
        RECT 77.695 192.750 83.430 192.890 ;
        RECT 77.695 192.705 77.985 192.750 ;
        RECT 74.935 192.550 75.225 192.595 ;
        RECT 77.770 192.550 77.910 192.705 ;
        RECT 74.935 192.410 77.910 192.550 ;
        RECT 74.935 192.365 75.225 192.410 ;
        RECT 78.140 192.350 78.460 192.610 ;
        RECT 80.440 192.550 80.760 192.610 ;
        RECT 81.360 192.550 81.680 192.610 ;
        RECT 81.910 192.595 82.050 192.750 ;
        RECT 80.440 192.410 81.680 192.550 ;
        RECT 80.440 192.350 80.760 192.410 ;
        RECT 81.360 192.350 81.680 192.410 ;
        RECT 81.835 192.365 82.125 192.595 ;
        RECT 82.740 192.550 83.060 192.610 ;
        RECT 82.370 192.410 83.060 192.550 ;
        RECT 76.315 192.210 76.605 192.255 ;
        RECT 76.760 192.210 77.080 192.270 ;
        RECT 78.230 192.210 78.370 192.350 ;
        RECT 76.315 192.070 77.080 192.210 ;
        RECT 76.315 192.025 76.605 192.070 ;
        RECT 76.760 192.010 77.080 192.070 ;
        RECT 77.310 192.070 78.370 192.210 ;
        RECT 77.310 191.590 77.450 192.070 ;
        RECT 80.900 192.010 81.220 192.270 ;
        RECT 82.370 192.255 82.510 192.410 ;
        RECT 82.740 192.350 83.060 192.410 ;
        RECT 82.295 192.025 82.585 192.255 ;
        RECT 83.290 192.210 83.430 192.750 ;
        RECT 86.880 192.550 87.200 192.610 ;
        RECT 87.355 192.550 87.645 192.595 ;
        RECT 89.885 192.550 90.025 193.090 ;
        RECT 93.320 193.030 93.640 193.090 ;
        RECT 94.240 193.230 94.560 193.290 ;
        RECT 104.820 193.230 105.140 193.290 ;
        RECT 105.755 193.230 106.045 193.275 ;
        RECT 94.240 193.090 102.750 193.230 ;
        RECT 94.240 193.030 94.560 193.090 ;
        RECT 90.560 192.690 90.880 192.950 ;
        RECT 92.875 192.890 93.165 192.935 ;
        RECT 93.410 192.890 93.550 193.030 ;
        RECT 92.875 192.750 93.550 192.890 ;
        RECT 94.715 192.890 95.005 192.935 ;
        RECT 95.620 192.890 95.940 192.950 ;
        RECT 94.715 192.750 95.940 192.890 ;
        RECT 92.875 192.705 93.165 192.750 ;
        RECT 94.715 192.705 95.005 192.750 ;
        RECT 95.620 192.690 95.940 192.750 ;
        RECT 96.080 192.890 96.400 192.950 ;
        RECT 98.395 192.890 98.685 192.935 ;
        RECT 99.300 192.890 99.620 192.950 ;
        RECT 96.080 192.750 99.620 192.890 ;
        RECT 96.080 192.690 96.400 192.750 ;
        RECT 98.395 192.705 98.685 192.750 ;
        RECT 99.300 192.690 99.620 192.750 ;
        RECT 100.695 192.705 100.985 192.935 ;
        RECT 86.880 192.410 90.025 192.550 ;
        RECT 86.880 192.350 87.200 192.410 ;
        RECT 87.355 192.365 87.645 192.410 ;
        RECT 91.020 192.350 91.340 192.610 ;
        RECT 93.320 192.550 93.640 192.610 ;
        RECT 97.000 192.550 97.320 192.610 ;
        RECT 100.770 192.550 100.910 192.705 ;
        RECT 102.610 192.595 102.750 193.090 ;
        RECT 104.820 193.090 106.045 193.230 ;
        RECT 104.820 193.030 105.140 193.090 ;
        RECT 105.755 193.045 106.045 193.090 ;
        RECT 106.200 193.230 106.520 193.290 ;
        RECT 110.800 193.230 111.120 193.290 ;
        RECT 106.200 193.090 111.120 193.230 ;
        RECT 106.200 193.030 106.520 193.090 ;
        RECT 107.135 192.890 107.425 192.935 ;
        RECT 107.580 192.890 107.900 192.950 ;
        RECT 108.590 192.935 108.730 193.090 ;
        RECT 110.800 193.030 111.120 193.090 ;
        RECT 111.720 193.230 112.040 193.290 ;
        RECT 113.575 193.230 113.865 193.275 ;
        RECT 111.720 193.090 113.865 193.230 ;
        RECT 111.720 193.030 112.040 193.090 ;
        RECT 113.575 193.045 113.865 193.090 ;
        RECT 114.020 193.230 114.340 193.290 ;
        RECT 128.740 193.230 129.060 193.290 ;
        RECT 114.020 193.090 129.060 193.230 ;
        RECT 114.020 193.030 114.340 193.090 ;
        RECT 128.740 193.030 129.060 193.090 ;
        RECT 129.660 193.230 129.980 193.290 ;
        RECT 130.595 193.230 130.885 193.275 ;
        RECT 129.660 193.090 130.885 193.230 ;
        RECT 129.660 193.030 129.980 193.090 ;
        RECT 130.595 193.045 130.885 193.090 ;
        RECT 137.065 193.230 137.355 193.275 ;
        RECT 137.065 193.090 138.630 193.230 ;
        RECT 137.065 193.045 137.355 193.090 ;
        RECT 104.910 192.750 107.900 192.890 ;
        RECT 104.910 192.595 105.050 192.750 ;
        RECT 107.135 192.705 107.425 192.750 ;
        RECT 107.580 192.690 107.900 192.750 ;
        RECT 108.515 192.705 108.805 192.935 ;
        RECT 108.975 192.890 109.265 192.935 ;
        RECT 108.975 192.750 114.250 192.890 ;
        RECT 108.975 192.705 109.265 192.750 ;
        RECT 93.320 192.410 95.390 192.550 ;
        RECT 93.320 192.350 93.640 192.410 ;
        RECT 85.975 192.210 86.265 192.255 ;
        RECT 82.830 192.070 86.265 192.210 ;
        RECT 82.830 191.590 82.970 192.070 ;
        RECT 85.975 192.025 86.265 192.070 ;
        RECT 88.275 192.210 88.565 192.255 ;
        RECT 89.195 192.210 89.485 192.255 ;
        RECT 92.400 192.210 92.720 192.270 ;
        RECT 94.255 192.210 94.545 192.255 ;
        RECT 88.275 192.070 94.545 192.210 ;
        RECT 88.275 192.025 88.565 192.070 ;
        RECT 89.195 192.025 89.485 192.070 ;
        RECT 92.400 192.010 92.720 192.070 ;
        RECT 94.255 192.025 94.545 192.070 ;
        RECT 89.655 191.870 89.945 191.915 ;
        RECT 93.795 191.870 94.085 191.915 ;
        RECT 89.655 191.730 94.085 191.870 ;
        RECT 95.250 191.870 95.390 192.410 ;
        RECT 97.000 192.410 100.910 192.550 ;
        RECT 97.000 192.350 97.320 192.410 ;
        RECT 102.535 192.365 102.825 192.595 ;
        RECT 102.995 192.365 103.285 192.595 ;
        RECT 104.835 192.365 105.125 192.595 ;
        RECT 109.420 192.550 109.740 192.610 ;
        RECT 105.370 192.410 109.740 192.550 ;
        RECT 97.935 192.210 98.225 192.255 ;
        RECT 99.760 192.210 100.080 192.270 ;
        RECT 97.935 192.070 100.080 192.210 ;
        RECT 97.935 192.025 98.225 192.070 ;
        RECT 99.760 192.010 100.080 192.070 ;
        RECT 102.060 192.210 102.380 192.270 ;
        RECT 103.070 192.210 103.210 192.365 ;
        RECT 102.060 192.070 103.210 192.210 ;
        RECT 102.060 192.010 102.380 192.070 ;
        RECT 100.695 191.870 100.985 191.915 ;
        RECT 105.370 191.870 105.510 192.410 ;
        RECT 109.420 192.350 109.740 192.410 ;
        RECT 109.880 192.550 110.200 192.610 ;
        RECT 110.815 192.550 111.105 192.595 ;
        RECT 109.880 192.410 111.105 192.550 ;
        RECT 109.880 192.350 110.200 192.410 ;
        RECT 110.815 192.365 111.105 192.410 ;
        RECT 112.775 192.550 113.065 192.595 ;
        RECT 113.560 192.550 113.880 192.610 ;
        RECT 112.775 192.410 113.880 192.550 ;
        RECT 112.775 192.365 113.065 192.410 ;
        RECT 113.560 192.350 113.880 192.410 ;
        RECT 111.260 192.265 111.580 192.270 ;
        RECT 112.210 192.265 112.470 192.300 ;
        RECT 111.260 192.255 112.470 192.265 ;
        RECT 106.215 192.210 106.505 192.255 ;
        RECT 107.135 192.210 107.425 192.255 ;
        RECT 111.260 192.210 112.485 192.255 ;
        RECT 106.215 192.070 112.485 192.210 ;
        RECT 106.215 192.025 106.505 192.070 ;
        RECT 107.135 192.025 107.425 192.070 ;
        RECT 111.260 192.010 111.580 192.070 ;
        RECT 112.195 192.025 112.485 192.070 ;
        RECT 112.210 191.980 112.470 192.025 ;
        RECT 95.250 191.730 105.510 191.870 ;
        RECT 107.595 191.870 107.885 191.915 ;
        RECT 111.735 191.870 112.025 191.915 ;
        RECT 107.595 191.730 112.025 191.870 ;
        RECT 114.110 191.870 114.250 192.750 ;
        RECT 119.630 192.750 122.990 192.890 ;
        RECT 115.400 192.350 115.720 192.610 ;
        RECT 117.700 192.550 118.020 192.610 ;
        RECT 119.630 192.595 119.770 192.750 ;
        RECT 119.555 192.550 119.845 192.595 ;
        RECT 117.700 192.410 119.845 192.550 ;
        RECT 117.700 192.350 118.020 192.410 ;
        RECT 119.555 192.365 119.845 192.410 ;
        RECT 120.920 192.350 121.240 192.610 ;
        RECT 122.850 192.595 122.990 192.750 ;
        RECT 127.360 192.690 127.680 192.950 ;
        RECT 138.490 192.890 138.630 193.090 ;
        RECT 140.560 192.890 140.850 192.935 ;
        RECT 138.490 192.750 140.850 192.890 ;
        RECT 140.560 192.705 140.850 192.750 ;
        RECT 122.775 192.550 123.065 192.595 ;
        RECT 124.600 192.550 124.920 192.610 ;
        RECT 122.775 192.410 124.920 192.550 ;
        RECT 127.450 192.545 127.590 192.690 ;
        RECT 128.295 192.550 128.585 192.595 ;
        RECT 129.660 192.550 129.980 192.610 ;
        RECT 122.775 192.365 123.065 192.410 ;
        RECT 124.600 192.350 124.920 192.410 ;
        RECT 127.375 192.315 127.665 192.545 ;
        RECT 128.295 192.410 129.980 192.550 ;
        RECT 128.295 192.365 128.585 192.410 ;
        RECT 129.660 192.350 129.980 192.410 ;
        RECT 131.975 192.365 132.265 192.595 ;
        RECT 136.575 192.550 136.865 192.595 ;
        RECT 137.020 192.550 137.340 192.610 ;
        RECT 136.575 192.410 137.340 192.550 ;
        RECT 136.575 192.365 136.865 192.410 ;
        RECT 120.475 192.210 120.765 192.255 ;
        RECT 122.300 192.210 122.620 192.270 ;
        RECT 125.980 192.210 126.300 192.270 ;
        RECT 130.580 192.210 130.900 192.270 ;
        RECT 132.050 192.210 132.190 192.365 ;
        RECT 137.020 192.350 137.340 192.410 ;
        RECT 137.480 192.350 137.800 192.610 ;
        RECT 137.940 192.350 138.260 192.610 ;
        RECT 139.335 192.550 139.625 192.595 ;
        RECT 139.780 192.550 140.100 192.610 ;
        RECT 147.600 192.550 147.920 192.610 ;
        RECT 139.335 192.410 140.100 192.550 ;
        RECT 139.335 192.365 139.625 192.410 ;
        RECT 120.475 192.070 122.620 192.210 ;
        RECT 120.475 192.025 120.765 192.070 ;
        RECT 122.300 192.010 122.620 192.070 ;
        RECT 122.850 192.070 126.300 192.210 ;
        RECT 116.335 191.870 116.625 191.915 ;
        RECT 116.780 191.870 117.100 191.930 ;
        RECT 114.110 191.730 117.100 191.870 ;
        RECT 89.655 191.685 89.945 191.730 ;
        RECT 93.795 191.685 94.085 191.730 ;
        RECT 100.695 191.685 100.985 191.730 ;
        RECT 107.595 191.685 107.885 191.730 ;
        RECT 111.735 191.685 112.025 191.730 ;
        RECT 116.335 191.685 116.625 191.730 ;
        RECT 116.780 191.670 117.100 191.730 ;
        RECT 117.240 191.870 117.560 191.930 ;
        RECT 118.635 191.870 118.925 191.915 ;
        RECT 122.850 191.870 122.990 192.070 ;
        RECT 125.980 192.010 126.300 192.070 ;
        RECT 128.370 192.070 130.350 192.210 ;
        RECT 128.370 191.870 128.510 192.070 ;
        RECT 117.240 191.730 118.925 191.870 ;
        RECT 117.240 191.670 117.560 191.730 ;
        RECT 118.635 191.685 118.925 191.730 ;
        RECT 120.550 191.730 122.990 191.870 ;
        RECT 123.310 191.730 128.510 191.870 ;
        RECT 75.395 191.530 75.685 191.575 ;
        RECT 77.220 191.530 77.540 191.590 ;
        RECT 75.395 191.390 77.540 191.530 ;
        RECT 75.395 191.345 75.685 191.390 ;
        RECT 77.220 191.330 77.540 191.390 ;
        RECT 82.740 191.330 83.060 191.590 ;
        RECT 90.115 191.530 90.405 191.575 ;
        RECT 91.495 191.530 91.785 191.575 ;
        RECT 90.115 191.390 91.785 191.530 ;
        RECT 90.115 191.345 90.405 191.390 ;
        RECT 91.495 191.345 91.785 191.390 ;
        RECT 92.415 191.530 92.705 191.575 ;
        RECT 94.715 191.530 95.005 191.575 ;
        RECT 92.415 191.390 95.005 191.530 ;
        RECT 92.415 191.345 92.705 191.390 ;
        RECT 94.715 191.345 95.005 191.390 ;
        RECT 95.620 191.330 95.940 191.590 ;
        RECT 97.000 191.330 97.320 191.590 ;
        RECT 104.835 191.530 105.125 191.575 ;
        RECT 107.120 191.530 107.440 191.590 ;
        RECT 104.835 191.390 107.440 191.530 ;
        RECT 104.835 191.345 105.125 191.390 ;
        RECT 107.120 191.330 107.440 191.390 ;
        RECT 108.055 191.530 108.345 191.575 ;
        RECT 109.435 191.530 109.725 191.575 ;
        RECT 108.055 191.390 109.725 191.530 ;
        RECT 108.055 191.345 108.345 191.390 ;
        RECT 109.435 191.345 109.725 191.390 ;
        RECT 110.355 191.530 110.645 191.575 ;
        RECT 112.655 191.530 112.945 191.575 ;
        RECT 110.355 191.390 112.945 191.530 ;
        RECT 116.870 191.530 117.010 191.670 ;
        RECT 120.550 191.530 120.690 191.730 ;
        RECT 123.310 191.590 123.450 191.730 ;
        RECT 128.755 191.685 129.045 191.915 ;
        RECT 130.210 191.870 130.350 192.070 ;
        RECT 130.580 192.070 132.190 192.210 ;
        RECT 132.420 192.210 132.740 192.270 ;
        RECT 139.410 192.210 139.550 192.365 ;
        RECT 139.780 192.350 140.100 192.410 ;
        RECT 146.310 192.410 147.920 192.550 ;
        RECT 132.420 192.070 139.550 192.210 ;
        RECT 140.215 192.210 140.505 192.255 ;
        RECT 141.405 192.210 141.695 192.255 ;
        RECT 143.925 192.210 144.215 192.255 ;
        RECT 140.215 192.070 144.215 192.210 ;
        RECT 130.580 192.010 130.900 192.070 ;
        RECT 132.420 192.010 132.740 192.070 ;
        RECT 140.215 192.025 140.505 192.070 ;
        RECT 141.405 192.025 141.695 192.070 ;
        RECT 143.925 192.025 144.215 192.070 ;
        RECT 132.895 191.870 133.185 191.915 ;
        RECT 137.940 191.870 138.260 191.930 ;
        RECT 146.310 191.915 146.450 192.410 ;
        RECT 147.600 192.350 147.920 192.410 ;
        RECT 130.210 191.730 138.260 191.870 ;
        RECT 132.895 191.685 133.185 191.730 ;
        RECT 116.870 191.390 120.690 191.530 ;
        RECT 110.355 191.345 110.645 191.390 ;
        RECT 112.655 191.345 112.945 191.390 ;
        RECT 120.920 191.330 121.240 191.590 ;
        RECT 123.220 191.330 123.540 191.590 ;
        RECT 123.680 191.530 124.000 191.590 ;
        RECT 125.520 191.530 125.840 191.590 ;
        RECT 123.680 191.390 125.840 191.530 ;
        RECT 123.680 191.330 124.000 191.390 ;
        RECT 125.520 191.330 125.840 191.390 ;
        RECT 126.440 191.330 126.760 191.590 ;
        RECT 126.900 191.530 127.220 191.590 ;
        RECT 128.830 191.530 128.970 191.685 ;
        RECT 137.940 191.670 138.260 191.730 ;
        RECT 139.820 191.870 140.110 191.915 ;
        RECT 141.920 191.870 142.210 191.915 ;
        RECT 143.490 191.870 143.780 191.915 ;
        RECT 139.820 191.730 143.780 191.870 ;
        RECT 139.820 191.685 140.110 191.730 ;
        RECT 141.920 191.685 142.210 191.730 ;
        RECT 143.490 191.685 143.780 191.730 ;
        RECT 146.235 191.685 146.525 191.915 ;
        RECT 146.680 191.870 147.000 191.930 ;
        RECT 148.060 191.870 148.380 191.930 ;
        RECT 146.680 191.730 148.380 191.870 ;
        RECT 146.680 191.670 147.000 191.730 ;
        RECT 148.060 191.670 148.380 191.730 ;
        RECT 126.900 191.390 128.970 191.530 ;
        RECT 130.120 191.530 130.440 191.590 ;
        RECT 130.595 191.530 130.885 191.575 ;
        RECT 130.120 191.390 130.885 191.530 ;
        RECT 126.900 191.330 127.220 191.390 ;
        RECT 130.120 191.330 130.440 191.390 ;
        RECT 130.595 191.345 130.885 191.390 ;
        RECT 131.500 191.330 131.820 191.590 ;
        RECT 70.710 190.710 156.270 191.190 ;
        RECT 85.040 190.510 85.360 190.570 ;
        RECT 86.895 190.510 87.185 190.555 ;
        RECT 85.040 190.370 87.185 190.510 ;
        RECT 85.040 190.310 85.360 190.370 ;
        RECT 86.895 190.325 87.185 190.370 ;
        RECT 91.955 190.510 92.245 190.555 ;
        RECT 92.860 190.510 93.180 190.570 ;
        RECT 91.955 190.370 93.180 190.510 ;
        RECT 91.955 190.325 92.245 190.370 ;
        RECT 92.860 190.310 93.180 190.370 ;
        RECT 94.700 190.310 95.020 190.570 ;
        RECT 97.000 190.510 97.320 190.570 ;
        RECT 95.710 190.370 97.320 190.510 ;
        RECT 77.220 190.170 77.540 190.230 ;
        RECT 80.915 190.170 81.205 190.215 ;
        RECT 77.220 190.030 81.205 190.170 ;
        RECT 77.220 189.970 77.540 190.030 ;
        RECT 80.915 189.985 81.205 190.030 ;
        RECT 86.050 190.030 91.250 190.170 ;
        RECT 86.050 189.890 86.190 190.030 ;
        RECT 80.440 189.830 80.760 189.890 ;
        RECT 82.755 189.830 83.045 189.875 ;
        RECT 80.440 189.690 83.045 189.830 ;
        RECT 80.440 189.630 80.760 189.690 ;
        RECT 82.755 189.645 83.045 189.690 ;
        RECT 85.960 189.630 86.280 189.890 ;
        RECT 88.735 189.830 89.025 189.875 ;
        RECT 89.640 189.830 89.960 189.890 ;
        RECT 88.735 189.690 89.960 189.830 ;
        RECT 88.735 189.645 89.025 189.690 ;
        RECT 89.640 189.630 89.960 189.690 ;
        RECT 80.900 189.490 81.220 189.550 ;
        RECT 81.835 189.490 82.125 189.535 ;
        RECT 80.900 189.350 82.125 189.490 ;
        RECT 80.900 189.290 81.220 189.350 ;
        RECT 81.835 189.305 82.125 189.350 ;
        RECT 84.135 189.490 84.425 189.535 ;
        RECT 85.515 189.490 85.805 189.535 ;
        RECT 86.050 189.490 86.190 189.630 ;
        RECT 84.135 189.350 86.190 189.490 ;
        RECT 84.135 189.305 84.425 189.350 ;
        RECT 85.515 189.305 85.805 189.350 ;
        RECT 86.420 189.290 86.740 189.550 ;
        RECT 87.340 189.490 87.660 189.550 ;
        RECT 86.970 189.350 87.660 189.490 ;
        RECT 85.975 189.150 86.265 189.195 ;
        RECT 86.970 189.150 87.110 189.350 ;
        RECT 87.340 189.290 87.660 189.350 ;
        RECT 87.800 189.290 88.120 189.550 ;
        RECT 88.260 189.290 88.580 189.550 ;
        RECT 89.180 189.490 89.500 189.550 ;
        RECT 89.180 189.350 89.695 189.490 ;
        RECT 89.180 189.290 89.500 189.350 ;
        RECT 90.115 189.305 90.405 189.535 ;
        RECT 85.975 189.010 87.110 189.150 ;
        RECT 85.975 188.965 86.265 189.010 ;
        RECT 85.055 188.810 85.345 188.855 ;
        RECT 88.350 188.810 88.490 189.290 ;
        RECT 90.190 189.150 90.330 189.305 ;
        RECT 89.270 189.010 90.330 189.150 ;
        RECT 91.110 189.150 91.250 190.030 ;
        RECT 94.790 189.830 94.930 190.310 ;
        RECT 92.950 189.690 94.930 189.830 ;
        RECT 91.495 189.490 91.785 189.535 ;
        RECT 91.940 189.490 92.260 189.550 ;
        RECT 92.950 189.535 93.090 189.690 ;
        RECT 91.495 189.350 92.260 189.490 ;
        RECT 91.495 189.305 91.785 189.350 ;
        RECT 91.940 189.290 92.260 189.350 ;
        RECT 92.875 189.305 93.165 189.535 ;
        RECT 94.240 189.290 94.560 189.550 ;
        RECT 95.710 189.535 95.850 190.370 ;
        RECT 97.000 190.310 97.320 190.370 ;
        RECT 101.140 190.310 101.460 190.570 ;
        RECT 102.060 190.310 102.380 190.570 ;
        RECT 103.900 190.310 104.220 190.570 ;
        RECT 104.835 190.325 105.125 190.555 ;
        RECT 108.040 190.510 108.360 190.570 ;
        RECT 114.020 190.510 114.340 190.570 ;
        RECT 108.040 190.370 114.340 190.510 ;
        RECT 100.220 190.170 100.540 190.230 ;
        RECT 97.550 190.030 100.540 190.170 ;
        RECT 102.150 190.170 102.290 190.310 ;
        RECT 104.910 190.170 105.050 190.325 ;
        RECT 108.040 190.310 108.360 190.370 ;
        RECT 109.895 190.170 110.185 190.215 ;
        RECT 102.150 190.030 105.050 190.170 ;
        RECT 109.050 190.030 110.185 190.170 ;
        RECT 97.550 189.830 97.690 190.030 ;
        RECT 100.220 189.970 100.540 190.030 ;
        RECT 109.050 189.890 109.190 190.030 ;
        RECT 109.895 189.985 110.185 190.030 ;
        RECT 96.630 189.690 97.690 189.830 ;
        RECT 98.380 189.830 98.700 189.890 ;
        RECT 98.855 189.830 99.145 189.875 ;
        RECT 98.380 189.690 99.145 189.830 ;
        RECT 95.635 189.305 95.925 189.535 ;
        RECT 96.095 189.490 96.385 189.535 ;
        RECT 96.630 189.490 96.770 189.690 ;
        RECT 98.380 189.630 98.700 189.690 ;
        RECT 98.855 189.645 99.145 189.690 ;
        RECT 99.390 189.690 102.750 189.830 ;
        RECT 99.390 189.550 99.530 189.690 ;
        RECT 99.300 189.490 99.620 189.550 ;
        RECT 102.610 189.535 102.750 189.690 ;
        RECT 104.360 189.630 104.680 189.890 ;
        RECT 108.960 189.830 109.280 189.890 ;
        RECT 104.910 189.690 109.280 189.830 ;
        RECT 96.095 189.350 96.770 189.490 ;
        RECT 99.105 189.350 99.620 189.490 ;
        RECT 96.095 189.305 96.385 189.350 ;
        RECT 99.300 189.290 99.620 189.350 ;
        RECT 101.155 189.305 101.445 189.535 ;
        RECT 102.535 189.305 102.825 189.535 ;
        RECT 104.450 189.490 104.590 189.630 ;
        RECT 104.910 189.550 105.050 189.690 ;
        RECT 108.960 189.630 109.280 189.690 ;
        RECT 109.420 189.830 109.740 189.890 ;
        RECT 111.720 189.830 112.040 189.890 ;
        RECT 109.420 189.690 112.040 189.830 ;
        RECT 109.420 189.630 109.740 189.690 ;
        RECT 111.720 189.630 112.040 189.690 ;
        RECT 103.070 189.350 104.590 189.490 ;
        RECT 99.760 189.150 100.080 189.210 ;
        RECT 101.230 189.150 101.370 189.305 ;
        RECT 91.110 189.010 98.610 189.150 ;
        RECT 89.270 188.870 89.410 189.010 ;
        RECT 85.055 188.670 88.490 188.810 ;
        RECT 85.055 188.625 85.345 188.670 ;
        RECT 89.180 188.610 89.500 188.870 ;
        RECT 91.035 188.810 91.325 188.855 ;
        RECT 97.920 188.810 98.240 188.870 ;
        RECT 91.035 188.670 98.240 188.810 ;
        RECT 98.470 188.810 98.610 189.010 ;
        RECT 99.760 189.010 101.370 189.150 ;
        RECT 99.760 188.950 100.080 189.010 ;
        RECT 99.850 188.810 99.990 188.950 ;
        RECT 98.470 188.670 99.990 188.810 ;
        RECT 102.075 188.810 102.365 188.855 ;
        RECT 103.070 188.810 103.210 189.350 ;
        RECT 104.820 189.290 105.140 189.550 ;
        RECT 106.660 189.290 106.980 189.550 ;
        RECT 107.135 189.490 107.425 189.535 ;
        RECT 107.580 189.490 107.900 189.550 ;
        RECT 112.270 189.535 112.410 190.370 ;
        RECT 114.020 190.310 114.340 190.370 ;
        RECT 115.875 190.510 116.165 190.555 ;
        RECT 117.255 190.510 117.545 190.555 ;
        RECT 115.875 190.370 117.545 190.510 ;
        RECT 115.875 190.325 116.165 190.370 ;
        RECT 117.255 190.325 117.545 190.370 ;
        RECT 118.175 190.510 118.465 190.555 ;
        RECT 120.475 190.510 120.765 190.555 ;
        RECT 118.175 190.370 120.765 190.510 ;
        RECT 118.175 190.325 118.465 190.370 ;
        RECT 120.475 190.325 120.765 190.370 ;
        RECT 120.920 190.510 121.240 190.570 ;
        RECT 123.235 190.510 123.525 190.555 ;
        RECT 126.900 190.510 127.220 190.570 ;
        RECT 127.835 190.510 128.125 190.555 ;
        RECT 136.115 190.510 136.405 190.555 ;
        RECT 136.560 190.510 136.880 190.570 ;
        RECT 120.920 190.370 128.125 190.510 ;
        RECT 120.920 190.310 121.240 190.370 ;
        RECT 123.235 190.325 123.525 190.370 ;
        RECT 126.900 190.310 127.220 190.370 ;
        RECT 127.835 190.325 128.125 190.370 ;
        RECT 128.370 190.370 135.870 190.510 ;
        RECT 115.415 190.170 115.705 190.215 ;
        RECT 119.555 190.170 119.845 190.215 ;
        RECT 115.415 190.030 119.845 190.170 ;
        RECT 115.415 189.985 115.705 190.030 ;
        RECT 119.555 189.985 119.845 190.030 ;
        RECT 121.395 190.170 121.685 190.215 ;
        RECT 122.760 190.170 123.080 190.230 ;
        RECT 121.395 190.030 123.080 190.170 ;
        RECT 121.395 189.985 121.685 190.030 ;
        RECT 122.760 189.970 123.080 190.030 ;
        RECT 124.140 190.170 124.460 190.230 ;
        RECT 128.370 190.170 128.510 190.370 ;
        RECT 124.140 190.030 128.510 190.170 ;
        RECT 124.140 189.970 124.460 190.030 ;
        RECT 128.740 189.970 129.060 190.230 ;
        RECT 129.200 189.970 129.520 190.230 ;
        RECT 114.035 189.830 114.325 189.875 ;
        RECT 114.955 189.830 115.245 189.875 ;
        RECT 120.015 189.830 120.305 189.875 ;
        RECT 125.995 189.830 126.285 189.875 ;
        RECT 128.280 189.830 128.600 189.890 ;
        RECT 114.035 189.690 120.305 189.830 ;
        RECT 114.035 189.645 114.325 189.690 ;
        RECT 114.955 189.645 115.245 189.690 ;
        RECT 115.490 189.550 115.630 189.690 ;
        RECT 120.015 189.645 120.305 189.690 ;
        RECT 121.470 189.690 122.530 189.830 ;
        RECT 110.815 189.490 111.105 189.535 ;
        RECT 107.135 189.350 107.900 189.490 ;
        RECT 107.135 189.305 107.425 189.350 ;
        RECT 102.075 188.670 103.210 188.810 ;
        RECT 103.455 188.810 103.745 188.855 ;
        RECT 107.210 188.810 107.350 189.305 ;
        RECT 107.580 189.290 107.900 189.350 ;
        RECT 109.970 189.350 111.105 189.490 ;
        RECT 109.970 189.150 110.110 189.350 ;
        RECT 110.815 189.305 111.105 189.350 ;
        RECT 112.195 189.305 112.485 189.535 ;
        RECT 115.400 189.290 115.720 189.550 ;
        RECT 115.860 189.490 116.180 189.550 ;
        RECT 116.795 189.490 117.085 189.535 ;
        RECT 115.860 189.350 117.085 189.490 ;
        RECT 115.860 189.290 116.180 189.350 ;
        RECT 116.795 189.305 117.085 189.350 ;
        RECT 113.560 189.150 113.880 189.210 ;
        RECT 109.970 189.010 113.880 189.150 ;
        RECT 109.970 188.870 110.110 189.010 ;
        RECT 113.560 188.950 113.880 189.010 ;
        RECT 116.320 188.950 116.640 189.210 ;
        RECT 118.160 189.150 118.480 189.210 ;
        RECT 118.635 189.150 118.925 189.195 ;
        RECT 121.470 189.150 121.610 189.690 ;
        RECT 122.390 189.490 122.530 189.690 ;
        RECT 125.995 189.690 128.600 189.830 ;
        RECT 125.995 189.645 126.285 189.690 ;
        RECT 128.280 189.630 128.600 189.690 ;
        RECT 122.390 189.350 127.130 189.490 ;
        RECT 123.220 189.195 123.540 189.210 ;
        RECT 118.160 189.010 118.925 189.150 ;
        RECT 118.160 188.950 118.480 189.010 ;
        RECT 118.635 188.965 118.925 189.010 ;
        RECT 120.550 189.010 121.610 189.150 ;
        RECT 103.455 188.670 107.350 188.810 ;
        RECT 91.035 188.625 91.325 188.670 ;
        RECT 97.920 188.610 98.240 188.670 ;
        RECT 102.075 188.625 102.365 188.670 ;
        RECT 103.455 188.625 103.745 188.670 ;
        RECT 109.880 188.610 110.200 188.870 ;
        RECT 111.720 188.810 112.040 188.870 ;
        RECT 113.115 188.810 113.405 188.855 ;
        RECT 114.955 188.810 115.245 188.855 ;
        RECT 111.720 188.670 115.245 188.810 ;
        RECT 116.410 188.810 116.550 188.950 ;
        RECT 117.240 188.810 117.560 188.870 ;
        RECT 116.410 188.670 117.560 188.810 ;
        RECT 111.720 188.610 112.040 188.670 ;
        RECT 113.115 188.625 113.405 188.670 ;
        RECT 114.955 188.625 115.245 188.670 ;
        RECT 117.240 188.610 117.560 188.670 ;
        RECT 119.080 188.810 119.400 188.870 ;
        RECT 120.550 188.855 120.690 189.010 ;
        RECT 123.155 188.965 123.540 189.195 ;
        RECT 124.155 189.150 124.445 189.195 ;
        RECT 124.600 189.150 124.920 189.210 ;
        RECT 124.155 189.010 124.920 189.150 ;
        RECT 124.155 188.965 124.445 189.010 ;
        RECT 123.220 188.950 123.540 188.965 ;
        RECT 124.600 188.950 124.920 189.010 ;
        RECT 125.075 189.150 125.365 189.195 ;
        RECT 125.980 189.150 126.300 189.210 ;
        RECT 125.075 189.010 126.300 189.150 ;
        RECT 126.990 189.150 127.130 189.350 ;
        RECT 127.360 189.290 127.680 189.550 ;
        RECT 128.830 189.535 128.970 189.970 ;
        RECT 129.290 189.535 129.430 189.970 ;
        RECT 135.730 189.875 135.870 190.370 ;
        RECT 136.115 190.370 136.880 190.510 ;
        RECT 136.115 190.325 136.405 190.370 ;
        RECT 136.560 190.310 136.880 190.370 ;
        RECT 137.495 190.510 137.785 190.555 ;
        RECT 138.400 190.510 138.720 190.570 ;
        RECT 137.495 190.370 138.720 190.510 ;
        RECT 137.495 190.325 137.785 190.370 ;
        RECT 138.400 190.310 138.720 190.370 ;
        RECT 137.940 190.170 138.260 190.230 ;
        RECT 136.650 190.030 138.260 190.170 ;
        RECT 136.650 189.875 136.790 190.030 ;
        RECT 137.940 189.970 138.260 190.030 ;
        RECT 140.280 190.170 140.570 190.215 ;
        RECT 142.380 190.170 142.670 190.215 ;
        RECT 143.950 190.170 144.240 190.215 ;
        RECT 140.280 190.030 144.240 190.170 ;
        RECT 140.280 189.985 140.570 190.030 ;
        RECT 142.380 189.985 142.670 190.030 ;
        RECT 143.950 189.985 144.240 190.030 ;
        RECT 146.695 190.170 146.985 190.215 ;
        RECT 146.695 190.030 147.370 190.170 ;
        RECT 146.695 189.985 146.985 190.030 ;
        RECT 132.435 189.830 132.725 189.875 ;
        RECT 131.130 189.690 132.725 189.830 ;
        RECT 131.130 189.550 131.270 189.690 ;
        RECT 132.435 189.645 132.725 189.690 ;
        RECT 135.655 189.645 135.945 189.875 ;
        RECT 136.575 189.645 136.865 189.875 ;
        RECT 137.480 189.830 137.800 189.890 ;
        RECT 140.675 189.830 140.965 189.875 ;
        RECT 141.865 189.830 142.155 189.875 ;
        RECT 144.385 189.830 144.675 189.875 ;
        RECT 137.480 189.690 140.470 189.830 ;
        RECT 137.480 189.630 137.800 189.690 ;
        RECT 128.755 189.305 129.045 189.535 ;
        RECT 129.215 189.305 129.505 189.535 ;
        RECT 130.580 189.290 130.900 189.550 ;
        RECT 131.040 189.290 131.360 189.550 ;
        RECT 131.515 189.490 131.805 189.535 ;
        RECT 133.815 189.490 134.105 189.535 ;
        RECT 137.035 189.490 137.325 189.535 ;
        RECT 137.570 189.490 137.710 189.630 ;
        RECT 131.515 189.350 136.790 189.490 ;
        RECT 131.515 189.305 131.805 189.350 ;
        RECT 133.815 189.305 134.105 189.350 ;
        RECT 136.650 189.150 136.790 189.350 ;
        RECT 137.035 189.350 137.710 189.490 ;
        RECT 137.035 189.305 137.325 189.350 ;
        RECT 139.780 189.290 140.100 189.550 ;
        RECT 126.990 189.010 133.110 189.150 ;
        RECT 136.650 189.010 137.710 189.150 ;
        RECT 125.075 188.965 125.365 189.010 ;
        RECT 125.980 188.950 126.300 189.010 ;
        RECT 120.475 188.810 120.765 188.855 ;
        RECT 119.080 188.670 120.765 188.810 ;
        RECT 119.080 188.610 119.400 188.670 ;
        RECT 120.475 188.625 120.765 188.670 ;
        RECT 120.920 188.810 121.240 188.870 ;
        RECT 122.315 188.810 122.605 188.855 ;
        RECT 120.920 188.670 122.605 188.810 ;
        RECT 124.690 188.810 124.830 188.950 ;
        RECT 126.455 188.810 126.745 188.855 ;
        RECT 124.690 188.670 126.745 188.810 ;
        RECT 120.920 188.610 121.240 188.670 ;
        RECT 122.315 188.625 122.605 188.670 ;
        RECT 126.455 188.625 126.745 188.670 ;
        RECT 130.120 188.610 130.440 188.870 ;
        RECT 132.970 188.855 133.110 189.010 ;
        RECT 132.895 188.810 133.185 188.855 ;
        RECT 137.020 188.810 137.340 188.870 ;
        RECT 132.895 188.670 137.340 188.810 ;
        RECT 137.570 188.810 137.710 189.010 ;
        RECT 138.400 188.950 138.720 189.210 ;
        RECT 139.335 188.965 139.625 189.195 ;
        RECT 140.330 189.150 140.470 189.690 ;
        RECT 140.675 189.690 144.675 189.830 ;
        RECT 140.675 189.645 140.965 189.690 ;
        RECT 141.865 189.645 142.155 189.690 ;
        RECT 144.385 189.645 144.675 189.690 ;
        RECT 141.130 189.490 141.420 189.535 ;
        RECT 146.680 189.490 147.000 189.550 ;
        RECT 141.130 189.350 147.000 189.490 ;
        RECT 147.230 189.490 147.370 190.030 ;
        RECT 147.600 189.970 147.920 190.230 ;
        RECT 151.295 190.170 151.585 190.215 ;
        RECT 153.580 190.170 153.900 190.230 ;
        RECT 149.070 190.030 153.900 190.170 ;
        RECT 147.690 189.830 147.830 189.970 ;
        RECT 149.070 189.890 149.210 190.030 ;
        RECT 151.295 189.985 151.585 190.030 ;
        RECT 153.580 189.970 153.900 190.030 ;
        RECT 148.535 189.830 148.825 189.875 ;
        RECT 147.690 189.690 148.825 189.830 ;
        RECT 148.535 189.645 148.825 189.690 ;
        RECT 148.980 189.630 149.300 189.890 ;
        RECT 149.900 189.630 150.220 189.890 ;
        RECT 148.075 189.490 148.365 189.535 ;
        RECT 151.740 189.490 152.060 189.550 ;
        RECT 147.230 189.350 152.060 189.490 ;
        RECT 141.130 189.305 141.420 189.350 ;
        RECT 146.680 189.290 147.000 189.350 ;
        RECT 148.075 189.305 148.365 189.350 ;
        RECT 151.740 189.290 152.060 189.350 ;
        RECT 152.200 189.290 152.520 189.550 ;
        RECT 153.595 189.490 153.885 189.535 ;
        RECT 153.210 189.350 153.885 189.490 ;
        RECT 153.210 189.210 153.350 189.350 ;
        RECT 153.595 189.305 153.885 189.350 ;
        RECT 141.620 189.150 141.940 189.210 ;
        RECT 140.330 189.010 141.940 189.150 ;
        RECT 139.410 188.810 139.550 188.965 ;
        RECT 141.620 188.950 141.940 189.010 ;
        RECT 153.120 188.950 153.440 189.210 ;
        RECT 152.675 188.810 152.965 188.855 ;
        RECT 154.960 188.810 155.280 188.870 ;
        RECT 137.570 188.670 155.280 188.810 ;
        RECT 132.895 188.625 133.185 188.670 ;
        RECT 137.020 188.610 137.340 188.670 ;
        RECT 152.675 188.625 152.965 188.670 ;
        RECT 154.960 188.610 155.280 188.670 ;
        RECT 70.710 187.990 156.270 188.470 ;
        RECT 78.600 187.790 78.920 187.850 ;
        RECT 84.595 187.790 84.885 187.835 ;
        RECT 85.500 187.790 85.820 187.850 ;
        RECT 78.600 187.650 83.430 187.790 ;
        RECT 78.600 187.590 78.920 187.650 ;
        RECT 80.900 187.250 81.220 187.510 ;
        RECT 83.290 187.495 83.430 187.650 ;
        RECT 84.595 187.650 85.820 187.790 ;
        RECT 84.595 187.605 84.885 187.650 ;
        RECT 85.500 187.590 85.820 187.650 ;
        RECT 85.960 187.590 86.280 187.850 ;
        RECT 87.355 187.790 87.645 187.835 ;
        RECT 87.800 187.790 88.120 187.850 ;
        RECT 87.355 187.650 88.120 187.790 ;
        RECT 87.355 187.605 87.645 187.650 ;
        RECT 87.800 187.590 88.120 187.650 ;
        RECT 89.640 187.590 89.960 187.850 ;
        RECT 97.015 187.790 97.305 187.835 ;
        RECT 102.520 187.790 102.840 187.850 ;
        RECT 106.200 187.790 106.520 187.850 ;
        RECT 96.170 187.650 101.370 187.790 ;
        RECT 82.215 187.450 82.505 187.495 ;
        RECT 82.215 187.265 82.510 187.450 ;
        RECT 83.215 187.265 83.505 187.495 ;
        RECT 89.195 187.450 89.485 187.495 ;
        RECT 89.730 187.450 89.870 187.590 ;
        RECT 86.510 187.310 89.870 187.450 ;
        RECT 74.000 187.155 74.320 187.170 ;
        RECT 73.970 186.925 74.320 187.155 ;
        RECT 80.990 187.075 81.130 187.250 ;
        RECT 74.000 186.910 74.320 186.925 ;
        RECT 80.915 186.845 81.205 187.075 ;
        RECT 72.160 186.770 72.480 186.830 ;
        RECT 72.635 186.770 72.925 186.815 ;
        RECT 72.160 186.630 72.925 186.770 ;
        RECT 72.160 186.570 72.480 186.630 ;
        RECT 72.635 186.585 72.925 186.630 ;
        RECT 73.515 186.770 73.805 186.815 ;
        RECT 74.705 186.770 74.995 186.815 ;
        RECT 77.225 186.770 77.515 186.815 ;
        RECT 73.515 186.630 77.515 186.770 ;
        RECT 73.515 186.585 73.805 186.630 ;
        RECT 74.705 186.585 74.995 186.630 ;
        RECT 77.225 186.585 77.515 186.630 ;
        RECT 73.120 186.430 73.410 186.475 ;
        RECT 75.220 186.430 75.510 186.475 ;
        RECT 76.790 186.430 77.080 186.475 ;
        RECT 82.370 186.430 82.510 187.265 ;
        RECT 83.290 187.110 83.430 187.265 ;
        RECT 83.675 187.110 83.965 187.155 ;
        RECT 83.290 186.970 83.965 187.110 ;
        RECT 83.675 186.925 83.965 186.970 ;
        RECT 85.055 186.925 85.345 187.155 ;
        RECT 85.130 186.430 85.270 186.925 ;
        RECT 73.120 186.290 77.080 186.430 ;
        RECT 73.120 186.245 73.410 186.290 ;
        RECT 75.220 186.245 75.510 186.290 ;
        RECT 76.790 186.245 77.080 186.290 ;
        RECT 79.610 186.290 85.270 186.430 ;
        RECT 79.610 186.150 79.750 186.290 ;
        RECT 79.520 185.890 79.840 186.150 ;
        RECT 79.980 185.890 80.300 186.150 ;
        RECT 80.440 186.090 80.760 186.150 ;
        RECT 81.375 186.090 81.665 186.135 ;
        RECT 80.440 185.950 81.665 186.090 ;
        RECT 80.440 185.890 80.760 185.950 ;
        RECT 81.375 185.905 81.665 185.950 ;
        RECT 82.295 186.090 82.585 186.135 ;
        RECT 84.120 186.090 84.440 186.150 ;
        RECT 86.510 186.090 86.650 187.310 ;
        RECT 89.195 187.265 89.485 187.310 ;
        RECT 96.170 187.170 96.310 187.650 ;
        RECT 97.015 187.605 97.305 187.650 ;
        RECT 99.760 187.450 100.080 187.510 ;
        RECT 100.695 187.450 100.985 187.495 ;
        RECT 99.760 187.310 100.985 187.450 ;
        RECT 101.230 187.450 101.370 187.650 ;
        RECT 102.520 187.650 106.520 187.790 ;
        RECT 102.520 187.590 102.840 187.650 ;
        RECT 106.200 187.590 106.520 187.650 ;
        RECT 113.560 187.790 113.880 187.850 ;
        RECT 115.415 187.790 115.705 187.835 ;
        RECT 113.560 187.650 115.705 187.790 ;
        RECT 113.560 187.590 113.880 187.650 ;
        RECT 115.415 187.605 115.705 187.650 ;
        RECT 116.335 187.790 116.625 187.835 ;
        RECT 118.160 187.790 118.480 187.850 ;
        RECT 116.335 187.650 118.480 187.790 ;
        RECT 116.335 187.605 116.625 187.650 ;
        RECT 118.160 187.590 118.480 187.650 ;
        RECT 121.395 187.790 121.685 187.835 ;
        RECT 122.300 187.790 122.620 187.850 ;
        RECT 121.395 187.650 122.620 187.790 ;
        RECT 121.395 187.605 121.685 187.650 ;
        RECT 122.300 187.590 122.620 187.650 ;
        RECT 128.280 187.790 128.600 187.850 ;
        RECT 128.280 187.650 131.730 187.790 ;
        RECT 128.280 187.590 128.600 187.650 ;
        RECT 102.060 187.450 102.380 187.510 ;
        RECT 101.230 187.310 102.380 187.450 ;
        RECT 99.760 187.250 100.080 187.310 ;
        RECT 100.695 187.265 100.985 187.310 ;
        RECT 102.060 187.250 102.380 187.310 ;
        RECT 104.375 187.450 104.665 187.495 ;
        RECT 104.820 187.450 105.140 187.510 ;
        RECT 104.375 187.310 105.140 187.450 ;
        RECT 104.375 187.265 104.665 187.310 ;
        RECT 104.820 187.250 105.140 187.310 ;
        RECT 107.580 187.450 107.900 187.510 ;
        RECT 108.975 187.450 109.265 187.495 ;
        RECT 109.880 187.450 110.200 187.510 ;
        RECT 107.580 187.310 108.730 187.450 ;
        RECT 107.580 187.250 107.900 187.310 ;
        RECT 88.275 186.925 88.565 187.155 ;
        RECT 89.640 187.110 89.960 187.170 ;
        RECT 90.575 187.110 90.865 187.155 ;
        RECT 89.640 186.970 90.865 187.110 ;
        RECT 88.350 186.770 88.490 186.925 ;
        RECT 89.640 186.910 89.960 186.970 ;
        RECT 90.575 186.925 90.865 186.970 ;
        RECT 91.020 186.910 91.340 187.170 ;
        RECT 92.400 187.110 92.720 187.170 ;
        RECT 92.400 186.970 95.390 187.110 ;
        RECT 92.400 186.910 92.720 186.970 ;
        RECT 91.110 186.770 91.250 186.910 ;
        RECT 88.350 186.630 91.250 186.770 ;
        RECT 94.700 186.570 95.020 186.830 ;
        RECT 95.250 186.770 95.390 186.970 ;
        RECT 96.080 186.910 96.400 187.170 ;
        RECT 97.935 187.110 98.225 187.155 ;
        RECT 98.380 187.110 98.700 187.170 ;
        RECT 102.520 187.110 102.840 187.170 ;
        RECT 97.935 186.970 98.700 187.110 ;
        RECT 97.935 186.925 98.225 186.970 ;
        RECT 98.380 186.910 98.700 186.970 ;
        RECT 98.930 186.970 102.840 187.110 ;
        RECT 108.590 187.110 108.730 187.310 ;
        RECT 108.975 187.310 110.200 187.450 ;
        RECT 108.975 187.265 109.265 187.310 ;
        RECT 109.880 187.250 110.200 187.310 ;
        RECT 114.495 187.450 114.785 187.495 ;
        RECT 115.860 187.450 116.180 187.510 ;
        RECT 119.080 187.450 119.400 187.510 ;
        RECT 131.040 187.450 131.360 187.510 ;
        RECT 114.495 187.310 115.170 187.450 ;
        RECT 114.495 187.265 114.785 187.310 ;
        RECT 115.030 187.170 115.170 187.310 ;
        RECT 115.860 187.310 118.390 187.450 ;
        RECT 115.860 187.250 116.180 187.310 ;
        RECT 110.355 187.110 110.645 187.155 ;
        RECT 108.590 186.970 110.645 187.110 ;
        RECT 98.930 186.770 99.070 186.970 ;
        RECT 102.520 186.910 102.840 186.970 ;
        RECT 110.355 186.925 110.645 186.970 ;
        RECT 110.800 186.910 111.120 187.170 ;
        RECT 111.260 187.110 111.580 187.170 ;
        RECT 112.655 187.110 112.945 187.155 ;
        RECT 111.260 186.970 112.945 187.110 ;
        RECT 111.260 186.910 111.580 186.970 ;
        RECT 112.655 186.925 112.945 186.970 ;
        RECT 114.940 186.910 115.260 187.170 ;
        RECT 117.255 186.925 117.545 187.155 ;
        RECT 95.250 186.630 99.070 186.770 ;
        RECT 99.775 186.770 100.065 186.815 ;
        RECT 100.695 186.770 100.985 186.815 ;
        RECT 105.755 186.770 106.045 186.815 ;
        RECT 107.120 186.770 107.440 186.830 ;
        RECT 99.775 186.630 107.440 186.770 ;
        RECT 99.775 186.585 100.065 186.630 ;
        RECT 100.695 186.585 100.985 186.630 ;
        RECT 105.755 186.585 106.045 186.630 ;
        RECT 107.120 186.570 107.440 186.630 ;
        RECT 108.055 186.770 108.345 186.815 ;
        RECT 108.975 186.770 109.265 186.815 ;
        RECT 114.035 186.770 114.325 186.815 ;
        RECT 116.780 186.770 117.100 186.830 ;
        RECT 108.055 186.630 117.100 186.770 ;
        RECT 108.055 186.585 108.345 186.630 ;
        RECT 108.975 186.585 109.265 186.630 ;
        RECT 114.035 186.585 114.325 186.630 ;
        RECT 116.780 186.570 117.100 186.630 ;
        RECT 92.860 186.430 93.180 186.490 ;
        RECT 96.540 186.430 96.860 186.490 ;
        RECT 92.860 186.290 96.860 186.430 ;
        RECT 92.860 186.230 93.180 186.290 ;
        RECT 96.540 186.230 96.860 186.290 ;
        RECT 101.155 186.430 101.445 186.475 ;
        RECT 105.295 186.430 105.585 186.475 ;
        RECT 101.155 186.290 105.585 186.430 ;
        RECT 101.155 186.245 101.445 186.290 ;
        RECT 105.295 186.245 105.585 186.290 ;
        RECT 109.435 186.430 109.725 186.475 ;
        RECT 113.575 186.430 113.865 186.475 ;
        RECT 109.435 186.290 113.865 186.430 ;
        RECT 109.435 186.245 109.725 186.290 ;
        RECT 113.575 186.245 113.865 186.290 ;
        RECT 116.320 186.430 116.640 186.490 ;
        RECT 117.330 186.430 117.470 186.925 ;
        RECT 118.250 186.815 118.390 187.310 ;
        RECT 118.710 187.310 119.400 187.450 ;
        RECT 118.710 187.155 118.850 187.310 ;
        RECT 119.080 187.250 119.400 187.310 ;
        RECT 120.550 187.310 131.360 187.450 ;
        RECT 131.590 187.450 131.730 187.650 ;
        RECT 131.960 187.590 132.280 187.850 ;
        RECT 132.420 187.790 132.740 187.850 ;
        RECT 133.340 187.790 133.660 187.850 ;
        RECT 132.420 187.650 133.660 187.790 ;
        RECT 132.420 187.590 132.740 187.650 ;
        RECT 133.340 187.590 133.660 187.650 ;
        RECT 134.350 187.650 136.790 187.790 ;
        RECT 134.350 187.450 134.490 187.650 ;
        RECT 131.590 187.310 134.490 187.450 ;
        RECT 120.550 187.155 120.690 187.310 ;
        RECT 131.040 187.250 131.360 187.310 ;
        RECT 134.720 187.250 135.040 187.510 ;
        RECT 136.650 187.495 136.790 187.650 ;
        RECT 146.680 187.590 147.000 187.850 ;
        RECT 152.215 187.605 152.505 187.835 ;
        RECT 136.575 187.265 136.865 187.495 ;
        RECT 137.940 187.450 138.260 187.510 ;
        RECT 140.255 187.450 140.545 187.495 ;
        RECT 152.290 187.450 152.430 187.605 ;
        RECT 153.580 187.590 153.900 187.850 ;
        RECT 137.940 187.310 152.430 187.450 ;
        RECT 137.940 187.250 138.260 187.310 ;
        RECT 140.255 187.265 140.545 187.310 ;
        RECT 145.850 187.170 145.990 187.310 ;
        RECT 118.635 186.925 118.925 187.155 ;
        RECT 120.475 186.925 120.765 187.155 ;
        RECT 120.920 187.110 121.240 187.170 ;
        RECT 123.695 187.110 123.985 187.155 ;
        RECT 120.920 186.970 123.985 187.110 ;
        RECT 120.920 186.910 121.240 186.970 ;
        RECT 123.695 186.925 123.985 186.970 ;
        RECT 124.600 186.910 124.920 187.170 ;
        RECT 125.520 187.110 125.840 187.170 ;
        RECT 128.740 187.110 129.060 187.170 ;
        RECT 133.430 187.110 134.490 187.140 ;
        RECT 136.115 187.110 136.405 187.155 ;
        RECT 125.520 187.000 136.405 187.110 ;
        RECT 125.520 186.970 133.570 187.000 ;
        RECT 134.350 186.970 136.405 187.000 ;
        RECT 125.520 186.910 125.840 186.970 ;
        RECT 128.740 186.910 129.060 186.970 ;
        RECT 136.115 186.925 136.405 186.970 ;
        RECT 137.020 187.110 137.340 187.170 ;
        RECT 138.415 187.110 138.705 187.155 ;
        RECT 142.540 187.110 142.860 187.170 ;
        RECT 137.020 186.970 142.860 187.110 ;
        RECT 137.020 186.910 137.340 186.970 ;
        RECT 138.415 186.925 138.705 186.970 ;
        RECT 142.540 186.910 142.860 186.970 ;
        RECT 145.760 186.910 146.080 187.170 ;
        RECT 147.600 186.910 147.920 187.170 ;
        RECT 148.060 187.110 148.380 187.170 ;
        RECT 149.455 187.110 149.745 187.155 ;
        RECT 148.060 186.970 149.745 187.110 ;
        RECT 148.060 186.910 148.380 186.970 ;
        RECT 149.455 186.925 149.745 186.970 ;
        RECT 149.900 187.110 150.220 187.170 ;
        RECT 149.900 186.970 151.050 187.110 ;
        RECT 149.900 186.910 150.220 186.970 ;
        RECT 118.175 186.585 118.465 186.815 ;
        RECT 125.060 186.770 125.380 186.830 ;
        RECT 133.815 186.770 134.105 186.815 ;
        RECT 134.735 186.770 135.025 186.815 ;
        RECT 139.795 186.770 140.085 186.815 ;
        RECT 119.630 186.630 123.450 186.770 ;
        RECT 119.630 186.490 119.770 186.630 ;
        RECT 119.080 186.430 119.400 186.490 ;
        RECT 116.320 186.290 119.400 186.430 ;
        RECT 116.320 186.230 116.640 186.290 ;
        RECT 119.080 186.230 119.400 186.290 ;
        RECT 119.540 186.230 119.860 186.490 ;
        RECT 122.775 186.430 123.065 186.475 ;
        RECT 121.470 186.290 123.065 186.430 ;
        RECT 121.470 186.150 121.610 186.290 ;
        RECT 122.775 186.245 123.065 186.290 ;
        RECT 82.295 185.950 86.650 186.090 ;
        RECT 91.495 186.090 91.785 186.135 ;
        RECT 93.780 186.090 94.100 186.150 ;
        RECT 91.495 185.950 94.100 186.090 ;
        RECT 82.295 185.905 82.585 185.950 ;
        RECT 84.120 185.890 84.440 185.950 ;
        RECT 91.495 185.905 91.785 185.950 ;
        RECT 93.780 185.890 94.100 185.950 ;
        RECT 101.615 186.090 101.905 186.135 ;
        RECT 102.995 186.090 103.285 186.135 ;
        RECT 101.615 185.950 103.285 186.090 ;
        RECT 101.615 185.905 101.905 185.950 ;
        RECT 102.995 185.905 103.285 185.950 ;
        RECT 103.915 186.090 104.205 186.135 ;
        RECT 106.215 186.090 106.505 186.135 ;
        RECT 103.915 185.950 106.505 186.090 ;
        RECT 103.915 185.905 104.205 185.950 ;
        RECT 106.215 185.905 106.505 185.950 ;
        RECT 107.135 186.090 107.425 186.135 ;
        RECT 107.580 186.090 107.900 186.150 ;
        RECT 107.135 185.950 107.900 186.090 ;
        RECT 107.135 185.905 107.425 185.950 ;
        RECT 107.580 185.890 107.900 185.950 ;
        RECT 109.895 186.090 110.185 186.135 ;
        RECT 111.275 186.090 111.565 186.135 ;
        RECT 109.895 185.950 111.565 186.090 ;
        RECT 109.895 185.905 110.185 185.950 ;
        RECT 111.275 185.905 111.565 185.950 ;
        RECT 112.195 186.090 112.485 186.135 ;
        RECT 114.495 186.090 114.785 186.135 ;
        RECT 112.195 185.950 114.785 186.090 ;
        RECT 112.195 185.905 112.485 185.950 ;
        RECT 114.495 185.905 114.785 185.950 ;
        RECT 117.240 186.090 117.560 186.150 ;
        RECT 120.015 186.090 120.305 186.135 ;
        RECT 120.920 186.090 121.240 186.150 ;
        RECT 117.240 185.950 121.240 186.090 ;
        RECT 117.240 185.890 117.560 185.950 ;
        RECT 120.015 185.905 120.305 185.950 ;
        RECT 120.920 185.890 121.240 185.950 ;
        RECT 121.380 185.890 121.700 186.150 ;
        RECT 123.310 186.090 123.450 186.630 ;
        RECT 125.060 186.630 140.085 186.770 ;
        RECT 125.060 186.570 125.380 186.630 ;
        RECT 133.815 186.585 134.105 186.630 ;
        RECT 134.735 186.585 135.025 186.630 ;
        RECT 139.795 186.585 140.085 186.630 ;
        RECT 140.700 186.770 141.020 186.830 ;
        RECT 142.095 186.770 142.385 186.815 ;
        RECT 140.700 186.630 142.385 186.770 ;
        RECT 140.700 186.570 141.020 186.630 ;
        RECT 142.095 186.585 142.385 186.630 ;
        RECT 143.475 186.585 143.765 186.815 ;
        RECT 150.375 186.585 150.665 186.815 ;
        RECT 150.910 186.770 151.050 186.970 ;
        RECT 151.740 186.910 152.060 187.170 ;
        RECT 153.135 187.110 153.425 187.155 ;
        RECT 153.670 187.110 153.810 187.590 ;
        RECT 153.135 186.970 153.810 187.110 ;
        RECT 153.135 186.925 153.425 186.970 ;
        RECT 154.515 186.925 154.805 187.155 ;
        RECT 154.590 186.770 154.730 186.925 ;
        RECT 150.910 186.630 154.730 186.770 ;
        RECT 135.195 186.430 135.485 186.475 ;
        RECT 139.335 186.430 139.625 186.475 ;
        RECT 135.195 186.290 139.625 186.430 ;
        RECT 135.195 186.245 135.485 186.290 ;
        RECT 139.335 186.245 139.625 186.290 ;
        RECT 141.620 186.430 141.940 186.490 ;
        RECT 143.550 186.430 143.690 186.585 ;
        RECT 141.620 186.290 143.690 186.430 ;
        RECT 144.380 186.430 144.700 186.490 ;
        RECT 150.450 186.430 150.590 186.585 ;
        RECT 150.835 186.430 151.125 186.475 ;
        RECT 144.380 186.290 151.125 186.430 ;
        RECT 141.620 186.230 141.940 186.290 ;
        RECT 144.380 186.230 144.700 186.290 ;
        RECT 150.835 186.245 151.125 186.290 ;
        RECT 133.800 186.090 134.120 186.150 ;
        RECT 123.310 185.950 134.120 186.090 ;
        RECT 133.800 185.890 134.120 185.950 ;
        RECT 135.655 186.090 135.945 186.135 ;
        RECT 137.035 186.090 137.325 186.135 ;
        RECT 135.655 185.950 137.325 186.090 ;
        RECT 135.655 185.905 135.945 185.950 ;
        RECT 137.035 185.905 137.325 185.950 ;
        RECT 137.955 186.090 138.245 186.135 ;
        RECT 140.255 186.090 140.545 186.135 ;
        RECT 137.955 185.950 140.545 186.090 ;
        RECT 137.955 185.905 138.245 185.950 ;
        RECT 140.255 185.905 140.545 185.950 ;
        RECT 141.175 186.090 141.465 186.135 ;
        RECT 144.840 186.090 145.160 186.150 ;
        RECT 141.175 185.950 145.160 186.090 ;
        RECT 141.175 185.905 141.465 185.950 ;
        RECT 144.840 185.890 145.160 185.950 ;
        RECT 146.680 186.090 147.000 186.150 ;
        RECT 148.535 186.090 148.825 186.135 ;
        RECT 146.680 185.950 148.825 186.090 ;
        RECT 146.680 185.890 147.000 185.950 ;
        RECT 148.535 185.905 148.825 185.950 ;
        RECT 153.580 185.890 153.900 186.150 ;
        RECT 70.710 185.270 156.270 185.750 ;
        RECT 74.000 185.070 74.320 185.130 ;
        RECT 74.475 185.070 74.765 185.115 ;
        RECT 74.000 184.930 74.765 185.070 ;
        RECT 74.000 184.870 74.320 184.930 ;
        RECT 74.475 184.885 74.765 184.930 ;
        RECT 76.760 184.870 77.080 185.130 ;
        RECT 82.280 184.870 82.600 185.130 ;
        RECT 94.700 185.070 95.020 185.130 ;
        RECT 84.210 184.930 95.020 185.070 ;
        RECT 76.300 184.730 76.620 184.790 ;
        RECT 75.470 184.590 76.620 184.730 ;
        RECT 75.470 184.095 75.610 184.590 ;
        RECT 76.300 184.530 76.620 184.590 ;
        RECT 75.855 184.390 76.145 184.435 ;
        RECT 76.850 184.390 76.990 184.870 ;
        RECT 84.210 184.390 84.350 184.930 ;
        RECT 94.700 184.870 95.020 184.930 ;
        RECT 97.460 185.070 97.780 185.130 ;
        RECT 98.395 185.070 98.685 185.115 ;
        RECT 97.460 184.930 98.685 185.070 ;
        RECT 97.460 184.870 97.780 184.930 ;
        RECT 98.395 184.885 98.685 184.930 ;
        RECT 102.980 185.070 103.300 185.130 ;
        RECT 103.455 185.070 103.745 185.115 ;
        RECT 102.980 184.930 103.745 185.070 ;
        RECT 102.980 184.870 103.300 184.930 ;
        RECT 103.455 184.885 103.745 184.930 ;
        RECT 109.880 185.070 110.200 185.130 ;
        RECT 115.400 185.070 115.720 185.130 ;
        RECT 109.880 184.930 115.720 185.070 ;
        RECT 109.880 184.870 110.200 184.930 ;
        RECT 115.400 184.870 115.720 184.930 ;
        RECT 116.320 184.870 116.640 185.130 ;
        RECT 118.635 185.070 118.925 185.115 ;
        RECT 120.015 185.070 120.305 185.115 ;
        RECT 118.635 184.930 120.305 185.070 ;
        RECT 118.635 184.885 118.925 184.930 ;
        RECT 120.015 184.885 120.305 184.930 ;
        RECT 120.935 185.070 121.225 185.115 ;
        RECT 123.235 185.070 123.525 185.115 ;
        RECT 127.835 185.070 128.125 185.115 ;
        RECT 134.260 185.070 134.580 185.130 ;
        RECT 140.700 185.070 141.020 185.130 ;
        RECT 120.935 184.930 123.525 185.070 ;
        RECT 120.935 184.885 121.225 184.930 ;
        RECT 123.235 184.885 123.525 184.930 ;
        RECT 125.150 184.930 132.650 185.070 ;
        RECT 84.620 184.730 84.910 184.775 ;
        RECT 86.720 184.730 87.010 184.775 ;
        RECT 88.290 184.730 88.580 184.775 ;
        RECT 84.620 184.590 88.580 184.730 ;
        RECT 84.620 184.545 84.910 184.590 ;
        RECT 86.720 184.545 87.010 184.590 ;
        RECT 88.290 184.545 88.580 184.590 ;
        RECT 91.020 184.730 91.340 184.790 ;
        RECT 116.410 184.730 116.550 184.870 ;
        RECT 91.020 184.590 101.960 184.730 ;
        RECT 91.020 184.530 91.340 184.590 ;
        RECT 75.855 184.250 76.990 184.390 ;
        RECT 77.310 184.250 84.350 184.390 ;
        RECT 85.015 184.390 85.305 184.435 ;
        RECT 86.205 184.390 86.495 184.435 ;
        RECT 88.725 184.390 89.015 184.435 ;
        RECT 85.015 184.250 89.015 184.390 ;
        RECT 75.855 184.205 76.145 184.250 ;
        RECT 74.475 183.865 74.765 184.095 ;
        RECT 75.395 183.865 75.685 184.095 ;
        RECT 74.550 183.710 74.690 183.865 ;
        RECT 75.855 183.710 76.145 183.755 ;
        RECT 74.550 183.570 76.145 183.710 ;
        RECT 76.390 183.710 76.530 184.250 ;
        RECT 76.760 183.850 77.080 184.110 ;
        RECT 77.310 184.095 77.450 184.250 ;
        RECT 85.015 184.205 85.305 184.250 ;
        RECT 86.205 184.205 86.495 184.250 ;
        RECT 88.725 184.205 89.015 184.250 ;
        RECT 93.780 184.190 94.100 184.450 ;
        RECT 100.680 184.190 101.000 184.450 ;
        RECT 101.140 184.190 101.460 184.450 ;
        RECT 101.820 184.390 101.960 184.590 ;
        RECT 116.180 184.590 116.550 184.730 ;
        RECT 118.175 184.730 118.465 184.775 ;
        RECT 122.315 184.730 122.605 184.775 ;
        RECT 118.175 184.590 122.605 184.730 ;
        RECT 116.180 184.390 116.320 184.590 ;
        RECT 118.175 184.545 118.465 184.590 ;
        RECT 122.315 184.545 122.605 184.590 ;
        RECT 116.810 184.435 117.070 184.480 ;
        RECT 125.150 184.450 125.290 184.930 ;
        RECT 127.835 184.885 128.125 184.930 ;
        RECT 126.900 184.530 127.220 184.790 ;
        RECT 127.375 184.730 127.665 184.775 ;
        RECT 127.375 184.590 131.270 184.730 ;
        RECT 127.375 184.545 127.665 184.590 ;
        RECT 101.820 184.250 116.320 184.390 ;
        RECT 116.795 184.390 117.085 184.435 ;
        RECT 117.715 184.390 118.005 184.435 ;
        RECT 122.775 184.390 123.065 184.435 ;
        RECT 116.795 184.250 123.065 184.390 ;
        RECT 116.795 184.205 117.085 184.250 ;
        RECT 117.715 184.205 118.005 184.250 ;
        RECT 122.775 184.205 123.065 184.250 ;
        RECT 116.810 184.160 117.070 184.205 ;
        RECT 125.060 184.190 125.380 184.450 ;
        RECT 77.235 183.865 77.525 184.095 ;
        RECT 77.680 184.050 78.000 184.110 ;
        RECT 79.980 184.050 80.300 184.110 ;
        RECT 80.455 184.050 80.745 184.095 ;
        RECT 77.680 183.910 80.745 184.050 ;
        RECT 77.680 183.850 78.000 183.910 ;
        RECT 79.980 183.850 80.300 183.910 ;
        RECT 80.455 183.865 80.745 183.910 ;
        RECT 84.135 184.050 84.425 184.095 ;
        RECT 84.135 183.910 86.190 184.050 ;
        RECT 84.135 183.865 84.425 183.910 ;
        RECT 86.050 183.770 86.190 183.910 ;
        RECT 93.320 183.850 93.640 184.110 ;
        RECT 95.175 183.865 95.465 184.095 ;
        RECT 99.300 184.050 99.620 184.110 ;
        RECT 100.235 184.050 100.525 184.095 ;
        RECT 102.535 184.050 102.825 184.095 ;
        RECT 103.440 184.050 103.760 184.110 ;
        RECT 109.880 184.050 110.200 184.110 ;
        RECT 99.300 183.910 100.525 184.050 ;
        RECT 80.900 183.710 81.220 183.770 ;
        RECT 85.500 183.755 85.820 183.770 ;
        RECT 76.390 183.570 85.270 183.710 ;
        RECT 75.855 183.525 76.145 183.570 ;
        RECT 80.900 183.510 81.220 183.570 ;
        RECT 81.820 183.370 82.140 183.430 ;
        RECT 82.295 183.370 82.585 183.415 ;
        RECT 82.740 183.370 83.060 183.430 ;
        RECT 81.820 183.230 83.060 183.370 ;
        RECT 81.820 183.170 82.140 183.230 ;
        RECT 82.295 183.185 82.585 183.230 ;
        RECT 82.740 183.170 83.060 183.230 ;
        RECT 83.200 183.170 83.520 183.430 ;
        RECT 85.130 183.370 85.270 183.570 ;
        RECT 85.470 183.525 85.820 183.755 ;
        RECT 85.500 183.510 85.820 183.525 ;
        RECT 85.960 183.510 86.280 183.770 ;
        RECT 88.720 183.510 89.040 183.770 ;
        RECT 88.810 183.370 88.950 183.510 ;
        RECT 85.130 183.230 88.950 183.370 ;
        RECT 92.400 183.170 92.720 183.430 ;
        RECT 95.250 183.370 95.390 183.865 ;
        RECT 99.300 183.850 99.620 183.910 ;
        RECT 100.235 183.865 100.525 183.910 ;
        RECT 101.230 183.910 110.200 184.050 ;
        RECT 98.840 183.710 99.160 183.770 ;
        RECT 101.230 183.710 101.370 183.910 ;
        RECT 102.535 183.865 102.825 183.910 ;
        RECT 103.440 183.850 103.760 183.910 ;
        RECT 109.880 183.850 110.200 183.910 ;
        RECT 115.860 184.050 116.180 184.110 ;
        RECT 116.335 184.050 116.625 184.095 ;
        RECT 121.380 184.050 121.700 184.110 ;
        RECT 115.860 183.910 116.625 184.050 ;
        RECT 115.860 183.850 116.180 183.910 ;
        RECT 116.335 183.865 116.625 183.910 ;
        RECT 117.330 183.910 121.700 184.050 ;
        RECT 98.840 183.570 101.370 183.710 ;
        RECT 98.840 183.510 99.160 183.570 ;
        RECT 101.600 183.510 101.920 183.770 ;
        RECT 102.060 183.710 102.380 183.770 ;
        RECT 109.420 183.710 109.740 183.770 ;
        RECT 110.815 183.710 111.105 183.755 ;
        RECT 114.940 183.710 115.260 183.770 ;
        RECT 117.330 183.710 117.470 183.910 ;
        RECT 121.380 183.850 121.700 183.910 ;
        RECT 123.355 184.050 123.645 184.095 ;
        RECT 126.455 184.050 126.745 184.095 ;
        RECT 126.990 184.050 127.130 184.530 ;
        RECT 127.820 184.190 128.140 184.450 ;
        RECT 128.740 184.190 129.060 184.450 ;
        RECT 130.135 184.390 130.425 184.435 ;
        RECT 130.580 184.390 130.900 184.450 ;
        RECT 130.135 184.250 130.900 184.390 ;
        RECT 130.135 184.205 130.425 184.250 ;
        RECT 130.580 184.190 130.900 184.250 ;
        RECT 123.355 183.910 127.130 184.050 ;
        RECT 123.355 183.865 123.645 183.910 ;
        RECT 126.455 183.865 126.745 183.910 ;
        RECT 102.060 183.570 109.740 183.710 ;
        RECT 102.060 183.510 102.380 183.570 ;
        RECT 109.420 183.510 109.740 183.570 ;
        RECT 109.970 183.570 117.470 183.710 ;
        RECT 101.690 183.370 101.830 183.510 ;
        RECT 102.980 183.370 103.300 183.430 ;
        RECT 95.250 183.230 103.300 183.370 ;
        RECT 102.980 183.170 103.300 183.230 ;
        RECT 107.120 183.370 107.440 183.430 ;
        RECT 109.970 183.370 110.110 183.570 ;
        RECT 110.815 183.525 111.105 183.570 ;
        RECT 114.940 183.510 115.260 183.570 ;
        RECT 117.700 183.510 118.020 183.770 ;
        RECT 119.095 183.525 119.385 183.755 ;
        RECT 107.120 183.230 110.110 183.370 ;
        RECT 110.355 183.370 110.645 183.415 ;
        RECT 111.260 183.370 111.580 183.430 ;
        RECT 113.560 183.370 113.880 183.430 ;
        RECT 110.355 183.230 113.880 183.370 ;
        RECT 107.120 183.170 107.440 183.230 ;
        RECT 110.355 183.185 110.645 183.230 ;
        RECT 111.260 183.170 111.580 183.230 ;
        RECT 113.560 183.170 113.880 183.230 ;
        RECT 115.400 183.370 115.720 183.430 ;
        RECT 119.170 183.370 119.310 183.525 ;
        RECT 119.540 183.510 119.860 183.770 ;
        RECT 122.300 183.710 122.620 183.770 ;
        RECT 127.910 183.710 128.050 184.190 ;
        RECT 128.830 183.975 128.970 184.190 ;
        RECT 131.130 184.110 131.270 184.590 ;
        RECT 131.960 184.190 132.280 184.450 ;
        RECT 132.510 184.435 132.650 184.930 ;
        RECT 134.260 184.930 141.020 185.070 ;
        RECT 134.260 184.870 134.580 184.930 ;
        RECT 140.700 184.870 141.020 184.930 ;
        RECT 152.200 185.070 152.520 185.130 ;
        RECT 154.040 185.070 154.360 185.130 ;
        RECT 152.200 184.930 154.360 185.070 ;
        RECT 152.200 184.870 152.520 184.930 ;
        RECT 154.040 184.870 154.360 184.930 ;
        RECT 147.640 184.730 147.930 184.775 ;
        RECT 149.740 184.730 150.030 184.775 ;
        RECT 151.310 184.730 151.600 184.775 ;
        RECT 147.640 184.590 151.600 184.730 ;
        RECT 147.640 184.545 147.930 184.590 ;
        RECT 149.740 184.545 150.030 184.590 ;
        RECT 151.310 184.545 151.600 184.590 ;
        RECT 132.435 184.205 132.725 184.435 ;
        RECT 143.475 184.390 143.765 184.435 ;
        RECT 132.970 184.250 143.765 184.390 ;
        RECT 128.755 183.745 129.045 183.975 ;
        RECT 131.040 183.850 131.360 184.110 ;
        RECT 131.515 183.865 131.805 184.095 ;
        RECT 131.590 183.710 131.730 183.865 ;
        RECT 132.970 183.710 133.110 184.250 ;
        RECT 143.475 184.205 143.765 184.250 ;
        RECT 148.035 184.390 148.325 184.435 ;
        RECT 149.225 184.390 149.515 184.435 ;
        RECT 151.745 184.390 152.035 184.435 ;
        RECT 148.035 184.250 152.035 184.390 ;
        RECT 148.035 184.205 148.325 184.250 ;
        RECT 149.225 184.205 149.515 184.250 ;
        RECT 151.745 184.205 152.035 184.250 ;
        RECT 136.560 183.850 136.880 184.110 ;
        RECT 137.035 184.050 137.325 184.095 ;
        RECT 137.940 184.050 138.260 184.110 ;
        RECT 137.035 183.910 138.260 184.050 ;
        RECT 137.035 183.865 137.325 183.910 ;
        RECT 137.940 183.850 138.260 183.910 ;
        RECT 138.415 184.050 138.705 184.095 ;
        RECT 139.320 184.050 139.640 184.110 ;
        RECT 138.415 183.910 139.640 184.050 ;
        RECT 138.415 183.865 138.705 183.910 ;
        RECT 139.320 183.850 139.640 183.910 ;
        RECT 142.095 184.050 142.385 184.095 ;
        RECT 142.540 184.050 142.860 184.110 ;
        RECT 142.095 183.910 142.860 184.050 ;
        RECT 142.095 183.865 142.385 183.910 ;
        RECT 142.540 183.850 142.860 183.910 ;
        RECT 143.920 184.050 144.240 184.110 ;
        RECT 147.155 184.050 147.445 184.095 ;
        RECT 143.920 183.910 147.445 184.050 ;
        RECT 143.920 183.850 144.240 183.910 ;
        RECT 147.155 183.865 147.445 183.910 ;
        RECT 148.490 184.050 148.780 184.095 ;
        RECT 153.580 184.050 153.900 184.110 ;
        RECT 148.490 183.910 153.900 184.050 ;
        RECT 148.490 183.865 148.780 183.910 ;
        RECT 153.580 183.850 153.900 183.910 ;
        RECT 122.300 183.570 128.050 183.710 ;
        RECT 131.130 183.570 133.110 183.710 ;
        RECT 133.340 183.710 133.660 183.770 ;
        RECT 138.860 183.710 139.180 183.770 ;
        RECT 144.380 183.710 144.700 183.770 ;
        RECT 133.340 183.570 144.700 183.710 ;
        RECT 122.300 183.510 122.620 183.570 ;
        RECT 131.130 183.430 131.270 183.570 ;
        RECT 133.340 183.510 133.660 183.570 ;
        RECT 138.860 183.510 139.180 183.570 ;
        RECT 144.380 183.510 144.700 183.570 ;
        RECT 145.300 183.710 145.620 183.770 ;
        RECT 149.900 183.710 150.220 183.770 ;
        RECT 145.300 183.570 150.220 183.710 ;
        RECT 145.300 183.510 145.620 183.570 ;
        RECT 149.900 183.510 150.220 183.570 ;
        RECT 115.400 183.230 119.310 183.370 ;
        RECT 124.155 183.370 124.445 183.415 ;
        RECT 126.900 183.370 127.220 183.430 ;
        RECT 124.155 183.230 127.220 183.370 ;
        RECT 115.400 183.170 115.720 183.230 ;
        RECT 124.155 183.185 124.445 183.230 ;
        RECT 126.900 183.170 127.220 183.230 ;
        RECT 131.040 183.170 131.360 183.430 ;
        RECT 131.960 183.370 132.280 183.430 ;
        RECT 135.655 183.370 135.945 183.415 ;
        RECT 136.100 183.370 136.420 183.430 ;
        RECT 131.960 183.230 136.420 183.370 ;
        RECT 131.960 183.170 132.280 183.230 ;
        RECT 135.655 183.185 135.945 183.230 ;
        RECT 136.100 183.170 136.420 183.230 ;
        RECT 142.080 183.370 142.400 183.430 ;
        RECT 147.600 183.370 147.920 183.430 ;
        RECT 142.080 183.230 147.920 183.370 ;
        RECT 142.080 183.170 142.400 183.230 ;
        RECT 147.600 183.170 147.920 183.230 ;
        RECT 70.710 182.550 156.270 183.030 ;
        RECT 82.740 182.150 83.060 182.410 ;
        RECT 83.675 182.350 83.965 182.395 ;
        RECT 85.500 182.350 85.820 182.410 ;
        RECT 83.675 182.210 85.820 182.350 ;
        RECT 83.675 182.165 83.965 182.210 ;
        RECT 85.500 182.150 85.820 182.210 ;
        RECT 85.975 182.165 86.265 182.395 ;
        RECT 88.720 182.350 89.040 182.410 ;
        RECT 90.345 182.350 90.635 182.395 ;
        RECT 102.060 182.350 102.380 182.410 ;
        RECT 88.720 182.210 102.380 182.350 ;
        RECT 82.830 182.010 82.970 182.150 ;
        RECT 86.050 182.010 86.190 182.165 ;
        RECT 88.720 182.150 89.040 182.210 ;
        RECT 90.345 182.165 90.635 182.210 ;
        RECT 102.060 182.150 102.380 182.210 ;
        RECT 107.580 182.150 107.900 182.410 ;
        RECT 109.880 182.150 110.200 182.410 ;
        RECT 130.580 182.350 130.900 182.410 ;
        RECT 134.260 182.350 134.580 182.410 ;
        RECT 130.580 182.210 134.580 182.350 ;
        RECT 130.580 182.150 130.900 182.210 ;
        RECT 134.260 182.150 134.580 182.210 ;
        RECT 137.035 182.350 137.325 182.395 ;
        RECT 137.035 182.210 141.390 182.350 ;
        RECT 137.035 182.165 137.325 182.210 ;
        RECT 82.830 181.870 92.170 182.010 ;
        RECT 73.540 181.715 73.860 181.730 ;
        RECT 73.510 181.485 73.860 181.715 ;
        RECT 73.540 181.470 73.860 181.485 ;
        RECT 82.740 181.470 83.060 181.730 ;
        RECT 92.030 181.715 92.170 181.870 ;
        RECT 96.540 181.810 96.860 182.070 ;
        RECT 100.220 182.010 100.540 182.070 ;
        RECT 105.755 182.010 106.045 182.055 ;
        RECT 98.010 181.870 99.530 182.010 ;
        RECT 85.515 181.485 85.805 181.715 ;
        RECT 86.895 181.670 87.185 181.715 ;
        RECT 86.895 181.530 91.710 181.670 ;
        RECT 86.895 181.485 87.185 181.530 ;
        RECT 72.160 181.130 72.480 181.390 ;
        RECT 73.055 181.330 73.345 181.375 ;
        RECT 74.245 181.330 74.535 181.375 ;
        RECT 76.765 181.330 77.055 181.375 ;
        RECT 73.055 181.190 77.055 181.330 ;
        RECT 73.055 181.145 73.345 181.190 ;
        RECT 74.245 181.145 74.535 181.190 ;
        RECT 76.765 181.145 77.055 181.190 ;
        RECT 79.060 181.130 79.380 181.390 ;
        RECT 85.590 181.330 85.730 181.485 ;
        RECT 89.180 181.330 89.500 181.390 ;
        RECT 91.570 181.375 91.710 181.530 ;
        RECT 91.955 181.485 92.245 181.715 ;
        RECT 96.630 181.670 96.770 181.810 ;
        RECT 98.010 181.715 98.150 181.870 ;
        RECT 97.935 181.670 98.225 181.715 ;
        RECT 96.630 181.530 98.225 181.670 ;
        RECT 97.935 181.485 98.225 181.530 ;
        RECT 98.840 181.470 99.160 181.730 ;
        RECT 99.390 181.715 99.530 181.870 ;
        RECT 100.220 181.870 106.045 182.010 ;
        RECT 100.220 181.810 100.540 181.870 ;
        RECT 105.755 181.825 106.045 181.870 ;
        RECT 106.445 182.010 106.735 182.055 ;
        RECT 109.420 182.010 109.740 182.070 ;
        RECT 124.140 182.010 124.460 182.070 ;
        RECT 136.100 182.010 136.420 182.070 ;
        RECT 137.955 182.010 138.245 182.055 ;
        RECT 140.700 182.010 141.020 182.070 ;
        RECT 106.445 181.870 109.190 182.010 ;
        RECT 106.445 181.825 106.735 181.870 ;
        RECT 99.315 181.485 99.605 181.715 ;
        RECT 101.600 181.670 101.920 181.730 ;
        RECT 103.915 181.670 104.205 181.715 ;
        RECT 101.600 181.530 104.205 181.670 ;
        RECT 101.600 181.470 101.920 181.530 ;
        RECT 103.915 181.485 104.205 181.530 ;
        RECT 104.360 181.670 104.680 181.730 ;
        RECT 104.835 181.670 105.125 181.715 ;
        RECT 104.360 181.530 105.125 181.670 ;
        RECT 104.360 181.470 104.680 181.530 ;
        RECT 104.835 181.485 105.125 181.530 ;
        RECT 105.295 181.485 105.585 181.715 ;
        RECT 108.515 181.670 108.805 181.715 ;
        RECT 107.670 181.530 108.805 181.670 ;
        RECT 109.050 181.670 109.190 181.870 ;
        RECT 109.420 181.870 124.460 182.010 ;
        RECT 109.420 181.810 109.740 181.870 ;
        RECT 124.140 181.810 124.460 181.870 ;
        RECT 125.150 181.870 135.870 182.010 ;
        RECT 110.815 181.670 111.105 181.715 ;
        RECT 114.480 181.670 114.800 181.730 ;
        RECT 109.050 181.530 109.650 181.670 ;
        RECT 85.590 181.190 89.500 181.330 ;
        RECT 89.180 181.130 89.500 181.190 ;
        RECT 91.495 181.145 91.785 181.375 ;
        RECT 93.335 181.330 93.625 181.375 ;
        RECT 100.695 181.330 100.985 181.375 ;
        RECT 101.140 181.330 101.460 181.390 ;
        RECT 93.335 181.190 100.450 181.330 ;
        RECT 93.335 181.145 93.625 181.190 ;
        RECT 72.660 180.990 72.950 181.035 ;
        RECT 74.760 180.990 75.050 181.035 ;
        RECT 76.330 180.990 76.620 181.035 ;
        RECT 72.660 180.850 76.620 180.990 ;
        RECT 79.150 180.990 79.290 181.130 ;
        RECT 91.570 180.990 91.710 181.145 ;
        RECT 92.860 180.990 93.180 181.050 ;
        RECT 97.015 180.990 97.305 181.035 ;
        RECT 79.150 180.850 85.685 180.990 ;
        RECT 91.570 180.850 97.305 180.990 ;
        RECT 100.310 180.990 100.450 181.190 ;
        RECT 100.695 181.190 101.460 181.330 ;
        RECT 100.695 181.145 100.985 181.190 ;
        RECT 101.140 181.130 101.460 181.190 ;
        RECT 103.440 180.990 103.760 181.050 ;
        RECT 100.310 180.850 103.760 180.990 ;
        RECT 105.370 180.990 105.510 181.485 ;
        RECT 107.120 181.130 107.440 181.390 ;
        RECT 107.670 180.990 107.810 181.530 ;
        RECT 108.515 181.485 108.805 181.530 ;
        RECT 109.510 181.390 109.650 181.530 ;
        RECT 110.815 181.530 114.800 181.670 ;
        RECT 110.815 181.485 111.105 181.530 ;
        RECT 109.420 181.130 109.740 181.390 ;
        RECT 110.890 181.330 111.030 181.485 ;
        RECT 114.480 181.470 114.800 181.530 ;
        RECT 122.760 181.670 123.080 181.730 ;
        RECT 125.150 181.715 125.290 181.870 ;
        RECT 126.440 181.715 126.760 181.730 ;
        RECT 125.075 181.670 125.365 181.715 ;
        RECT 122.760 181.530 125.365 181.670 ;
        RECT 122.760 181.470 123.080 181.530 ;
        RECT 125.075 181.485 125.365 181.530 ;
        RECT 126.410 181.485 126.760 181.715 ;
        RECT 126.440 181.470 126.760 181.485 ;
        RECT 109.970 181.190 111.030 181.330 ;
        RECT 125.955 181.330 126.245 181.375 ;
        RECT 127.145 181.330 127.435 181.375 ;
        RECT 129.665 181.330 129.955 181.375 ;
        RECT 125.955 181.190 129.955 181.330 ;
        RECT 105.370 180.850 107.810 180.990 ;
        RECT 72.660 180.805 72.950 180.850 ;
        RECT 74.760 180.805 75.050 180.850 ;
        RECT 76.330 180.805 76.620 180.850 ;
        RECT 78.600 180.650 78.920 180.710 ;
        RECT 79.075 180.650 79.365 180.695 ;
        RECT 78.600 180.510 79.365 180.650 ;
        RECT 78.600 180.450 78.920 180.510 ;
        RECT 79.075 180.465 79.365 180.510 ;
        RECT 85.040 180.450 85.360 180.710 ;
        RECT 85.545 180.650 85.685 180.850 ;
        RECT 92.860 180.790 93.180 180.850 ;
        RECT 97.015 180.805 97.305 180.850 ;
        RECT 103.440 180.790 103.760 180.850 ;
        RECT 107.670 180.710 107.810 180.850 ;
        RECT 108.500 180.990 108.820 181.050 ;
        RECT 109.970 180.990 110.110 181.190 ;
        RECT 125.955 181.145 126.245 181.190 ;
        RECT 127.145 181.145 127.435 181.190 ;
        RECT 129.665 181.145 129.955 181.190 ;
        RECT 108.500 180.850 110.110 180.990 ;
        RECT 110.800 180.990 111.120 181.050 ;
        RECT 112.640 180.990 112.960 181.050 ;
        RECT 110.800 180.850 112.960 180.990 ;
        RECT 108.500 180.790 108.820 180.850 ;
        RECT 110.800 180.790 111.120 180.850 ;
        RECT 112.640 180.790 112.960 180.850 ;
        RECT 114.940 180.990 115.260 181.050 ;
        RECT 125.560 180.990 125.850 181.035 ;
        RECT 127.660 180.990 127.950 181.035 ;
        RECT 129.230 180.990 129.520 181.035 ;
        RECT 114.940 180.850 125.290 180.990 ;
        RECT 114.940 180.790 115.260 180.850 ;
        RECT 92.400 180.650 92.720 180.710 ;
        RECT 100.680 180.650 101.000 180.710 ;
        RECT 85.545 180.510 101.000 180.650 ;
        RECT 92.400 180.450 92.720 180.510 ;
        RECT 100.680 180.450 101.000 180.510 ;
        RECT 103.900 180.650 104.220 180.710 ;
        RECT 106.660 180.650 106.980 180.710 ;
        RECT 103.900 180.510 106.980 180.650 ;
        RECT 103.900 180.450 104.220 180.510 ;
        RECT 106.660 180.450 106.980 180.510 ;
        RECT 107.580 180.450 107.900 180.710 ;
        RECT 110.340 180.650 110.660 180.710 ;
        RECT 124.600 180.650 124.920 180.710 ;
        RECT 110.340 180.510 124.920 180.650 ;
        RECT 125.150 180.650 125.290 180.850 ;
        RECT 125.560 180.850 129.520 180.990 ;
        RECT 125.560 180.805 125.850 180.850 ;
        RECT 127.660 180.805 127.950 180.850 ;
        RECT 129.230 180.805 129.520 180.850 ;
        RECT 130.580 180.650 130.900 180.710 ;
        RECT 125.150 180.510 130.900 180.650 ;
        RECT 110.340 180.450 110.660 180.510 ;
        RECT 124.600 180.450 124.920 180.510 ;
        RECT 130.580 180.450 130.900 180.510 ;
        RECT 131.960 180.450 132.280 180.710 ;
        RECT 135.730 180.650 135.870 181.870 ;
        RECT 136.100 181.870 141.020 182.010 ;
        RECT 141.250 182.010 141.390 182.210 ;
        RECT 145.300 182.150 145.620 182.410 ;
        RECT 152.660 182.350 152.980 182.410 ;
        RECT 154.040 182.350 154.360 182.410 ;
        RECT 152.660 182.210 154.360 182.350 ;
        RECT 152.660 182.150 152.980 182.210 ;
        RECT 154.040 182.150 154.360 182.210 ;
        RECT 141.940 182.010 142.230 182.055 ;
        RECT 141.250 181.870 142.230 182.010 ;
        RECT 136.100 181.810 136.420 181.870 ;
        RECT 137.955 181.825 138.245 181.870 ;
        RECT 140.700 181.810 141.020 181.870 ;
        RECT 141.940 181.825 142.230 181.870 ;
        RECT 136.575 181.670 136.865 181.715 ;
        RECT 137.020 181.670 137.340 181.730 ;
        RECT 136.575 181.530 137.340 181.670 ;
        RECT 136.575 181.485 136.865 181.530 ;
        RECT 137.020 181.470 137.340 181.530 ;
        RECT 137.480 181.470 137.800 181.730 ;
        RECT 145.390 181.670 145.530 182.150 ;
        RECT 151.370 181.870 154.270 182.010 ;
        RECT 151.370 181.715 151.510 181.870 ;
        RECT 154.130 181.715 154.270 181.870 ;
        RECT 151.295 181.670 151.585 181.715 ;
        RECT 140.330 181.530 145.530 181.670 ;
        RECT 147.690 181.530 151.585 181.670 ;
        RECT 140.330 181.375 140.470 181.530 ;
        RECT 140.255 181.145 140.545 181.375 ;
        RECT 140.715 181.145 141.005 181.375 ;
        RECT 141.595 181.330 141.885 181.375 ;
        RECT 142.785 181.330 143.075 181.375 ;
        RECT 145.305 181.330 145.595 181.375 ;
        RECT 141.595 181.190 145.595 181.330 ;
        RECT 141.595 181.145 141.885 181.190 ;
        RECT 142.785 181.145 143.075 181.190 ;
        RECT 145.305 181.145 145.595 181.190 ;
        RECT 139.320 180.790 139.640 181.050 ;
        RECT 140.790 180.650 140.930 181.145 ;
        RECT 141.200 180.990 141.490 181.035 ;
        RECT 143.300 180.990 143.590 181.035 ;
        RECT 144.870 180.990 145.160 181.035 ;
        RECT 141.200 180.850 145.160 180.990 ;
        RECT 141.200 180.805 141.490 180.850 ;
        RECT 143.300 180.805 143.590 180.850 ;
        RECT 144.870 180.805 145.160 180.850 ;
        RECT 142.540 180.650 142.860 180.710 ;
        RECT 135.730 180.510 142.860 180.650 ;
        RECT 142.540 180.450 142.860 180.510 ;
        RECT 143.920 180.650 144.240 180.710 ;
        RECT 147.690 180.695 147.830 181.530 ;
        RECT 151.295 181.485 151.585 181.530 ;
        RECT 153.595 181.485 153.885 181.715 ;
        RECT 154.055 181.485 154.345 181.715 ;
        RECT 151.755 181.330 152.045 181.375 ;
        RECT 153.120 181.330 153.440 181.390 ;
        RECT 151.755 181.190 153.440 181.330 ;
        RECT 153.670 181.330 153.810 181.485 ;
        RECT 154.960 181.330 155.280 181.390 ;
        RECT 153.670 181.190 155.280 181.330 ;
        RECT 151.755 181.145 152.045 181.190 ;
        RECT 153.120 181.130 153.440 181.190 ;
        RECT 154.960 181.130 155.280 181.190 ;
        RECT 147.615 180.650 147.905 180.695 ;
        RECT 143.920 180.510 147.905 180.650 ;
        RECT 143.920 180.450 144.240 180.510 ;
        RECT 147.615 180.465 147.905 180.510 ;
        RECT 148.980 180.650 149.300 180.710 ;
        RECT 149.455 180.650 149.745 180.695 ;
        RECT 148.980 180.510 149.745 180.650 ;
        RECT 148.980 180.450 149.300 180.510 ;
        RECT 149.455 180.465 149.745 180.510 ;
        RECT 152.660 180.450 152.980 180.710 ;
        RECT 70.710 179.830 156.270 180.310 ;
        RECT 73.540 179.630 73.860 179.690 ;
        RECT 74.935 179.630 75.225 179.675 ;
        RECT 73.540 179.490 75.225 179.630 ;
        RECT 73.540 179.430 73.860 179.490 ;
        RECT 74.935 179.445 75.225 179.490 ;
        RECT 76.760 179.430 77.080 179.690 ;
        RECT 77.695 179.630 77.985 179.675 ;
        RECT 81.360 179.630 81.680 179.690 ;
        RECT 77.695 179.490 81.680 179.630 ;
        RECT 77.695 179.445 77.985 179.490 ;
        RECT 81.360 179.430 81.680 179.490 ;
        RECT 83.660 179.630 83.980 179.690 ;
        RECT 87.815 179.630 88.105 179.675 ;
        RECT 83.660 179.490 88.105 179.630 ;
        RECT 83.660 179.430 83.980 179.490 ;
        RECT 87.815 179.445 88.105 179.490 ;
        RECT 104.360 179.430 104.680 179.690 ;
        RECT 107.120 179.630 107.440 179.690 ;
        RECT 108.055 179.630 108.345 179.675 ;
        RECT 110.815 179.630 111.105 179.675 ;
        RECT 107.120 179.490 108.345 179.630 ;
        RECT 107.120 179.430 107.440 179.490 ;
        RECT 108.055 179.445 108.345 179.490 ;
        RECT 108.590 179.490 111.105 179.630 ;
        RECT 74.935 178.425 75.225 178.655 ;
        RECT 75.855 178.610 76.145 178.655 ;
        RECT 76.850 178.610 76.990 179.430 ;
        RECT 80.900 179.290 81.220 179.350 ;
        RECT 79.150 179.150 81.220 179.290 ;
        RECT 79.150 178.995 79.290 179.150 ;
        RECT 80.900 179.090 81.220 179.150 ;
        RECT 84.580 179.290 84.900 179.350 ;
        RECT 98.840 179.290 99.160 179.350 ;
        RECT 104.450 179.290 104.590 179.430 ;
        RECT 108.590 179.290 108.730 179.490 ;
        RECT 110.815 179.445 111.105 179.490 ;
        RECT 113.115 179.630 113.405 179.675 ;
        RECT 114.940 179.630 115.260 179.690 ;
        RECT 113.115 179.490 115.260 179.630 ;
        RECT 113.115 179.445 113.405 179.490 ;
        RECT 114.940 179.430 115.260 179.490 ;
        RECT 123.695 179.630 123.985 179.675 ;
        RECT 124.615 179.630 124.905 179.675 ;
        RECT 123.695 179.490 124.905 179.630 ;
        RECT 123.695 179.445 123.985 179.490 ;
        RECT 124.615 179.445 124.905 179.490 ;
        RECT 126.440 179.630 126.760 179.690 ;
        RECT 127.375 179.630 127.665 179.675 ;
        RECT 126.440 179.490 127.665 179.630 ;
        RECT 126.440 179.430 126.760 179.490 ;
        RECT 127.375 179.445 127.665 179.490 ;
        RECT 132.895 179.630 133.185 179.675 ;
        RECT 133.340 179.630 133.660 179.690 ;
        RECT 137.495 179.630 137.785 179.675 ;
        RECT 132.895 179.490 133.660 179.630 ;
        RECT 132.895 179.445 133.185 179.490 ;
        RECT 133.340 179.430 133.660 179.490 ;
        RECT 137.110 179.490 137.785 179.630 ;
        RECT 84.580 179.150 97.690 179.290 ;
        RECT 84.580 179.090 84.900 179.150 ;
        RECT 79.075 178.765 79.365 178.995 ;
        RECT 75.855 178.470 76.990 178.610 ;
        RECT 78.140 178.610 78.460 178.670 ;
        RECT 78.140 178.470 78.830 178.610 ;
        RECT 75.855 178.425 76.145 178.470 ;
        RECT 75.010 178.270 75.150 178.425 ;
        RECT 78.140 178.410 78.460 178.470 ;
        RECT 78.690 178.315 78.830 178.470 ;
        RECT 79.980 178.410 80.300 178.670 ;
        RECT 80.455 178.425 80.745 178.655 ;
        RECT 85.590 178.610 85.730 179.150 ;
        RECT 97.550 179.010 97.690 179.150 ;
        RECT 98.840 179.150 104.130 179.290 ;
        RECT 104.450 179.150 108.730 179.290 ;
        RECT 113.575 179.290 113.865 179.335 ;
        RECT 114.480 179.290 114.800 179.350 ;
        RECT 128.755 179.290 129.045 179.335 ;
        RECT 133.800 179.290 134.120 179.350 ;
        RECT 135.655 179.290 135.945 179.335 ;
        RECT 113.575 179.150 114.800 179.290 ;
        RECT 98.840 179.090 99.160 179.150 ;
        RECT 85.960 178.950 86.280 179.010 ;
        RECT 91.035 178.950 91.325 178.995 ;
        RECT 85.960 178.810 91.325 178.950 ;
        RECT 85.960 178.750 86.280 178.810 ;
        RECT 91.035 178.765 91.325 178.810 ;
        RECT 97.460 178.750 97.780 179.010 ;
        RECT 99.760 178.950 100.080 179.010 ;
        RECT 101.140 178.950 101.460 179.010 ;
        RECT 99.760 178.810 101.460 178.950 ;
        RECT 103.990 178.950 104.130 179.150 ;
        RECT 113.575 179.105 113.865 179.150 ;
        RECT 114.480 179.090 114.800 179.150 ;
        RECT 126.530 179.150 128.510 179.290 ;
        RECT 112.655 178.950 112.945 178.995 ;
        RECT 119.080 178.950 119.400 179.010 ;
        RECT 126.530 178.950 126.670 179.150 ;
        RECT 103.990 178.810 105.970 178.950 ;
        RECT 99.760 178.750 100.080 178.810 ;
        RECT 101.140 178.750 101.460 178.810 ;
        RECT 87.355 178.610 87.645 178.655 ;
        RECT 85.590 178.470 87.645 178.610 ;
        RECT 87.355 178.425 87.645 178.470 ;
        RECT 87.800 178.610 88.120 178.670 ;
        RECT 88.735 178.610 89.025 178.655 ;
        RECT 87.800 178.470 89.025 178.610 ;
        RECT 78.615 178.270 78.905 178.315 ;
        RECT 80.530 178.270 80.670 178.425 ;
        RECT 87.800 178.410 88.120 178.470 ;
        RECT 88.735 178.425 89.025 178.470 ;
        RECT 89.640 178.410 89.960 178.670 ;
        RECT 90.575 178.610 90.865 178.655 ;
        RECT 91.940 178.610 92.260 178.670 ;
        RECT 100.220 178.610 100.540 178.670 ;
        RECT 90.575 178.470 92.260 178.610 ;
        RECT 90.575 178.425 90.865 178.470 ;
        RECT 91.940 178.410 92.260 178.470 ;
        RECT 95.250 178.470 100.540 178.610 ;
        RECT 75.010 178.130 78.370 178.270 ;
        RECT 77.680 177.975 78.000 177.990 ;
        RECT 77.615 177.745 78.000 177.975 ;
        RECT 78.230 177.930 78.370 178.130 ;
        RECT 78.615 178.130 80.670 178.270 ;
        RECT 85.040 178.270 85.360 178.330 ;
        RECT 89.195 178.270 89.485 178.315 ;
        RECT 95.250 178.270 95.390 178.470 ;
        RECT 100.220 178.410 100.540 178.470 ;
        RECT 102.980 178.610 103.300 178.670 ;
        RECT 105.830 178.655 105.970 178.810 ;
        RECT 109.050 178.810 112.945 178.950 ;
        RECT 104.835 178.610 105.125 178.655 ;
        RECT 102.980 178.470 105.125 178.610 ;
        RECT 102.980 178.410 103.300 178.470 ;
        RECT 104.835 178.425 105.125 178.470 ;
        RECT 105.755 178.425 106.045 178.655 ;
        RECT 106.200 178.410 106.520 178.670 ;
        RECT 106.660 178.410 106.980 178.670 ;
        RECT 107.135 178.610 107.425 178.655 ;
        RECT 108.040 178.610 108.360 178.670 ;
        RECT 107.135 178.470 108.360 178.610 ;
        RECT 107.135 178.425 107.425 178.470 ;
        RECT 108.040 178.410 108.360 178.470 ;
        RECT 85.040 178.130 95.390 178.270 ;
        RECT 98.840 178.270 99.160 178.330 ;
        RECT 99.775 178.270 100.065 178.315 ;
        RECT 98.840 178.130 100.065 178.270 ;
        RECT 78.615 178.085 78.905 178.130 ;
        RECT 85.040 178.070 85.360 178.130 ;
        RECT 89.195 178.085 89.485 178.130 ;
        RECT 98.840 178.070 99.160 178.130 ;
        RECT 99.775 178.085 100.065 178.130 ;
        RECT 79.075 177.930 79.365 177.975 ;
        RECT 78.230 177.790 79.365 177.930 ;
        RECT 79.075 177.745 79.365 177.790 ;
        RECT 86.435 177.930 86.725 177.975 ;
        RECT 88.720 177.930 89.040 177.990 ;
        RECT 86.435 177.790 89.040 177.930 ;
        RECT 86.435 177.745 86.725 177.790 ;
        RECT 77.680 177.730 78.000 177.745 ;
        RECT 88.720 177.730 89.040 177.790 ;
        RECT 92.860 177.930 93.180 177.990 ;
        RECT 94.700 177.930 95.020 177.990 ;
        RECT 92.860 177.790 95.020 177.930 ;
        RECT 92.860 177.730 93.180 177.790 ;
        RECT 94.700 177.730 95.020 177.790 ;
        RECT 104.820 177.930 105.140 177.990 ;
        RECT 109.050 177.930 109.190 178.810 ;
        RECT 112.655 178.765 112.945 178.810 ;
        RECT 114.570 178.810 118.390 178.950 ;
        RECT 111.735 178.590 112.025 178.655 ;
        RECT 111.735 178.450 112.410 178.590 ;
        RECT 111.735 178.425 112.025 178.450 ;
        RECT 112.270 178.270 112.410 178.450 ;
        RECT 113.100 178.410 113.420 178.670 ;
        RECT 114.570 178.655 114.710 178.810 ;
        RECT 114.495 178.610 114.785 178.655 ;
        RECT 114.110 178.470 114.785 178.610 ;
        RECT 113.560 178.270 113.880 178.330 ;
        RECT 114.110 178.270 114.250 178.470 ;
        RECT 114.495 178.425 114.785 178.470 ;
        RECT 114.940 178.410 115.260 178.670 ;
        RECT 115.400 178.610 115.720 178.670 ;
        RECT 117.255 178.610 117.545 178.655 ;
        RECT 117.700 178.610 118.020 178.670 ;
        RECT 118.250 178.655 118.390 178.810 ;
        RECT 119.080 178.810 121.150 178.950 ;
        RECT 119.080 178.750 119.400 178.810 ;
        RECT 121.010 178.655 121.150 178.810 ;
        RECT 126.070 178.810 126.670 178.950 ;
        RECT 115.400 178.470 117.010 178.610 ;
        RECT 115.400 178.410 115.720 178.470 ;
        RECT 112.270 178.130 114.250 178.270 ;
        RECT 113.560 178.070 113.880 178.130 ;
        RECT 115.860 178.070 116.180 178.330 ;
        RECT 116.870 178.270 117.010 178.470 ;
        RECT 117.255 178.470 118.020 178.610 ;
        RECT 117.255 178.425 117.545 178.470 ;
        RECT 117.700 178.410 118.020 178.470 ;
        RECT 118.175 178.425 118.465 178.655 ;
        RECT 118.635 178.610 118.925 178.655 ;
        RECT 120.935 178.610 121.225 178.655 ;
        RECT 123.695 178.610 123.985 178.655 ;
        RECT 118.635 178.470 120.690 178.610 ;
        RECT 118.635 178.425 118.925 178.470 ;
        RECT 120.550 178.315 120.690 178.470 ;
        RECT 120.935 178.470 123.985 178.610 ;
        RECT 120.935 178.425 121.225 178.470 ;
        RECT 123.695 178.425 123.985 178.470 ;
        RECT 124.140 178.610 124.460 178.670 ;
        RECT 126.070 178.655 126.210 178.810 ;
        RECT 127.835 178.765 128.125 178.995 ;
        RECT 128.370 178.950 128.510 179.150 ;
        RECT 128.755 179.150 135.945 179.290 ;
        RECT 128.755 179.105 129.045 179.150 ;
        RECT 133.800 179.090 134.120 179.150 ;
        RECT 135.655 179.105 135.945 179.150 ;
        RECT 137.110 179.010 137.250 179.490 ;
        RECT 137.495 179.445 137.785 179.490 ;
        RECT 138.415 179.630 138.705 179.675 ;
        RECT 139.795 179.630 140.085 179.675 ;
        RECT 145.760 179.630 146.080 179.690 ;
        RECT 151.295 179.630 151.585 179.675 ;
        RECT 138.415 179.490 139.550 179.630 ;
        RECT 138.415 179.445 138.705 179.490 ;
        RECT 139.410 179.290 139.550 179.490 ;
        RECT 139.795 179.490 151.585 179.630 ;
        RECT 139.795 179.445 140.085 179.490 ;
        RECT 145.760 179.430 146.080 179.490 ;
        RECT 151.295 179.445 151.585 179.490 ;
        RECT 142.080 179.290 142.400 179.350 ;
        RECT 139.410 179.150 142.400 179.290 ;
        RECT 142.080 179.090 142.400 179.150 ;
        RECT 144.880 179.290 145.170 179.335 ;
        RECT 146.980 179.290 147.270 179.335 ;
        RECT 148.550 179.290 148.840 179.335 ;
        RECT 144.880 179.150 148.840 179.290 ;
        RECT 144.880 179.105 145.170 179.150 ;
        RECT 146.980 179.105 147.270 179.150 ;
        RECT 148.550 179.105 148.840 179.150 ;
        RECT 131.960 178.950 132.280 179.010 ;
        RECT 128.370 178.810 130.120 178.950 ;
        RECT 125.995 178.610 126.285 178.655 ;
        RECT 124.140 178.470 126.285 178.610 ;
        RECT 124.140 178.410 124.460 178.470 ;
        RECT 125.995 178.425 126.285 178.470 ;
        RECT 126.440 178.410 126.760 178.670 ;
        RECT 127.375 178.425 127.665 178.655 ;
        RECT 127.910 178.610 128.050 178.765 ;
        RECT 127.910 178.470 128.510 178.610 ;
        RECT 120.475 178.270 120.765 178.315 ;
        RECT 127.450 178.270 127.590 178.425 ;
        RECT 128.370 178.330 128.510 178.470 ;
        RECT 129.215 178.425 129.505 178.655 ;
        RECT 129.980 178.610 130.120 178.810 ;
        RECT 130.670 178.810 134.030 178.950 ;
        RECT 130.670 178.610 130.810 178.810 ;
        RECT 131.960 178.750 132.280 178.810 ;
        RECT 129.980 178.470 130.810 178.610 ;
        RECT 131.515 178.610 131.805 178.655 ;
        RECT 133.340 178.610 133.660 178.670 ;
        RECT 131.515 178.470 133.660 178.610 ;
        RECT 131.515 178.425 131.805 178.470 ;
        RECT 127.835 178.270 128.125 178.315 ;
        RECT 116.870 178.130 118.850 178.270 ;
        RECT 118.710 177.990 118.850 178.130 ;
        RECT 120.475 178.130 123.450 178.270 ;
        RECT 127.450 178.130 128.125 178.270 ;
        RECT 120.475 178.085 120.765 178.130 ;
        RECT 123.310 177.990 123.450 178.130 ;
        RECT 127.835 178.085 128.125 178.130 ;
        RECT 128.280 178.070 128.600 178.330 ;
        RECT 104.820 177.790 109.190 177.930 ;
        RECT 104.820 177.730 105.140 177.790 ;
        RECT 116.320 177.730 116.640 177.990 ;
        RECT 118.620 177.730 118.940 177.990 ;
        RECT 123.220 177.730 123.540 177.990 ;
        RECT 125.075 177.930 125.365 177.975 ;
        RECT 125.520 177.930 125.840 177.990 ;
        RECT 129.290 177.930 129.430 178.425 ;
        RECT 133.340 178.410 133.660 178.470 ;
        RECT 133.890 178.315 134.030 178.810 ;
        RECT 137.020 178.750 137.340 179.010 ;
        RECT 145.275 178.950 145.565 178.995 ;
        RECT 146.465 178.950 146.755 178.995 ;
        RECT 148.985 178.950 149.275 178.995 ;
        RECT 145.275 178.810 149.275 178.950 ;
        RECT 145.275 178.765 145.565 178.810 ;
        RECT 146.465 178.765 146.755 178.810 ;
        RECT 148.985 178.765 149.275 178.810 ;
        RECT 141.175 178.610 141.465 178.655 ;
        RECT 137.140 178.470 141.465 178.610 ;
        RECT 130.210 178.130 132.190 178.270 ;
        RECT 125.075 177.790 129.430 177.930 ;
        RECT 129.660 177.930 129.980 177.990 ;
        RECT 130.210 177.930 130.350 178.130 ;
        RECT 129.660 177.790 130.350 177.930 ;
        RECT 130.595 177.930 130.885 177.975 ;
        RECT 131.500 177.930 131.820 177.990 ;
        RECT 132.050 177.975 132.190 178.130 ;
        RECT 133.815 178.085 134.105 178.315 ;
        RECT 130.595 177.790 131.820 177.930 ;
        RECT 125.075 177.745 125.365 177.790 ;
        RECT 125.520 177.730 125.840 177.790 ;
        RECT 129.660 177.730 129.980 177.790 ;
        RECT 130.595 177.745 130.885 177.790 ;
        RECT 131.500 177.730 131.820 177.790 ;
        RECT 131.975 177.745 132.265 177.975 ;
        RECT 132.815 177.930 133.105 177.975 ;
        RECT 136.560 177.930 136.880 177.990 ;
        RECT 137.140 177.930 137.280 178.470 ;
        RECT 141.175 178.425 141.465 178.470 ;
        RECT 141.620 178.610 141.940 178.670 ;
        RECT 142.095 178.610 142.385 178.655 ;
        RECT 141.620 178.470 142.385 178.610 ;
        RECT 141.620 178.410 141.940 178.470 ;
        RECT 142.095 178.425 142.385 178.470 ;
        RECT 142.540 178.610 142.860 178.670 ;
        RECT 144.395 178.610 144.685 178.655 ;
        RECT 142.540 178.470 144.685 178.610 ;
        RECT 142.540 178.410 142.860 178.470 ;
        RECT 144.395 178.425 144.685 178.470 ;
        RECT 137.495 178.270 137.785 178.315 ;
        RECT 140.715 178.270 141.005 178.315 ;
        RECT 143.460 178.270 143.780 178.330 ;
        RECT 137.495 178.130 140.470 178.270 ;
        RECT 137.495 178.085 137.785 178.130 ;
        RECT 139.780 177.975 140.100 177.990 ;
        RECT 138.875 177.930 139.165 177.975 ;
        RECT 132.815 177.790 139.165 177.930 ;
        RECT 132.815 177.745 133.105 177.790 ;
        RECT 136.560 177.730 136.880 177.790 ;
        RECT 138.875 177.745 139.165 177.790 ;
        RECT 139.690 177.745 140.100 177.975 ;
        RECT 140.330 177.930 140.470 178.130 ;
        RECT 140.715 178.130 143.780 178.270 ;
        RECT 140.715 178.085 141.005 178.130 ;
        RECT 143.460 178.070 143.780 178.130 ;
        RECT 145.730 178.270 146.020 178.315 ;
        RECT 148.520 178.270 148.840 178.330 ;
        RECT 145.730 178.130 148.840 178.270 ;
        RECT 145.730 178.085 146.020 178.130 ;
        RECT 148.520 178.070 148.840 178.130 ;
        RECT 143.015 177.930 143.305 177.975 ;
        RECT 140.330 177.790 143.305 177.930 ;
        RECT 143.015 177.745 143.305 177.790 ;
        RECT 139.780 177.730 140.100 177.745 ;
        RECT 70.710 177.110 156.270 177.590 ;
        RECT 76.315 176.910 76.605 176.955 ;
        RECT 76.760 176.910 77.080 176.970 ;
        RECT 79.980 176.910 80.300 176.970 ;
        RECT 76.315 176.770 80.300 176.910 ;
        RECT 76.315 176.725 76.605 176.770 ;
        RECT 76.760 176.710 77.080 176.770 ;
        RECT 79.980 176.710 80.300 176.770 ;
        RECT 89.195 176.910 89.485 176.955 ;
        RECT 89.640 176.910 89.960 176.970 ;
        RECT 91.035 176.910 91.325 176.955 ;
        RECT 91.940 176.910 92.260 176.970 ;
        RECT 89.195 176.770 90.790 176.910 ;
        RECT 89.195 176.725 89.485 176.770 ;
        RECT 89.640 176.710 89.960 176.770 ;
        RECT 72.160 176.570 72.480 176.630 ;
        RECT 82.250 176.570 82.540 176.615 ;
        RECT 88.260 176.570 88.580 176.630 ;
        RECT 72.160 176.430 81.130 176.570 ;
        RECT 72.160 176.370 72.480 176.430 ;
        RECT 77.235 176.230 77.525 176.275 ;
        RECT 77.680 176.230 78.000 176.290 ;
        RECT 80.990 176.275 81.130 176.430 ;
        RECT 82.250 176.430 88.580 176.570 ;
        RECT 82.250 176.385 82.540 176.430 ;
        RECT 88.260 176.370 88.580 176.430 ;
        RECT 88.720 176.570 89.040 176.630 ;
        RECT 90.650 176.570 90.790 176.770 ;
        RECT 91.035 176.770 92.260 176.910 ;
        RECT 91.035 176.725 91.325 176.770 ;
        RECT 91.940 176.710 92.260 176.770 ;
        RECT 102.520 176.910 102.840 176.970 ;
        RECT 106.675 176.910 106.965 176.955 ;
        RECT 107.580 176.910 107.900 176.970 ;
        RECT 102.520 176.770 105.050 176.910 ;
        RECT 102.520 176.710 102.840 176.770 ;
        RECT 104.910 176.570 105.050 176.770 ;
        RECT 106.675 176.770 107.900 176.910 ;
        RECT 106.675 176.725 106.965 176.770 ;
        RECT 107.580 176.710 107.900 176.770 ;
        RECT 108.040 176.710 108.360 176.970 ;
        RECT 109.880 176.910 110.200 176.970 ;
        RECT 110.800 176.910 111.120 176.970 ;
        RECT 109.880 176.770 111.120 176.910 ;
        RECT 109.880 176.710 110.200 176.770 ;
        RECT 110.800 176.710 111.120 176.770 ;
        RECT 111.275 176.910 111.565 176.955 ;
        RECT 113.100 176.910 113.420 176.970 ;
        RECT 111.275 176.770 113.420 176.910 ;
        RECT 111.275 176.725 111.565 176.770 ;
        RECT 113.100 176.710 113.420 176.770 ;
        RECT 114.035 176.910 114.325 176.955 ;
        RECT 115.860 176.910 116.180 176.970 ;
        RECT 114.035 176.770 116.180 176.910 ;
        RECT 114.035 176.725 114.325 176.770 ;
        RECT 115.860 176.710 116.180 176.770 ;
        RECT 119.080 176.710 119.400 176.970 ;
        RECT 124.140 176.710 124.460 176.970 ;
        RECT 126.440 176.910 126.760 176.970 ;
        RECT 129.660 176.910 129.980 176.970 ;
        RECT 126.440 176.770 129.980 176.910 ;
        RECT 126.440 176.710 126.760 176.770 ;
        RECT 129.660 176.710 129.980 176.770 ;
        RECT 132.420 176.910 132.740 176.970 ;
        RECT 133.340 176.910 133.660 176.970 ;
        RECT 132.420 176.770 133.660 176.910 ;
        RECT 132.420 176.710 132.740 176.770 ;
        RECT 133.340 176.710 133.660 176.770 ;
        RECT 137.480 176.910 137.800 176.970 ;
        RECT 146.235 176.910 146.525 176.955 ;
        RECT 137.480 176.770 146.525 176.910 ;
        RECT 137.480 176.710 137.800 176.770 ;
        RECT 146.235 176.725 146.525 176.770 ;
        RECT 148.520 176.710 148.840 176.970 ;
        RECT 148.980 176.710 149.300 176.970 ;
        RECT 152.660 176.710 152.980 176.970 ;
        RECT 108.130 176.570 108.270 176.710 ;
        RECT 88.720 176.430 90.330 176.570 ;
        RECT 90.650 176.430 93.550 176.570 ;
        RECT 88.720 176.370 89.040 176.430 ;
        RECT 77.235 176.090 78.000 176.230 ;
        RECT 77.235 176.045 77.525 176.090 ;
        RECT 77.680 176.030 78.000 176.090 ;
        RECT 78.155 176.230 78.445 176.275 ;
        RECT 78.615 176.230 78.905 176.275 ;
        RECT 80.915 176.230 81.205 176.275 ;
        RECT 85.960 176.230 86.280 176.290 ;
        RECT 90.190 176.275 90.330 176.430 ;
        RECT 93.410 176.290 93.550 176.430 ;
        RECT 93.870 176.430 100.910 176.570 ;
        RECT 78.155 176.090 80.670 176.230 ;
        RECT 78.155 176.045 78.445 176.090 ;
        RECT 78.615 176.045 78.905 176.090 ;
        RECT 77.770 175.550 77.910 176.030 ;
        RECT 79.520 175.890 79.840 175.950 ;
        RECT 79.995 175.890 80.285 175.935 ;
        RECT 79.520 175.750 80.285 175.890 ;
        RECT 79.520 175.690 79.840 175.750 ;
        RECT 79.995 175.705 80.285 175.750 ;
        RECT 79.075 175.550 79.365 175.595 ;
        RECT 77.770 175.410 79.365 175.550 ;
        RECT 79.075 175.365 79.365 175.410 ;
        RECT 79.520 175.010 79.840 175.270 ;
        RECT 80.530 175.210 80.670 176.090 ;
        RECT 80.915 176.090 86.280 176.230 ;
        RECT 80.915 176.045 81.205 176.090 ;
        RECT 85.960 176.030 86.280 176.090 ;
        RECT 89.655 176.045 89.945 176.275 ;
        RECT 90.115 176.230 90.405 176.275 ;
        RECT 91.940 176.230 92.260 176.290 ;
        RECT 90.115 176.090 92.260 176.230 ;
        RECT 90.115 176.045 90.405 176.090 ;
        RECT 81.795 175.890 82.085 175.935 ;
        RECT 82.985 175.890 83.275 175.935 ;
        RECT 85.505 175.890 85.795 175.935 ;
        RECT 81.795 175.750 85.795 175.890 ;
        RECT 81.795 175.705 82.085 175.750 ;
        RECT 82.985 175.705 83.275 175.750 ;
        RECT 85.505 175.705 85.795 175.750 ;
        RECT 88.720 175.890 89.040 175.950 ;
        RECT 89.730 175.890 89.870 176.045 ;
        RECT 91.940 176.030 92.260 176.090 ;
        RECT 92.860 176.030 93.180 176.290 ;
        RECT 93.320 176.030 93.640 176.290 ;
        RECT 93.870 176.275 94.010 176.430 ;
        RECT 93.795 176.045 94.085 176.275 ;
        RECT 94.255 176.045 94.545 176.275 ;
        RECT 97.000 176.230 97.320 176.290 ;
        RECT 95.710 176.090 97.320 176.230 ;
        RECT 94.330 175.890 94.470 176.045 ;
        RECT 88.720 175.750 89.870 175.890 ;
        RECT 93.870 175.750 94.470 175.890 ;
        RECT 88.720 175.690 89.040 175.750 ;
        RECT 93.870 175.610 94.010 175.750 ;
        RECT 81.400 175.550 81.690 175.595 ;
        RECT 83.500 175.550 83.790 175.595 ;
        RECT 85.070 175.550 85.360 175.595 ;
        RECT 81.400 175.410 85.360 175.550 ;
        RECT 81.400 175.365 81.690 175.410 ;
        RECT 83.500 175.365 83.790 175.410 ;
        RECT 85.070 175.365 85.360 175.410 ;
        RECT 87.815 175.550 88.105 175.595 ;
        RECT 88.275 175.550 88.565 175.595 ;
        RECT 93.780 175.550 94.100 175.610 ;
        RECT 87.815 175.410 94.100 175.550 ;
        RECT 87.815 175.365 88.105 175.410 ;
        RECT 88.275 175.365 88.565 175.410 ;
        RECT 93.780 175.350 94.100 175.410 ;
        RECT 95.710 175.270 95.850 176.090 ;
        RECT 97.000 176.030 97.320 176.090 ;
        RECT 96.540 175.890 96.860 175.950 ;
        RECT 99.760 175.890 100.080 175.950 ;
        RECT 96.540 175.750 100.080 175.890 ;
        RECT 100.770 175.890 100.910 176.430 ;
        RECT 101.230 176.430 104.590 176.570 ;
        RECT 104.910 176.430 106.890 176.570 ;
        RECT 108.130 176.430 116.090 176.570 ;
        RECT 101.230 176.290 101.370 176.430 ;
        RECT 101.140 176.030 101.460 176.290 ;
        RECT 101.600 176.030 101.920 176.290 ;
        RECT 102.060 176.230 102.380 176.290 ;
        RECT 102.995 176.230 103.285 176.275 ;
        RECT 102.060 176.090 103.285 176.230 ;
        RECT 104.450 176.230 104.590 176.430 ;
        RECT 104.820 176.230 105.140 176.290 ;
        RECT 104.450 176.090 105.140 176.230 ;
        RECT 102.060 176.030 102.380 176.090 ;
        RECT 102.995 176.045 103.285 176.090 ;
        RECT 104.820 176.030 105.140 176.090 ;
        RECT 105.295 176.045 105.585 176.275 ;
        RECT 106.750 176.220 106.890 176.430 ;
        RECT 107.135 176.220 107.425 176.275 ;
        RECT 106.750 176.080 107.425 176.220 ;
        RECT 107.135 176.045 107.425 176.080 ;
        RECT 108.040 176.230 108.360 176.290 ;
        RECT 112.195 176.230 112.485 176.275 ;
        RECT 108.040 176.090 112.485 176.230 ;
        RECT 105.370 175.890 105.510 176.045 ;
        RECT 108.040 176.030 108.360 176.090 ;
        RECT 112.195 176.045 112.485 176.090 ;
        RECT 113.575 176.230 113.865 176.275 ;
        RECT 114.020 176.230 114.340 176.290 ;
        RECT 115.950 176.275 116.090 176.430 ;
        RECT 113.575 176.090 114.340 176.230 ;
        RECT 113.575 176.045 113.865 176.090 ;
        RECT 114.020 176.030 114.340 176.090 ;
        RECT 115.875 176.045 116.165 176.275 ;
        RECT 119.170 176.230 119.310 176.710 ;
        RECT 120.935 176.230 121.225 176.275 ;
        RECT 119.170 176.090 121.225 176.230 ;
        RECT 120.935 176.045 121.225 176.090 ;
        RECT 121.855 176.230 122.145 176.275 ;
        RECT 124.230 176.230 124.370 176.710 ;
        RECT 124.600 176.570 124.920 176.630 ;
        RECT 130.135 176.570 130.425 176.615 ;
        RECT 141.620 176.570 141.940 176.630 ;
        RECT 124.600 176.430 130.425 176.570 ;
        RECT 124.600 176.370 124.920 176.430 ;
        RECT 130.135 176.385 130.425 176.430 ;
        RECT 138.490 176.430 141.940 176.570 ;
        RECT 149.070 176.570 149.210 176.710 ;
        RECT 149.070 176.430 150.590 176.570 ;
        RECT 138.490 176.290 138.630 176.430 ;
        RECT 141.620 176.370 141.940 176.430 ;
        RECT 121.855 176.090 124.370 176.230 ;
        RECT 121.855 176.045 122.145 176.090 ;
        RECT 125.980 176.030 126.300 176.290 ;
        RECT 131.500 176.230 131.820 176.290 ;
        RECT 138.400 176.230 138.720 176.290 ;
        RECT 131.500 176.090 138.720 176.230 ;
        RECT 131.500 176.030 131.820 176.090 ;
        RECT 138.400 176.030 138.720 176.090 ;
        RECT 138.875 176.230 139.165 176.275 ;
        RECT 142.540 176.230 142.860 176.290 ;
        RECT 138.875 176.090 142.860 176.230 ;
        RECT 138.875 176.045 139.165 176.090 ;
        RECT 142.540 176.030 142.860 176.090 ;
        RECT 143.460 176.230 143.780 176.290 ;
        RECT 145.775 176.230 146.065 176.275 ;
        RECT 147.615 176.230 147.905 176.275 ;
        RECT 143.460 176.090 146.065 176.230 ;
        RECT 143.460 176.030 143.780 176.090 ;
        RECT 145.775 176.045 146.065 176.090 ;
        RECT 146.770 176.090 147.905 176.230 ;
        RECT 108.500 175.890 108.820 175.950 ;
        RECT 100.770 175.750 104.590 175.890 ;
        RECT 105.370 175.750 108.820 175.890 ;
        RECT 96.540 175.690 96.860 175.750 ;
        RECT 99.760 175.690 100.080 175.750 ;
        RECT 104.450 175.595 104.590 175.750 ;
        RECT 108.500 175.690 108.820 175.750 ;
        RECT 113.115 175.705 113.405 175.935 ;
        RECT 114.480 175.890 114.800 175.950 ;
        RECT 115.415 175.890 115.705 175.935 ;
        RECT 114.480 175.750 115.705 175.890 ;
        RECT 102.075 175.550 102.365 175.595 ;
        RECT 103.915 175.550 104.205 175.595 ;
        RECT 102.075 175.410 104.205 175.550 ;
        RECT 102.075 175.365 102.365 175.410 ;
        RECT 103.915 175.365 104.205 175.410 ;
        RECT 104.375 175.550 104.665 175.595 ;
        RECT 110.800 175.550 111.120 175.610 ;
        RECT 104.375 175.410 111.120 175.550 ;
        RECT 113.190 175.550 113.330 175.705 ;
        RECT 114.480 175.690 114.800 175.750 ;
        RECT 115.415 175.705 115.705 175.750 ;
        RECT 117.700 175.890 118.020 175.950 ;
        RECT 120.015 175.890 120.305 175.935 ;
        RECT 117.700 175.750 120.305 175.890 ;
        RECT 117.700 175.690 118.020 175.750 ;
        RECT 120.015 175.705 120.305 175.750 ;
        RECT 123.220 175.890 123.540 175.950 ;
        RECT 125.075 175.890 125.365 175.935 ;
        RECT 123.220 175.750 125.365 175.890 ;
        RECT 123.220 175.690 123.540 175.750 ;
        RECT 125.075 175.705 125.365 175.750 ;
        RECT 129.200 175.690 129.520 175.950 ;
        RECT 140.700 175.890 141.020 175.950 ;
        RECT 143.000 175.890 143.320 175.950 ;
        RECT 140.700 175.750 143.320 175.890 ;
        RECT 140.700 175.690 141.020 175.750 ;
        RECT 143.000 175.690 143.320 175.750 ;
        RECT 146.235 175.705 146.525 175.935 ;
        RECT 136.100 175.550 136.420 175.610 ;
        RECT 113.190 175.410 136.420 175.550 ;
        RECT 104.375 175.365 104.665 175.410 ;
        RECT 84.580 175.210 84.900 175.270 ;
        RECT 80.530 175.070 84.900 175.210 ;
        RECT 84.580 175.010 84.900 175.070 ;
        RECT 86.420 175.210 86.740 175.270 ;
        RECT 91.495 175.210 91.785 175.255 ;
        RECT 86.420 175.070 91.785 175.210 ;
        RECT 86.420 175.010 86.740 175.070 ;
        RECT 91.495 175.025 91.785 175.070 ;
        RECT 92.875 175.210 93.165 175.255 ;
        RECT 94.700 175.210 95.020 175.270 ;
        RECT 92.875 175.070 95.020 175.210 ;
        RECT 92.875 175.025 93.165 175.070 ;
        RECT 94.700 175.010 95.020 175.070 ;
        RECT 95.175 175.210 95.465 175.255 ;
        RECT 95.620 175.210 95.940 175.270 ;
        RECT 95.175 175.070 95.940 175.210 ;
        RECT 95.175 175.025 95.465 175.070 ;
        RECT 95.620 175.010 95.940 175.070 ;
        RECT 97.935 175.210 98.225 175.255 ;
        RECT 100.220 175.210 100.540 175.270 ;
        RECT 101.600 175.210 101.920 175.270 ;
        RECT 97.935 175.070 101.920 175.210 ;
        RECT 103.990 175.210 104.130 175.365 ;
        RECT 110.800 175.350 111.120 175.410 ;
        RECT 136.100 175.350 136.420 175.410 ;
        RECT 139.320 175.550 139.640 175.610 ;
        RECT 146.310 175.550 146.450 175.705 ;
        RECT 139.320 175.410 146.450 175.550 ;
        RECT 139.320 175.350 139.640 175.410 ;
        RECT 112.195 175.210 112.485 175.255 ;
        RECT 103.990 175.070 112.485 175.210 ;
        RECT 97.935 175.025 98.225 175.070 ;
        RECT 100.220 175.010 100.540 175.070 ;
        RECT 101.600 175.010 101.920 175.070 ;
        RECT 112.195 175.025 112.485 175.070 ;
        RECT 115.860 175.010 116.180 175.270 ;
        RECT 118.620 175.210 118.940 175.270 ;
        RECT 123.680 175.210 124.000 175.270 ;
        RECT 118.620 175.070 124.000 175.210 ;
        RECT 118.620 175.010 118.940 175.070 ;
        RECT 123.680 175.010 124.000 175.070 ;
        RECT 126.475 175.210 126.765 175.255 ;
        RECT 127.395 175.210 127.685 175.255 ;
        RECT 126.475 175.070 127.685 175.210 ;
        RECT 126.475 175.025 126.765 175.070 ;
        RECT 127.395 175.025 127.685 175.070 ;
        RECT 128.280 175.210 128.600 175.270 ;
        RECT 139.410 175.210 139.550 175.350 ;
        RECT 128.280 175.070 139.550 175.210 ;
        RECT 140.700 175.210 141.020 175.270 ;
        RECT 144.625 175.210 144.915 175.255 ;
        RECT 146.770 175.210 146.910 176.090 ;
        RECT 147.615 176.045 147.905 176.090 ;
        RECT 149.440 176.030 149.760 176.290 ;
        RECT 150.450 176.275 150.590 176.430 ;
        RECT 150.375 176.045 150.665 176.275 ;
        RECT 150.820 176.030 151.140 176.290 ;
        RECT 151.755 176.230 152.045 176.275 ;
        RECT 152.750 176.230 152.890 176.710 ;
        RECT 151.755 176.090 152.890 176.230 ;
        RECT 151.755 176.045 152.045 176.090 ;
        RECT 152.675 175.550 152.965 175.595 ;
        RECT 155.420 175.550 155.740 175.610 ;
        RECT 152.675 175.410 155.740 175.550 ;
        RECT 152.675 175.365 152.965 175.410 ;
        RECT 155.420 175.350 155.740 175.410 ;
        RECT 140.700 175.070 146.910 175.210 ;
        RECT 128.280 175.010 128.600 175.070 ;
        RECT 140.700 175.010 141.020 175.070 ;
        RECT 144.625 175.025 144.915 175.070 ;
        RECT 147.140 175.010 147.460 175.270 ;
        RECT 70.710 174.390 156.270 174.870 ;
        RECT 89.180 174.190 89.500 174.250 ;
        RECT 90.575 174.190 90.865 174.235 ;
        RECT 89.180 174.050 90.865 174.190 ;
        RECT 89.180 173.990 89.500 174.050 ;
        RECT 90.575 174.005 90.865 174.050 ;
        RECT 93.335 174.190 93.625 174.235 ;
        RECT 97.000 174.190 97.320 174.250 ;
        RECT 93.335 174.050 97.320 174.190 ;
        RECT 93.335 174.005 93.625 174.050 ;
        RECT 97.000 173.990 97.320 174.050 ;
        RECT 102.520 173.990 102.840 174.250 ;
        RECT 102.980 173.990 103.300 174.250 ;
        RECT 107.135 174.005 107.425 174.235 ;
        RECT 108.040 174.190 108.360 174.250 ;
        RECT 114.940 174.190 115.260 174.250 ;
        RECT 108.040 174.050 115.260 174.190 ;
        RECT 89.640 173.650 89.960 173.910 ;
        RECT 95.175 173.850 95.465 173.895 ;
        RECT 100.220 173.850 100.540 173.910 ;
        RECT 95.175 173.710 100.540 173.850 ;
        RECT 95.175 173.665 95.465 173.710 ;
        RECT 100.220 173.650 100.540 173.710 ;
        RECT 100.680 173.850 101.000 173.910 ;
        RECT 102.610 173.850 102.750 173.990 ;
        RECT 107.210 173.850 107.350 174.005 ;
        RECT 108.040 173.990 108.360 174.050 ;
        RECT 114.940 173.990 115.260 174.050 ;
        RECT 115.860 174.190 116.180 174.250 ;
        RECT 131.960 174.190 132.280 174.250 ;
        RECT 115.860 174.050 132.280 174.190 ;
        RECT 115.860 173.990 116.180 174.050 ;
        RECT 131.960 173.990 132.280 174.050 ;
        RECT 133.800 174.190 134.120 174.250 ;
        RECT 135.655 174.190 135.945 174.235 ;
        RECT 133.800 174.050 135.945 174.190 ;
        RECT 133.800 173.990 134.120 174.050 ;
        RECT 135.655 174.005 135.945 174.050 ;
        RECT 137.480 174.190 137.800 174.250 ;
        RECT 141.635 174.190 141.925 174.235 ;
        RECT 142.080 174.190 142.400 174.250 ;
        RECT 137.480 174.050 142.400 174.190 ;
        RECT 137.480 173.990 137.800 174.050 ;
        RECT 141.635 174.005 141.925 174.050 ;
        RECT 142.080 173.990 142.400 174.050 ;
        RECT 142.555 174.190 142.845 174.235 ;
        RECT 149.440 174.190 149.760 174.250 ;
        RECT 142.555 174.050 149.760 174.190 ;
        RECT 142.555 174.005 142.845 174.050 ;
        RECT 149.440 173.990 149.760 174.050 ;
        RECT 100.680 173.650 101.040 173.850 ;
        RECT 88.260 173.510 88.580 173.570 ;
        RECT 89.730 173.510 89.870 173.650 ;
        RECT 88.260 173.370 89.870 173.510 ;
        RECT 92.415 173.510 92.705 173.555 ;
        RECT 94.240 173.510 94.560 173.570 ;
        RECT 97.935 173.510 98.225 173.555 ;
        RECT 99.760 173.510 100.080 173.570 ;
        RECT 92.415 173.370 94.560 173.510 ;
        RECT 88.260 173.310 88.580 173.370 ;
        RECT 92.415 173.325 92.705 173.370 ;
        RECT 94.240 173.310 94.560 173.370 ;
        RECT 94.790 173.370 96.770 173.510 ;
        RECT 75.395 172.985 75.685 173.215 ;
        RECT 76.315 173.170 76.605 173.215 ;
        RECT 76.760 173.170 77.080 173.230 ;
        RECT 76.315 173.030 77.080 173.170 ;
        RECT 76.315 172.985 76.605 173.030 ;
        RECT 75.470 172.830 75.610 172.985 ;
        RECT 76.760 172.970 77.080 173.030 ;
        RECT 79.520 172.970 79.840 173.230 ;
        RECT 89.655 173.170 89.945 173.215 ;
        RECT 89.270 173.030 89.945 173.170 ;
        RECT 79.610 172.830 79.750 172.970 ;
        RECT 75.470 172.690 79.750 172.830 ;
        RECT 89.270 172.550 89.410 173.030 ;
        RECT 89.655 172.985 89.945 173.030 ;
        RECT 91.020 173.170 91.340 173.230 ;
        RECT 91.495 173.170 91.785 173.215 ;
        RECT 91.020 173.030 91.785 173.170 ;
        RECT 91.020 172.970 91.340 173.030 ;
        RECT 91.495 172.985 91.785 173.030 ;
        RECT 93.320 173.170 93.640 173.230 ;
        RECT 94.790 173.170 94.930 173.370 ;
        RECT 96.095 173.170 96.385 173.215 ;
        RECT 93.320 173.030 94.930 173.170 ;
        RECT 95.710 173.030 96.385 173.170 ;
        RECT 96.630 173.170 96.770 173.370 ;
        RECT 97.935 173.370 100.080 173.510 ;
        RECT 97.935 173.325 98.225 173.370 ;
        RECT 99.760 173.310 100.080 173.370 ;
        RECT 98.395 173.170 98.685 173.215 ;
        RECT 96.630 173.030 98.685 173.170 ;
        RECT 93.320 172.970 93.640 173.030 ;
        RECT 93.795 172.830 94.085 172.875 ;
        RECT 94.240 172.830 94.560 172.890 ;
        RECT 95.710 172.830 95.850 173.030 ;
        RECT 96.095 172.985 96.385 173.030 ;
        RECT 98.395 172.985 98.685 173.030 ;
        RECT 99.315 172.985 99.605 173.215 ;
        RECT 97.015 172.830 97.305 172.875 ;
        RECT 93.795 172.690 95.850 172.830 ;
        RECT 96.170 172.690 97.305 172.830 ;
        RECT 93.795 172.645 94.085 172.690 ;
        RECT 94.240 172.630 94.560 172.690 ;
        RECT 75.840 172.290 76.160 172.550 ;
        RECT 89.180 172.290 89.500 172.550 ;
        RECT 94.700 172.490 95.020 172.550 ;
        RECT 96.170 172.490 96.310 172.690 ;
        RECT 97.015 172.645 97.305 172.690 ;
        RECT 99.390 172.550 99.530 172.985 ;
        RECT 99.760 172.630 100.080 172.890 ;
        RECT 100.220 172.630 100.540 172.890 ;
        RECT 100.900 172.875 101.040 173.650 ;
        RECT 102.610 173.710 107.350 173.850 ;
        RECT 107.580 173.850 107.900 173.910 ;
        RECT 110.800 173.850 111.120 173.910 ;
        RECT 107.580 173.710 111.120 173.850 ;
        RECT 101.615 173.510 101.905 173.555 ;
        RECT 102.610 173.510 102.750 173.710 ;
        RECT 103.440 173.510 103.760 173.570 ;
        RECT 101.615 173.370 102.750 173.510 ;
        RECT 103.070 173.370 103.760 173.510 ;
        RECT 101.615 173.325 101.905 173.370 ;
        RECT 102.060 172.970 102.380 173.230 ;
        RECT 103.070 173.140 103.210 173.370 ;
        RECT 103.440 173.310 103.760 173.370 ;
        RECT 105.370 173.230 105.510 173.710 ;
        RECT 107.580 173.650 107.900 173.710 ;
        RECT 110.800 173.650 111.120 173.710 ;
        RECT 113.100 173.850 113.420 173.910 ;
        RECT 124.140 173.850 124.460 173.910 ;
        RECT 113.100 173.710 124.460 173.850 ;
        RECT 113.100 173.650 113.420 173.710 ;
        RECT 124.140 173.650 124.460 173.710 ;
        RECT 124.600 173.850 124.920 173.910 ;
        RECT 139.795 173.850 140.085 173.895 ;
        RECT 143.920 173.850 144.240 173.910 ;
        RECT 147.140 173.850 147.460 173.910 ;
        RECT 124.600 173.710 139.550 173.850 ;
        RECT 124.600 173.650 124.920 173.710 ;
        RECT 108.500 173.510 108.820 173.570 ;
        RECT 131.500 173.510 131.820 173.570 ;
        RECT 132.895 173.510 133.185 173.555 ;
        RECT 137.940 173.510 138.260 173.570 ;
        RECT 106.290 173.370 108.820 173.510 ;
        RECT 103.915 173.140 104.205 173.215 ;
        RECT 103.070 173.000 104.205 173.140 ;
        RECT 103.915 172.985 104.205 173.000 ;
        RECT 105.280 172.970 105.600 173.230 ;
        RECT 106.290 173.215 106.430 173.370 ;
        RECT 108.500 173.310 108.820 173.370 ;
        RECT 116.180 173.370 122.990 173.510 ;
        RECT 105.755 172.985 106.045 173.215 ;
        RECT 106.215 172.985 106.505 173.215 ;
        RECT 116.180 173.170 116.320 173.370 ;
        RECT 109.280 173.030 116.320 173.170 ;
        RECT 119.095 173.170 119.385 173.215 ;
        RECT 122.300 173.170 122.620 173.230 ;
        RECT 119.095 173.030 122.620 173.170 ;
        RECT 122.850 173.170 122.990 173.370 ;
        RECT 131.500 173.370 132.650 173.510 ;
        RECT 131.500 173.310 131.820 173.370 ;
        RECT 126.440 173.170 126.760 173.230 ;
        RECT 122.850 173.030 126.760 173.170 ;
        RECT 100.900 172.830 101.215 172.875 ;
        RECT 101.600 172.830 101.920 172.890 ;
        RECT 100.900 172.690 101.920 172.830 ;
        RECT 102.150 172.830 102.290 172.970 ;
        RECT 104.375 172.830 104.665 172.875 ;
        RECT 102.150 172.690 104.665 172.830 ;
        RECT 100.925 172.645 101.215 172.690 ;
        RECT 101.600 172.630 101.920 172.690 ;
        RECT 104.375 172.645 104.665 172.690 ;
        RECT 104.820 172.630 105.140 172.890 ;
        RECT 94.700 172.350 96.310 172.490 ;
        RECT 94.700 172.290 95.020 172.350 ;
        RECT 96.540 172.290 96.860 172.550 ;
        RECT 99.300 172.290 99.620 172.550 ;
        RECT 103.440 172.490 103.760 172.550 ;
        RECT 105.830 172.490 105.970 172.985 ;
        RECT 103.440 172.350 105.970 172.490 ;
        RECT 106.200 172.490 106.520 172.550 ;
        RECT 109.280 172.490 109.420 173.030 ;
        RECT 119.095 172.985 119.385 173.030 ;
        RECT 122.300 172.970 122.620 173.030 ;
        RECT 126.440 172.970 126.760 173.030 ;
        RECT 131.975 172.985 132.265 173.215 ;
        RECT 132.510 173.170 132.650 173.370 ;
        RECT 132.895 173.370 138.260 173.510 ;
        RECT 139.410 173.510 139.550 173.710 ;
        RECT 139.795 173.710 147.460 173.850 ;
        RECT 139.795 173.665 140.085 173.710 ;
        RECT 143.920 173.650 144.240 173.710 ;
        RECT 147.140 173.650 147.460 173.710 ;
        RECT 144.380 173.510 144.700 173.570 ;
        RECT 139.410 173.370 144.700 173.510 ;
        RECT 132.895 173.325 133.185 173.370 ;
        RECT 137.940 173.310 138.260 173.370 ;
        RECT 144.380 173.310 144.700 173.370 ;
        RECT 145.760 173.310 146.080 173.570 ;
        RECT 148.980 173.510 149.300 173.570 ;
        RECT 149.915 173.510 150.205 173.555 ;
        RECT 148.980 173.370 150.205 173.510 ;
        RECT 148.980 173.310 149.300 173.370 ;
        RECT 149.915 173.325 150.205 173.370 ;
        RECT 133.355 173.170 133.645 173.215 ;
        RECT 132.510 173.030 133.645 173.170 ;
        RECT 133.355 172.985 133.645 173.030 ;
        RECT 134.275 173.170 134.565 173.215 ;
        RECT 134.720 173.170 135.040 173.230 ;
        RECT 134.275 173.030 135.040 173.170 ;
        RECT 134.275 172.985 134.565 173.030 ;
        RECT 111.275 172.830 111.565 172.875 ;
        RECT 110.430 172.690 111.565 172.830 ;
        RECT 110.430 172.550 110.570 172.690 ;
        RECT 111.275 172.645 111.565 172.690 ;
        RECT 113.100 172.830 113.420 172.890 ;
        RECT 132.050 172.830 132.190 172.985 ;
        RECT 134.720 172.970 135.040 173.030 ;
        RECT 136.575 173.170 136.865 173.215 ;
        RECT 137.020 173.170 137.340 173.230 ;
        RECT 136.575 173.030 137.340 173.170 ;
        RECT 136.575 172.985 136.865 173.030 ;
        RECT 137.020 172.970 137.340 173.030 ;
        RECT 137.495 173.170 137.785 173.215 ;
        RECT 138.400 173.170 138.720 173.230 ;
        RECT 144.855 173.170 145.145 173.215 ;
        RECT 137.495 173.030 138.720 173.170 ;
        RECT 137.495 172.985 137.785 173.030 ;
        RECT 138.400 172.970 138.720 173.030 ;
        RECT 141.710 173.030 145.145 173.170 ;
        RECT 145.850 173.170 145.990 173.310 ;
        RECT 146.235 173.170 146.525 173.215 ;
        RECT 147.140 173.170 147.460 173.230 ;
        RECT 150.375 173.170 150.665 173.215 ;
        RECT 145.850 173.030 147.460 173.170 ;
        RECT 133.815 172.830 134.105 172.875 ;
        RECT 139.780 172.830 140.100 172.890 ;
        RECT 141.710 172.875 141.850 173.030 ;
        RECT 144.855 172.985 145.145 173.030 ;
        RECT 146.235 172.985 146.525 173.030 ;
        RECT 147.140 172.970 147.460 173.030 ;
        RECT 149.070 173.030 150.665 173.170 ;
        RECT 113.100 172.690 130.120 172.830 ;
        RECT 132.050 172.690 140.100 172.830 ;
        RECT 113.100 172.630 113.420 172.690 ;
        RECT 106.200 172.350 109.420 172.490 ;
        RECT 103.440 172.290 103.760 172.350 ;
        RECT 106.200 172.290 106.520 172.350 ;
        RECT 110.340 172.290 110.660 172.550 ;
        RECT 110.800 172.490 111.120 172.550 ;
        RECT 119.080 172.490 119.400 172.550 ;
        RECT 110.800 172.350 119.400 172.490 ;
        RECT 129.980 172.490 130.120 172.690 ;
        RECT 133.815 172.645 134.105 172.690 ;
        RECT 139.780 172.630 140.100 172.690 ;
        RECT 141.635 172.645 141.925 172.875 ;
        RECT 143.015 172.645 143.305 172.875 ;
        RECT 143.460 172.830 143.780 172.890 ;
        RECT 143.935 172.830 144.225 172.875 ;
        RECT 143.460 172.690 144.225 172.830 ;
        RECT 131.055 172.490 131.345 172.535 ;
        RECT 129.980 172.350 131.345 172.490 ;
        RECT 110.800 172.290 111.120 172.350 ;
        RECT 119.080 172.290 119.400 172.350 ;
        RECT 131.055 172.305 131.345 172.350 ;
        RECT 135.640 172.490 135.960 172.550 ;
        RECT 143.090 172.490 143.230 172.645 ;
        RECT 143.460 172.630 143.780 172.690 ;
        RECT 143.935 172.645 144.225 172.690 ;
        RECT 135.640 172.350 143.230 172.490 ;
        RECT 144.010 172.490 144.150 172.645 ;
        RECT 149.070 172.550 149.210 173.030 ;
        RECT 150.375 172.985 150.665 173.030 ;
        RECT 145.315 172.490 145.605 172.535 ;
        RECT 144.010 172.350 145.605 172.490 ;
        RECT 135.640 172.290 135.960 172.350 ;
        RECT 145.315 172.305 145.605 172.350 ;
        RECT 148.980 172.290 149.300 172.550 ;
        RECT 152.215 172.490 152.505 172.535 ;
        RECT 152.660 172.490 152.980 172.550 ;
        RECT 152.215 172.350 152.980 172.490 ;
        RECT 152.215 172.305 152.505 172.350 ;
        RECT 152.660 172.290 152.980 172.350 ;
        RECT 70.710 171.670 156.270 172.150 ;
        RECT 86.895 171.470 87.185 171.515 ;
        RECT 87.800 171.470 88.120 171.530 ;
        RECT 86.895 171.330 88.120 171.470 ;
        RECT 86.895 171.285 87.185 171.330 ;
        RECT 87.800 171.270 88.120 171.330 ;
        RECT 88.720 171.270 89.040 171.530 ;
        RECT 89.655 171.470 89.945 171.515 ;
        RECT 91.480 171.470 91.800 171.530 ;
        RECT 89.655 171.330 91.800 171.470 ;
        RECT 89.655 171.285 89.945 171.330 ;
        RECT 91.480 171.270 91.800 171.330 ;
        RECT 92.415 171.470 92.705 171.515 ;
        RECT 92.860 171.470 93.180 171.530 ;
        RECT 92.415 171.330 93.180 171.470 ;
        RECT 92.415 171.285 92.705 171.330 ;
        RECT 92.860 171.270 93.180 171.330 ;
        RECT 93.320 171.270 93.640 171.530 ;
        RECT 94.700 171.470 95.020 171.530 ;
        RECT 95.175 171.470 95.465 171.515 ;
        RECT 94.700 171.330 95.465 171.470 ;
        RECT 94.700 171.270 95.020 171.330 ;
        RECT 95.175 171.285 95.465 171.330 ;
        RECT 97.460 171.470 97.780 171.530 ;
        RECT 98.015 171.470 98.305 171.515 ;
        RECT 97.460 171.330 98.305 171.470 ;
        RECT 97.460 171.270 97.780 171.330 ;
        RECT 98.015 171.285 98.305 171.330 ;
        RECT 99.760 171.470 100.080 171.530 ;
        RECT 102.535 171.470 102.825 171.515 ;
        RECT 107.595 171.470 107.885 171.515 ;
        RECT 99.760 171.330 102.825 171.470 ;
        RECT 99.760 171.270 100.080 171.330 ;
        RECT 102.535 171.285 102.825 171.330 ;
        RECT 103.070 171.330 107.885 171.470 ;
        RECT 80.870 171.130 81.160 171.175 ;
        RECT 93.410 171.130 93.550 171.270 ;
        RECT 97.015 171.130 97.305 171.175 ;
        RECT 103.070 171.130 103.210 171.330 ;
        RECT 107.595 171.285 107.885 171.330 ;
        RECT 113.560 171.470 113.880 171.530 ;
        RECT 114.495 171.470 114.785 171.515 ;
        RECT 119.095 171.470 119.385 171.515 ;
        RECT 113.560 171.330 119.385 171.470 ;
        RECT 113.560 171.270 113.880 171.330 ;
        RECT 114.495 171.285 114.785 171.330 ;
        RECT 119.095 171.285 119.385 171.330 ;
        RECT 120.000 171.470 120.320 171.530 ;
        RECT 124.600 171.470 124.920 171.530 ;
        RECT 120.000 171.330 124.920 171.470 ;
        RECT 120.000 171.270 120.320 171.330 ;
        RECT 124.600 171.270 124.920 171.330 ;
        RECT 129.660 171.470 129.980 171.530 ;
        RECT 130.580 171.470 130.900 171.530 ;
        RECT 131.515 171.470 131.805 171.515 ;
        RECT 129.660 171.270 130.120 171.470 ;
        RECT 130.580 171.330 131.805 171.470 ;
        RECT 130.580 171.270 130.900 171.330 ;
        RECT 131.515 171.285 131.805 171.330 ;
        RECT 131.960 171.470 132.280 171.530 ;
        RECT 136.115 171.470 136.405 171.515 ;
        RECT 137.020 171.470 137.340 171.530 ;
        RECT 131.960 171.330 137.340 171.470 ;
        RECT 131.960 171.270 132.280 171.330 ;
        RECT 136.115 171.285 136.405 171.330 ;
        RECT 137.020 171.270 137.340 171.330 ;
        RECT 139.795 171.470 140.085 171.515 ;
        RECT 143.920 171.470 144.240 171.530 ;
        RECT 139.795 171.330 144.240 171.470 ;
        RECT 139.795 171.285 140.085 171.330 ;
        RECT 143.920 171.270 144.240 171.330 ;
        RECT 144.380 171.470 144.700 171.530 ;
        RECT 151.295 171.470 151.585 171.515 ;
        RECT 155.880 171.470 156.200 171.530 ;
        RECT 144.380 171.330 150.130 171.470 ;
        RECT 144.380 171.270 144.700 171.330 ;
        RECT 72.250 170.990 79.750 171.130 ;
        RECT 72.250 170.510 72.390 170.990 ;
        RECT 73.510 170.790 73.800 170.835 ;
        RECT 75.840 170.790 76.160 170.850 ;
        RECT 79.610 170.835 79.750 170.990 ;
        RECT 80.870 170.990 93.550 171.130 ;
        RECT 93.870 170.990 97.305 171.130 ;
        RECT 80.870 170.945 81.160 170.990 ;
        RECT 73.510 170.650 76.160 170.790 ;
        RECT 73.510 170.605 73.800 170.650 ;
        RECT 75.840 170.590 76.160 170.650 ;
        RECT 79.535 170.605 79.825 170.835 ;
        RECT 87.340 170.790 87.660 170.850 ;
        RECT 87.815 170.790 88.105 170.835 ;
        RECT 87.340 170.650 88.105 170.790 ;
        RECT 87.340 170.590 87.660 170.650 ;
        RECT 87.815 170.605 88.105 170.650 ;
        RECT 88.260 170.590 88.580 170.850 ;
        RECT 90.575 170.790 90.865 170.835 ;
        RECT 91.940 170.790 92.260 170.850 ;
        RECT 90.575 170.650 92.260 170.790 ;
        RECT 90.575 170.605 90.865 170.650 ;
        RECT 91.940 170.590 92.260 170.650 ;
        RECT 93.320 170.590 93.640 170.850 ;
        RECT 72.160 170.250 72.480 170.510 ;
        RECT 73.055 170.450 73.345 170.495 ;
        RECT 74.245 170.450 74.535 170.495 ;
        RECT 76.765 170.450 77.055 170.495 ;
        RECT 73.055 170.310 77.055 170.450 ;
        RECT 73.055 170.265 73.345 170.310 ;
        RECT 74.245 170.265 74.535 170.310 ;
        RECT 76.765 170.265 77.055 170.310 ;
        RECT 80.415 170.450 80.705 170.495 ;
        RECT 81.605 170.450 81.895 170.495 ;
        RECT 84.125 170.450 84.415 170.495 ;
        RECT 80.415 170.310 84.415 170.450 ;
        RECT 80.415 170.265 80.705 170.310 ;
        RECT 81.605 170.265 81.895 170.310 ;
        RECT 84.125 170.265 84.415 170.310 ;
        RECT 89.640 170.450 89.960 170.510 ;
        RECT 90.115 170.450 90.405 170.495 ;
        RECT 89.640 170.310 90.405 170.450 ;
        RECT 89.640 170.250 89.960 170.310 ;
        RECT 90.115 170.265 90.405 170.310 ;
        RECT 91.035 170.450 91.325 170.495 ;
        RECT 93.870 170.450 94.010 170.990 ;
        RECT 97.015 170.945 97.305 170.990 ;
        RECT 97.550 170.990 103.210 171.130 ;
        RECT 103.455 171.130 103.745 171.175 ;
        RECT 105.280 171.130 105.600 171.190 ;
        RECT 120.935 171.130 121.225 171.175 ;
        RECT 103.455 170.990 105.970 171.130 ;
        RECT 94.240 170.590 94.560 170.850 ;
        RECT 94.715 170.790 95.005 170.835 ;
        RECT 96.540 170.790 96.860 170.850 ;
        RECT 97.550 170.790 97.690 170.990 ;
        RECT 103.455 170.945 103.745 170.990 ;
        RECT 105.280 170.930 105.600 170.990 ;
        RECT 94.715 170.650 97.690 170.790 ;
        RECT 100.235 170.790 100.525 170.835 ;
        RECT 102.060 170.790 102.380 170.850 ;
        RECT 100.235 170.650 102.380 170.790 ;
        RECT 94.715 170.605 95.005 170.650 ;
        RECT 96.540 170.590 96.860 170.650 ;
        RECT 100.235 170.605 100.525 170.650 ;
        RECT 102.060 170.590 102.380 170.650 ;
        RECT 103.900 170.790 104.220 170.850 ;
        RECT 105.830 170.835 105.970 170.990 ;
        RECT 109.050 170.990 116.090 171.130 ;
        RECT 109.050 170.835 109.190 170.990 ;
        RECT 112.730 170.835 112.870 170.990 ;
        RECT 104.375 170.790 104.665 170.835 ;
        RECT 104.835 170.790 105.125 170.835 ;
        RECT 103.900 170.650 105.125 170.790 ;
        RECT 103.900 170.590 104.220 170.650 ;
        RECT 104.375 170.605 104.665 170.650 ;
        RECT 104.835 170.605 105.125 170.650 ;
        RECT 105.755 170.605 106.045 170.835 ;
        RECT 108.975 170.605 109.265 170.835 ;
        RECT 109.665 170.790 109.955 170.835 ;
        RECT 109.665 170.650 112.410 170.790 ;
        RECT 109.665 170.605 109.955 170.650 ;
        RECT 91.035 170.310 94.010 170.450 ;
        RECT 96.095 170.450 96.385 170.495 ;
        RECT 98.380 170.450 98.700 170.510 ;
        RECT 96.095 170.310 98.700 170.450 ;
        RECT 91.035 170.265 91.325 170.310 ;
        RECT 96.095 170.265 96.385 170.310 ;
        RECT 72.660 170.110 72.950 170.155 ;
        RECT 74.760 170.110 75.050 170.155 ;
        RECT 76.330 170.110 76.620 170.155 ;
        RECT 72.660 169.970 76.620 170.110 ;
        RECT 72.660 169.925 72.950 169.970 ;
        RECT 74.760 169.925 75.050 169.970 ;
        RECT 76.330 169.925 76.620 169.970 ;
        RECT 80.020 170.110 80.310 170.155 ;
        RECT 82.120 170.110 82.410 170.155 ;
        RECT 83.690 170.110 83.980 170.155 ;
        RECT 80.020 169.970 83.980 170.110 ;
        RECT 80.020 169.925 80.310 169.970 ;
        RECT 82.120 169.925 82.410 169.970 ;
        RECT 83.690 169.925 83.980 169.970 ;
        RECT 86.435 170.110 86.725 170.155 ;
        RECT 89.180 170.110 89.500 170.170 ;
        RECT 91.110 170.110 91.250 170.265 ;
        RECT 98.380 170.250 98.700 170.310 ;
        RECT 99.300 170.450 99.620 170.510 ;
        RECT 100.695 170.450 100.985 170.495 ;
        RECT 105.295 170.450 105.585 170.495 ;
        RECT 99.300 170.310 105.585 170.450 ;
        RECT 99.300 170.250 99.620 170.310 ;
        RECT 100.695 170.265 100.985 170.310 ;
        RECT 105.295 170.265 105.585 170.310 ;
        RECT 108.500 170.250 108.820 170.510 ;
        RECT 110.355 170.265 110.645 170.495 ;
        RECT 86.435 169.970 91.250 170.110 ;
        RECT 93.780 170.110 94.100 170.170 ;
        RECT 98.855 170.110 99.145 170.155 ;
        RECT 110.430 170.110 110.570 170.265 ;
        RECT 110.800 170.250 111.120 170.510 ;
        RECT 93.780 169.970 98.150 170.110 ;
        RECT 86.435 169.925 86.725 169.970 ;
        RECT 89.180 169.910 89.500 169.970 ;
        RECT 93.780 169.910 94.100 169.970 ;
        RECT 79.075 169.770 79.365 169.815 ;
        RECT 81.360 169.770 81.680 169.830 ;
        RECT 79.075 169.630 81.680 169.770 ;
        RECT 79.075 169.585 79.365 169.630 ;
        RECT 81.360 169.570 81.680 169.630 ;
        RECT 88.720 169.770 89.040 169.830 ;
        RECT 90.575 169.770 90.865 169.815 ;
        RECT 91.940 169.770 92.260 169.830 ;
        RECT 98.010 169.815 98.150 169.970 ;
        RECT 98.855 169.970 110.570 170.110 ;
        RECT 112.270 170.110 112.410 170.650 ;
        RECT 112.655 170.605 112.945 170.835 ;
        RECT 114.020 170.590 114.340 170.850 ;
        RECT 115.415 170.790 115.705 170.835 ;
        RECT 115.950 170.790 116.090 170.990 ;
        RECT 119.630 170.990 121.225 171.130 ;
        RECT 119.630 170.850 119.770 170.990 ;
        RECT 120.935 170.945 121.225 170.990 ;
        RECT 121.840 171.130 122.160 171.190 ;
        RECT 124.000 171.130 124.290 171.175 ;
        RECT 121.840 170.990 124.290 171.130 ;
        RECT 121.840 170.930 122.160 170.990 ;
        RECT 124.000 170.945 124.290 170.990 ;
        RECT 125.980 171.130 126.300 171.190 ;
        RECT 129.980 171.130 130.120 171.270 ;
        RECT 149.990 171.130 150.130 171.330 ;
        RECT 151.295 171.330 156.200 171.470 ;
        RECT 151.295 171.285 151.585 171.330 ;
        RECT 155.880 171.270 156.200 171.330 ;
        RECT 152.215 171.130 152.505 171.175 ;
        RECT 125.980 170.990 128.510 171.130 ;
        RECT 129.980 170.990 149.670 171.130 ;
        RECT 149.990 170.990 152.505 171.130 ;
        RECT 125.980 170.930 126.300 170.990 ;
        RECT 116.335 170.790 116.625 170.835 ;
        RECT 115.415 170.650 116.625 170.790 ;
        RECT 115.415 170.605 115.705 170.650 ;
        RECT 116.335 170.605 116.625 170.650 ;
        RECT 116.780 170.590 117.100 170.850 ;
        RECT 117.700 170.790 118.020 170.850 ;
        RECT 118.175 170.790 118.465 170.835 ;
        RECT 117.700 170.650 118.465 170.790 ;
        RECT 117.700 170.590 118.020 170.650 ;
        RECT 118.175 170.605 118.465 170.650 ;
        RECT 119.540 170.590 119.860 170.850 ;
        RECT 120.000 170.790 120.320 170.850 ;
        RECT 120.475 170.790 120.765 170.835 ;
        RECT 120.000 170.650 120.765 170.790 ;
        RECT 120.000 170.590 120.320 170.650 ;
        RECT 120.475 170.605 120.765 170.650 ;
        RECT 121.380 170.590 121.700 170.850 ;
        RECT 122.760 170.590 123.080 170.850 ;
        RECT 128.370 170.790 128.510 170.990 ;
        RECT 132.510 170.835 132.650 170.990 ;
        RECT 131.055 170.790 131.345 170.835 ;
        RECT 123.310 170.650 128.050 170.790 ;
        RECT 128.370 170.650 131.345 170.790 ;
        RECT 113.560 170.250 113.880 170.510 ;
        RECT 114.110 170.450 114.250 170.590 ;
        RECT 123.310 170.450 123.450 170.650 ;
        RECT 114.110 170.310 123.450 170.450 ;
        RECT 123.655 170.450 123.945 170.495 ;
        RECT 124.845 170.450 125.135 170.495 ;
        RECT 127.365 170.450 127.655 170.495 ;
        RECT 123.655 170.310 127.655 170.450 ;
        RECT 127.910 170.450 128.050 170.650 ;
        RECT 131.055 170.605 131.345 170.650 ;
        RECT 132.435 170.605 132.725 170.835 ;
        RECT 135.195 170.605 135.485 170.835 ;
        RECT 135.640 170.790 135.960 170.850 ;
        RECT 138.875 170.790 139.165 170.835 ;
        RECT 135.640 170.650 139.165 170.790 ;
        RECT 135.270 170.450 135.410 170.605 ;
        RECT 135.640 170.590 135.960 170.650 ;
        RECT 138.875 170.605 139.165 170.650 ;
        RECT 140.240 170.790 140.560 170.850 ;
        RECT 144.380 170.790 144.700 170.850 ;
        RECT 144.930 170.835 145.070 170.990 ;
        RECT 140.240 170.650 144.700 170.790 ;
        RECT 140.240 170.590 140.560 170.650 ;
        RECT 144.380 170.590 144.700 170.650 ;
        RECT 144.855 170.605 145.145 170.835 ;
        RECT 146.235 170.790 146.525 170.835 ;
        RECT 146.680 170.790 147.000 170.850 ;
        RECT 149.530 170.835 149.670 170.990 ;
        RECT 152.215 170.945 152.505 170.990 ;
        RECT 146.235 170.650 147.000 170.790 ;
        RECT 146.235 170.605 146.525 170.650 ;
        RECT 146.680 170.590 147.000 170.650 ;
        RECT 147.155 170.605 147.445 170.835 ;
        RECT 147.615 170.790 147.905 170.835 ;
        RECT 147.615 170.650 148.290 170.790 ;
        RECT 147.615 170.605 147.905 170.650 ;
        RECT 137.480 170.450 137.800 170.510 ;
        RECT 127.910 170.310 137.800 170.450 ;
        RECT 123.655 170.265 123.945 170.310 ;
        RECT 124.845 170.265 125.135 170.310 ;
        RECT 127.365 170.265 127.655 170.310 ;
        RECT 137.480 170.250 137.800 170.310 ;
        RECT 137.955 170.450 138.245 170.495 ;
        RECT 141.620 170.450 141.940 170.510 ;
        RECT 143.460 170.450 143.780 170.510 ;
        RECT 147.230 170.450 147.370 170.605 ;
        RECT 148.150 170.510 148.290 170.650 ;
        RECT 149.455 170.605 149.745 170.835 ;
        RECT 151.740 170.590 152.060 170.850 ;
        RECT 152.675 170.605 152.965 170.835 ;
        RECT 137.955 170.310 143.780 170.450 ;
        RECT 137.955 170.265 138.245 170.310 ;
        RECT 141.620 170.250 141.940 170.310 ;
        RECT 143.460 170.250 143.780 170.310 ;
        RECT 144.470 170.310 147.370 170.450 ;
        RECT 148.060 170.450 148.380 170.510 ;
        RECT 148.995 170.450 149.285 170.495 ;
        RECT 148.060 170.310 149.285 170.450 ;
        RECT 152.750 170.450 152.890 170.605 ;
        RECT 153.120 170.590 153.440 170.850 ;
        RECT 152.750 170.310 153.810 170.450 ;
        RECT 123.260 170.110 123.550 170.155 ;
        RECT 125.360 170.110 125.650 170.155 ;
        RECT 126.930 170.110 127.220 170.155 ;
        RECT 129.660 170.110 129.980 170.170 ;
        RECT 144.470 170.155 144.610 170.310 ;
        RECT 148.060 170.250 148.380 170.310 ;
        RECT 148.995 170.265 149.285 170.310 ;
        RECT 144.395 170.110 144.685 170.155 ;
        RECT 112.270 169.970 122.990 170.110 ;
        RECT 98.855 169.925 99.145 169.970 ;
        RECT 88.720 169.630 92.260 169.770 ;
        RECT 88.720 169.570 89.040 169.630 ;
        RECT 90.575 169.585 90.865 169.630 ;
        RECT 91.940 169.570 92.260 169.630 ;
        RECT 97.935 169.585 98.225 169.815 ;
        RECT 101.615 169.770 101.905 169.815 ;
        RECT 103.440 169.770 103.760 169.830 ;
        RECT 101.615 169.630 103.760 169.770 ;
        RECT 101.615 169.585 101.905 169.630 ;
        RECT 103.440 169.570 103.760 169.630 ;
        RECT 107.580 169.770 107.900 169.830 ;
        RECT 111.735 169.770 112.025 169.815 ;
        RECT 107.580 169.630 112.025 169.770 ;
        RECT 112.270 169.770 112.410 169.970 ;
        RECT 112.655 169.770 112.945 169.815 ;
        RECT 112.270 169.630 112.945 169.770 ;
        RECT 107.580 169.570 107.900 169.630 ;
        RECT 111.735 169.585 112.025 169.630 ;
        RECT 112.655 169.585 112.945 169.630 ;
        RECT 116.320 169.770 116.640 169.830 ;
        RECT 117.700 169.770 118.020 169.830 ;
        RECT 116.320 169.630 118.020 169.770 ;
        RECT 116.320 169.570 116.640 169.630 ;
        RECT 117.700 169.570 118.020 169.630 ;
        RECT 118.160 169.570 118.480 169.830 ;
        RECT 120.000 169.770 120.320 169.830 ;
        RECT 121.840 169.770 122.160 169.830 ;
        RECT 120.000 169.630 122.160 169.770 ;
        RECT 122.850 169.770 122.990 169.970 ;
        RECT 123.260 169.970 127.220 170.110 ;
        RECT 123.260 169.925 123.550 169.970 ;
        RECT 125.360 169.925 125.650 169.970 ;
        RECT 126.930 169.925 127.220 169.970 ;
        RECT 127.450 169.970 144.685 170.110 ;
        RECT 127.450 169.770 127.590 169.970 ;
        RECT 129.660 169.910 129.980 169.970 ;
        RECT 144.395 169.925 144.685 169.970 ;
        RECT 153.670 169.830 153.810 170.310 ;
        RECT 122.850 169.630 127.590 169.770 ;
        RECT 120.000 169.570 120.320 169.630 ;
        RECT 121.840 169.570 122.160 169.630 ;
        RECT 130.120 169.570 130.440 169.830 ;
        RECT 145.300 169.570 145.620 169.830 ;
        RECT 153.580 169.570 153.900 169.830 ;
        RECT 70.710 168.950 156.270 169.430 ;
        RECT 88.720 168.550 89.040 168.810 ;
        RECT 89.195 168.750 89.485 168.795 ;
        RECT 94.240 168.750 94.560 168.810 ;
        RECT 89.195 168.610 94.560 168.750 ;
        RECT 89.195 168.565 89.485 168.610 ;
        RECT 94.240 168.550 94.560 168.610 ;
        RECT 97.000 168.750 97.320 168.810 ;
        RECT 116.780 168.750 117.100 168.810 ;
        RECT 125.980 168.750 126.300 168.810 ;
        RECT 127.375 168.750 127.665 168.795 ;
        RECT 97.000 168.610 127.665 168.750 ;
        RECT 97.000 168.550 97.320 168.610 ;
        RECT 116.780 168.550 117.100 168.610 ;
        RECT 125.980 168.550 126.300 168.610 ;
        RECT 127.375 168.565 127.665 168.610 ;
        RECT 129.660 168.750 129.980 168.810 ;
        RECT 130.135 168.750 130.425 168.795 ;
        RECT 129.660 168.610 130.425 168.750 ;
        RECT 129.660 168.550 129.980 168.610 ;
        RECT 130.135 168.565 130.425 168.610 ;
        RECT 133.815 168.565 134.105 168.795 ;
        RECT 137.480 168.750 137.800 168.810 ;
        RECT 137.480 168.610 155.190 168.750 ;
        RECT 72.660 168.410 72.950 168.455 ;
        RECT 74.760 168.410 75.050 168.455 ;
        RECT 76.330 168.410 76.620 168.455 ;
        RECT 80.455 168.410 80.745 168.455 ;
        RECT 87.340 168.410 87.660 168.470 ;
        RECT 72.660 168.270 76.620 168.410 ;
        RECT 72.660 168.225 72.950 168.270 ;
        RECT 74.760 168.225 75.050 168.270 ;
        RECT 76.330 168.225 76.620 168.270 ;
        RECT 77.770 168.270 87.660 168.410 ;
        RECT 77.770 168.130 77.910 168.270 ;
        RECT 80.455 168.225 80.745 168.270 ;
        RECT 87.340 168.210 87.660 168.270 ;
        RECT 87.815 168.410 88.105 168.455 ;
        RECT 88.810 168.410 88.950 168.550 ;
        RECT 87.815 168.270 88.950 168.410 ;
        RECT 96.540 168.410 96.860 168.470 ;
        RECT 101.140 168.410 101.460 168.470 ;
        RECT 96.540 168.270 101.460 168.410 ;
        RECT 87.815 168.225 88.105 168.270 ;
        RECT 96.540 168.210 96.860 168.270 ;
        RECT 101.140 168.210 101.460 168.270 ;
        RECT 102.060 168.410 102.380 168.470 ;
        RECT 103.900 168.410 104.220 168.470 ;
        RECT 102.060 168.270 104.220 168.410 ;
        RECT 102.060 168.210 102.380 168.270 ;
        RECT 103.900 168.210 104.220 168.270 ;
        RECT 113.560 168.410 113.880 168.470 ;
        RECT 119.080 168.410 119.400 168.470 ;
        RECT 113.560 168.270 119.400 168.410 ;
        RECT 113.560 168.210 113.880 168.270 ;
        RECT 119.080 168.210 119.400 168.270 ;
        RECT 120.000 168.210 120.320 168.470 ;
        RECT 120.960 168.410 121.250 168.455 ;
        RECT 123.060 168.410 123.350 168.455 ;
        RECT 124.630 168.410 124.920 168.455 ;
        RECT 133.890 168.410 134.030 168.565 ;
        RECT 137.480 168.550 137.800 168.610 ;
        RECT 120.960 168.270 124.920 168.410 ;
        RECT 120.960 168.225 121.250 168.270 ;
        RECT 123.060 168.225 123.350 168.270 ;
        RECT 124.630 168.225 124.920 168.270 ;
        RECT 133.460 168.270 134.030 168.410 ;
        RECT 73.055 168.070 73.345 168.115 ;
        RECT 74.245 168.070 74.535 168.115 ;
        RECT 76.765 168.070 77.055 168.115 ;
        RECT 73.055 167.930 77.055 168.070 ;
        RECT 73.055 167.885 73.345 167.930 ;
        RECT 74.245 167.885 74.535 167.930 ;
        RECT 76.765 167.885 77.055 167.930 ;
        RECT 77.680 167.870 78.000 168.130 ;
        RECT 79.060 168.070 79.380 168.130 ;
        RECT 81.375 168.070 81.665 168.115 ;
        RECT 85.500 168.070 85.820 168.130 ;
        RECT 93.780 168.070 94.100 168.130 ;
        RECT 102.535 168.070 102.825 168.115 ;
        RECT 79.060 167.930 85.820 168.070 ;
        RECT 79.060 167.870 79.380 167.930 ;
        RECT 81.375 167.885 81.665 167.930 ;
        RECT 85.500 167.870 85.820 167.930 ;
        RECT 86.970 167.930 94.100 168.070 ;
        RECT 86.970 167.790 87.110 167.930 ;
        RECT 93.780 167.870 94.100 167.930 ;
        RECT 99.850 167.930 102.825 168.070 ;
        RECT 99.850 167.790 99.990 167.930 ;
        RECT 102.535 167.885 102.825 167.930 ;
        RECT 114.480 168.070 114.800 168.130 ;
        RECT 117.700 168.070 118.020 168.130 ;
        RECT 121.355 168.070 121.645 168.115 ;
        RECT 122.545 168.070 122.835 168.115 ;
        RECT 125.065 168.070 125.355 168.115 ;
        RECT 133.460 168.070 133.600 168.270 ;
        RECT 139.320 168.210 139.640 168.470 ;
        RECT 142.580 168.410 142.870 168.455 ;
        RECT 144.680 168.410 144.970 168.455 ;
        RECT 146.250 168.410 146.540 168.455 ;
        RECT 142.580 168.270 146.540 168.410 ;
        RECT 142.580 168.225 142.870 168.270 ;
        RECT 144.680 168.225 144.970 168.270 ;
        RECT 146.250 168.225 146.540 168.270 ;
        RECT 148.995 168.410 149.285 168.455 ;
        RECT 153.120 168.410 153.440 168.470 ;
        RECT 148.995 168.270 153.440 168.410 ;
        RECT 148.995 168.225 149.285 168.270 ;
        RECT 153.120 168.210 153.440 168.270 ;
        RECT 114.480 167.930 118.390 168.070 ;
        RECT 114.480 167.870 114.800 167.930 ;
        RECT 117.700 167.870 118.020 167.930 ;
        RECT 72.160 167.530 72.480 167.790 ;
        RECT 79.535 167.730 79.825 167.775 ;
        RECT 80.915 167.730 81.205 167.775 ;
        RECT 79.535 167.590 81.205 167.730 ;
        RECT 79.535 167.545 79.825 167.590 ;
        RECT 80.915 167.545 81.205 167.590 ;
        RECT 73.510 167.390 73.800 167.435 ;
        RECT 77.220 167.390 77.540 167.450 ;
        RECT 73.510 167.250 77.540 167.390 ;
        RECT 73.510 167.205 73.800 167.250 ;
        RECT 77.220 167.190 77.540 167.250 ;
        RECT 79.075 167.050 79.365 167.095 ;
        RECT 80.990 167.050 81.130 167.545 ;
        RECT 86.880 167.530 87.200 167.790 ;
        RECT 88.260 167.530 88.580 167.790 ;
        RECT 88.720 167.730 89.040 167.790 ;
        RECT 89.195 167.730 89.485 167.775 ;
        RECT 88.720 167.590 89.485 167.730 ;
        RECT 88.720 167.530 89.040 167.590 ;
        RECT 89.195 167.545 89.485 167.590 ;
        RECT 90.560 167.730 90.880 167.790 ;
        RECT 94.240 167.730 94.560 167.790 ;
        RECT 90.560 167.590 94.560 167.730 ;
        RECT 90.560 167.530 90.880 167.590 ;
        RECT 87.340 167.390 87.660 167.450 ;
        RECT 91.020 167.390 91.340 167.450 ;
        RECT 87.340 167.250 91.340 167.390 ;
        RECT 87.340 167.190 87.660 167.250 ;
        RECT 91.020 167.190 91.340 167.250 ;
        RECT 91.570 167.050 91.710 167.590 ;
        RECT 94.240 167.530 94.560 167.590 ;
        RECT 98.840 167.530 99.160 167.790 ;
        RECT 99.760 167.530 100.080 167.790 ;
        RECT 100.220 167.530 100.540 167.790 ;
        RECT 101.140 167.730 101.460 167.790 ;
        RECT 113.100 167.730 113.420 167.790 ;
        RECT 113.575 167.730 113.865 167.775 ;
        RECT 101.140 167.590 113.865 167.730 ;
        RECT 101.140 167.530 101.460 167.590 ;
        RECT 113.100 167.530 113.420 167.590 ;
        RECT 113.575 167.545 113.865 167.590 ;
        RECT 116.780 167.530 117.100 167.790 ;
        RECT 118.250 167.775 118.390 167.930 ;
        RECT 121.355 167.930 125.355 168.070 ;
        RECT 121.355 167.885 121.645 167.930 ;
        RECT 122.545 167.885 122.835 167.930 ;
        RECT 125.065 167.885 125.355 167.930 ;
        RECT 129.750 167.930 133.600 168.070 ;
        RECT 134.260 168.070 134.580 168.130 ;
        RECT 139.410 168.070 139.550 168.210 ;
        RECT 155.050 168.130 155.190 168.610 ;
        RECT 134.260 167.930 135.870 168.070 ;
        RECT 118.175 167.545 118.465 167.775 ;
        RECT 118.620 167.530 118.940 167.790 ;
        RECT 119.095 167.730 119.385 167.775 ;
        RECT 119.540 167.730 119.860 167.790 ;
        RECT 119.095 167.590 119.860 167.730 ;
        RECT 119.095 167.545 119.385 167.590 ;
        RECT 119.540 167.530 119.860 167.590 ;
        RECT 120.475 167.730 120.765 167.775 ;
        RECT 123.220 167.730 123.540 167.790 ;
        RECT 120.475 167.590 123.540 167.730 ;
        RECT 120.475 167.545 120.765 167.590 ;
        RECT 123.220 167.530 123.540 167.590 ;
        RECT 126.440 167.730 126.760 167.790 ;
        RECT 129.200 167.730 129.520 167.790 ;
        RECT 129.750 167.775 129.890 167.930 ;
        RECT 134.260 167.870 134.580 167.930 ;
        RECT 126.440 167.590 129.520 167.730 ;
        RECT 126.440 167.530 126.760 167.590 ;
        RECT 129.200 167.530 129.520 167.590 ;
        RECT 129.675 167.545 129.965 167.775 ;
        RECT 131.960 167.730 132.280 167.790 ;
        RECT 135.730 167.775 135.870 167.930 ;
        RECT 138.490 167.930 139.550 168.070 ;
        RECT 142.975 168.070 143.265 168.115 ;
        RECT 144.165 168.070 144.455 168.115 ;
        RECT 146.685 168.070 146.975 168.115 ;
        RECT 151.755 168.070 152.045 168.115 ;
        RECT 142.975 167.930 146.975 168.070 ;
        RECT 138.490 167.775 138.630 167.930 ;
        RECT 142.975 167.885 143.265 167.930 ;
        RECT 144.165 167.885 144.455 167.930 ;
        RECT 146.685 167.885 146.975 167.930 ;
        RECT 149.070 167.930 152.045 168.070 ;
        RECT 149.070 167.790 149.210 167.930 ;
        RECT 151.755 167.885 152.045 167.930 ;
        RECT 154.960 167.870 155.280 168.130 ;
        RECT 134.735 167.730 135.025 167.775 ;
        RECT 101.600 167.435 101.920 167.450 ;
        RECT 100.695 167.390 100.985 167.435 ;
        RECT 98.930 167.250 100.985 167.390 ;
        RECT 98.930 167.110 99.070 167.250 ;
        RECT 100.695 167.205 100.985 167.250 ;
        RECT 101.600 167.205 102.035 167.435 ;
        RECT 117.585 167.390 117.875 167.435 ;
        RECT 102.610 167.250 119.310 167.390 ;
        RECT 101.600 167.190 101.920 167.205 ;
        RECT 102.610 167.110 102.750 167.250 ;
        RECT 117.585 167.205 117.875 167.250 ;
        RECT 119.170 167.110 119.310 167.250 ;
        RECT 121.755 167.205 122.045 167.435 ;
        RECT 79.075 166.910 91.710 167.050 ;
        RECT 79.075 166.865 79.365 166.910 ;
        RECT 92.400 166.850 92.720 167.110 ;
        RECT 98.840 166.850 99.160 167.110 ;
        RECT 99.300 166.850 99.620 167.110 ;
        RECT 101.140 167.050 101.460 167.110 ;
        RECT 102.520 167.050 102.840 167.110 ;
        RECT 101.140 166.910 102.840 167.050 ;
        RECT 101.140 166.850 101.460 166.910 ;
        RECT 102.520 166.850 102.840 166.910 ;
        RECT 104.360 167.050 104.680 167.110 ;
        RECT 114.480 167.050 114.800 167.110 ;
        RECT 104.360 166.910 114.800 167.050 ;
        RECT 104.360 166.850 104.680 166.910 ;
        RECT 114.480 166.850 114.800 166.910 ;
        RECT 119.080 166.850 119.400 167.110 ;
        RECT 121.885 167.050 122.025 167.205 ;
        RECT 129.750 167.110 129.890 167.545 ;
        RECT 131.055 167.450 131.345 167.655 ;
        RECT 131.960 167.590 135.025 167.730 ;
        RECT 131.960 167.530 132.280 167.590 ;
        RECT 134.735 167.545 135.025 167.590 ;
        RECT 135.655 167.545 135.945 167.775 ;
        RECT 138.415 167.545 138.705 167.775 ;
        RECT 139.320 167.530 139.640 167.790 ;
        RECT 139.780 167.530 140.100 167.790 ;
        RECT 140.240 167.530 140.560 167.790 ;
        RECT 142.095 167.730 142.385 167.775 ;
        RECT 142.540 167.730 142.860 167.790 ;
        RECT 142.095 167.590 142.860 167.730 ;
        RECT 142.095 167.545 142.385 167.590 ;
        RECT 142.540 167.530 142.860 167.590 ;
        RECT 148.980 167.530 149.300 167.790 ;
        RECT 150.375 167.545 150.665 167.775 ;
        RECT 130.595 167.205 130.885 167.435 ;
        RECT 123.220 167.050 123.540 167.110 ;
        RECT 121.885 166.910 123.540 167.050 ;
        RECT 123.220 166.850 123.540 166.910 ;
        RECT 123.680 167.050 124.000 167.110 ;
        RECT 128.295 167.050 128.585 167.095 ;
        RECT 123.680 166.910 128.585 167.050 ;
        RECT 123.680 166.850 124.000 166.910 ;
        RECT 128.295 166.865 128.585 166.910 ;
        RECT 129.660 166.850 129.980 167.110 ;
        RECT 130.120 167.050 130.440 167.110 ;
        RECT 130.670 167.050 130.810 167.205 ;
        RECT 131.040 167.190 131.360 167.450 ;
        RECT 136.575 167.390 136.865 167.435 ;
        RECT 132.050 167.250 136.865 167.390 ;
        RECT 132.050 167.110 132.190 167.250 ;
        RECT 136.575 167.205 136.865 167.250 ;
        RECT 141.635 167.390 141.925 167.435 ;
        RECT 143.320 167.390 143.610 167.435 ;
        RECT 141.635 167.250 143.610 167.390 ;
        RECT 150.450 167.390 150.590 167.545 ;
        RECT 150.450 167.250 152.430 167.390 ;
        RECT 141.635 167.205 141.925 167.250 ;
        RECT 143.320 167.205 143.610 167.250 ;
        RECT 152.290 167.110 152.430 167.250 ;
        RECT 130.120 166.910 130.810 167.050 ;
        RECT 130.120 166.850 130.440 166.910 ;
        RECT 131.960 166.850 132.280 167.110 ;
        RECT 137.495 167.050 137.785 167.095 ;
        RECT 137.940 167.050 138.260 167.110 ;
        RECT 137.495 166.910 138.260 167.050 ;
        RECT 137.495 166.865 137.785 166.910 ;
        RECT 137.940 166.850 138.260 166.910 ;
        RECT 139.780 167.050 140.100 167.110 ;
        RECT 140.700 167.050 141.020 167.110 ;
        RECT 139.780 166.910 141.020 167.050 ;
        RECT 139.780 166.850 140.100 166.910 ;
        RECT 140.700 166.850 141.020 166.910 ;
        RECT 152.200 166.850 152.520 167.110 ;
        RECT 70.710 166.230 156.270 166.710 ;
        RECT 83.675 166.030 83.965 166.075 ;
        RECT 88.720 166.030 89.040 166.090 ;
        RECT 83.675 165.890 89.040 166.030 ;
        RECT 83.675 165.845 83.965 165.890 ;
        RECT 88.720 165.830 89.040 165.890 ;
        RECT 92.400 165.830 92.720 166.090 ;
        RECT 98.840 165.830 99.160 166.090 ;
        RECT 100.220 166.030 100.540 166.090 ;
        RECT 105.295 166.030 105.585 166.075 ;
        RECT 100.220 165.890 105.585 166.030 ;
        RECT 100.220 165.830 100.540 165.890 ;
        RECT 105.295 165.845 105.585 165.890 ;
        RECT 117.700 165.830 118.020 166.090 ;
        RECT 118.620 166.030 118.940 166.090 ;
        RECT 121.395 166.030 121.685 166.075 ;
        RECT 123.220 166.030 123.540 166.090 ;
        RECT 118.620 165.890 121.150 166.030 ;
        RECT 118.620 165.830 118.940 165.890 ;
        RECT 76.850 165.550 91.250 165.690 ;
        RECT 72.160 165.350 72.480 165.410 ;
        RECT 76.850 165.395 76.990 165.550 ;
        RECT 76.775 165.350 77.065 165.395 ;
        RECT 72.160 165.210 77.065 165.350 ;
        RECT 72.160 165.150 72.480 165.210 ;
        RECT 76.775 165.165 77.065 165.210 ;
        RECT 78.110 165.350 78.400 165.395 ;
        RECT 80.900 165.350 81.220 165.410 ;
        RECT 86.880 165.350 87.200 165.410 ;
        RECT 91.110 165.395 91.250 165.550 ;
        RECT 78.110 165.210 81.220 165.350 ;
        RECT 78.110 165.165 78.400 165.210 ;
        RECT 80.900 165.150 81.220 165.210 ;
        RECT 86.050 165.210 87.200 165.350 ;
        RECT 77.655 165.010 77.945 165.055 ;
        RECT 78.845 165.010 79.135 165.055 ;
        RECT 81.365 165.010 81.655 165.055 ;
        RECT 77.655 164.870 81.655 165.010 ;
        RECT 77.655 164.825 77.945 164.870 ;
        RECT 78.845 164.825 79.135 164.870 ;
        RECT 81.365 164.825 81.655 164.870 ;
        RECT 77.260 164.670 77.550 164.715 ;
        RECT 79.360 164.670 79.650 164.715 ;
        RECT 80.930 164.670 81.220 164.715 ;
        RECT 77.260 164.530 81.220 164.670 ;
        RECT 77.260 164.485 77.550 164.530 ;
        RECT 79.360 164.485 79.650 164.530 ;
        RECT 80.930 164.485 81.220 164.530 ;
        RECT 84.135 164.670 84.425 164.715 ;
        RECT 86.050 164.670 86.190 165.210 ;
        RECT 86.880 165.150 87.200 165.210 ;
        RECT 89.755 165.350 90.045 165.395 ;
        RECT 91.035 165.350 91.325 165.395 ;
        RECT 92.490 165.350 92.630 165.830 ;
        RECT 102.995 165.690 103.285 165.735 ;
        RECT 104.360 165.690 104.680 165.750 ;
        RECT 98.470 165.550 102.290 165.690 ;
        RECT 89.755 165.210 90.790 165.350 ;
        RECT 89.755 165.165 90.045 165.210 ;
        RECT 86.445 165.010 86.735 165.055 ;
        RECT 88.965 165.010 89.255 165.055 ;
        RECT 90.155 165.010 90.445 165.055 ;
        RECT 86.445 164.870 90.445 165.010 ;
        RECT 90.650 165.010 90.790 165.210 ;
        RECT 91.035 165.210 92.630 165.350 ;
        RECT 95.620 165.350 95.940 165.410 ;
        RECT 98.470 165.395 98.610 165.550 ;
        RECT 102.150 165.410 102.290 165.550 ;
        RECT 102.995 165.550 104.680 165.690 ;
        RECT 102.995 165.505 103.285 165.550 ;
        RECT 104.360 165.490 104.680 165.550 ;
        RECT 112.640 165.490 112.960 165.750 ;
        RECT 113.560 165.690 113.880 165.750 ;
        RECT 117.790 165.690 117.930 165.830 ;
        RECT 121.010 165.690 121.150 165.890 ;
        RECT 121.395 165.890 123.540 166.030 ;
        RECT 121.395 165.845 121.685 165.890 ;
        RECT 123.220 165.830 123.540 165.890 ;
        RECT 137.020 166.030 137.340 166.090 ;
        RECT 139.320 166.030 139.640 166.090 ;
        RECT 143.475 166.030 143.765 166.075 ;
        RECT 137.020 165.890 139.090 166.030 ;
        RECT 137.020 165.830 137.340 165.890 ;
        RECT 122.775 165.690 123.065 165.735 ;
        RECT 123.750 165.690 124.040 165.735 ;
        RECT 113.560 165.550 116.090 165.690 ;
        RECT 117.790 165.550 119.310 165.690 ;
        RECT 121.010 165.550 123.065 165.690 ;
        RECT 113.560 165.490 113.880 165.550 ;
        RECT 97.475 165.350 97.765 165.395 ;
        RECT 95.620 165.210 97.765 165.350 ;
        RECT 91.035 165.165 91.325 165.210 ;
        RECT 95.620 165.150 95.940 165.210 ;
        RECT 97.475 165.165 97.765 165.210 ;
        RECT 98.395 165.165 98.685 165.395 ;
        RECT 91.495 165.010 91.785 165.055 ;
        RECT 91.940 165.010 92.260 165.070 ;
        RECT 90.650 164.870 91.250 165.010 ;
        RECT 86.445 164.825 86.735 164.870 ;
        RECT 88.965 164.825 89.255 164.870 ;
        RECT 90.155 164.825 90.445 164.870 ;
        RECT 84.135 164.530 86.190 164.670 ;
        RECT 86.880 164.670 87.170 164.715 ;
        RECT 88.450 164.670 88.740 164.715 ;
        RECT 90.550 164.670 90.840 164.715 ;
        RECT 86.880 164.530 90.840 164.670 ;
        RECT 91.110 164.670 91.250 164.870 ;
        RECT 91.495 164.870 92.260 165.010 ;
        RECT 91.495 164.825 91.785 164.870 ;
        RECT 91.940 164.810 92.260 164.870 ;
        RECT 92.875 165.010 93.165 165.055 ;
        RECT 93.780 165.010 94.100 165.070 ;
        RECT 92.875 164.870 94.100 165.010 ;
        RECT 97.550 165.010 97.690 165.165 ;
        RECT 99.760 165.150 100.080 165.410 ;
        RECT 100.695 165.350 100.985 165.395 ;
        RECT 101.600 165.350 101.920 165.410 ;
        RECT 100.695 165.210 101.920 165.350 ;
        RECT 100.695 165.165 100.985 165.210 ;
        RECT 101.600 165.150 101.920 165.210 ;
        RECT 102.060 165.150 102.380 165.410 ;
        RECT 102.520 165.150 102.840 165.410 ;
        RECT 103.585 165.350 103.875 165.395 ;
        RECT 103.070 165.210 103.875 165.350 ;
        RECT 101.140 165.010 101.460 165.070 ;
        RECT 103.070 165.010 103.210 165.210 ;
        RECT 103.585 165.165 103.875 165.210 ;
        RECT 104.835 165.165 105.125 165.395 ;
        RECT 107.120 165.350 107.440 165.410 ;
        RECT 108.055 165.350 108.345 165.395 ;
        RECT 107.120 165.210 108.345 165.350 ;
        RECT 97.550 164.870 99.990 165.010 ;
        RECT 92.875 164.825 93.165 164.870 ;
        RECT 93.780 164.810 94.100 164.870 ;
        RECT 99.300 164.670 99.620 164.730 ;
        RECT 91.110 164.530 99.620 164.670 ;
        RECT 99.850 164.670 99.990 164.870 ;
        RECT 101.140 164.870 103.210 165.010 ;
        RECT 101.140 164.810 101.460 164.870 ;
        RECT 104.360 164.810 104.680 165.070 ;
        RECT 103.440 164.670 103.760 164.730 ;
        RECT 104.910 164.670 105.050 165.165 ;
        RECT 107.120 165.150 107.440 165.210 ;
        RECT 108.055 165.165 108.345 165.210 ;
        RECT 114.035 165.165 114.325 165.395 ;
        RECT 109.435 165.010 109.725 165.055 ;
        RECT 114.110 165.010 114.250 165.165 ;
        RECT 114.480 165.150 114.800 165.410 ;
        RECT 115.950 165.395 116.090 165.550 ;
        RECT 114.955 165.165 115.245 165.395 ;
        RECT 115.875 165.350 116.165 165.395 ;
        RECT 115.875 165.210 117.930 165.350 ;
        RECT 115.875 165.165 116.165 165.210 ;
        RECT 115.030 165.010 115.170 165.165 ;
        RECT 116.780 165.010 117.100 165.070 ;
        RECT 109.435 164.870 110.570 165.010 ;
        RECT 114.110 164.870 114.710 165.010 ;
        RECT 115.030 164.870 117.100 165.010 ;
        RECT 117.790 165.010 117.930 165.210 ;
        RECT 118.160 165.340 118.480 165.410 ;
        RECT 118.735 165.350 119.025 165.395 ;
        RECT 118.710 165.340 119.025 165.350 ;
        RECT 118.160 165.200 119.025 165.340 ;
        RECT 119.170 165.350 119.310 165.550 ;
        RECT 122.775 165.505 123.065 165.550 ;
        RECT 123.430 165.550 124.040 165.690 ;
        RECT 119.555 165.350 119.845 165.395 ;
        RECT 119.170 165.210 119.845 165.350 ;
        RECT 118.160 165.150 118.480 165.200 ;
        RECT 118.735 165.165 119.025 165.200 ;
        RECT 119.555 165.165 119.845 165.210 ;
        RECT 120.000 165.150 120.320 165.410 ;
        RECT 120.460 165.150 120.780 165.410 ;
        RECT 121.840 165.350 122.160 165.410 ;
        RECT 123.430 165.350 123.570 165.550 ;
        RECT 123.750 165.505 124.040 165.550 ;
        RECT 124.600 165.690 124.920 165.750 ;
        RECT 125.835 165.690 126.125 165.735 ;
        RECT 124.600 165.550 126.125 165.690 ;
        RECT 124.600 165.490 124.920 165.550 ;
        RECT 125.835 165.505 126.125 165.550 ;
        RECT 126.440 165.690 126.760 165.750 ;
        RECT 126.915 165.690 127.205 165.735 ;
        RECT 130.120 165.690 130.440 165.750 ;
        RECT 126.440 165.550 127.205 165.690 ;
        RECT 126.440 165.490 126.760 165.550 ;
        RECT 126.915 165.505 127.205 165.550 ;
        RECT 129.750 165.550 130.440 165.690 ;
        RECT 128.280 165.350 128.600 165.410 ;
        RECT 129.750 165.395 129.890 165.550 ;
        RECT 130.120 165.490 130.440 165.550 ;
        RECT 133.800 165.690 134.120 165.750 ;
        RECT 137.480 165.690 137.800 165.750 ;
        RECT 133.800 165.550 138.630 165.690 ;
        RECT 121.840 165.210 123.570 165.350 ;
        RECT 124.075 165.270 128.600 165.350 ;
        RECT 123.770 165.210 128.600 165.270 ;
        RECT 121.840 165.150 122.160 165.210 ;
        RECT 123.770 165.130 124.215 165.210 ;
        RECT 128.280 165.150 128.600 165.210 ;
        RECT 129.675 165.165 129.965 165.395 ;
        RECT 130.595 165.350 130.885 165.395 ;
        RECT 131.500 165.350 131.820 165.410 ;
        RECT 130.595 165.210 131.820 165.350 ;
        RECT 131.960 165.350 132.280 165.530 ;
        RECT 133.800 165.490 134.120 165.550 ;
        RECT 137.480 165.490 137.800 165.550 ;
        RECT 132.435 165.350 132.725 165.395 ;
        RECT 137.020 165.350 137.340 165.410 ;
        RECT 138.490 165.395 138.630 165.550 ;
        RECT 131.960 165.270 137.340 165.350 ;
        RECT 132.050 165.210 137.340 165.270 ;
        RECT 130.595 165.165 130.885 165.210 ;
        RECT 123.770 165.010 123.910 165.130 ;
        RECT 130.670 165.010 130.810 165.165 ;
        RECT 131.500 165.150 131.820 165.210 ;
        RECT 132.435 165.165 132.725 165.210 ;
        RECT 137.020 165.150 137.340 165.210 ;
        RECT 138.415 165.165 138.705 165.395 ;
        RECT 138.950 165.350 139.090 165.890 ;
        RECT 139.320 165.890 143.765 166.030 ;
        RECT 139.320 165.830 139.640 165.890 ;
        RECT 143.475 165.845 143.765 165.890 ;
        RECT 147.155 166.030 147.445 166.075 ;
        RECT 151.740 166.030 152.060 166.090 ;
        RECT 147.155 165.890 152.060 166.030 ;
        RECT 147.155 165.845 147.445 165.890 ;
        RECT 151.740 165.830 152.060 165.890 ;
        RECT 153.120 165.830 153.440 166.090 ;
        RECT 140.700 165.350 141.020 165.410 ;
        RECT 141.635 165.350 141.925 165.395 ;
        RECT 143.895 165.350 144.185 165.395 ;
        RECT 138.950 165.210 141.925 165.350 ;
        RECT 140.700 165.150 141.020 165.210 ;
        RECT 141.635 165.165 141.925 165.210 ;
        RECT 143.550 165.210 144.185 165.350 ;
        RECT 117.790 164.870 123.910 165.010 ;
        RECT 124.690 164.870 130.810 165.010 ;
        RECT 131.960 165.010 132.280 165.070 ;
        RECT 133.815 165.010 134.105 165.055 ;
        RECT 131.960 164.870 134.105 165.010 ;
        RECT 109.435 164.825 109.725 164.870 ;
        RECT 110.430 164.730 110.570 164.870 ;
        RECT 99.850 164.530 101.830 164.670 ;
        RECT 84.135 164.485 84.425 164.530 ;
        RECT 86.880 164.485 87.170 164.530 ;
        RECT 88.450 164.485 88.740 164.530 ;
        RECT 90.550 164.485 90.840 164.530 ;
        RECT 99.300 164.470 99.620 164.530 ;
        RECT 98.380 164.130 98.700 164.390 ;
        RECT 100.220 164.330 100.540 164.390 ;
        RECT 101.155 164.330 101.445 164.375 ;
        RECT 100.220 164.190 101.445 164.330 ;
        RECT 101.690 164.330 101.830 164.530 ;
        RECT 103.440 164.530 105.050 164.670 ;
        RECT 103.440 164.470 103.760 164.530 ;
        RECT 110.340 164.470 110.660 164.730 ;
        RECT 114.570 164.670 114.710 164.870 ;
        RECT 116.780 164.810 117.100 164.870 ;
        RECT 124.690 164.670 124.830 164.870 ;
        RECT 131.960 164.810 132.280 164.870 ;
        RECT 133.815 164.825 134.105 164.870 ;
        RECT 114.570 164.530 124.830 164.670 ;
        RECT 129.200 164.670 129.520 164.730 ;
        RECT 130.595 164.670 130.885 164.715 ;
        RECT 140.240 164.670 140.560 164.730 ;
        RECT 142.555 164.670 142.845 164.715 ;
        RECT 129.200 164.530 140.010 164.670 ;
        RECT 114.570 164.330 114.710 164.530 ;
        RECT 129.200 164.470 129.520 164.530 ;
        RECT 130.595 164.485 130.885 164.530 ;
        RECT 101.690 164.190 114.710 164.330 ;
        RECT 116.320 164.330 116.640 164.390 ;
        RECT 125.075 164.330 125.365 164.375 ;
        RECT 116.320 164.190 125.365 164.330 ;
        RECT 100.220 164.130 100.540 164.190 ;
        RECT 101.155 164.145 101.445 164.190 ;
        RECT 116.320 164.130 116.640 164.190 ;
        RECT 125.075 164.145 125.365 164.190 ;
        RECT 125.995 164.330 126.285 164.375 ;
        RECT 131.040 164.330 131.360 164.390 ;
        RECT 125.995 164.190 131.360 164.330 ;
        RECT 139.870 164.330 140.010 164.530 ;
        RECT 140.240 164.530 142.845 164.670 ;
        RECT 140.240 164.470 140.560 164.530 ;
        RECT 142.555 164.485 142.845 164.530 ;
        RECT 143.550 164.330 143.690 165.210 ;
        RECT 143.895 165.165 144.185 165.210 ;
        RECT 146.680 165.150 147.000 165.410 ;
        RECT 147.615 165.350 147.905 165.395 ;
        RECT 152.200 165.350 152.520 165.410 ;
        RECT 153.210 165.395 153.350 165.830 ;
        RECT 147.615 165.210 152.520 165.350 ;
        RECT 147.615 165.165 147.905 165.210 ;
        RECT 152.200 165.150 152.520 165.210 ;
        RECT 153.135 165.165 153.425 165.395 ;
        RECT 146.770 165.010 146.910 165.150 ;
        RECT 148.060 165.010 148.380 165.070 ;
        RECT 151.295 165.010 151.585 165.055 ;
        RECT 146.770 164.870 151.585 165.010 ;
        RECT 148.060 164.810 148.380 164.870 ;
        RECT 151.295 164.825 151.585 164.870 ;
        RECT 152.675 165.010 152.965 165.055 ;
        RECT 153.580 165.010 153.900 165.070 ;
        RECT 152.675 164.870 153.900 165.010 ;
        RECT 152.675 164.825 152.965 164.870 ;
        RECT 153.580 164.810 153.900 164.870 ;
        RECT 143.920 164.330 144.240 164.390 ;
        RECT 139.870 164.190 144.240 164.330 ;
        RECT 125.995 164.145 126.285 164.190 ;
        RECT 131.040 164.130 131.360 164.190 ;
        RECT 143.920 164.130 144.240 164.190 ;
        RECT 153.580 164.330 153.900 164.390 ;
        RECT 154.055 164.330 154.345 164.375 ;
        RECT 154.960 164.330 155.280 164.390 ;
        RECT 153.580 164.190 155.280 164.330 ;
        RECT 153.580 164.130 153.900 164.190 ;
        RECT 154.055 164.145 154.345 164.190 ;
        RECT 154.960 164.130 155.280 164.190 ;
        RECT 70.710 163.510 156.270 163.990 ;
        RECT 72.175 163.310 72.465 163.355 ;
        RECT 83.660 163.310 83.980 163.370 ;
        RECT 72.175 163.170 83.980 163.310 ;
        RECT 72.175 163.125 72.465 163.170 ;
        RECT 83.660 163.110 83.980 163.170 ;
        RECT 91.495 163.310 91.785 163.355 ;
        RECT 92.415 163.310 92.705 163.355 ;
        RECT 91.495 163.170 92.705 163.310 ;
        RECT 91.495 163.125 91.785 163.170 ;
        RECT 92.415 163.125 92.705 163.170 ;
        RECT 95.620 163.110 95.940 163.370 ;
        RECT 96.540 163.110 96.860 163.370 ;
        RECT 98.380 163.310 98.700 163.370 ;
        RECT 99.315 163.310 99.605 163.355 ;
        RECT 98.380 163.170 99.605 163.310 ;
        RECT 98.380 163.110 98.700 163.170 ;
        RECT 99.315 163.125 99.605 163.170 ;
        RECT 102.060 163.110 102.380 163.370 ;
        RECT 102.520 163.310 102.840 163.370 ;
        RECT 106.215 163.310 106.505 163.355 ;
        RECT 102.520 163.170 106.505 163.310 ;
        RECT 102.520 163.110 102.840 163.170 ;
        RECT 106.215 163.125 106.505 163.170 ;
        RECT 107.120 163.110 107.440 163.370 ;
        RECT 114.480 163.310 114.800 163.370 ;
        RECT 115.415 163.310 115.705 163.355 ;
        RECT 114.480 163.170 115.705 163.310 ;
        RECT 114.480 163.110 114.800 163.170 ;
        RECT 115.415 163.125 115.705 163.170 ;
        RECT 116.780 163.110 117.100 163.370 ;
        RECT 129.660 163.310 129.980 163.370 ;
        RECT 133.800 163.310 134.120 163.370 ;
        RECT 129.660 163.170 134.120 163.310 ;
        RECT 129.660 163.110 129.980 163.170 ;
        RECT 133.800 163.110 134.120 163.170 ;
        RECT 152.200 163.310 152.520 163.370 ;
        RECT 154.515 163.310 154.805 163.355 ;
        RECT 152.200 163.170 154.805 163.310 ;
        RECT 152.200 163.110 152.520 163.170 ;
        RECT 154.515 163.125 154.805 163.170 ;
        RECT 74.920 162.970 75.210 163.015 ;
        RECT 76.490 162.970 76.780 163.015 ;
        RECT 78.590 162.970 78.880 163.015 ;
        RECT 97.460 162.970 97.780 163.030 ;
        RECT 74.920 162.830 78.880 162.970 ;
        RECT 74.920 162.785 75.210 162.830 ;
        RECT 76.490 162.785 76.780 162.830 ;
        RECT 78.590 162.785 78.880 162.830 ;
        RECT 81.680 162.830 97.230 162.970 ;
        RECT 72.160 162.430 72.480 162.690 ;
        RECT 74.485 162.630 74.775 162.675 ;
        RECT 77.005 162.630 77.295 162.675 ;
        RECT 78.195 162.630 78.485 162.675 ;
        RECT 74.485 162.490 78.485 162.630 ;
        RECT 74.485 162.445 74.775 162.490 ;
        RECT 77.005 162.445 77.295 162.490 ;
        RECT 78.195 162.445 78.485 162.490 ;
        RECT 72.250 162.290 72.390 162.430 ;
        RECT 79.075 162.290 79.365 162.335 ;
        RECT 72.250 162.150 79.365 162.290 ;
        RECT 79.075 162.105 79.365 162.150 ;
        RECT 77.850 161.950 78.140 161.995 ;
        RECT 81.680 161.950 81.820 162.830 ;
        RECT 87.800 162.630 88.120 162.690 ;
        RECT 97.090 162.675 97.230 162.830 ;
        RECT 97.460 162.830 100.910 162.970 ;
        RECT 97.460 162.770 97.780 162.830 ;
        RECT 93.335 162.630 93.625 162.675 ;
        RECT 87.800 162.490 93.625 162.630 ;
        RECT 87.800 162.430 88.120 162.490 ;
        RECT 93.335 162.445 93.625 162.490 ;
        RECT 97.015 162.445 97.305 162.675 ;
        RECT 100.235 162.630 100.525 162.675 ;
        RECT 98.010 162.490 100.525 162.630 ;
        RECT 87.340 162.290 87.660 162.350 ;
        RECT 88.735 162.290 89.025 162.335 ;
        RECT 91.495 162.290 91.785 162.335 ;
        RECT 87.340 162.150 91.785 162.290 ;
        RECT 87.340 162.090 87.660 162.150 ;
        RECT 88.735 162.105 89.025 162.150 ;
        RECT 91.495 162.105 91.785 162.150 ;
        RECT 91.955 162.105 92.245 162.335 ;
        RECT 93.795 162.105 94.085 162.335 ;
        RECT 95.635 162.290 95.925 162.335 ;
        RECT 96.080 162.290 96.400 162.350 ;
        RECT 97.460 162.290 97.780 162.350 ;
        RECT 98.010 162.335 98.150 162.490 ;
        RECT 100.235 162.445 100.525 162.490 ;
        RECT 95.635 162.150 97.780 162.290 ;
        RECT 95.635 162.105 95.925 162.150 ;
        RECT 77.850 161.810 81.820 161.950 ;
        RECT 77.850 161.765 78.140 161.810 ;
        RECT 86.880 161.750 87.200 162.010 ;
        RECT 92.030 161.950 92.170 162.105 ;
        RECT 93.870 161.950 94.010 162.105 ;
        RECT 96.080 162.090 96.400 162.150 ;
        RECT 97.460 162.090 97.780 162.150 ;
        RECT 97.935 162.105 98.225 162.335 ;
        RECT 98.395 162.105 98.685 162.335 ;
        RECT 99.775 162.290 100.065 162.335 ;
        RECT 100.770 162.290 100.910 162.830 ;
        RECT 101.155 162.785 101.445 163.015 ;
        RECT 102.150 162.970 102.290 163.110 ;
        RECT 103.455 162.970 103.745 163.015 ;
        RECT 102.150 162.830 104.590 162.970 ;
        RECT 103.455 162.785 103.745 162.830 ;
        RECT 99.775 162.150 100.910 162.290 ;
        RECT 99.775 162.105 100.065 162.150 ;
        RECT 92.030 161.810 94.010 161.950 ;
        RECT 98.470 161.950 98.610 162.105 ;
        RECT 100.680 161.950 101.000 162.010 ;
        RECT 98.470 161.810 101.000 161.950 ;
        RECT 101.230 161.950 101.370 162.785 ;
        RECT 101.600 162.630 101.920 162.690 ;
        RECT 102.535 162.630 102.825 162.675 ;
        RECT 101.600 162.490 102.825 162.630 ;
        RECT 101.600 162.430 101.920 162.490 ;
        RECT 102.535 162.445 102.825 162.490 ;
        RECT 102.980 162.090 103.300 162.350 ;
        RECT 104.450 162.335 104.590 162.830 ;
        RECT 104.820 162.430 105.140 162.690 ;
        RECT 107.210 162.630 107.350 163.110 ;
        RECT 121.840 162.970 122.160 163.030 ;
        RECT 125.060 162.970 125.380 163.030 ;
        RECT 121.840 162.830 125.380 162.970 ;
        RECT 121.840 162.770 122.160 162.830 ;
        RECT 125.060 162.770 125.380 162.830 ;
        RECT 148.100 162.970 148.390 163.015 ;
        RECT 150.200 162.970 150.490 163.015 ;
        RECT 151.770 162.970 152.060 163.015 ;
        RECT 148.100 162.830 152.060 162.970 ;
        RECT 148.100 162.785 148.390 162.830 ;
        RECT 150.200 162.785 150.490 162.830 ;
        RECT 151.770 162.785 152.060 162.830 ;
        RECT 110.355 162.630 110.645 162.675 ;
        RECT 116.320 162.630 116.640 162.690 ;
        RECT 119.540 162.630 119.860 162.690 ;
        RECT 129.200 162.630 129.520 162.690 ;
        RECT 107.210 162.490 110.645 162.630 ;
        RECT 104.375 162.105 104.665 162.335 ;
        RECT 105.280 162.090 105.600 162.350 ;
        RECT 107.120 162.300 107.440 162.350 ;
        RECT 106.750 162.290 107.440 162.300 ;
        RECT 106.290 162.160 107.440 162.290 ;
        RECT 106.290 162.150 106.890 162.160 ;
        RECT 104.820 161.950 105.140 162.010 ;
        RECT 106.290 161.950 106.430 162.150 ;
        RECT 107.120 162.090 107.440 162.160 ;
        RECT 101.230 161.810 104.590 161.950 ;
        RECT 93.870 161.670 94.010 161.810 ;
        RECT 100.680 161.750 101.000 161.810 ;
        RECT 93.780 161.410 94.100 161.670 ;
        RECT 104.450 161.610 104.590 161.810 ;
        RECT 104.820 161.810 106.430 161.950 ;
        RECT 104.820 161.750 105.140 161.810 ;
        RECT 107.670 161.610 107.810 162.490 ;
        RECT 110.355 162.445 110.645 162.490 ;
        RECT 111.350 162.490 116.640 162.630 ;
        RECT 108.500 162.290 108.820 162.350 ;
        RECT 111.350 162.290 111.490 162.490 ;
        RECT 108.500 162.150 111.490 162.290 ;
        RECT 111.735 162.290 112.025 162.335 ;
        RECT 113.560 162.290 113.880 162.350 ;
        RECT 115.950 162.335 116.090 162.490 ;
        RECT 116.320 162.430 116.640 162.490 ;
        RECT 118.250 162.490 119.860 162.630 ;
        RECT 118.250 162.350 118.390 162.490 ;
        RECT 119.540 162.430 119.860 162.490 ;
        RECT 120.090 162.490 129.520 162.630 ;
        RECT 111.735 162.150 113.880 162.290 ;
        RECT 108.500 162.090 108.820 162.150 ;
        RECT 111.735 162.105 112.025 162.150 ;
        RECT 113.560 162.090 113.880 162.150 ;
        RECT 114.955 162.105 115.245 162.335 ;
        RECT 115.875 162.105 116.165 162.335 ;
        RECT 108.040 161.950 108.360 162.010 ;
        RECT 115.030 161.950 115.170 162.105 ;
        RECT 117.700 162.090 118.020 162.350 ;
        RECT 118.160 162.090 118.480 162.350 ;
        RECT 120.090 162.335 120.230 162.490 ;
        RECT 129.200 162.430 129.520 162.490 ;
        RECT 137.020 162.430 137.340 162.690 ;
        RECT 142.540 162.630 142.860 162.690 ;
        RECT 147.615 162.630 147.905 162.675 ;
        RECT 142.540 162.490 147.905 162.630 ;
        RECT 142.540 162.430 142.860 162.490 ;
        RECT 147.615 162.445 147.905 162.490 ;
        RECT 148.495 162.630 148.785 162.675 ;
        RECT 149.685 162.630 149.975 162.675 ;
        RECT 152.205 162.630 152.495 162.675 ;
        RECT 148.495 162.490 152.495 162.630 ;
        RECT 148.495 162.445 148.785 162.490 ;
        RECT 149.685 162.445 149.975 162.490 ;
        RECT 152.205 162.445 152.495 162.490 ;
        RECT 120.015 162.105 120.305 162.335 ;
        RECT 126.440 162.290 126.760 162.350 ;
        RECT 126.440 162.150 127.590 162.290 ;
        RECT 126.440 162.090 126.760 162.150 ;
        RECT 117.790 161.950 117.930 162.090 ;
        RECT 127.450 162.010 127.590 162.150 ;
        RECT 135.655 162.105 135.945 162.335 ;
        RECT 136.575 162.290 136.865 162.335 ;
        RECT 137.495 162.290 137.785 162.335 ;
        RECT 136.190 162.150 136.865 162.290 ;
        RECT 119.080 161.950 119.400 162.010 ;
        RECT 108.040 161.810 117.930 161.950 ;
        RECT 118.710 161.810 119.400 161.950 ;
        RECT 108.040 161.750 108.360 161.810 ;
        RECT 118.710 161.655 118.850 161.810 ;
        RECT 119.080 161.750 119.400 161.810 ;
        RECT 124.155 161.765 124.445 161.995 ;
        RECT 118.635 161.610 118.925 161.655 ;
        RECT 104.450 161.470 107.810 161.610 ;
        RECT 118.525 161.470 118.925 161.610 ;
        RECT 118.635 161.425 118.925 161.470 ;
        RECT 119.555 161.610 119.845 161.655 ;
        RECT 122.760 161.610 123.080 161.670 ;
        RECT 119.555 161.470 123.080 161.610 ;
        RECT 119.555 161.425 119.845 161.470 ;
        RECT 122.760 161.410 123.080 161.470 ;
        RECT 123.220 161.410 123.540 161.670 ;
        RECT 124.230 161.610 124.370 161.765 ;
        RECT 125.060 161.750 125.380 162.010 ;
        RECT 127.360 161.750 127.680 162.010 ;
        RECT 135.730 161.670 135.870 162.105 ;
        RECT 136.190 161.670 136.330 162.150 ;
        RECT 136.575 162.105 136.865 162.150 ;
        RECT 137.110 162.150 137.785 162.290 ;
        RECT 137.110 161.670 137.250 162.150 ;
        RECT 137.495 162.105 137.785 162.150 ;
        RECT 138.415 162.290 138.705 162.335 ;
        RECT 138.860 162.290 139.180 162.350 ;
        RECT 138.415 162.150 139.180 162.290 ;
        RECT 138.415 162.105 138.705 162.150 ;
        RECT 138.860 162.090 139.180 162.150 ;
        RECT 148.950 161.950 149.240 161.995 ;
        RECT 151.740 161.950 152.060 162.010 ;
        RECT 138.950 161.810 140.010 161.950 ;
        RECT 138.950 161.670 139.090 161.810 ;
        RECT 139.870 161.670 140.010 161.810 ;
        RECT 148.950 161.810 152.060 161.950 ;
        RECT 148.950 161.765 149.240 161.810 ;
        RECT 151.740 161.750 152.060 161.810 ;
        RECT 125.535 161.610 125.825 161.655 ;
        RECT 128.740 161.610 129.060 161.670 ;
        RECT 124.230 161.470 129.060 161.610 ;
        RECT 125.535 161.425 125.825 161.470 ;
        RECT 128.740 161.410 129.060 161.470 ;
        RECT 135.640 161.410 135.960 161.670 ;
        RECT 136.100 161.410 136.420 161.670 ;
        RECT 137.020 161.410 137.340 161.670 ;
        RECT 138.860 161.410 139.180 161.670 ;
        RECT 139.320 161.410 139.640 161.670 ;
        RECT 139.780 161.410 140.100 161.670 ;
        RECT 70.710 160.790 156.270 161.270 ;
        RECT 79.060 160.390 79.380 160.650 ;
        RECT 81.360 160.390 81.680 160.650 ;
        RECT 84.120 160.390 84.440 160.650 ;
        RECT 89.180 160.390 89.500 160.650 ;
        RECT 98.525 160.590 98.815 160.635 ;
        RECT 101.615 160.590 101.905 160.635 ;
        RECT 102.980 160.590 103.300 160.650 ;
        RECT 98.525 160.450 103.300 160.590 ;
        RECT 98.525 160.405 98.815 160.450 ;
        RECT 101.615 160.405 101.905 160.450 ;
        RECT 102.980 160.390 103.300 160.450 ;
        RECT 118.620 160.590 118.940 160.650 ;
        RECT 137.020 160.590 137.340 160.650 ;
        RECT 118.620 160.450 129.430 160.590 ;
        RECT 118.620 160.390 118.940 160.450 ;
        RECT 79.150 160.250 79.290 160.390 ;
        RECT 78.690 160.110 79.290 160.250 ;
        RECT 81.450 160.250 81.590 160.390 ;
        RECT 81.450 160.110 83.430 160.250 ;
        RECT 75.855 159.910 76.145 159.955 ;
        RECT 77.680 159.910 78.000 159.970 ;
        RECT 78.690 159.955 78.830 160.110 ;
        RECT 75.855 159.770 78.000 159.910 ;
        RECT 75.855 159.725 76.145 159.770 ;
        RECT 77.680 159.710 78.000 159.770 ;
        RECT 78.615 159.725 78.905 159.955 ;
        RECT 79.060 159.710 79.380 159.970 ;
        RECT 79.520 159.910 79.840 159.970 ;
        RECT 80.900 159.910 81.220 159.970 ;
        RECT 83.290 159.955 83.430 160.110 ;
        RECT 81.835 159.910 82.125 159.955 ;
        RECT 79.520 159.770 82.125 159.910 ;
        RECT 79.520 159.710 79.840 159.770 ;
        RECT 80.900 159.710 81.220 159.770 ;
        RECT 81.835 159.725 82.125 159.770 ;
        RECT 82.755 159.725 83.045 159.955 ;
        RECT 83.215 159.725 83.505 159.955 ;
        RECT 83.660 159.910 83.980 159.970 ;
        RECT 88.260 159.910 88.580 159.970 ;
        RECT 83.660 159.770 88.580 159.910 ;
        RECT 89.270 159.910 89.410 160.390 ;
        RECT 91.035 160.250 91.325 160.295 ;
        RECT 93.780 160.250 94.100 160.310 ;
        RECT 91.035 160.110 94.100 160.250 ;
        RECT 91.035 160.065 91.325 160.110 ;
        RECT 93.780 160.050 94.100 160.110 ;
        RECT 97.460 160.050 97.780 160.310 ;
        RECT 99.775 160.250 100.065 160.295 ;
        RECT 98.470 160.110 100.065 160.250 ;
        RECT 89.640 159.910 89.960 159.970 ;
        RECT 89.270 159.770 89.960 159.910 ;
        RECT 77.220 159.370 77.540 159.630 ;
        RECT 78.155 159.385 78.445 159.615 ;
        RECT 79.150 159.570 79.290 159.710 ;
        RECT 82.830 159.570 82.970 159.725 ;
        RECT 83.660 159.710 83.980 159.770 ;
        RECT 88.260 159.710 88.580 159.770 ;
        RECT 89.640 159.710 89.960 159.770 ;
        RECT 92.400 159.910 92.720 159.970 ;
        RECT 93.335 159.910 93.625 159.955 ;
        RECT 92.400 159.770 93.625 159.910 ;
        RECT 92.400 159.710 92.720 159.770 ;
        RECT 93.335 159.725 93.625 159.770 ;
        RECT 94.240 159.910 94.560 159.970 ;
        RECT 94.715 159.910 95.005 159.955 ;
        RECT 94.240 159.770 95.005 159.910 ;
        RECT 94.240 159.710 94.560 159.770 ;
        RECT 94.715 159.725 95.005 159.770 ;
        RECT 95.620 159.710 95.940 159.970 ;
        RECT 92.875 159.570 93.165 159.615 ;
        RECT 95.710 159.570 95.850 159.710 ;
        RECT 98.470 159.630 98.610 160.110 ;
        RECT 99.775 160.065 100.065 160.110 ;
        RECT 100.855 160.250 101.145 160.295 ;
        RECT 108.500 160.250 108.820 160.310 ;
        RECT 100.855 160.110 108.820 160.250 ;
        RECT 100.855 160.065 101.145 160.110 ;
        RECT 108.500 160.050 108.820 160.110 ;
        RECT 109.420 160.250 109.740 160.310 ;
        RECT 114.020 160.250 114.340 160.310 ;
        RECT 129.290 160.250 129.430 160.450 ;
        RECT 137.020 160.450 141.390 160.590 ;
        RECT 137.020 160.390 137.340 160.450 ;
        RECT 109.420 160.110 114.340 160.250 ;
        RECT 109.420 160.050 109.740 160.110 ;
        RECT 114.020 160.050 114.340 160.110 ;
        RECT 121.930 160.110 128.970 160.250 ;
        RECT 108.040 159.910 108.360 159.970 ;
        RECT 121.930 159.955 122.070 160.110 ;
        RECT 128.830 159.970 128.970 160.110 ;
        RECT 129.290 160.110 140.470 160.250 ;
        RECT 108.040 159.770 108.730 159.910 ;
        RECT 108.040 159.710 108.360 159.770 ;
        RECT 79.150 159.430 82.970 159.570 ;
        RECT 90.650 159.430 95.850 159.570 ;
        RECT 76.315 159.230 76.605 159.275 ;
        RECT 77.680 159.230 78.000 159.290 ;
        RECT 78.230 159.230 78.370 159.385 ;
        RECT 76.315 159.090 78.370 159.230 ;
        RECT 80.455 159.230 80.745 159.275 ;
        RECT 85.500 159.230 85.820 159.290 ;
        RECT 80.455 159.090 85.820 159.230 ;
        RECT 76.315 159.045 76.605 159.090 ;
        RECT 77.680 159.030 78.000 159.090 ;
        RECT 80.455 159.045 80.745 159.090 ;
        RECT 85.500 159.030 85.820 159.090 ;
        RECT 87.800 159.230 88.120 159.290 ;
        RECT 90.650 159.275 90.790 159.430 ;
        RECT 92.875 159.385 93.165 159.430 ;
        RECT 98.380 159.370 98.700 159.630 ;
        RECT 108.590 159.615 108.730 159.770 ;
        RECT 119.555 159.725 119.845 159.955 ;
        RECT 120.475 159.910 120.765 159.955 ;
        RECT 121.855 159.910 122.145 159.955 ;
        RECT 120.475 159.770 122.145 159.910 ;
        RECT 120.475 159.725 120.765 159.770 ;
        RECT 121.855 159.725 122.145 159.770 ;
        RECT 123.695 159.910 123.985 159.955 ;
        RECT 124.140 159.910 124.460 159.970 ;
        RECT 123.695 159.770 124.460 159.910 ;
        RECT 123.695 159.725 123.985 159.770 ;
        RECT 108.515 159.385 108.805 159.615 ;
        RECT 109.895 159.570 110.185 159.615 ;
        RECT 119.630 159.570 119.770 159.725 ;
        RECT 124.140 159.710 124.460 159.770 ;
        RECT 125.075 159.910 125.365 159.955 ;
        RECT 126.455 159.910 126.745 159.955 ;
        RECT 125.075 159.770 126.745 159.910 ;
        RECT 125.075 159.725 125.365 159.770 ;
        RECT 126.455 159.725 126.745 159.770 ;
        RECT 127.375 159.725 127.665 159.955 ;
        RECT 125.520 159.570 125.840 159.630 ;
        RECT 127.450 159.570 127.590 159.725 ;
        RECT 128.740 159.710 129.060 159.970 ;
        RECT 129.290 159.955 129.430 160.110 ;
        RECT 136.190 159.970 136.330 160.110 ;
        RECT 129.215 159.725 129.505 159.955 ;
        RECT 130.135 159.725 130.425 159.955 ;
        RECT 109.895 159.430 110.570 159.570 ;
        RECT 119.630 159.430 122.070 159.570 ;
        RECT 109.895 159.385 110.185 159.430 ;
        RECT 90.575 159.230 90.865 159.275 ;
        RECT 95.635 159.230 95.925 159.275 ;
        RECT 98.470 159.230 98.610 159.370 ;
        RECT 87.800 159.090 90.865 159.230 ;
        RECT 87.800 159.030 88.120 159.090 ;
        RECT 90.575 159.045 90.865 159.090 ;
        RECT 93.410 159.090 98.610 159.230 ;
        RECT 99.315 159.230 99.605 159.275 ;
        RECT 103.440 159.230 103.760 159.290 ;
        RECT 99.315 159.090 103.760 159.230 ;
        RECT 76.760 158.690 77.080 158.950 ;
        RECT 80.900 158.690 81.220 158.950 ;
        RECT 89.195 158.890 89.485 158.935 ;
        RECT 92.860 158.890 93.180 158.950 ;
        RECT 93.410 158.935 93.550 159.090 ;
        RECT 95.635 159.045 95.925 159.090 ;
        RECT 99.315 159.045 99.605 159.090 ;
        RECT 103.440 159.030 103.760 159.090 ;
        RECT 110.430 158.950 110.570 159.430 ;
        RECT 121.930 159.290 122.070 159.430 ;
        RECT 125.520 159.430 127.590 159.570 ;
        RECT 125.520 159.370 125.840 159.430 ;
        RECT 128.295 159.385 128.585 159.615 ;
        RECT 130.210 159.570 130.350 159.725 ;
        RECT 130.580 159.710 130.900 159.970 ;
        RECT 133.800 159.710 134.120 159.970 ;
        RECT 135.195 159.910 135.485 159.955 ;
        RECT 135.640 159.910 135.960 159.970 ;
        RECT 135.195 159.770 135.960 159.910 ;
        RECT 135.195 159.725 135.485 159.770 ;
        RECT 135.640 159.710 135.960 159.770 ;
        RECT 136.100 159.955 136.420 159.970 ;
        RECT 136.100 159.725 136.425 159.955 ;
        RECT 136.100 159.710 136.420 159.725 ;
        RECT 137.020 159.710 137.340 159.970 ;
        RECT 137.955 159.910 138.245 159.955 ;
        RECT 138.860 159.910 139.180 159.970 ;
        RECT 140.330 159.955 140.470 160.110 ;
        RECT 137.955 159.770 139.180 159.910 ;
        RECT 137.955 159.725 138.245 159.770 ;
        RECT 138.860 159.710 139.180 159.770 ;
        RECT 139.335 159.725 139.625 159.955 ;
        RECT 140.255 159.725 140.545 159.955 ;
        RECT 133.890 159.570 134.030 159.710 ;
        RECT 136.575 159.570 136.865 159.615 ;
        RECT 130.210 159.430 131.730 159.570 ;
        RECT 133.890 159.430 136.865 159.570 ;
        RECT 120.935 159.230 121.225 159.275 ;
        RECT 118.250 159.090 121.225 159.230 ;
        RECT 118.250 158.950 118.390 159.090 ;
        RECT 120.935 159.045 121.225 159.090 ;
        RECT 121.840 159.030 122.160 159.290 ;
        RECT 126.440 159.230 126.760 159.290 ;
        RECT 124.230 159.090 126.760 159.230 ;
        RECT 89.195 158.750 93.180 158.890 ;
        RECT 89.195 158.705 89.485 158.750 ;
        RECT 92.860 158.690 93.180 158.750 ;
        RECT 93.335 158.705 93.625 158.935 ;
        RECT 94.240 158.690 94.560 158.950 ;
        RECT 95.160 158.890 95.480 158.950 ;
        RECT 98.395 158.890 98.685 158.935 ;
        RECT 95.160 158.750 98.685 158.890 ;
        RECT 95.160 158.690 95.480 158.750 ;
        RECT 98.395 158.705 98.685 158.750 ;
        RECT 100.680 158.890 101.000 158.950 ;
        RECT 110.340 158.890 110.660 158.950 ;
        RECT 100.680 158.750 110.660 158.890 ;
        RECT 100.680 158.690 101.000 158.750 ;
        RECT 110.340 158.690 110.660 158.750 ;
        RECT 118.160 158.690 118.480 158.950 ;
        RECT 120.000 158.690 120.320 158.950 ;
        RECT 121.380 158.890 121.700 158.950 ;
        RECT 124.230 158.935 124.370 159.090 ;
        RECT 126.440 159.030 126.760 159.090 ;
        RECT 124.155 158.890 124.445 158.935 ;
        RECT 121.380 158.750 124.445 158.890 ;
        RECT 121.380 158.690 121.700 158.750 ;
        RECT 124.155 158.705 124.445 158.750 ;
        RECT 125.980 158.690 126.300 158.950 ;
        RECT 128.370 158.890 128.510 159.385 ;
        RECT 131.590 159.275 131.730 159.430 ;
        RECT 136.575 159.385 136.865 159.430 ;
        RECT 131.515 159.230 131.805 159.275 ;
        RECT 135.640 159.230 135.960 159.290 ;
        RECT 139.410 159.230 139.550 159.725 ;
        RECT 140.700 159.710 141.020 159.970 ;
        RECT 141.250 159.955 141.390 160.450 ;
        RECT 143.920 160.390 144.240 160.650 ;
        RECT 144.395 160.590 144.685 160.635 ;
        RECT 149.535 160.590 149.825 160.635 ;
        RECT 144.395 160.450 149.825 160.590 ;
        RECT 144.395 160.405 144.685 160.450 ;
        RECT 149.535 160.405 149.825 160.450 ;
        RECT 150.835 160.590 151.125 160.635 ;
        RECT 151.740 160.590 152.060 160.650 ;
        RECT 150.835 160.450 152.060 160.590 ;
        RECT 150.835 160.405 151.125 160.450 ;
        RECT 151.740 160.390 152.060 160.450 ;
        RECT 144.010 160.250 144.150 160.390 ;
        RECT 145.315 160.250 145.605 160.295 ;
        RECT 144.010 160.110 145.605 160.250 ;
        RECT 141.175 159.725 141.465 159.955 ;
        RECT 141.620 159.910 141.940 159.970 ;
        RECT 142.095 159.910 142.385 159.955 ;
        RECT 142.540 159.910 142.860 159.970 ;
        RECT 141.620 159.770 142.860 159.910 ;
        RECT 141.620 159.710 141.940 159.770 ;
        RECT 142.095 159.725 142.385 159.770 ;
        RECT 142.540 159.710 142.860 159.770 ;
        RECT 143.920 159.710 144.240 159.970 ;
        RECT 144.930 159.955 145.070 160.110 ;
        RECT 145.315 160.065 145.605 160.110 ;
        RECT 146.680 160.250 147.000 160.310 ;
        RECT 148.535 160.250 148.825 160.295 ;
        RECT 146.680 160.110 148.825 160.250 ;
        RECT 146.680 160.050 147.000 160.110 ;
        RECT 148.535 160.065 148.825 160.110 ;
        RECT 144.855 159.725 145.145 159.955 ;
        RECT 146.235 159.725 146.525 159.955 ;
        RECT 151.755 159.910 152.045 159.955 ;
        RECT 150.450 159.770 152.045 159.910 ;
        RECT 131.515 159.090 139.550 159.230 ;
        RECT 141.160 159.230 141.480 159.290 ;
        RECT 146.310 159.230 146.450 159.725 ;
        RECT 150.450 159.275 150.590 159.770 ;
        RECT 151.755 159.725 152.045 159.770 ;
        RECT 141.160 159.090 146.450 159.230 ;
        RECT 131.515 159.045 131.805 159.090 ;
        RECT 135.640 159.030 135.960 159.090 ;
        RECT 141.160 159.030 141.480 159.090 ;
        RECT 150.375 159.045 150.665 159.275 ;
        RECT 129.660 158.890 129.980 158.950 ;
        RECT 137.020 158.890 137.340 158.950 ;
        RECT 128.370 158.750 137.340 158.890 ;
        RECT 129.660 158.690 129.980 158.750 ;
        RECT 137.020 158.690 137.340 158.750 ;
        RECT 138.875 158.890 139.165 158.935 ;
        RECT 142.540 158.890 142.860 158.950 ;
        RECT 138.875 158.750 142.860 158.890 ;
        RECT 138.875 158.705 139.165 158.750 ;
        RECT 142.540 158.690 142.860 158.750 ;
        RECT 143.000 158.690 143.320 158.950 ;
        RECT 147.155 158.890 147.445 158.935 ;
        RECT 149.455 158.890 149.745 158.935 ;
        RECT 147.155 158.750 149.745 158.890 ;
        RECT 147.155 158.705 147.445 158.750 ;
        RECT 149.455 158.705 149.745 158.750 ;
        RECT 70.710 158.070 156.270 158.550 ;
        RECT 77.220 157.670 77.540 157.930 ;
        RECT 77.680 157.870 78.000 157.930 ;
        RECT 78.155 157.870 78.445 157.915 ;
        RECT 77.680 157.730 78.445 157.870 ;
        RECT 77.680 157.670 78.000 157.730 ;
        RECT 78.155 157.685 78.445 157.730 ;
        RECT 80.900 157.670 81.220 157.930 ;
        RECT 89.180 157.870 89.500 157.930 ;
        RECT 89.655 157.870 89.945 157.915 ;
        RECT 91.035 157.870 91.325 157.915 ;
        RECT 89.180 157.730 89.945 157.870 ;
        RECT 89.180 157.670 89.500 157.730 ;
        RECT 89.655 157.685 89.945 157.730 ;
        RECT 90.650 157.730 91.325 157.870 ;
        RECT 77.310 157.530 77.450 157.670 ;
        RECT 79.535 157.530 79.825 157.575 ;
        RECT 77.310 157.390 79.825 157.530 ;
        RECT 77.310 156.850 77.450 157.390 ;
        RECT 79.535 157.345 79.825 157.390 ;
        RECT 80.990 157.190 81.130 157.670 ;
        RECT 88.720 157.330 89.040 157.590 ;
        RECT 78.690 157.050 81.130 157.190 ;
        RECT 86.435 157.190 86.725 157.235 ;
        RECT 90.115 157.190 90.405 157.235 ;
        RECT 90.650 157.190 90.790 157.730 ;
        RECT 91.035 157.685 91.325 157.730 ;
        RECT 92.860 157.870 93.180 157.930 ;
        RECT 93.795 157.870 94.085 157.915 ;
        RECT 95.160 157.870 95.480 157.930 ;
        RECT 92.860 157.730 95.480 157.870 ;
        RECT 92.860 157.670 93.180 157.730 ;
        RECT 93.795 157.685 94.085 157.730 ;
        RECT 95.160 157.670 95.480 157.730 ;
        RECT 95.635 157.870 95.925 157.915 ;
        RECT 97.000 157.870 97.320 157.930 ;
        RECT 95.635 157.730 97.320 157.870 ;
        RECT 95.635 157.685 95.925 157.730 ;
        RECT 97.000 157.670 97.320 157.730 ;
        RECT 97.460 157.870 97.780 157.930 ;
        RECT 98.395 157.870 98.685 157.915 ;
        RECT 97.460 157.730 98.685 157.870 ;
        RECT 97.460 157.670 97.780 157.730 ;
        RECT 98.395 157.685 98.685 157.730 ;
        RECT 100.220 157.870 100.540 157.930 ;
        RECT 115.400 157.870 115.720 157.930 ;
        RECT 100.220 157.730 115.720 157.870 ;
        RECT 100.220 157.670 100.540 157.730 ;
        RECT 115.400 157.670 115.720 157.730 ;
        RECT 116.320 157.870 116.640 157.930 ;
        RECT 116.320 157.730 118.390 157.870 ;
        RECT 116.320 157.670 116.640 157.730 ;
        RECT 94.240 157.530 94.560 157.590 ;
        RECT 107.580 157.530 107.900 157.590 ;
        RECT 116.780 157.530 117.100 157.590 ;
        RECT 94.240 157.390 107.900 157.530 ;
        RECT 94.240 157.330 94.560 157.390 ;
        RECT 107.580 157.330 107.900 157.390 ;
        RECT 111.350 157.390 117.100 157.530 ;
        RECT 118.250 157.530 118.390 157.730 ;
        RECT 118.620 157.670 118.940 157.930 ;
        RECT 120.000 157.670 120.320 157.930 ;
        RECT 121.380 157.670 121.700 157.930 ;
        RECT 125.980 157.670 126.300 157.930 ;
        RECT 126.440 157.670 126.760 157.930 ;
        RECT 128.295 157.870 128.585 157.915 ;
        RECT 128.740 157.870 129.060 157.930 ;
        RECT 128.295 157.730 129.060 157.870 ;
        RECT 128.295 157.685 128.585 157.730 ;
        RECT 128.740 157.670 129.060 157.730 ;
        RECT 129.660 157.670 129.980 157.930 ;
        RECT 130.120 157.870 130.440 157.930 ;
        RECT 132.420 157.870 132.740 157.930 ;
        RECT 130.120 157.730 132.740 157.870 ;
        RECT 130.120 157.670 130.440 157.730 ;
        RECT 132.420 157.670 132.740 157.730 ;
        RECT 137.020 157.870 137.340 157.930 ;
        RECT 141.620 157.870 141.940 157.930 ;
        RECT 137.020 157.730 141.940 157.870 ;
        RECT 137.020 157.670 137.340 157.730 ;
        RECT 141.620 157.670 141.940 157.730 ;
        RECT 119.540 157.530 119.860 157.590 ;
        RECT 118.250 157.390 119.860 157.530 ;
        RECT 120.090 157.530 120.230 157.670 ;
        RECT 120.090 157.390 124.830 157.530 ;
        RECT 86.435 157.050 90.790 157.190 ;
        RECT 93.780 157.190 94.100 157.250 ;
        RECT 93.780 157.050 97.690 157.190 ;
        RECT 78.690 156.895 78.830 157.050 ;
        RECT 86.435 157.005 86.725 157.050 ;
        RECT 90.115 157.005 90.405 157.050 ;
        RECT 93.780 156.990 94.100 157.050 ;
        RECT 77.695 156.850 77.985 156.895 ;
        RECT 77.310 156.710 77.985 156.850 ;
        RECT 77.695 156.665 77.985 156.710 ;
        RECT 78.615 156.665 78.905 156.895 ;
        RECT 79.075 156.850 79.365 156.895 ;
        RECT 79.520 156.850 79.840 156.910 ;
        RECT 79.075 156.710 79.840 156.850 ;
        RECT 79.075 156.665 79.365 156.710 ;
        RECT 79.520 156.650 79.840 156.710 ;
        RECT 79.995 156.665 80.285 156.895 ;
        RECT 76.760 156.170 77.080 156.230 ;
        RECT 78.140 156.170 78.460 156.230 ;
        RECT 76.760 156.030 78.460 156.170 ;
        RECT 76.760 155.970 77.080 156.030 ;
        RECT 78.140 155.970 78.460 156.030 ;
        RECT 79.060 156.170 79.380 156.230 ;
        RECT 80.070 156.170 80.210 156.665 ;
        RECT 80.440 156.650 80.760 156.910 ;
        RECT 81.360 156.650 81.680 156.910 ;
        RECT 82.295 156.850 82.585 156.895 ;
        RECT 86.895 156.850 87.185 156.895 ;
        RECT 82.295 156.710 87.185 156.850 ;
        RECT 82.295 156.665 82.585 156.710 ;
        RECT 86.895 156.665 87.185 156.710 ;
        RECT 84.120 156.310 84.440 156.570 ;
        RECT 86.970 156.510 87.110 156.665 ;
        RECT 87.800 156.650 88.120 156.910 ;
        RECT 90.575 156.850 90.865 156.895 ;
        RECT 88.350 156.710 90.865 156.850 ;
        RECT 87.340 156.510 87.660 156.570 ;
        RECT 88.350 156.510 88.490 156.710 ;
        RECT 90.575 156.665 90.865 156.710 ;
        RECT 91.035 156.665 91.325 156.895 ;
        RECT 91.955 156.665 92.245 156.895 ;
        RECT 92.400 156.850 92.720 156.910 ;
        RECT 92.875 156.850 93.165 156.895 ;
        RECT 94.715 156.850 95.005 156.895 ;
        RECT 92.400 156.710 95.005 156.850 ;
        RECT 86.970 156.370 88.490 156.510 ;
        RECT 89.195 156.510 89.485 156.555 ;
        RECT 89.640 156.510 89.960 156.570 ;
        RECT 89.195 156.370 89.960 156.510 ;
        RECT 87.340 156.310 87.660 156.370 ;
        RECT 89.195 156.325 89.485 156.370 ;
        RECT 89.640 156.310 89.960 156.370 ;
        RECT 79.060 156.030 80.210 156.170 ;
        RECT 84.210 156.170 84.350 156.310 ;
        RECT 91.110 156.170 91.250 156.665 ;
        RECT 92.030 156.510 92.170 156.665 ;
        RECT 92.400 156.650 92.720 156.710 ;
        RECT 92.875 156.665 93.165 156.710 ;
        RECT 94.715 156.665 95.005 156.710 ;
        RECT 95.620 156.850 95.940 156.910 ;
        RECT 97.550 156.895 97.690 157.050 ;
        RECT 97.920 156.990 98.240 157.250 ;
        RECT 100.680 156.990 101.000 157.250 ;
        RECT 96.095 156.850 96.385 156.895 ;
        RECT 95.620 156.710 96.385 156.850 ;
        RECT 95.620 156.650 95.940 156.710 ;
        RECT 96.095 156.665 96.385 156.710 ;
        RECT 97.475 156.665 97.765 156.895 ;
        RECT 98.010 156.850 98.150 156.990 ;
        RECT 99.775 156.850 100.065 156.895 ;
        RECT 98.010 156.710 100.065 156.850 ;
        RECT 99.775 156.665 100.065 156.710 ;
        RECT 100.770 156.510 100.910 156.990 ;
        RECT 102.060 156.650 102.380 156.910 ;
        RECT 108.500 156.850 108.820 156.910 ;
        RECT 110.815 156.850 111.105 156.895 ;
        RECT 108.500 156.710 111.105 156.850 ;
        RECT 111.350 156.850 111.490 157.390 ;
        RECT 116.780 157.330 117.100 157.390 ;
        RECT 119.540 157.330 119.860 157.390 ;
        RECT 123.220 157.190 123.540 157.250 ;
        RECT 124.690 157.235 124.830 157.390 ;
        RECT 124.155 157.190 124.445 157.235 ;
        RECT 113.190 157.050 116.320 157.190 ;
        RECT 113.190 156.930 113.330 157.050 ;
        RECT 112.730 156.895 113.330 156.930 ;
        RECT 111.735 156.850 112.025 156.895 ;
        RECT 111.350 156.710 112.025 156.850 ;
        RECT 108.500 156.650 108.820 156.710 ;
        RECT 110.815 156.665 111.105 156.710 ;
        RECT 111.735 156.665 112.025 156.710 ;
        RECT 112.195 156.665 112.485 156.895 ;
        RECT 112.655 156.790 113.330 156.895 ;
        RECT 112.655 156.665 112.945 156.790 ;
        RECT 92.030 156.370 92.630 156.510 ;
        RECT 92.490 156.230 92.630 156.370 ;
        RECT 97.090 156.370 100.910 156.510 ;
        RECT 102.150 156.510 102.290 156.650 ;
        RECT 111.810 156.510 111.950 156.665 ;
        RECT 102.150 156.370 111.950 156.510 ;
        RECT 84.210 156.030 91.250 156.170 ;
        RECT 79.060 155.970 79.380 156.030 ;
        RECT 92.400 155.970 92.720 156.230 ;
        RECT 93.780 156.170 94.100 156.230 ;
        RECT 97.090 156.215 97.230 156.370 ;
        RECT 97.015 156.170 97.305 156.215 ;
        RECT 93.780 156.030 97.305 156.170 ;
        RECT 93.780 155.970 94.100 156.030 ;
        RECT 97.015 155.985 97.305 156.030 ;
        RECT 99.760 156.170 100.080 156.230 ;
        RECT 100.695 156.170 100.985 156.215 ;
        RECT 103.440 156.170 103.760 156.230 ;
        RECT 99.760 156.030 103.760 156.170 ;
        RECT 99.760 155.970 100.080 156.030 ;
        RECT 100.695 155.985 100.985 156.030 ;
        RECT 103.440 155.970 103.760 156.030 ;
        RECT 109.895 156.170 110.185 156.215 ;
        RECT 110.800 156.170 111.120 156.230 ;
        RECT 109.895 156.030 111.120 156.170 ;
        RECT 112.270 156.170 112.410 156.665 ;
        RECT 112.730 156.510 112.870 156.665 ;
        RECT 113.560 156.650 113.880 156.910 ;
        RECT 114.020 156.650 114.340 156.910 ;
        RECT 114.495 156.665 114.785 156.895 ;
        RECT 114.570 156.510 114.710 156.665 ;
        RECT 115.400 156.650 115.720 156.910 ;
        RECT 116.180 156.850 116.320 157.050 ;
        RECT 123.220 157.050 124.445 157.190 ;
        RECT 123.220 156.990 123.540 157.050 ;
        RECT 124.155 157.005 124.445 157.050 ;
        RECT 124.615 157.005 124.905 157.235 ;
        RECT 125.535 157.190 125.825 157.235 ;
        RECT 126.070 157.190 126.210 157.670 ;
        RECT 126.530 157.530 126.670 157.670 ;
        RECT 137.955 157.530 138.245 157.575 ;
        RECT 140.715 157.530 141.005 157.575 ;
        RECT 144.855 157.530 145.145 157.575 ;
        RECT 126.530 157.390 145.145 157.530 ;
        RECT 137.955 157.345 138.245 157.390 ;
        RECT 140.715 157.345 141.005 157.390 ;
        RECT 144.855 157.345 145.145 157.390 ;
        RECT 145.760 157.530 146.080 157.590 ;
        RECT 146.680 157.530 147.000 157.590 ;
        RECT 145.760 157.390 147.000 157.530 ;
        RECT 145.760 157.330 146.080 157.390 ;
        RECT 146.680 157.330 147.000 157.390 ;
        RECT 125.535 157.050 126.210 157.190 ;
        RECT 127.820 157.190 128.140 157.250 ;
        RECT 137.495 157.190 137.785 157.235 ;
        RECT 127.820 157.050 137.785 157.190 ;
        RECT 125.535 157.005 125.825 157.050 ;
        RECT 127.820 156.990 128.140 157.050 ;
        RECT 137.495 157.005 137.785 157.050 ;
        RECT 139.780 157.190 140.100 157.250 ;
        RECT 140.255 157.190 140.545 157.235 ;
        RECT 139.780 157.050 140.545 157.190 ;
        RECT 139.780 156.990 140.100 157.050 ;
        RECT 140.255 157.005 140.545 157.050 ;
        RECT 142.540 156.990 142.860 157.250 ;
        RECT 143.000 156.990 143.320 157.250 ;
        RECT 117.715 156.850 118.005 156.895 ;
        RECT 119.095 156.850 119.385 156.895 ;
        RECT 116.180 156.710 119.385 156.850 ;
        RECT 117.715 156.665 118.005 156.710 ;
        RECT 119.095 156.665 119.385 156.710 ;
        RECT 120.015 156.665 120.305 156.895 ;
        RECT 120.090 156.510 120.230 156.665 ;
        RECT 120.460 156.650 120.780 156.910 ;
        RECT 125.075 156.850 125.365 156.895 ;
        RECT 125.980 156.850 126.300 156.910 ;
        RECT 122.850 156.590 123.910 156.730 ;
        RECT 125.075 156.710 126.300 156.850 ;
        RECT 125.075 156.665 125.365 156.710 ;
        RECT 125.980 156.650 126.300 156.710 ;
        RECT 129.215 156.665 129.505 156.895 ;
        RECT 129.660 156.850 129.980 156.910 ;
        RECT 130.595 156.850 130.885 156.895 ;
        RECT 132.420 156.850 132.740 156.910 ;
        RECT 129.660 156.710 132.740 156.850 ;
        RECT 122.850 156.510 122.990 156.590 ;
        RECT 112.730 156.370 113.790 156.510 ;
        RECT 114.570 156.370 118.850 156.510 ;
        RECT 120.090 156.370 122.990 156.510 ;
        RECT 123.770 156.510 123.910 156.590 ;
        RECT 129.290 156.510 129.430 156.665 ;
        RECT 129.660 156.650 129.980 156.710 ;
        RECT 130.595 156.665 130.885 156.710 ;
        RECT 132.420 156.650 132.740 156.710 ;
        RECT 138.875 156.850 139.165 156.895 ;
        RECT 139.320 156.850 139.640 156.910 ;
        RECT 138.875 156.710 139.640 156.850 ;
        RECT 138.875 156.665 139.165 156.710 ;
        RECT 139.320 156.650 139.640 156.710 ;
        RECT 141.635 156.850 141.925 156.895 ;
        RECT 142.630 156.850 142.770 156.990 ;
        RECT 141.635 156.710 142.770 156.850 ;
        RECT 143.090 156.850 143.230 156.990 ;
        RECT 143.935 156.850 144.225 156.895 ;
        RECT 143.090 156.710 144.225 156.850 ;
        RECT 141.635 156.665 141.925 156.710 ;
        RECT 143.935 156.665 144.225 156.710 ;
        RECT 144.840 156.850 145.160 156.910 ;
        RECT 145.315 156.850 145.605 156.895 ;
        RECT 145.760 156.850 146.080 156.910 ;
        RECT 144.840 156.710 146.080 156.850 ;
        RECT 144.840 156.650 145.160 156.710 ;
        RECT 145.315 156.665 145.605 156.710 ;
        RECT 145.760 156.650 146.080 156.710 ;
        RECT 146.220 156.850 146.540 156.910 ;
        RECT 148.980 156.850 149.300 156.910 ;
        RECT 151.295 156.850 151.585 156.895 ;
        RECT 146.220 156.710 151.585 156.850 ;
        RECT 146.220 156.650 146.540 156.710 ;
        RECT 148.980 156.650 149.300 156.710 ;
        RECT 151.295 156.665 151.585 156.710 ;
        RECT 152.215 156.850 152.505 156.895 ;
        RECT 154.040 156.850 154.360 156.910 ;
        RECT 152.215 156.710 154.360 156.850 ;
        RECT 152.215 156.665 152.505 156.710 ;
        RECT 154.040 156.650 154.360 156.710 ;
        RECT 151.755 156.510 152.045 156.555 ;
        RECT 123.770 156.370 152.045 156.510 ;
        RECT 113.650 156.230 113.790 156.370 ;
        RECT 118.710 156.230 118.850 156.370 ;
        RECT 151.755 156.325 152.045 156.370 ;
        RECT 113.100 156.170 113.420 156.230 ;
        RECT 112.270 156.030 113.420 156.170 ;
        RECT 109.895 155.985 110.185 156.030 ;
        RECT 110.800 155.970 111.120 156.030 ;
        RECT 113.100 155.970 113.420 156.030 ;
        RECT 113.560 155.970 113.880 156.230 ;
        RECT 114.480 156.170 114.800 156.230 ;
        RECT 116.335 156.170 116.625 156.215 ;
        RECT 114.480 156.030 116.625 156.170 ;
        RECT 114.480 155.970 114.800 156.030 ;
        RECT 116.335 155.985 116.625 156.030 ;
        RECT 118.620 156.170 118.940 156.230 ;
        RECT 119.555 156.170 119.845 156.215 ;
        RECT 118.620 156.030 119.845 156.170 ;
        RECT 118.620 155.970 118.940 156.030 ;
        RECT 119.555 155.985 119.845 156.030 ;
        RECT 123.220 155.970 123.540 156.230 ;
        RECT 133.800 156.170 134.120 156.230 ;
        RECT 139.795 156.170 140.085 156.215 ;
        RECT 133.800 156.030 140.085 156.170 ;
        RECT 133.800 155.970 134.120 156.030 ;
        RECT 139.795 155.985 140.085 156.030 ;
        RECT 142.540 155.970 142.860 156.230 ;
        RECT 143.000 155.970 143.320 156.230 ;
        RECT 70.710 155.350 156.270 155.830 ;
        RECT 87.340 155.150 87.660 155.210 ;
        RECT 89.640 155.150 89.960 155.210 ;
        RECT 87.340 155.010 89.960 155.150 ;
        RECT 87.340 154.950 87.660 155.010 ;
        RECT 89.640 154.950 89.960 155.010 ;
        RECT 97.920 155.150 98.240 155.210 ;
        RECT 113.100 155.150 113.420 155.210 ;
        RECT 97.920 155.010 113.420 155.150 ;
        RECT 97.920 154.950 98.240 155.010 ;
        RECT 85.500 154.810 85.820 154.870 ;
        RECT 88.720 154.810 89.040 154.870 ;
        RECT 94.240 154.810 94.560 154.870 ;
        RECT 102.980 154.810 103.300 154.870 ;
        RECT 85.500 154.670 88.490 154.810 ;
        RECT 85.500 154.610 85.820 154.670 ;
        RECT 73.510 154.470 73.800 154.515 ;
        RECT 77.220 154.470 77.540 154.530 ;
        RECT 80.440 154.470 80.760 154.530 ;
        RECT 86.050 154.515 86.190 154.670 ;
        RECT 81.375 154.470 81.665 154.515 ;
        RECT 73.510 154.330 77.540 154.470 ;
        RECT 73.510 154.285 73.800 154.330 ;
        RECT 77.220 154.270 77.540 154.330 ;
        RECT 79.150 154.330 81.665 154.470 ;
        RECT 72.160 153.930 72.480 154.190 ;
        RECT 73.055 154.130 73.345 154.175 ;
        RECT 74.245 154.130 74.535 154.175 ;
        RECT 76.765 154.130 77.055 154.175 ;
        RECT 73.055 153.990 77.055 154.130 ;
        RECT 73.055 153.945 73.345 153.990 ;
        RECT 74.245 153.945 74.535 153.990 ;
        RECT 76.765 153.945 77.055 153.990 ;
        RECT 79.150 153.835 79.290 154.330 ;
        RECT 80.440 154.270 80.760 154.330 ;
        RECT 81.375 154.285 81.665 154.330 ;
        RECT 85.975 154.285 86.265 154.515 ;
        RECT 86.895 154.470 87.185 154.515 ;
        RECT 87.340 154.470 87.660 154.530 ;
        RECT 86.895 154.330 87.660 154.470 ;
        RECT 86.895 154.285 87.185 154.330 ;
        RECT 87.340 154.270 87.660 154.330 ;
        RECT 87.815 154.285 88.105 154.515 ;
        RECT 88.350 154.470 88.490 154.670 ;
        RECT 88.720 154.670 91.710 154.810 ;
        RECT 88.720 154.610 89.040 154.670 ;
        RECT 89.195 154.470 89.485 154.515 ;
        RECT 88.350 154.330 89.485 154.470 ;
        RECT 89.195 154.285 89.485 154.330 ;
        RECT 87.890 154.130 88.030 154.285 ;
        RECT 89.640 154.270 89.960 154.530 ;
        RECT 91.570 154.515 91.710 154.670 ;
        RECT 94.240 154.670 103.300 154.810 ;
        RECT 94.240 154.610 94.560 154.670 ;
        RECT 102.980 154.610 103.300 154.670 ;
        RECT 103.900 154.810 104.220 154.870 ;
        RECT 108.500 154.810 108.820 154.870 ;
        RECT 103.900 154.670 109.190 154.810 ;
        RECT 103.900 154.610 104.220 154.670 ;
        RECT 108.500 154.610 108.820 154.670 ;
        RECT 91.495 154.285 91.785 154.515 ;
        RECT 92.415 154.285 92.705 154.515 ;
        RECT 104.360 154.470 104.680 154.530 ;
        RECT 104.360 154.330 106.890 154.470 ;
        RECT 92.490 154.130 92.630 154.285 ;
        RECT 104.360 154.270 104.680 154.330 ;
        RECT 106.750 154.190 106.890 154.330 ;
        RECT 107.135 154.285 107.425 154.515 ;
        RECT 108.055 154.285 108.345 154.515 ;
        RECT 109.050 154.470 109.190 154.670 ;
        RECT 109.970 154.515 110.110 155.010 ;
        RECT 113.100 154.950 113.420 155.010 ;
        RECT 122.760 155.150 123.080 155.210 ;
        RECT 143.920 155.150 144.240 155.210 ;
        RECT 144.840 155.150 145.160 155.210 ;
        RECT 122.760 155.010 145.160 155.150 ;
        RECT 122.760 154.950 123.080 155.010 ;
        RECT 143.920 154.950 144.240 155.010 ;
        RECT 144.840 154.950 145.160 155.010 ;
        RECT 110.800 154.810 111.120 154.870 ;
        RECT 115.400 154.810 115.720 154.870 ;
        RECT 127.360 154.810 127.680 154.870 ;
        RECT 110.800 154.670 115.720 154.810 ;
        RECT 110.800 154.610 111.120 154.670 ;
        RECT 115.400 154.610 115.720 154.670 ;
        RECT 118.250 154.670 121.150 154.810 ;
        RECT 118.250 154.530 118.390 154.670 ;
        RECT 108.590 154.330 109.190 154.470 ;
        RECT 87.890 153.990 89.410 154.130 ;
        RECT 72.660 153.790 72.950 153.835 ;
        RECT 74.760 153.790 75.050 153.835 ;
        RECT 76.330 153.790 76.620 153.835 ;
        RECT 72.660 153.650 76.620 153.790 ;
        RECT 72.660 153.605 72.950 153.650 ;
        RECT 74.760 153.605 75.050 153.650 ;
        RECT 76.330 153.605 76.620 153.650 ;
        RECT 79.075 153.605 79.365 153.835 ;
        RECT 87.815 153.790 88.105 153.835 ;
        RECT 88.260 153.790 88.580 153.850 ;
        RECT 87.815 153.650 88.580 153.790 ;
        RECT 87.815 153.605 88.105 153.650 ;
        RECT 88.260 153.590 88.580 153.650 ;
        RECT 89.270 153.790 89.410 153.990 ;
        RECT 90.650 153.990 92.630 154.130 ;
        RECT 90.650 153.790 90.790 153.990 ;
        RECT 102.980 153.930 103.300 154.190 ;
        RECT 103.440 153.930 103.760 154.190 ;
        RECT 103.915 154.130 104.205 154.175 ;
        RECT 105.280 154.130 105.600 154.190 ;
        RECT 103.915 153.990 105.600 154.130 ;
        RECT 103.915 153.945 104.205 153.990 ;
        RECT 105.280 153.930 105.600 153.990 ;
        RECT 106.660 153.930 106.980 154.190 ;
        RECT 107.210 154.130 107.350 154.285 ;
        RECT 107.580 154.130 107.900 154.190 ;
        RECT 107.210 153.990 107.900 154.130 ;
        RECT 89.270 153.650 90.790 153.790 ;
        RECT 91.035 153.790 91.325 153.835 ;
        RECT 91.940 153.790 92.260 153.850 ;
        RECT 107.210 153.790 107.350 153.990 ;
        RECT 107.580 153.930 107.900 153.990 ;
        RECT 91.035 153.650 92.260 153.790 ;
        RECT 89.270 153.510 89.410 153.650 ;
        RECT 91.035 153.605 91.325 153.650 ;
        RECT 91.940 153.590 92.260 153.650 ;
        RECT 100.770 153.650 107.350 153.790 ;
        RECT 100.770 153.510 100.910 153.650 ;
        RECT 82.295 153.450 82.585 153.495 ;
        RECT 85.960 153.450 86.280 153.510 ;
        RECT 82.295 153.310 86.280 153.450 ;
        RECT 82.295 153.265 82.585 153.310 ;
        RECT 85.960 153.250 86.280 153.310 ;
        RECT 89.180 153.250 89.500 153.510 ;
        RECT 89.640 153.450 89.960 153.510 ;
        RECT 91.495 153.450 91.785 153.495 ;
        RECT 89.640 153.310 91.785 153.450 ;
        RECT 89.640 153.250 89.960 153.310 ;
        RECT 91.495 153.265 91.785 153.310 ;
        RECT 100.680 153.250 101.000 153.510 ;
        RECT 105.295 153.450 105.585 153.495 ;
        RECT 107.580 153.450 107.900 153.510 ;
        RECT 105.295 153.310 107.900 153.450 ;
        RECT 108.130 153.450 108.270 154.285 ;
        RECT 108.590 154.175 108.730 154.330 ;
        RECT 109.895 154.285 110.185 154.515 ;
        RECT 113.560 154.470 113.880 154.530 ;
        RECT 116.795 154.470 117.085 154.515 ;
        RECT 113.560 154.330 117.085 154.470 ;
        RECT 113.560 154.270 113.880 154.330 ;
        RECT 116.795 154.285 117.085 154.330 ;
        RECT 118.160 154.270 118.480 154.530 ;
        RECT 118.620 154.270 118.940 154.530 ;
        RECT 121.010 154.515 121.150 154.670 ;
        RECT 123.770 154.670 127.680 154.810 ;
        RECT 120.935 154.285 121.225 154.515 ;
        RECT 122.760 154.270 123.080 154.530 ;
        RECT 123.770 154.515 123.910 154.670 ;
        RECT 127.360 154.610 127.680 154.670 ;
        RECT 134.260 154.610 134.580 154.870 ;
        RECT 138.400 154.810 138.720 154.870 ;
        RECT 139.780 154.810 140.100 154.870 ;
        RECT 138.400 154.670 140.100 154.810 ;
        RECT 138.400 154.610 138.720 154.670 ;
        RECT 139.780 154.610 140.100 154.670 ;
        RECT 141.160 154.610 141.480 154.870 ;
        RECT 148.980 154.810 149.300 154.870 ;
        RECT 150.360 154.810 150.680 154.870 ;
        RECT 150.835 154.810 151.125 154.855 ;
        RECT 148.980 154.670 151.125 154.810 ;
        RECT 148.980 154.610 149.300 154.670 ;
        RECT 150.360 154.610 150.680 154.670 ;
        RECT 150.835 154.625 151.125 154.670 ;
        RECT 124.600 154.515 124.920 154.530 ;
        RECT 123.695 154.285 123.985 154.515 ;
        RECT 124.385 154.285 124.920 154.515 ;
        RECT 125.535 154.285 125.825 154.515 ;
        RECT 126.455 154.285 126.745 154.515 ;
        RECT 134.350 154.470 134.490 154.610 ;
        RECT 137.035 154.470 137.325 154.515 ;
        RECT 134.350 154.330 137.325 154.470 ;
        RECT 137.035 154.285 137.325 154.330 ;
        RECT 124.600 154.270 124.920 154.285 ;
        RECT 108.515 153.945 108.805 154.175 ;
        RECT 108.975 153.945 109.265 154.175 ;
        RECT 109.050 153.790 109.190 153.945 ;
        RECT 110.800 153.930 111.120 154.190 ;
        RECT 114.020 154.130 114.340 154.190 ;
        RECT 114.955 154.130 115.245 154.175 ;
        RECT 115.400 154.130 115.720 154.190 ;
        RECT 114.020 153.990 115.720 154.130 ;
        RECT 114.020 153.930 114.340 153.990 ;
        RECT 114.955 153.945 115.245 153.990 ;
        RECT 115.400 153.930 115.720 153.990 ;
        RECT 116.335 154.130 116.625 154.175 ;
        RECT 118.710 154.130 118.850 154.270 ;
        RECT 116.335 153.990 118.850 154.130 ;
        RECT 119.095 154.130 119.385 154.175 ;
        RECT 119.540 154.130 119.860 154.190 ;
        RECT 119.095 153.990 119.860 154.130 ;
        RECT 116.335 153.945 116.625 153.990 ;
        RECT 119.095 153.945 119.385 153.990 ;
        RECT 119.540 153.930 119.860 153.990 ;
        RECT 120.000 153.930 120.320 154.190 ;
        RECT 120.460 153.930 120.780 154.190 ;
        RECT 121.395 154.130 121.685 154.175 ;
        RECT 123.220 154.130 123.540 154.190 ;
        RECT 121.395 153.990 123.540 154.130 ;
        RECT 121.395 153.945 121.685 153.990 ;
        RECT 123.220 153.930 123.540 153.990 ;
        RECT 125.060 153.930 125.380 154.190 ;
        RECT 116.780 153.790 117.100 153.850 ;
        RECT 109.050 153.650 117.100 153.790 ;
        RECT 116.780 153.590 117.100 153.650 ;
        RECT 110.340 153.450 110.660 153.510 ;
        RECT 117.715 153.450 118.005 153.495 ;
        RECT 125.610 153.450 125.750 154.285 ;
        RECT 126.530 153.850 126.670 154.285 ;
        RECT 141.250 154.130 141.390 154.610 ;
        RECT 147.600 154.470 147.920 154.530 ;
        RECT 148.520 154.470 148.840 154.530 ;
        RECT 149.915 154.470 150.205 154.515 ;
        RECT 147.600 154.330 150.205 154.470 ;
        RECT 147.600 154.270 147.920 154.330 ;
        RECT 148.520 154.270 148.840 154.330 ;
        RECT 149.915 154.285 150.205 154.330 ;
        RECT 138.030 153.990 141.390 154.130 ;
        RECT 142.540 154.130 142.860 154.190 ;
        RECT 148.995 154.130 149.285 154.175 ;
        RECT 142.540 153.990 149.285 154.130 ;
        RECT 126.440 153.590 126.760 153.850 ;
        RECT 138.030 153.835 138.170 153.990 ;
        RECT 142.540 153.930 142.860 153.990 ;
        RECT 148.995 153.945 149.285 153.990 ;
        RECT 137.955 153.605 138.245 153.835 ;
        RECT 139.780 153.790 140.100 153.850 ;
        RECT 142.080 153.790 142.400 153.850 ;
        RECT 139.780 153.650 142.400 153.790 ;
        RECT 139.780 153.590 140.100 153.650 ;
        RECT 142.080 153.590 142.400 153.650 ;
        RECT 128.740 153.450 129.060 153.510 ;
        RECT 108.130 153.310 129.060 153.450 ;
        RECT 105.295 153.265 105.585 153.310 ;
        RECT 107.580 153.250 107.900 153.310 ;
        RECT 110.340 153.250 110.660 153.310 ;
        RECT 117.715 153.265 118.005 153.310 ;
        RECT 128.740 153.250 129.060 153.310 ;
        RECT 130.580 153.450 130.900 153.510 ;
        RECT 133.340 153.450 133.660 153.510 ;
        RECT 130.580 153.310 133.660 153.450 ;
        RECT 130.580 153.250 130.900 153.310 ;
        RECT 133.340 153.250 133.660 153.310 ;
        RECT 70.710 152.630 156.270 153.110 ;
        RECT 86.420 152.430 86.740 152.490 ;
        RECT 100.220 152.430 100.540 152.490 ;
        RECT 86.420 152.290 100.540 152.430 ;
        RECT 86.420 152.230 86.740 152.290 ;
        RECT 100.220 152.230 100.540 152.290 ;
        RECT 102.980 152.430 103.300 152.490 ;
        RECT 109.895 152.430 110.185 152.475 ;
        RECT 102.980 152.290 110.185 152.430 ;
        RECT 102.980 152.230 103.300 152.290 ;
        RECT 109.895 152.245 110.185 152.290 ;
        RECT 110.800 152.230 111.120 152.490 ;
        RECT 111.735 152.245 112.025 152.475 ;
        RECT 97.000 152.090 97.320 152.150 ;
        RECT 99.300 152.090 99.620 152.150 ;
        RECT 107.135 152.090 107.425 152.135 ;
        RECT 97.000 151.950 98.610 152.090 ;
        RECT 97.000 151.890 97.320 151.950 ;
        RECT 98.470 151.795 98.610 151.950 ;
        RECT 99.300 151.950 107.425 152.090 ;
        RECT 99.300 151.890 99.620 151.950 ;
        RECT 107.135 151.905 107.425 151.950 ;
        RECT 98.395 151.565 98.685 151.795 ;
        RECT 102.060 151.750 102.380 151.810 ;
        RECT 99.390 151.610 102.380 151.750 ;
        RECT 80.900 151.410 81.220 151.470 ;
        RECT 81.835 151.410 82.125 151.455 ;
        RECT 79.150 151.270 82.125 151.410 ;
        RECT 79.150 151.130 79.290 151.270 ;
        RECT 80.900 151.210 81.220 151.270 ;
        RECT 81.835 151.225 82.125 151.270 ;
        RECT 97.935 151.410 98.225 151.455 ;
        RECT 99.390 151.410 99.530 151.610 ;
        RECT 102.060 151.550 102.380 151.610 ;
        RECT 103.440 151.750 103.760 151.810 ;
        RECT 105.295 151.750 105.585 151.795 ;
        RECT 103.440 151.610 105.585 151.750 ;
        RECT 103.440 151.550 103.760 151.610 ;
        RECT 105.295 151.565 105.585 151.610 ;
        RECT 106.290 151.610 108.730 151.750 ;
        RECT 103.900 151.410 104.220 151.470 ;
        RECT 97.935 151.270 99.530 151.410 ;
        RECT 99.850 151.270 104.220 151.410 ;
        RECT 97.935 151.225 98.225 151.270 ;
        RECT 79.060 150.870 79.380 151.130 ;
        RECT 99.850 151.070 99.990 151.270 ;
        RECT 103.900 151.210 104.220 151.270 ;
        RECT 104.820 151.210 105.140 151.470 ;
        RECT 105.755 151.410 106.045 151.455 ;
        RECT 106.290 151.410 106.430 151.610 ;
        RECT 108.590 151.470 108.730 151.610 ;
        RECT 105.755 151.270 106.430 151.410 ;
        RECT 105.755 151.225 106.045 151.270 ;
        RECT 80.070 150.930 99.990 151.070 ;
        RECT 78.140 150.730 78.460 150.790 ;
        RECT 80.070 150.730 80.210 150.930 ;
        RECT 102.980 150.870 103.300 151.130 ;
        RECT 106.290 151.070 106.430 151.270 ;
        RECT 106.675 151.225 106.965 151.455 ;
        RECT 108.055 151.225 108.345 151.455 ;
        RECT 103.530 150.930 106.430 151.070 ;
        RECT 78.140 150.590 80.210 150.730 ;
        RECT 80.440 150.730 80.760 150.790 ;
        RECT 80.915 150.730 81.205 150.775 ;
        RECT 80.440 150.590 81.205 150.730 ;
        RECT 78.140 150.530 78.460 150.590 ;
        RECT 80.440 150.530 80.760 150.590 ;
        RECT 80.915 150.545 81.205 150.590 ;
        RECT 96.540 150.730 96.860 150.790 ;
        RECT 98.840 150.730 99.160 150.790 ;
        RECT 96.540 150.590 99.160 150.730 ;
        RECT 96.540 150.530 96.860 150.590 ;
        RECT 98.840 150.530 99.160 150.590 ;
        RECT 99.545 150.730 99.835 150.775 ;
        RECT 103.530 150.730 103.670 150.930 ;
        RECT 99.545 150.590 103.670 150.730 ;
        RECT 103.900 150.730 104.220 150.790 ;
        RECT 106.750 150.730 106.890 151.225 ;
        RECT 108.130 151.070 108.270 151.225 ;
        RECT 108.500 151.210 108.820 151.470 ;
        RECT 110.890 151.455 111.030 152.230 ;
        RECT 111.810 152.090 111.950 152.245 ;
        RECT 113.560 152.230 113.880 152.490 ;
        RECT 114.940 152.230 115.260 152.490 ;
        RECT 116.780 152.230 117.100 152.490 ;
        RECT 123.220 152.230 123.540 152.490 ;
        RECT 124.140 152.430 124.460 152.490 ;
        RECT 125.075 152.430 125.365 152.475 ;
        RECT 129.200 152.430 129.520 152.490 ;
        RECT 140.255 152.430 140.545 152.475 ;
        RECT 145.760 152.430 146.080 152.490 ;
        RECT 124.140 152.290 125.365 152.430 ;
        RECT 124.140 152.230 124.460 152.290 ;
        RECT 125.075 152.245 125.365 152.290 ;
        RECT 125.750 152.290 129.520 152.430 ;
        RECT 112.640 152.090 112.960 152.150 ;
        RECT 115.030 152.090 115.170 152.230 ;
        RECT 111.810 151.950 115.170 152.090 ;
        RECT 116.870 152.090 117.010 152.230 ;
        RECT 124.600 152.090 124.920 152.150 ;
        RECT 125.750 152.090 125.890 152.290 ;
        RECT 129.200 152.230 129.520 152.290 ;
        RECT 132.970 152.290 137.250 152.430 ;
        RECT 132.970 152.090 133.110 152.290 ;
        RECT 116.870 151.950 125.890 152.090 ;
        RECT 126.070 151.950 133.110 152.090 ;
        RECT 137.110 152.090 137.250 152.290 ;
        RECT 140.255 152.290 146.080 152.430 ;
        RECT 140.255 152.245 140.545 152.290 ;
        RECT 145.760 152.230 146.080 152.290 ;
        RECT 147.140 152.430 147.460 152.490 ;
        RECT 148.980 152.430 149.300 152.490 ;
        RECT 147.140 152.290 149.300 152.430 ;
        RECT 147.140 152.230 147.460 152.290 ;
        RECT 148.980 152.230 149.300 152.290 ;
        RECT 149.915 152.090 150.205 152.135 ;
        RECT 137.110 151.950 150.205 152.090 ;
        RECT 112.640 151.890 112.960 151.950 ;
        RECT 124.600 151.890 124.920 151.950 ;
        RECT 112.195 151.750 112.485 151.795 ;
        RECT 125.060 151.750 125.380 151.810 ;
        RECT 125.535 151.750 125.825 151.795 ;
        RECT 112.195 151.610 125.825 151.750 ;
        RECT 112.195 151.565 112.485 151.610 ;
        RECT 110.815 151.225 111.105 151.455 ;
        RECT 111.260 151.410 111.580 151.470 ;
        RECT 112.270 151.410 112.410 151.565 ;
        RECT 125.060 151.550 125.380 151.610 ;
        RECT 125.535 151.565 125.825 151.610 ;
        RECT 111.260 151.270 112.410 151.410 ;
        RECT 111.260 151.210 111.580 151.270 ;
        RECT 112.655 151.225 112.945 151.455 ;
        RECT 117.700 151.410 118.020 151.470 ;
        RECT 119.540 151.410 119.860 151.470 ;
        RECT 117.700 151.270 119.860 151.410 ;
        RECT 112.730 151.070 112.870 151.225 ;
        RECT 117.700 151.210 118.020 151.270 ;
        RECT 119.540 151.210 119.860 151.270 ;
        RECT 122.760 151.410 123.080 151.470 ;
        RECT 124.155 151.410 124.445 151.455 ;
        RECT 122.760 151.270 124.445 151.410 ;
        RECT 122.760 151.210 123.080 151.270 ;
        RECT 124.155 151.225 124.445 151.270 ;
        RECT 126.070 151.070 126.210 151.950 ;
        RECT 149.915 151.905 150.205 151.950 ;
        RECT 128.370 151.610 135.870 151.750 ;
        RECT 126.900 151.410 127.220 151.470 ;
        RECT 127.375 151.410 127.665 151.455 ;
        RECT 126.900 151.270 127.665 151.410 ;
        RECT 126.900 151.210 127.220 151.270 ;
        RECT 127.375 151.225 127.665 151.270 ;
        RECT 108.130 150.930 126.210 151.070 ;
        RECT 103.900 150.590 106.890 150.730 ;
        RECT 108.040 150.730 108.360 150.790 ;
        RECT 126.440 150.730 126.760 150.790 ;
        RECT 128.370 150.775 128.510 151.610 ;
        RECT 129.200 151.410 129.520 151.470 ;
        RECT 131.960 151.410 132.280 151.470 ;
        RECT 135.730 151.455 135.870 151.610 ;
        RECT 137.020 151.550 137.340 151.810 ;
        RECT 139.335 151.750 139.625 151.795 ;
        RECT 142.080 151.750 142.400 151.810 ;
        RECT 143.475 151.750 143.765 151.795 ;
        RECT 151.295 151.750 151.585 151.795 ;
        RECT 139.335 151.610 141.390 151.750 ;
        RECT 139.335 151.565 139.625 151.610 ;
        RECT 129.200 151.270 132.280 151.410 ;
        RECT 129.200 151.210 129.520 151.270 ;
        RECT 131.960 151.210 132.280 151.270 ;
        RECT 135.655 151.225 135.945 151.455 ;
        RECT 136.575 151.225 136.865 151.455 ;
        RECT 137.495 151.410 137.785 151.455 ;
        RECT 137.495 151.270 138.170 151.410 ;
        RECT 137.495 151.225 137.785 151.270 ;
        RECT 128.740 151.070 129.060 151.130 ;
        RECT 136.650 151.070 136.790 151.225 ;
        RECT 128.740 150.930 136.790 151.070 ;
        RECT 128.740 150.870 129.060 150.930 ;
        RECT 128.295 150.730 128.585 150.775 ;
        RECT 108.040 150.590 128.585 150.730 ;
        RECT 99.545 150.545 99.835 150.590 ;
        RECT 103.900 150.530 104.220 150.590 ;
        RECT 108.040 150.530 108.360 150.590 ;
        RECT 126.440 150.530 126.760 150.590 ;
        RECT 128.295 150.545 128.585 150.590 ;
        RECT 129.200 150.730 129.520 150.790 ;
        RECT 131.055 150.730 131.345 150.775 ;
        RECT 138.030 150.730 138.170 151.270 ;
        RECT 138.415 151.225 138.705 151.455 ;
        RECT 138.860 151.410 139.180 151.470 ;
        RECT 139.795 151.410 140.085 151.455 ;
        RECT 138.860 151.270 140.085 151.410 ;
        RECT 138.490 151.070 138.630 151.225 ;
        RECT 138.860 151.210 139.180 151.270 ;
        RECT 139.795 151.225 140.085 151.270 ;
        RECT 140.700 151.210 141.020 151.470 ;
        RECT 141.250 151.455 141.390 151.610 ;
        RECT 142.080 151.610 143.765 151.750 ;
        RECT 142.080 151.550 142.400 151.610 ;
        RECT 143.475 151.565 143.765 151.610 ;
        RECT 144.470 151.610 151.585 151.750 ;
        RECT 141.175 151.225 141.465 151.455 ;
        RECT 140.790 151.070 140.930 151.210 ;
        RECT 138.490 150.930 140.930 151.070 ;
        RECT 143.920 151.070 144.240 151.130 ;
        RECT 144.470 151.070 144.610 151.610 ;
        RECT 144.855 151.225 145.145 151.455 ;
        RECT 145.760 151.410 146.080 151.470 ;
        RECT 148.075 151.410 148.365 151.455 ;
        RECT 145.760 151.270 148.365 151.410 ;
        RECT 143.920 150.930 144.610 151.070 ;
        RECT 144.930 151.070 145.070 151.225 ;
        RECT 145.760 151.210 146.080 151.270 ;
        RECT 148.075 151.225 148.365 151.270 ;
        RECT 148.520 151.410 148.840 151.470 ;
        RECT 150.450 151.455 150.590 151.610 ;
        RECT 151.295 151.565 151.585 151.610 ;
        RECT 148.995 151.410 149.285 151.455 ;
        RECT 149.455 151.410 149.745 151.455 ;
        RECT 148.520 151.270 149.745 151.410 ;
        RECT 148.520 151.210 148.840 151.270 ;
        RECT 148.995 151.225 149.285 151.270 ;
        RECT 149.455 151.225 149.745 151.270 ;
        RECT 150.375 151.225 150.665 151.455 ;
        RECT 150.820 151.210 151.140 151.470 ;
        RECT 153.135 151.410 153.425 151.455 ;
        RECT 154.040 151.410 154.360 151.470 ;
        RECT 153.135 151.270 154.360 151.410 ;
        RECT 153.135 151.225 153.425 151.270 ;
        RECT 154.040 151.210 154.360 151.270 ;
        RECT 144.930 150.930 145.990 151.070 ;
        RECT 143.920 150.870 144.240 150.930 ;
        RECT 145.850 150.790 145.990 150.930 ;
        RECT 129.200 150.590 138.170 150.730 ;
        RECT 129.200 150.530 129.520 150.590 ;
        RECT 131.055 150.545 131.345 150.590 ;
        RECT 142.080 150.530 142.400 150.790 ;
        RECT 145.760 150.530 146.080 150.790 ;
        RECT 148.520 150.530 148.840 150.790 ;
        RECT 152.200 150.530 152.520 150.790 ;
        RECT 70.710 149.910 156.270 150.390 ;
        RECT 77.220 149.710 77.540 149.770 ;
        RECT 80.915 149.710 81.205 149.755 ;
        RECT 77.220 149.570 81.205 149.710 ;
        RECT 77.220 149.510 77.540 149.570 ;
        RECT 80.915 149.525 81.205 149.570 ;
        RECT 82.295 149.710 82.585 149.755 ;
        RECT 84.580 149.710 84.900 149.770 ;
        RECT 82.295 149.570 84.900 149.710 ;
        RECT 82.295 149.525 82.585 149.570 ;
        RECT 84.580 149.510 84.900 149.570 ;
        RECT 87.800 149.710 88.120 149.770 ;
        RECT 89.425 149.710 89.715 149.755 ;
        RECT 103.440 149.710 103.760 149.770 ;
        RECT 104.360 149.710 104.680 149.770 ;
        RECT 87.800 149.570 99.530 149.710 ;
        RECT 87.800 149.510 88.120 149.570 ;
        RECT 89.425 149.525 89.715 149.570 ;
        RECT 86.435 149.370 86.725 149.415 ;
        RECT 96.080 149.370 96.400 149.430 ;
        RECT 99.390 149.370 99.530 149.570 ;
        RECT 103.440 149.570 104.680 149.710 ;
        RECT 103.440 149.510 103.760 149.570 ;
        RECT 104.360 149.510 104.680 149.570 ;
        RECT 104.820 149.710 105.140 149.770 ;
        RECT 109.880 149.710 110.200 149.770 ;
        RECT 145.760 149.710 146.080 149.770 ;
        RECT 104.820 149.570 146.080 149.710 ;
        RECT 104.820 149.510 105.140 149.570 ;
        RECT 109.880 149.510 110.200 149.570 ;
        RECT 145.760 149.510 146.080 149.570 ;
        RECT 148.060 149.510 148.380 149.770 ;
        RECT 148.520 149.510 148.840 149.770 ;
        RECT 148.980 149.710 149.300 149.770 ;
        RECT 148.980 149.570 149.750 149.710 ;
        RECT 148.980 149.510 149.300 149.570 ;
        RECT 117.255 149.370 117.545 149.415 ;
        RECT 143.920 149.370 144.240 149.430 ;
        RECT 81.450 149.230 86.725 149.370 ;
        RECT 81.450 149.075 81.590 149.230 ;
        RECT 86.435 149.185 86.725 149.230 ;
        RECT 87.430 149.230 88.490 149.370 ;
        RECT 73.510 149.030 73.800 149.075 ;
        RECT 73.510 148.890 78.370 149.030 ;
        RECT 73.510 148.845 73.800 148.890 ;
        RECT 72.160 148.490 72.480 148.750 ;
        RECT 73.055 148.690 73.345 148.735 ;
        RECT 74.245 148.690 74.535 148.735 ;
        RECT 76.765 148.690 77.055 148.735 ;
        RECT 73.055 148.550 77.055 148.690 ;
        RECT 73.055 148.505 73.345 148.550 ;
        RECT 74.245 148.505 74.535 148.550 ;
        RECT 76.765 148.505 77.055 148.550 ;
        RECT 72.660 148.350 72.950 148.395 ;
        RECT 74.760 148.350 75.050 148.395 ;
        RECT 76.330 148.350 76.620 148.395 ;
        RECT 72.660 148.210 76.620 148.350 ;
        RECT 78.230 148.350 78.370 148.890 ;
        RECT 80.455 148.845 80.745 149.075 ;
        RECT 81.375 148.845 81.665 149.075 ;
        RECT 81.835 149.030 82.125 149.075 ;
        RECT 81.835 148.890 82.235 149.030 ;
        RECT 81.835 148.845 82.125 148.890 ;
        RECT 79.980 148.690 80.300 148.750 ;
        RECT 80.530 148.690 80.670 148.845 ;
        RECT 81.910 148.690 82.050 148.845 ;
        RECT 83.200 148.830 83.520 149.090 ;
        RECT 85.055 148.845 85.345 149.075 ;
        RECT 85.960 149.030 86.280 149.090 ;
        RECT 87.430 149.030 87.570 149.230 ;
        RECT 85.960 148.890 87.570 149.030 ;
        RECT 79.980 148.550 84.350 148.690 ;
        RECT 79.980 148.490 80.300 148.550 ;
        RECT 83.215 148.350 83.505 148.395 ;
        RECT 78.230 148.210 83.505 148.350 ;
        RECT 72.660 148.165 72.950 148.210 ;
        RECT 74.760 148.165 75.050 148.210 ;
        RECT 76.330 148.165 76.620 148.210 ;
        RECT 83.215 148.165 83.505 148.210 ;
        RECT 84.210 148.070 84.350 148.550 ;
        RECT 85.130 148.350 85.270 148.845 ;
        RECT 85.960 148.830 86.280 148.890 ;
        RECT 87.800 148.830 88.120 149.090 ;
        RECT 85.500 148.690 85.820 148.750 ;
        RECT 86.420 148.690 86.740 148.750 ;
        RECT 88.350 148.735 88.490 149.230 ;
        RECT 96.080 149.230 98.610 149.370 ;
        RECT 99.390 149.230 116.090 149.370 ;
        RECT 96.080 149.170 96.400 149.230 ;
        RECT 97.935 148.845 98.225 149.075 ;
        RECT 98.470 149.030 98.610 149.230 ;
        RECT 115.950 149.090 116.090 149.230 ;
        RECT 117.255 149.230 119.770 149.370 ;
        RECT 117.255 149.185 117.545 149.230 ;
        RECT 99.315 149.030 99.605 149.075 ;
        RECT 98.470 148.890 99.605 149.030 ;
        RECT 99.315 148.845 99.605 148.890 ;
        RECT 85.500 148.550 86.740 148.690 ;
        RECT 85.500 148.490 85.820 148.550 ;
        RECT 86.420 148.490 86.740 148.550 ;
        RECT 87.355 148.505 87.645 148.735 ;
        RECT 88.275 148.690 88.565 148.735 ;
        RECT 92.400 148.690 92.720 148.750 ;
        RECT 95.620 148.690 95.940 148.750 ;
        RECT 88.275 148.550 95.940 148.690 ;
        RECT 88.275 148.505 88.565 148.550 ;
        RECT 85.960 148.350 86.280 148.410 ;
        RECT 87.430 148.350 87.570 148.505 ;
        RECT 92.400 148.490 92.720 148.550 ;
        RECT 95.620 148.490 95.940 148.550 ;
        RECT 94.240 148.350 94.560 148.410 ;
        RECT 85.130 148.210 94.560 148.350 ;
        RECT 98.010 148.350 98.150 148.845 ;
        RECT 99.760 148.830 100.080 149.090 ;
        RECT 100.680 148.830 101.000 149.090 ;
        RECT 102.980 149.030 103.300 149.090 ;
        RECT 103.455 149.030 103.745 149.075 ;
        RECT 114.955 149.030 115.245 149.075 ;
        RECT 102.980 148.890 103.745 149.030 ;
        RECT 102.980 148.830 103.300 148.890 ;
        RECT 103.455 148.845 103.745 148.890 ;
        RECT 103.990 148.890 115.245 149.030 ;
        RECT 98.840 148.490 99.160 148.750 ;
        RECT 102.060 148.690 102.380 148.750 ;
        RECT 103.990 148.690 104.130 148.890 ;
        RECT 114.955 148.845 115.245 148.890 ;
        RECT 115.860 148.830 116.180 149.090 ;
        RECT 119.630 149.075 119.770 149.230 ;
        RECT 129.750 149.230 135.410 149.370 ;
        RECT 118.175 148.845 118.465 149.075 ;
        RECT 119.555 148.845 119.845 149.075 ;
        RECT 124.600 149.030 124.920 149.090 ;
        RECT 127.835 149.030 128.125 149.075 ;
        RECT 124.600 148.890 128.125 149.030 ;
        RECT 102.060 148.550 104.130 148.690 ;
        RECT 104.360 148.690 104.680 148.750 ;
        RECT 104.835 148.690 105.125 148.735 ;
        RECT 104.360 148.550 105.125 148.690 ;
        RECT 102.060 148.490 102.380 148.550 ;
        RECT 104.360 148.490 104.680 148.550 ;
        RECT 104.835 148.505 105.125 148.550 ;
        RECT 110.800 148.690 111.120 148.750 ;
        RECT 113.575 148.690 113.865 148.735 ;
        RECT 118.250 148.690 118.390 148.845 ;
        RECT 110.800 148.550 118.390 148.690 ;
        RECT 119.630 148.690 119.770 148.845 ;
        RECT 124.600 148.830 124.920 148.890 ;
        RECT 127.835 148.845 128.125 148.890 ;
        RECT 128.755 148.845 129.045 149.075 ;
        RECT 128.830 148.690 128.970 148.845 ;
        RECT 129.200 148.830 129.520 149.090 ;
        RECT 129.750 149.075 129.890 149.230 ;
        RECT 129.675 148.845 129.965 149.075 ;
        RECT 131.960 149.030 132.280 149.090 ;
        RECT 132.435 149.030 132.725 149.075 ;
        RECT 131.960 148.890 132.725 149.030 ;
        RECT 131.960 148.830 132.280 148.890 ;
        RECT 132.435 148.845 132.725 148.890 ;
        RECT 132.895 148.845 133.185 149.075 ;
        RECT 131.515 148.690 131.805 148.735 ;
        RECT 132.970 148.690 133.110 148.845 ;
        RECT 134.260 148.830 134.580 149.090 ;
        RECT 119.630 148.550 127.130 148.690 ;
        RECT 128.830 148.550 131.805 148.690 ;
        RECT 110.800 148.490 111.120 148.550 ;
        RECT 113.575 148.505 113.865 148.550 ;
        RECT 115.030 148.410 115.170 148.550 ;
        RECT 126.990 148.410 127.130 148.550 ;
        RECT 131.515 148.505 131.805 148.550 ;
        RECT 132.050 148.550 133.110 148.690 ;
        RECT 135.270 148.690 135.410 149.230 ;
        RECT 135.730 149.230 140.930 149.370 ;
        RECT 135.730 149.075 135.870 149.230 ;
        RECT 140.790 149.090 140.930 149.230 ;
        RECT 143.550 149.230 144.240 149.370 ;
        RECT 135.655 148.845 135.945 149.075 ;
        RECT 136.100 148.830 136.420 149.090 ;
        RECT 137.020 149.030 137.340 149.090 ;
        RECT 137.495 149.030 137.785 149.075 ;
        RECT 137.020 148.890 137.785 149.030 ;
        RECT 137.020 148.830 137.340 148.890 ;
        RECT 137.495 148.845 137.785 148.890 ;
        RECT 136.190 148.690 136.330 148.830 ;
        RECT 135.270 148.550 136.330 148.690 ;
        RECT 111.260 148.350 111.580 148.410 ;
        RECT 98.010 148.210 111.580 148.350 ;
        RECT 85.960 148.150 86.280 148.210 ;
        RECT 94.240 148.150 94.560 148.210 ;
        RECT 111.260 148.150 111.580 148.210 ;
        RECT 112.640 148.150 112.960 148.410 ;
        RECT 114.940 148.150 115.260 148.410 ;
        RECT 115.875 148.350 116.165 148.395 ;
        RECT 119.080 148.350 119.400 148.410 ;
        RECT 115.875 148.210 119.400 148.350 ;
        RECT 115.875 148.165 116.165 148.210 ;
        RECT 119.080 148.150 119.400 148.210 ;
        RECT 126.900 148.350 127.220 148.410 ;
        RECT 132.050 148.350 132.190 148.550 ;
        RECT 126.900 148.210 132.190 148.350 ;
        RECT 126.900 148.150 127.220 148.210 ;
        RECT 132.420 148.150 132.740 148.410 ;
        RECT 132.970 148.350 133.110 148.550 ;
        RECT 135.640 148.350 135.960 148.410 ;
        RECT 132.970 148.210 135.960 148.350 ;
        RECT 137.570 148.350 137.710 148.845 ;
        RECT 140.700 148.830 141.020 149.090 ;
        RECT 143.550 149.075 143.690 149.230 ;
        RECT 143.920 149.170 144.240 149.230 ;
        RECT 145.850 149.075 145.990 149.510 ;
        RECT 148.150 149.370 148.290 149.510 ;
        RECT 146.310 149.230 148.290 149.370 ;
        RECT 142.095 149.030 142.385 149.075 ;
        RECT 143.475 149.030 143.765 149.075 ;
        RECT 142.095 148.890 143.765 149.030 ;
        RECT 142.095 148.845 142.385 148.890 ;
        RECT 143.475 148.845 143.765 148.890 ;
        RECT 144.855 148.845 145.145 149.075 ;
        RECT 145.775 148.845 146.065 149.075 ;
        RECT 141.175 148.350 141.465 148.395 ;
        RECT 137.570 148.210 141.465 148.350 ;
        RECT 144.930 148.350 145.070 148.845 ;
        RECT 146.310 148.735 146.450 149.230 ;
        RECT 146.680 148.830 147.000 149.090 ;
        RECT 147.615 149.030 147.905 149.075 ;
        RECT 148.610 149.030 148.750 149.510 ;
        RECT 149.610 149.370 149.750 149.570 ;
        RECT 149.610 149.230 151.510 149.370 ;
        RECT 149.610 149.075 149.750 149.230 ;
        RECT 147.615 148.890 148.750 149.030 ;
        RECT 149.455 148.890 149.750 149.075 ;
        RECT 149.900 149.030 150.220 149.090 ;
        RECT 151.370 149.075 151.510 149.230 ;
        RECT 150.375 149.030 150.665 149.075 ;
        RECT 149.900 148.890 150.665 149.030 ;
        RECT 147.615 148.845 147.905 148.890 ;
        RECT 149.455 148.845 149.745 148.890 ;
        RECT 149.900 148.830 150.220 148.890 ;
        RECT 150.375 148.845 150.665 148.890 ;
        RECT 151.295 148.845 151.585 149.075 ;
        RECT 152.675 148.845 152.965 149.075 ;
        RECT 146.235 148.505 146.525 148.735 ;
        RECT 152.750 148.690 152.890 148.845 ;
        RECT 153.580 148.830 153.900 149.090 ;
        RECT 149.070 148.550 152.890 148.690 ;
        RECT 149.070 148.395 149.210 148.550 ;
        RECT 148.995 148.350 149.285 148.395 ;
        RECT 144.930 148.210 149.285 148.350 ;
        RECT 135.640 148.150 135.960 148.210 ;
        RECT 141.175 148.165 141.465 148.210 ;
        RECT 148.995 148.165 149.285 148.210 ;
        RECT 151.740 148.150 152.060 148.410 ;
        RECT 79.060 147.810 79.380 148.070 ;
        RECT 84.120 147.810 84.440 148.070 ;
        RECT 97.015 148.010 97.305 148.055 ;
        RECT 98.840 148.010 99.160 148.070 ;
        RECT 97.015 147.870 99.160 148.010 ;
        RECT 97.015 147.825 97.305 147.870 ;
        RECT 98.840 147.810 99.160 147.870 ;
        RECT 100.220 148.010 100.540 148.070 ;
        RECT 102.535 148.010 102.825 148.055 ;
        RECT 100.220 147.870 102.825 148.010 ;
        RECT 100.220 147.810 100.540 147.870 ;
        RECT 102.535 147.825 102.825 147.870 ;
        RECT 104.375 148.010 104.665 148.055 ;
        RECT 112.730 148.010 112.870 148.150 ;
        RECT 104.375 147.870 112.870 148.010 ;
        RECT 104.375 147.825 104.665 147.870 ;
        RECT 114.020 147.810 114.340 148.070 ;
        RECT 115.400 148.010 115.720 148.070 ;
        RECT 116.335 148.010 116.625 148.055 ;
        RECT 115.400 147.870 116.625 148.010 ;
        RECT 115.400 147.810 115.720 147.870 ;
        RECT 116.335 147.825 116.625 147.870 ;
        RECT 118.160 148.010 118.480 148.070 ;
        RECT 118.635 148.010 118.925 148.055 ;
        RECT 118.160 147.870 118.925 148.010 ;
        RECT 118.160 147.810 118.480 147.870 ;
        RECT 118.635 147.825 118.925 147.870 ;
        RECT 121.840 148.010 122.160 148.070 ;
        RECT 124.140 148.010 124.460 148.070 ;
        RECT 121.840 147.870 124.460 148.010 ;
        RECT 121.840 147.810 122.160 147.870 ;
        RECT 124.140 147.810 124.460 147.870 ;
        RECT 126.440 148.010 126.760 148.070 ;
        RECT 127.820 148.010 128.140 148.070 ;
        RECT 126.440 147.870 128.140 148.010 ;
        RECT 126.440 147.810 126.760 147.870 ;
        RECT 127.820 147.810 128.140 147.870 ;
        RECT 130.580 148.010 130.900 148.070 ;
        RECT 131.055 148.010 131.345 148.055 ;
        RECT 130.580 147.870 131.345 148.010 ;
        RECT 132.510 148.010 132.650 148.150 ;
        RECT 133.815 148.010 134.105 148.055 ;
        RECT 132.510 147.870 134.105 148.010 ;
        RECT 130.580 147.810 130.900 147.870 ;
        RECT 131.055 147.825 131.345 147.870 ;
        RECT 133.815 147.825 134.105 147.870 ;
        RECT 134.260 148.010 134.580 148.070 ;
        RECT 134.735 148.010 135.025 148.055 ;
        RECT 134.260 147.870 135.025 148.010 ;
        RECT 134.260 147.810 134.580 147.870 ;
        RECT 134.735 147.825 135.025 147.870 ;
        RECT 137.035 148.010 137.325 148.055 ;
        RECT 138.400 148.010 138.720 148.070 ;
        RECT 137.035 147.870 138.720 148.010 ;
        RECT 137.035 147.825 137.325 147.870 ;
        RECT 138.400 147.810 138.720 147.870 ;
        RECT 138.860 148.010 139.180 148.070 ;
        RECT 142.555 148.010 142.845 148.055 ;
        RECT 138.860 147.870 142.845 148.010 ;
        RECT 138.860 147.810 139.180 147.870 ;
        RECT 142.555 147.825 142.845 147.870 ;
        RECT 143.920 147.810 144.240 148.070 ;
        RECT 152.660 147.810 152.980 148.070 ;
        RECT 70.710 147.190 156.270 147.670 ;
        RECT 72.635 146.990 72.925 147.035 ;
        RECT 78.155 146.990 78.445 147.035 ;
        RECT 72.635 146.850 78.445 146.990 ;
        RECT 72.635 146.805 72.925 146.850 ;
        RECT 78.155 146.805 78.445 146.850 ;
        RECT 82.295 146.990 82.585 147.035 ;
        RECT 85.055 146.990 85.345 147.035 ;
        RECT 82.295 146.850 85.345 146.990 ;
        RECT 82.295 146.805 82.585 146.850 ;
        RECT 85.055 146.805 85.345 146.850 ;
        RECT 96.095 146.990 96.385 147.035 ;
        RECT 102.060 146.990 102.380 147.050 ;
        RECT 96.095 146.850 102.380 146.990 ;
        RECT 96.095 146.805 96.385 146.850 ;
        RECT 102.060 146.790 102.380 146.850 ;
        RECT 105.755 146.990 106.045 147.035 ;
        RECT 108.500 146.990 108.820 147.050 ;
        RECT 110.800 146.990 111.120 147.050 ;
        RECT 116.780 146.990 117.100 147.050 ;
        RECT 131.960 146.990 132.280 147.050 ;
        RECT 136.115 146.990 136.405 147.035 ;
        RECT 105.755 146.850 111.120 146.990 ;
        RECT 105.755 146.805 106.045 146.850 ;
        RECT 108.500 146.790 108.820 146.850 ;
        RECT 110.800 146.790 111.120 146.850 ;
        RECT 111.350 146.850 131.730 146.990 ;
        RECT 79.995 146.650 80.285 146.695 ;
        RECT 89.195 146.650 89.485 146.695 ;
        RECT 100.680 146.650 101.000 146.710 ;
        RECT 111.350 146.650 111.490 146.850 ;
        RECT 116.780 146.790 117.100 146.850 ;
        RECT 75.010 146.510 80.285 146.650 ;
        RECT 75.010 146.310 75.150 146.510 ;
        RECT 79.995 146.465 80.285 146.510 ;
        RECT 87.890 146.510 101.000 146.650 ;
        RECT 78.140 146.310 78.460 146.370 ;
        RECT 72.250 146.170 75.150 146.310 ;
        RECT 72.250 146.015 72.390 146.170 ;
        RECT 75.010 146.015 75.150 146.170 ;
        RECT 75.470 146.170 78.460 146.310 ;
        RECT 80.070 146.310 80.210 146.465 ;
        RECT 84.580 146.310 84.900 146.370 ;
        RECT 86.895 146.310 87.185 146.355 ;
        RECT 87.890 146.310 88.030 146.510 ;
        RECT 89.195 146.465 89.485 146.510 ;
        RECT 100.680 146.450 101.000 146.510 ;
        RECT 103.070 146.510 111.490 146.650 ;
        RECT 111.720 146.650 112.040 146.710 ;
        RECT 112.195 146.650 112.485 146.695 ;
        RECT 111.720 146.510 112.485 146.650 ;
        RECT 80.070 146.170 81.590 146.310 ;
        RECT 72.175 145.785 72.465 146.015 ;
        RECT 73.095 145.970 73.385 146.015 ;
        RECT 73.095 145.830 74.230 145.970 ;
        RECT 73.095 145.785 73.385 145.830 ;
        RECT 74.090 145.335 74.230 145.830 ;
        RECT 74.475 145.785 74.765 146.015 ;
        RECT 74.935 145.785 75.225 146.015 ;
        RECT 74.550 145.630 74.690 145.785 ;
        RECT 75.470 145.690 75.610 146.170 ;
        RECT 78.140 146.110 78.460 146.170 ;
        RECT 79.535 145.970 79.825 146.015 ;
        RECT 79.980 145.970 80.300 146.030 ;
        RECT 79.535 145.830 80.300 145.970 ;
        RECT 79.535 145.785 79.825 145.830 ;
        RECT 79.980 145.770 80.300 145.830 ;
        RECT 80.900 145.770 81.220 146.030 ;
        RECT 75.380 145.630 75.700 145.690 ;
        RECT 74.550 145.490 75.700 145.630 ;
        RECT 75.380 145.430 75.700 145.490 ;
        RECT 75.855 145.445 76.145 145.675 ;
        RECT 76.775 145.630 77.065 145.675 ;
        RECT 77.995 145.630 78.285 145.675 ;
        RECT 76.775 145.490 78.285 145.630 ;
        RECT 76.775 145.445 77.065 145.490 ;
        RECT 77.995 145.445 78.285 145.490 ;
        RECT 78.600 145.630 78.920 145.690 ;
        RECT 79.075 145.630 79.365 145.675 ;
        RECT 78.600 145.490 79.365 145.630 ;
        RECT 74.015 145.290 74.305 145.335 ;
        RECT 75.930 145.290 76.070 145.445 ;
        RECT 78.600 145.430 78.920 145.490 ;
        RECT 79.075 145.445 79.365 145.490 ;
        RECT 80.455 145.630 80.745 145.675 ;
        RECT 81.450 145.630 81.590 146.170 ;
        RECT 84.580 146.170 88.030 146.310 ;
        RECT 84.580 146.110 84.900 146.170 ;
        RECT 86.895 146.125 87.185 146.170 ;
        RECT 93.780 146.110 94.100 146.370 ;
        RECT 94.255 146.310 94.545 146.355 ;
        RECT 97.000 146.310 97.320 146.370 ;
        RECT 94.255 146.170 97.320 146.310 ;
        RECT 94.255 146.125 94.545 146.170 ;
        RECT 97.000 146.110 97.320 146.170 ;
        RECT 97.920 146.310 98.240 146.370 ;
        RECT 98.855 146.310 99.145 146.355 ;
        RECT 99.300 146.310 99.620 146.370 ;
        RECT 97.920 146.170 99.620 146.310 ;
        RECT 97.920 146.110 98.240 146.170 ;
        RECT 98.855 146.125 99.145 146.170 ;
        RECT 99.300 146.110 99.620 146.170 ;
        RECT 99.760 146.310 100.080 146.370 ;
        RECT 100.235 146.310 100.525 146.355 ;
        RECT 103.070 146.310 103.210 146.510 ;
        RECT 111.720 146.450 112.040 146.510 ;
        RECT 112.195 146.465 112.485 146.510 ;
        RECT 114.940 146.450 115.260 146.710 ;
        RECT 116.320 146.650 116.640 146.710 ;
        RECT 124.615 146.650 124.905 146.695 ;
        RECT 116.180 146.450 116.640 146.650 ;
        RECT 117.330 146.510 129.890 146.650 ;
        RECT 99.760 146.170 103.210 146.310 ;
        RECT 108.040 146.310 108.360 146.370 ;
        RECT 111.810 146.310 111.950 146.450 ;
        RECT 116.180 146.310 116.320 146.450 ;
        RECT 108.040 146.170 111.950 146.310 ;
        RECT 112.730 146.170 114.710 146.310 ;
        RECT 99.760 146.110 100.080 146.170 ;
        RECT 100.235 146.125 100.525 146.170 ;
        RECT 108.040 146.110 108.360 146.170 ;
        RECT 85.960 145.770 86.280 146.030 ;
        RECT 86.435 145.785 86.725 146.015 ;
        RECT 82.135 145.630 82.425 145.675 ;
        RECT 80.455 145.490 81.130 145.630 ;
        RECT 81.450 145.490 82.425 145.630 ;
        RECT 80.455 145.445 80.745 145.490 ;
        RECT 80.990 145.350 81.130 145.490 ;
        RECT 82.135 145.445 82.425 145.490 ;
        RECT 83.215 145.630 83.505 145.675 ;
        RECT 85.500 145.630 85.820 145.690 ;
        RECT 83.215 145.490 85.820 145.630 ;
        RECT 86.510 145.630 86.650 145.785 ;
        RECT 87.340 145.770 87.660 146.030 ;
        RECT 88.275 145.785 88.565 146.015 ;
        RECT 87.800 145.630 88.120 145.690 ;
        RECT 86.510 145.490 88.120 145.630 ;
        RECT 83.215 145.445 83.505 145.490 ;
        RECT 85.500 145.430 85.820 145.490 ;
        RECT 87.800 145.430 88.120 145.490 ;
        RECT 74.015 145.150 76.070 145.290 ;
        RECT 74.015 145.105 74.305 145.150 ;
        RECT 77.220 145.090 77.540 145.350 ;
        RECT 80.900 145.090 81.220 145.350 ;
        RECT 81.360 145.090 81.680 145.350 ;
        RECT 82.740 145.290 83.060 145.350 ;
        RECT 87.340 145.290 87.660 145.350 ;
        RECT 82.740 145.150 87.660 145.290 ;
        RECT 88.350 145.290 88.490 145.785 ;
        RECT 92.400 145.770 92.720 146.030 ;
        RECT 93.335 145.785 93.625 146.015 ;
        RECT 95.175 145.970 95.465 146.015 ;
        RECT 95.620 145.970 95.940 146.030 ;
        RECT 95.175 145.830 95.940 145.970 ;
        RECT 95.175 145.785 95.465 145.830 ;
        RECT 93.410 145.630 93.550 145.785 ;
        RECT 95.620 145.770 95.940 145.830 ;
        RECT 96.540 145.970 96.860 146.030 ;
        RECT 104.375 145.970 104.665 146.015 ;
        RECT 96.540 145.830 104.665 145.970 ;
        RECT 96.540 145.770 96.860 145.830 ;
        RECT 104.375 145.785 104.665 145.830 ;
        RECT 104.820 145.770 105.140 146.030 ;
        RECT 105.740 145.970 106.060 146.030 ;
        RECT 106.215 145.970 106.505 146.015 ;
        RECT 105.740 145.830 106.505 145.970 ;
        RECT 105.740 145.770 106.060 145.830 ;
        RECT 106.215 145.785 106.505 145.830 ;
        RECT 109.880 145.770 110.200 146.030 ;
        RECT 110.340 145.970 110.660 146.030 ;
        RECT 110.815 145.970 111.105 146.015 ;
        RECT 110.340 145.830 111.105 145.970 ;
        RECT 110.340 145.770 110.660 145.830 ;
        RECT 110.815 145.785 111.105 145.830 ;
        RECT 111.260 145.770 111.580 146.030 ;
        RECT 112.730 146.015 112.870 146.170 ;
        RECT 112.655 145.785 112.945 146.015 ;
        RECT 113.100 145.770 113.420 146.030 ;
        RECT 114.570 146.015 114.710 146.170 ;
        RECT 115.490 146.170 116.320 146.310 ;
        RECT 114.495 145.970 114.785 146.015 ;
        RECT 115.490 145.970 115.630 146.170 ;
        RECT 117.330 146.030 117.470 146.510 ;
        RECT 124.615 146.465 124.905 146.510 ;
        RECT 120.935 146.310 121.225 146.355 ;
        RECT 118.250 146.170 121.225 146.310 ;
        RECT 118.250 146.030 118.390 146.170 ;
        RECT 120.935 146.125 121.225 146.170 ;
        RECT 121.840 146.110 122.160 146.370 ;
        RECT 125.075 146.310 125.365 146.355 ;
        RECT 125.520 146.310 125.840 146.370 ;
        RECT 125.075 146.170 125.840 146.310 ;
        RECT 125.075 146.125 125.365 146.170 ;
        RECT 125.520 146.110 125.840 146.170 ;
        RECT 126.530 146.170 128.050 146.310 ;
        RECT 114.495 145.830 115.630 145.970 ;
        RECT 114.495 145.785 114.785 145.830 ;
        RECT 115.860 145.770 116.180 146.030 ;
        RECT 116.335 145.970 116.625 146.015 ;
        RECT 116.780 145.970 117.100 146.030 ;
        RECT 116.335 145.830 117.100 145.970 ;
        RECT 116.335 145.785 116.625 145.830 ;
        RECT 116.780 145.770 117.100 145.830 ;
        RECT 117.240 145.770 117.560 146.030 ;
        RECT 118.160 145.770 118.480 146.030 ;
        RECT 118.620 145.970 118.940 146.030 ;
        RECT 119.555 145.970 119.845 146.015 ;
        RECT 118.620 145.830 119.845 145.970 ;
        RECT 118.620 145.770 118.940 145.830 ;
        RECT 119.555 145.785 119.845 145.830 ;
        RECT 120.475 145.785 120.765 146.015 ;
        RECT 121.395 145.970 121.685 146.015 ;
        RECT 121.930 145.970 122.070 146.110 ;
        RECT 121.395 145.830 122.070 145.970 ;
        RECT 122.315 145.970 122.605 146.015 ;
        RECT 122.775 145.970 123.065 146.015 ;
        RECT 122.315 145.830 123.065 145.970 ;
        RECT 121.395 145.785 121.685 145.830 ;
        RECT 122.315 145.785 122.605 145.830 ;
        RECT 122.775 145.785 123.065 145.830 ;
        RECT 123.695 145.970 123.985 146.015 ;
        RECT 124.140 145.970 124.460 146.030 ;
        RECT 123.695 145.830 124.460 145.970 ;
        RECT 123.695 145.785 123.985 145.830 ;
        RECT 97.920 145.630 98.240 145.690 ;
        RECT 104.910 145.630 105.050 145.770 ;
        RECT 108.500 145.630 108.820 145.690 ;
        RECT 118.250 145.630 118.390 145.770 ;
        RECT 93.410 145.490 98.240 145.630 ;
        RECT 97.920 145.430 98.240 145.490 ;
        RECT 98.470 145.490 104.590 145.630 ;
        RECT 104.910 145.490 118.390 145.630 ;
        RECT 120.550 145.630 120.690 145.785 ;
        RECT 124.140 145.770 124.460 145.830 ;
        RECT 120.550 145.490 122.070 145.630 ;
        RECT 88.720 145.290 89.040 145.350 ;
        RECT 98.470 145.290 98.610 145.490 ;
        RECT 104.450 145.350 104.590 145.490 ;
        RECT 108.500 145.430 108.820 145.490 ;
        RECT 121.930 145.350 122.070 145.490 ;
        RECT 88.350 145.150 98.610 145.290 ;
        RECT 102.520 145.290 102.840 145.350 ;
        RECT 103.455 145.290 103.745 145.335 ;
        RECT 102.520 145.150 103.745 145.290 ;
        RECT 82.740 145.090 83.060 145.150 ;
        RECT 87.340 145.090 87.660 145.150 ;
        RECT 88.720 145.090 89.040 145.150 ;
        RECT 102.520 145.090 102.840 145.150 ;
        RECT 103.455 145.105 103.745 145.150 ;
        RECT 104.360 145.290 104.680 145.350 ;
        RECT 110.340 145.290 110.660 145.350 ;
        RECT 104.360 145.150 110.660 145.290 ;
        RECT 104.360 145.090 104.680 145.150 ;
        RECT 110.340 145.090 110.660 145.150 ;
        RECT 114.035 145.290 114.325 145.335 ;
        RECT 116.320 145.290 116.640 145.350 ;
        RECT 114.035 145.150 116.640 145.290 ;
        RECT 114.035 145.105 114.325 145.150 ;
        RECT 116.320 145.090 116.640 145.150 ;
        RECT 117.255 145.290 117.545 145.335 ;
        RECT 118.160 145.290 118.480 145.350 ;
        RECT 117.255 145.150 118.480 145.290 ;
        RECT 117.255 145.105 117.545 145.150 ;
        RECT 118.160 145.090 118.480 145.150 ;
        RECT 118.620 145.090 118.940 145.350 ;
        RECT 121.840 145.290 122.160 145.350 ;
        RECT 126.530 145.290 126.670 146.170 ;
        RECT 127.360 145.770 127.680 146.030 ;
        RECT 127.910 145.980 128.050 146.170 ;
        RECT 128.740 146.110 129.060 146.370 ;
        RECT 128.295 145.980 128.585 146.015 ;
        RECT 127.910 145.840 128.585 145.980 ;
        RECT 128.295 145.785 128.585 145.840 ;
        RECT 129.215 145.970 129.505 146.015 ;
        RECT 129.750 145.970 129.890 146.510 ;
        RECT 131.590 146.310 131.730 146.850 ;
        RECT 131.960 146.850 136.405 146.990 ;
        RECT 131.960 146.790 132.280 146.850 ;
        RECT 136.115 146.805 136.405 146.850 ;
        RECT 132.420 146.650 132.740 146.710 ;
        RECT 146.680 146.650 147.000 146.710 ;
        RECT 132.420 146.510 147.000 146.650 ;
        RECT 132.420 146.450 132.740 146.510 ;
        RECT 146.680 146.450 147.000 146.510 ;
        RECT 131.590 146.170 137.710 146.310 ;
        RECT 129.215 145.830 129.890 145.970 ;
        RECT 129.215 145.785 129.505 145.830 ;
        RECT 128.740 145.630 129.060 145.690 ;
        RECT 129.750 145.630 129.890 145.830 ;
        RECT 130.135 145.970 130.425 146.015 ;
        RECT 130.135 145.830 132.190 145.970 ;
        RECT 130.135 145.785 130.425 145.830 ;
        RECT 128.740 145.490 129.890 145.630 ;
        RECT 128.740 145.430 129.060 145.490 ;
        RECT 131.040 145.430 131.360 145.690 ;
        RECT 132.050 145.630 132.190 145.830 ;
        RECT 132.420 145.770 132.740 146.030 ;
        RECT 134.720 145.970 135.040 146.030 ;
        RECT 135.655 145.970 135.945 146.015 ;
        RECT 136.560 145.970 136.880 146.030 ;
        RECT 137.570 146.015 137.710 146.170 ;
        RECT 138.400 146.110 138.720 146.370 ;
        RECT 140.700 146.310 141.020 146.370 ;
        RECT 138.950 146.170 141.020 146.310 ;
        RECT 134.720 145.830 136.880 145.970 ;
        RECT 134.720 145.770 135.040 145.830 ;
        RECT 135.655 145.785 135.945 145.830 ;
        RECT 136.560 145.770 136.880 145.830 ;
        RECT 137.035 145.785 137.325 146.015 ;
        RECT 137.495 145.970 137.785 146.015 ;
        RECT 138.950 145.970 139.090 146.170 ;
        RECT 140.700 146.110 141.020 146.170 ;
        RECT 137.495 145.830 139.090 145.970 ;
        RECT 137.495 145.785 137.785 145.830 ;
        RECT 137.110 145.630 137.250 145.785 ;
        RECT 139.320 145.770 139.640 146.030 ;
        RECT 139.410 145.630 139.550 145.770 ;
        RECT 132.050 145.490 139.550 145.630 ;
        RECT 131.515 145.290 131.805 145.335 ;
        RECT 121.840 145.150 131.805 145.290 ;
        RECT 121.840 145.090 122.160 145.150 ;
        RECT 131.515 145.105 131.805 145.150 ;
        RECT 70.710 144.470 156.270 144.950 ;
        RECT 75.380 144.270 75.700 144.330 ;
        RECT 76.315 144.270 76.605 144.315 ;
        RECT 75.380 144.130 76.605 144.270 ;
        RECT 75.380 144.070 75.700 144.130 ;
        RECT 76.315 144.085 76.605 144.130 ;
        RECT 77.220 144.070 77.540 144.330 ;
        RECT 81.360 144.070 81.680 144.330 ;
        RECT 83.200 144.070 83.520 144.330 ;
        RECT 97.000 144.270 97.320 144.330 ;
        RECT 94.330 144.130 98.610 144.270 ;
        RECT 77.310 143.930 77.450 144.070 ;
        RECT 75.010 143.790 77.450 143.930 ;
        RECT 81.450 143.930 81.590 144.070 ;
        RECT 81.450 143.790 85.270 143.930 ;
        RECT 75.010 143.635 75.150 143.790 ;
        RECT 74.935 143.405 75.225 143.635 ;
        RECT 76.760 143.390 77.080 143.650 ;
        RECT 84.580 143.390 84.900 143.650 ;
        RECT 85.130 143.635 85.270 143.790 ;
        RECT 92.950 143.790 94.010 143.930 ;
        RECT 92.950 143.650 93.090 143.790 ;
        RECT 85.055 143.405 85.345 143.635 ;
        RECT 92.400 143.390 92.720 143.650 ;
        RECT 92.860 143.390 93.180 143.650 ;
        RECT 93.870 143.635 94.010 143.790 ;
        RECT 94.330 143.635 94.470 144.130 ;
        RECT 97.000 144.070 97.320 144.130 ;
        RECT 93.335 143.405 93.625 143.635 ;
        RECT 93.795 143.405 94.085 143.635 ;
        RECT 94.255 143.405 94.545 143.635 ;
        RECT 83.215 143.065 83.505 143.295 ;
        RECT 83.290 142.910 83.430 143.065 ;
        RECT 84.120 143.050 84.440 143.310 ;
        RECT 85.500 143.250 85.820 143.310 ;
        RECT 84.670 143.110 85.820 143.250 ;
        RECT 93.410 143.250 93.550 143.405 ;
        RECT 95.160 143.390 95.480 143.650 ;
        RECT 97.015 143.455 97.305 143.685 ;
        RECT 97.090 143.310 97.230 143.455 ;
        RECT 97.920 143.390 98.240 143.650 ;
        RECT 98.470 143.590 98.610 144.130 ;
        RECT 104.360 144.070 104.680 144.330 ;
        RECT 110.340 144.270 110.660 144.330 ;
        RECT 111.260 144.270 111.580 144.330 ;
        RECT 123.220 144.270 123.540 144.330 ;
        RECT 124.600 144.270 124.920 144.330 ;
        RECT 107.670 144.130 108.730 144.270 ;
        RECT 104.450 143.930 104.590 144.070 ;
        RECT 107.670 143.930 107.810 144.130 ;
        RECT 99.850 143.790 104.590 143.930 ;
        RECT 107.210 143.790 107.810 143.930 ;
        RECT 108.590 143.930 108.730 144.130 ;
        RECT 110.340 144.130 111.580 144.270 ;
        RECT 110.340 144.070 110.660 144.130 ;
        RECT 111.260 144.070 111.580 144.130 ;
        RECT 118.250 144.130 118.950 144.270 ;
        RECT 115.400 143.930 115.720 143.990 ;
        RECT 118.250 143.930 118.390 144.130 ;
        RECT 108.590 143.790 109.420 143.930 ;
        RECT 99.850 143.635 99.990 143.790 ;
        RECT 98.855 143.590 99.145 143.635 ;
        RECT 98.470 143.450 99.145 143.590 ;
        RECT 98.855 143.405 99.145 143.450 ;
        RECT 99.775 143.405 100.065 143.635 ;
        RECT 100.680 143.590 101.000 143.650 ;
        RECT 102.535 143.590 102.825 143.635 ;
        RECT 100.680 143.450 102.825 143.590 ;
        RECT 100.680 143.390 101.000 143.450 ;
        RECT 102.535 143.405 102.825 143.450 ;
        RECT 103.900 143.390 104.220 143.650 ;
        RECT 104.360 143.590 104.680 143.650 ;
        RECT 105.740 143.590 106.060 143.650 ;
        RECT 104.360 143.580 106.060 143.590 ;
        RECT 106.215 143.580 106.505 143.635 ;
        RECT 107.210 143.590 107.350 143.790 ;
        RECT 104.360 143.450 106.505 143.580 ;
        RECT 104.360 143.390 104.680 143.450 ;
        RECT 105.740 143.440 106.505 143.450 ;
        RECT 105.740 143.390 106.060 143.440 ;
        RECT 106.215 143.405 106.505 143.440 ;
        RECT 106.750 143.450 107.350 143.590 ;
        RECT 93.410 143.110 94.010 143.250 ;
        RECT 84.670 142.910 84.810 143.110 ;
        RECT 85.500 143.050 85.820 143.110 ;
        RECT 91.480 142.910 91.800 142.970 ;
        RECT 83.290 142.770 84.810 142.910 ;
        RECT 85.130 142.770 91.800 142.910 ;
        RECT 93.870 142.910 94.010 143.110 ;
        RECT 97.000 143.050 97.320 143.310 ;
        RECT 98.010 142.910 98.150 143.390 ;
        RECT 98.380 143.050 98.700 143.310 ;
        RECT 102.980 143.050 103.300 143.310 ;
        RECT 104.835 143.250 105.125 143.295 ;
        RECT 106.750 143.250 106.890 143.450 ;
        RECT 108.040 143.390 108.360 143.650 ;
        RECT 109.280 143.635 109.420 143.790 ;
        RECT 115.400 143.790 118.390 143.930 ;
        RECT 115.400 143.730 115.720 143.790 ;
        RECT 109.035 143.450 109.420 143.635 ;
        RECT 109.035 143.405 109.325 143.450 ;
        RECT 110.340 143.390 110.660 143.650 ;
        RECT 113.190 143.450 115.630 143.590 ;
        RECT 104.835 143.110 106.890 143.250 ;
        RECT 104.835 143.065 105.125 143.110 ;
        RECT 107.135 143.065 107.425 143.295 ;
        RECT 107.595 143.210 107.885 143.295 ;
        RECT 108.500 143.210 108.820 143.310 ;
        RECT 107.595 143.070 108.820 143.210 ;
        RECT 107.595 143.065 107.885 143.070 ;
        RECT 93.870 142.770 98.150 142.910 ;
        RECT 101.140 142.910 101.460 142.970 ;
        RECT 107.210 142.910 107.350 143.065 ;
        RECT 108.500 143.050 108.820 143.070 ;
        RECT 110.430 142.910 110.570 143.390 ;
        RECT 113.190 143.310 113.330 143.450 ;
        RECT 113.100 143.050 113.420 143.310 ;
        RECT 114.940 143.050 115.260 143.310 ;
        RECT 115.490 143.250 115.630 143.450 ;
        RECT 115.860 143.390 116.180 143.650 ;
        RECT 116.320 143.590 116.640 143.650 ;
        RECT 118.810 143.635 118.950 144.130 ;
        RECT 123.220 144.130 124.920 144.270 ;
        RECT 123.220 144.070 123.540 144.130 ;
        RECT 124.600 144.070 124.920 144.130 ;
        RECT 127.360 144.270 127.680 144.330 ;
        RECT 127.835 144.270 128.125 144.315 ;
        RECT 127.360 144.130 128.125 144.270 ;
        RECT 127.360 144.070 127.680 144.130 ;
        RECT 127.835 144.085 128.125 144.130 ;
        RECT 128.280 144.070 128.600 144.330 ;
        RECT 128.740 144.070 129.060 144.330 ;
        RECT 125.995 143.930 126.285 143.975 ;
        RECT 126.440 143.930 126.760 143.990 ;
        RECT 125.995 143.790 126.760 143.930 ;
        RECT 125.995 143.745 126.285 143.790 ;
        RECT 126.440 143.730 126.760 143.790 ;
        RECT 126.900 143.730 127.220 143.990 ;
        RECT 117.255 143.600 117.545 143.635 ;
        RECT 116.870 143.590 117.545 143.600 ;
        RECT 116.320 143.460 117.545 143.590 ;
        RECT 116.320 143.450 117.010 143.460 ;
        RECT 116.320 143.390 116.640 143.450 ;
        RECT 117.255 143.405 117.545 143.460 ;
        RECT 117.775 143.405 118.065 143.635 ;
        RECT 118.635 143.450 118.950 143.635 ;
        RECT 125.520 143.590 125.840 143.650 ;
        RECT 128.370 143.590 128.510 144.070 ;
        RECT 125.520 143.450 128.510 143.590 ;
        RECT 128.830 143.590 128.970 144.070 ;
        RECT 140.240 143.930 140.560 143.990 ;
        RECT 141.175 143.930 141.465 143.975 ;
        RECT 140.240 143.790 142.770 143.930 ;
        RECT 140.240 143.730 140.560 143.790 ;
        RECT 141.175 143.745 141.465 143.790 ;
        RECT 129.675 143.590 129.965 143.635 ;
        RECT 128.830 143.450 129.965 143.590 ;
        RECT 118.635 143.405 118.925 143.450 ;
        RECT 116.795 143.250 117.085 143.295 ;
        RECT 115.490 143.110 117.085 143.250 ;
        RECT 116.795 143.065 117.085 143.110 ;
        RECT 117.790 143.250 117.930 143.405 ;
        RECT 125.520 143.390 125.840 143.450 ;
        RECT 129.675 143.405 129.965 143.450 ;
        RECT 133.800 143.590 134.120 143.650 ;
        RECT 142.630 143.635 142.770 143.790 ;
        RECT 146.220 143.730 146.540 143.990 ;
        RECT 136.575 143.590 136.865 143.635 ;
        RECT 133.800 143.450 136.865 143.590 ;
        RECT 133.800 143.390 134.120 143.450 ;
        RECT 136.575 143.405 136.865 143.450 ;
        RECT 142.095 143.405 142.385 143.635 ;
        RECT 142.555 143.405 142.845 143.635 ;
        RECT 121.840 143.250 122.160 143.310 ;
        RECT 117.790 143.110 122.160 143.250 ;
        RECT 116.320 142.910 116.640 142.970 ;
        RECT 101.140 142.770 105.510 142.910 ;
        RECT 107.210 142.770 109.420 142.910 ;
        RECT 110.430 142.770 116.640 142.910 ;
        RECT 116.870 142.910 117.010 143.065 ;
        RECT 117.240 142.910 117.560 142.970 ;
        RECT 116.870 142.770 117.560 142.910 ;
        RECT 74.000 142.370 74.320 142.630 ;
        RECT 76.300 142.570 76.620 142.630 ;
        RECT 85.130 142.570 85.270 142.770 ;
        RECT 91.480 142.710 91.800 142.770 ;
        RECT 101.140 142.710 101.460 142.770 ;
        RECT 76.300 142.430 85.270 142.570 ;
        RECT 85.500 142.570 85.820 142.630 ;
        RECT 85.975 142.570 86.265 142.615 ;
        RECT 85.500 142.430 86.265 142.570 ;
        RECT 76.300 142.370 76.620 142.430 ;
        RECT 85.500 142.370 85.820 142.430 ;
        RECT 85.975 142.385 86.265 142.430 ;
        RECT 96.095 142.570 96.385 142.615 ;
        RECT 99.300 142.570 99.620 142.630 ;
        RECT 96.095 142.430 99.620 142.570 ;
        RECT 96.095 142.385 96.385 142.430 ;
        RECT 99.300 142.370 99.620 142.430 ;
        RECT 100.695 142.570 100.985 142.615 ;
        RECT 102.520 142.570 102.840 142.630 ;
        RECT 105.370 142.615 105.510 142.770 ;
        RECT 100.695 142.430 102.840 142.570 ;
        RECT 100.695 142.385 100.985 142.430 ;
        RECT 102.520 142.370 102.840 142.430 ;
        RECT 105.295 142.385 105.585 142.615 ;
        RECT 109.280 142.570 109.420 142.770 ;
        RECT 116.320 142.710 116.640 142.770 ;
        RECT 117.240 142.710 117.560 142.770 ;
        RECT 117.790 142.570 117.930 143.110 ;
        RECT 121.840 143.050 122.160 143.110 ;
        RECT 128.295 143.250 128.585 143.295 ;
        RECT 129.200 143.250 129.520 143.310 ;
        RECT 128.295 143.110 129.520 143.250 ;
        RECT 128.295 143.065 128.585 143.110 ;
        RECT 129.200 143.050 129.520 143.110 ;
        RECT 131.500 143.250 131.820 143.310 ;
        RECT 137.035 143.250 137.325 143.295 ;
        RECT 131.500 143.110 137.325 143.250 ;
        RECT 131.500 143.050 131.820 143.110 ;
        RECT 137.035 143.065 137.325 143.110 ;
        RECT 137.480 143.050 137.800 143.310 ;
        RECT 137.940 143.050 138.260 143.310 ;
        RECT 142.170 143.250 142.310 143.405 ;
        RECT 143.460 143.390 143.780 143.650 ;
        RECT 146.310 143.250 146.450 143.730 ;
        RECT 150.835 143.590 151.125 143.635 ;
        RECT 151.740 143.590 152.060 143.650 ;
        RECT 150.835 143.450 152.060 143.590 ;
        RECT 150.835 143.405 151.125 143.450 ;
        RECT 151.740 143.390 152.060 143.450 ;
        RECT 142.170 143.110 146.450 143.250 ;
        RECT 151.295 143.250 151.585 143.295 ;
        RECT 152.200 143.250 152.520 143.310 ;
        RECT 153.120 143.250 153.440 143.310 ;
        RECT 151.295 143.110 153.440 143.250 ;
        RECT 151.295 143.065 151.585 143.110 ;
        RECT 152.200 143.050 152.520 143.110 ;
        RECT 153.120 143.050 153.440 143.110 ;
        RECT 109.280 142.430 117.930 142.570 ;
        RECT 138.860 142.370 139.180 142.630 ;
        RECT 140.240 142.370 140.560 142.630 ;
        RECT 141.160 142.570 141.480 142.630 ;
        RECT 143.015 142.570 143.305 142.615 ;
        RECT 141.160 142.430 143.305 142.570 ;
        RECT 141.160 142.370 141.480 142.430 ;
        RECT 143.015 142.385 143.305 142.430 ;
        RECT 148.980 142.370 149.300 142.630 ;
        RECT 70.710 141.750 156.270 142.230 ;
        RECT 88.720 141.550 89.040 141.610 ;
        RECT 91.035 141.550 91.325 141.595 ;
        RECT 95.160 141.550 95.480 141.610 ;
        RECT 88.720 141.410 95.480 141.550 ;
        RECT 88.720 141.350 89.040 141.410 ;
        RECT 91.035 141.365 91.325 141.410 ;
        RECT 95.160 141.350 95.480 141.410 ;
        RECT 98.855 141.550 99.145 141.595 ;
        RECT 103.900 141.550 104.220 141.610 ;
        RECT 124.140 141.550 124.460 141.610 ;
        RECT 125.075 141.550 125.365 141.595 ;
        RECT 135.655 141.550 135.945 141.595 ;
        RECT 98.855 141.410 103.670 141.550 ;
        RECT 98.855 141.365 99.145 141.410 ;
        RECT 72.660 141.210 72.950 141.255 ;
        RECT 74.760 141.210 75.050 141.255 ;
        RECT 76.330 141.210 76.620 141.255 ;
        RECT 72.660 141.070 76.620 141.210 ;
        RECT 72.660 141.025 72.950 141.070 ;
        RECT 74.760 141.025 75.050 141.070 ;
        RECT 76.330 141.025 76.620 141.070 ;
        RECT 84.620 141.210 84.910 141.255 ;
        RECT 86.720 141.210 87.010 141.255 ;
        RECT 88.290 141.210 88.580 141.255 ;
        RECT 84.620 141.070 88.580 141.210 ;
        RECT 84.620 141.025 84.910 141.070 ;
        RECT 86.720 141.025 87.010 141.070 ;
        RECT 88.290 141.025 88.580 141.070 ;
        RECT 91.480 141.210 91.800 141.270 ;
        RECT 93.780 141.210 94.100 141.270 ;
        RECT 100.680 141.210 101.000 141.270 ;
        RECT 91.480 141.070 94.100 141.210 ;
        RECT 91.480 141.010 91.800 141.070 ;
        RECT 93.780 141.010 94.100 141.070 ;
        RECT 96.630 141.070 101.000 141.210 ;
        RECT 103.530 141.210 103.670 141.410 ;
        RECT 103.900 141.410 125.365 141.550 ;
        RECT 103.900 141.350 104.220 141.410 ;
        RECT 124.140 141.350 124.460 141.410 ;
        RECT 105.755 141.210 106.045 141.255 ;
        RECT 108.040 141.210 108.360 141.270 ;
        RECT 103.530 141.070 106.045 141.210 ;
        RECT 73.055 140.870 73.345 140.915 ;
        RECT 74.245 140.870 74.535 140.915 ;
        RECT 76.765 140.870 77.055 140.915 ;
        RECT 84.135 140.870 84.425 140.915 ;
        RECT 73.055 140.730 77.055 140.870 ;
        RECT 73.055 140.685 73.345 140.730 ;
        RECT 74.245 140.685 74.535 140.730 ;
        RECT 76.765 140.685 77.055 140.730 ;
        RECT 77.310 140.730 84.425 140.870 ;
        RECT 72.160 140.530 72.480 140.590 ;
        RECT 77.310 140.530 77.450 140.730 ;
        RECT 84.135 140.685 84.425 140.730 ;
        RECT 85.015 140.870 85.305 140.915 ;
        RECT 86.205 140.870 86.495 140.915 ;
        RECT 88.725 140.870 89.015 140.915 ;
        RECT 85.015 140.730 89.015 140.870 ;
        RECT 85.015 140.685 85.305 140.730 ;
        RECT 86.205 140.685 86.495 140.730 ;
        RECT 88.725 140.685 89.015 140.730 ;
        RECT 72.160 140.390 77.450 140.530 ;
        RECT 79.520 140.530 79.840 140.590 ;
        RECT 85.500 140.575 85.820 140.590 ;
        RECT 80.455 140.530 80.745 140.575 ;
        RECT 79.520 140.390 80.745 140.530 ;
        RECT 72.160 140.330 72.480 140.390 ;
        RECT 79.520 140.330 79.840 140.390 ;
        RECT 80.455 140.345 80.745 140.390 ;
        RECT 81.375 140.345 81.665 140.575 ;
        RECT 85.470 140.530 85.820 140.575 ;
        RECT 85.305 140.390 85.820 140.530 ;
        RECT 85.470 140.345 85.820 140.390 ;
        RECT 73.510 140.190 73.800 140.235 ;
        RECT 74.000 140.190 74.320 140.250 ;
        RECT 73.510 140.050 74.320 140.190 ;
        RECT 73.510 140.005 73.800 140.050 ;
        RECT 74.000 139.990 74.320 140.050 ;
        RECT 81.450 139.910 81.590 140.345 ;
        RECT 85.500 140.330 85.820 140.345 ;
        RECT 87.340 140.530 87.660 140.590 ;
        RECT 96.080 140.530 96.400 140.590 ;
        RECT 96.630 140.575 96.770 141.070 ;
        RECT 100.680 141.010 101.000 141.070 ;
        RECT 105.755 141.025 106.045 141.070 ;
        RECT 106.290 141.070 108.360 141.210 ;
        RECT 102.060 140.870 102.380 140.930 ;
        RECT 97.090 140.730 102.380 140.870 ;
        RECT 97.090 140.575 97.230 140.730 ;
        RECT 102.060 140.670 102.380 140.730 ;
        RECT 87.340 140.390 96.400 140.530 ;
        RECT 87.340 140.330 87.660 140.390 ;
        RECT 96.080 140.330 96.400 140.390 ;
        RECT 96.555 140.345 96.845 140.575 ;
        RECT 97.015 140.345 97.305 140.575 ;
        RECT 97.920 140.330 98.240 140.590 ;
        RECT 98.395 140.345 98.685 140.575 ;
        RECT 99.300 140.530 99.620 140.590 ;
        RECT 99.775 140.530 100.065 140.575 ;
        RECT 99.300 140.390 100.065 140.530 ;
        RECT 82.295 140.190 82.585 140.235 ;
        RECT 95.620 140.190 95.940 140.250 ;
        RECT 98.470 140.190 98.610 140.345 ;
        RECT 99.300 140.330 99.620 140.390 ;
        RECT 99.775 140.345 100.065 140.390 ;
        RECT 102.520 140.530 102.840 140.590 ;
        RECT 104.835 140.530 105.125 140.575 ;
        RECT 102.520 140.390 105.125 140.530 ;
        RECT 102.520 140.330 102.840 140.390 ;
        RECT 104.835 140.345 105.125 140.390 ;
        RECT 82.295 140.050 95.940 140.190 ;
        RECT 82.295 140.005 82.585 140.050 ;
        RECT 95.620 139.990 95.940 140.050 ;
        RECT 96.630 140.050 98.610 140.190 ;
        RECT 105.830 140.190 105.970 141.025 ;
        RECT 106.290 140.915 106.430 141.070 ;
        RECT 108.040 141.010 108.360 141.070 ;
        RECT 110.340 141.210 110.660 141.270 ;
        RECT 123.220 141.210 123.540 141.270 ;
        RECT 110.340 141.070 123.540 141.210 ;
        RECT 110.340 141.010 110.660 141.070 ;
        RECT 123.220 141.010 123.540 141.070 ;
        RECT 106.215 140.685 106.505 140.915 ;
        RECT 108.500 140.870 108.820 140.930 ;
        RECT 122.760 140.870 123.080 140.930 ;
        RECT 124.690 140.915 124.830 141.410 ;
        RECT 125.075 141.365 125.365 141.410 ;
        RECT 132.970 141.410 135.945 141.550 ;
        RECT 108.500 140.730 123.450 140.870 ;
        RECT 108.500 140.670 108.820 140.730 ;
        RECT 122.760 140.670 123.080 140.730 ;
        RECT 106.660 140.530 106.980 140.590 ;
        RECT 113.100 140.530 113.420 140.590 ;
        RECT 115.875 140.530 116.165 140.575 ;
        RECT 106.660 140.390 116.165 140.530 ;
        RECT 106.660 140.330 106.980 140.390 ;
        RECT 113.100 140.330 113.420 140.390 ;
        RECT 115.875 140.345 116.165 140.390 ;
        RECT 116.780 140.330 117.100 140.590 ;
        RECT 117.240 140.530 117.560 140.590 ;
        RECT 118.160 140.530 118.480 140.590 ;
        RECT 123.310 140.575 123.450 140.730 ;
        RECT 124.615 140.685 124.905 140.915 ;
        RECT 129.200 140.870 129.520 140.930 ;
        RECT 131.055 140.870 131.345 140.915 ;
        RECT 129.200 140.730 131.345 140.870 ;
        RECT 129.200 140.670 129.520 140.730 ;
        RECT 131.055 140.685 131.345 140.730 ;
        RECT 131.960 140.670 132.280 140.930 ;
        RECT 132.435 140.870 132.725 140.915 ;
        RECT 132.970 140.870 133.110 141.410 ;
        RECT 135.655 141.365 135.945 141.410 ;
        RECT 137.940 141.550 138.260 141.610 ;
        RECT 139.780 141.550 140.100 141.610 ;
        RECT 137.940 141.410 140.100 141.550 ;
        RECT 137.940 141.350 138.260 141.410 ;
        RECT 139.780 141.350 140.100 141.410 ;
        RECT 140.700 141.350 141.020 141.610 ;
        RECT 143.460 141.350 143.780 141.610 ;
        RECT 146.220 141.350 146.540 141.610 ;
        RECT 138.030 141.210 138.170 141.350 ;
        RECT 135.730 141.070 138.170 141.210 ;
        RECT 135.730 140.870 135.870 141.070 ;
        RECT 140.255 140.870 140.545 140.915 ;
        RECT 132.435 140.730 133.110 140.870 ;
        RECT 133.430 140.730 135.870 140.870 ;
        RECT 136.190 140.730 140.545 140.870 ;
        RECT 140.790 140.870 140.930 141.350 ;
        RECT 141.175 140.870 141.465 140.915 ;
        RECT 140.790 140.730 141.465 140.870 ;
        RECT 132.435 140.685 132.725 140.730 ;
        RECT 117.240 140.390 118.480 140.530 ;
        RECT 117.240 140.330 117.560 140.390 ;
        RECT 118.160 140.330 118.480 140.390 ;
        RECT 123.235 140.345 123.525 140.575 ;
        RECT 125.520 140.530 125.840 140.590 ;
        RECT 125.995 140.530 126.285 140.575 ;
        RECT 125.520 140.390 126.285 140.530 ;
        RECT 125.520 140.330 125.840 140.390 ;
        RECT 125.995 140.345 126.285 140.390 ;
        RECT 129.675 140.345 129.965 140.575 ;
        RECT 132.050 140.530 132.190 140.670 ;
        RECT 133.430 140.575 133.570 140.730 ;
        RECT 132.895 140.530 133.185 140.575 ;
        RECT 132.050 140.390 133.185 140.530 ;
        RECT 132.895 140.345 133.185 140.390 ;
        RECT 133.355 140.345 133.645 140.575 ;
        RECT 133.800 140.530 134.120 140.590 ;
        RECT 136.190 140.530 136.330 140.730 ;
        RECT 140.255 140.685 140.545 140.730 ;
        RECT 141.175 140.685 141.465 140.730 ;
        RECT 141.635 140.870 141.925 140.915 ;
        RECT 142.080 140.870 142.400 140.930 ;
        RECT 141.635 140.730 142.400 140.870 ;
        RECT 141.635 140.685 141.925 140.730 ;
        RECT 142.080 140.670 142.400 140.730 ;
        RECT 133.800 140.390 136.330 140.530 ;
        RECT 114.020 140.190 114.340 140.250 ;
        RECT 105.830 140.050 114.340 140.190 ;
        RECT 96.630 139.910 96.770 140.050 ;
        RECT 114.020 139.990 114.340 140.050 ;
        RECT 116.320 140.190 116.640 140.250 ;
        RECT 129.750 140.190 129.890 140.345 ;
        RECT 133.800 140.330 134.120 140.390 ;
        RECT 137.020 140.330 137.340 140.590 ;
        RECT 137.495 140.345 137.785 140.575 ;
        RECT 137.955 140.530 138.245 140.575 ;
        RECT 138.400 140.530 138.720 140.590 ;
        RECT 137.955 140.390 138.720 140.530 ;
        RECT 137.955 140.345 138.245 140.390 ;
        RECT 135.180 140.190 135.500 140.250 ;
        RECT 137.570 140.190 137.710 140.345 ;
        RECT 138.400 140.330 138.720 140.390 ;
        RECT 138.875 140.345 139.165 140.575 ;
        RECT 140.715 140.530 141.005 140.575 ;
        RECT 143.550 140.530 143.690 141.350 ;
        RECT 143.920 140.870 144.240 140.930 ;
        RECT 146.310 140.870 146.450 141.350 ;
        RECT 148.535 141.210 148.825 141.255 ;
        RECT 151.740 141.210 152.060 141.270 ;
        RECT 148.535 141.070 152.060 141.210 ;
        RECT 148.535 141.025 148.825 141.070 ;
        RECT 151.740 141.010 152.060 141.070 ;
        RECT 148.995 140.870 149.285 140.915 ;
        RECT 143.920 140.730 145.070 140.870 ;
        RECT 146.310 140.730 148.290 140.870 ;
        RECT 143.920 140.670 144.240 140.730 ;
        RECT 144.930 140.575 145.070 140.730 ;
        RECT 148.150 140.575 148.290 140.730 ;
        RECT 148.995 140.730 152.890 140.870 ;
        RECT 148.995 140.685 149.285 140.730 ;
        RECT 152.750 140.590 152.890 140.730 ;
        RECT 140.715 140.390 143.690 140.530 ;
        RECT 140.715 140.345 141.005 140.390 ;
        RECT 144.395 140.345 144.685 140.575 ;
        RECT 144.855 140.345 145.145 140.575 ;
        RECT 146.235 140.530 146.525 140.575 ;
        RECT 147.155 140.530 147.445 140.575 ;
        RECT 146.235 140.390 147.445 140.530 ;
        RECT 146.235 140.345 146.525 140.390 ;
        RECT 147.155 140.345 147.445 140.390 ;
        RECT 148.075 140.345 148.365 140.575 ;
        RECT 148.520 140.530 148.840 140.590 ;
        RECT 149.455 140.530 149.745 140.575 ;
        RECT 148.520 140.390 149.745 140.530 ;
        RECT 116.320 140.050 137.710 140.190 ;
        RECT 116.320 139.990 116.640 140.050 ;
        RECT 135.180 139.990 135.500 140.050 ;
        RECT 76.760 139.850 77.080 139.910 ;
        RECT 79.075 139.850 79.365 139.895 ;
        RECT 76.760 139.710 79.365 139.850 ;
        RECT 76.760 139.650 77.080 139.710 ;
        RECT 79.075 139.665 79.365 139.710 ;
        RECT 79.520 139.650 79.840 139.910 ;
        RECT 81.360 139.650 81.680 139.910 ;
        RECT 82.755 139.850 83.045 139.895 ;
        RECT 85.040 139.850 85.360 139.910 ;
        RECT 92.400 139.850 92.720 139.910 ;
        RECT 82.755 139.710 92.720 139.850 ;
        RECT 82.755 139.665 83.045 139.710 ;
        RECT 85.040 139.650 85.360 139.710 ;
        RECT 92.400 139.650 92.720 139.710 ;
        RECT 94.700 139.650 95.020 139.910 ;
        RECT 96.540 139.650 96.860 139.910 ;
        RECT 99.760 139.850 100.080 139.910 ;
        RECT 100.695 139.850 100.985 139.895 ;
        RECT 99.760 139.710 100.985 139.850 ;
        RECT 99.760 139.650 100.080 139.710 ;
        RECT 100.695 139.665 100.985 139.710 ;
        RECT 103.900 139.650 104.220 139.910 ;
        RECT 116.795 139.850 117.085 139.895 ;
        RECT 118.160 139.850 118.480 139.910 ;
        RECT 116.795 139.710 118.480 139.850 ;
        RECT 116.795 139.665 117.085 139.710 ;
        RECT 118.160 139.650 118.480 139.710 ;
        RECT 134.720 139.650 135.040 139.910 ;
        RECT 135.640 139.850 135.960 139.910 ;
        RECT 138.950 139.850 139.090 140.345 ;
        RECT 144.470 140.190 144.610 140.345 ;
        RECT 148.520 140.330 148.840 140.390 ;
        RECT 149.455 140.345 149.745 140.390 ;
        RECT 151.740 140.330 152.060 140.590 ;
        RECT 152.660 140.330 152.980 140.590 ;
        RECT 154.500 140.330 154.820 140.590 ;
        RECT 140.790 140.050 144.610 140.190 ;
        RECT 146.695 140.190 146.985 140.235 ;
        RECT 152.200 140.190 152.520 140.250 ;
        RECT 154.055 140.190 154.345 140.235 ;
        RECT 146.695 140.050 154.345 140.190 ;
        RECT 140.790 139.910 140.930 140.050 ;
        RECT 146.695 140.005 146.985 140.050 ;
        RECT 152.200 139.990 152.520 140.050 ;
        RECT 154.055 140.005 154.345 140.050 ;
        RECT 135.640 139.710 139.090 139.850 ;
        RECT 135.640 139.650 135.960 139.710 ;
        RECT 139.320 139.650 139.640 139.910 ;
        RECT 140.700 139.650 141.020 139.910 ;
        RECT 142.080 139.850 142.400 139.910 ;
        RECT 143.475 139.850 143.765 139.895 ;
        RECT 142.080 139.710 143.765 139.850 ;
        RECT 142.080 139.650 142.400 139.710 ;
        RECT 143.475 139.665 143.765 139.710 ;
        RECT 70.710 139.030 156.270 139.510 ;
        RECT 79.075 138.830 79.365 138.875 ;
        RECT 77.770 138.690 79.365 138.830 ;
        RECT 77.770 137.470 77.910 138.690 ;
        RECT 79.075 138.645 79.365 138.690 ;
        RECT 79.520 138.630 79.840 138.890 ;
        RECT 81.835 138.830 82.125 138.875 ;
        RECT 82.280 138.830 82.600 138.890 ;
        RECT 95.160 138.830 95.480 138.890 ;
        RECT 81.835 138.690 95.480 138.830 ;
        RECT 81.835 138.645 82.125 138.690 ;
        RECT 82.280 138.630 82.600 138.690 ;
        RECT 95.160 138.630 95.480 138.690 ;
        RECT 97.920 138.830 98.240 138.890 ;
        RECT 108.500 138.830 108.820 138.890 ;
        RECT 113.560 138.830 113.880 138.890 ;
        RECT 97.920 138.690 108.820 138.830 ;
        RECT 97.920 138.630 98.240 138.690 ;
        RECT 108.500 138.630 108.820 138.690 ;
        RECT 112.730 138.690 113.880 138.830 ;
        RECT 79.610 138.490 79.750 138.630 ;
        RECT 81.360 138.490 81.680 138.550 ;
        RECT 78.230 138.350 79.750 138.490 ;
        RECT 80.990 138.350 87.110 138.490 ;
        RECT 78.230 138.195 78.370 138.350 ;
        RECT 78.155 137.965 78.445 138.195 ;
        RECT 78.600 138.150 78.920 138.210 ;
        RECT 79.535 138.150 79.825 138.195 ;
        RECT 78.600 138.010 79.825 138.150 ;
        RECT 78.600 137.950 78.920 138.010 ;
        RECT 79.535 137.965 79.825 138.010 ;
        RECT 79.980 137.950 80.300 138.210 ;
        RECT 80.990 138.195 81.130 138.350 ;
        RECT 81.360 138.290 81.680 138.350 ;
        RECT 80.915 137.965 81.205 138.195 ;
        RECT 82.295 138.150 82.585 138.195 ;
        RECT 83.660 138.150 83.980 138.210 ;
        RECT 86.970 138.195 87.110 138.350 ;
        RECT 92.860 138.290 93.180 138.550 ;
        RECT 94.240 138.290 94.560 138.550 ;
        RECT 97.460 138.490 97.780 138.550 ;
        RECT 98.395 138.490 98.685 138.535 ;
        RECT 97.460 138.350 98.685 138.490 ;
        RECT 97.460 138.290 97.780 138.350 ;
        RECT 98.395 138.305 98.685 138.350 ;
        RECT 99.315 138.490 99.605 138.535 ;
        RECT 109.880 138.490 110.200 138.550 ;
        RECT 112.730 138.535 112.870 138.690 ;
        RECT 113.560 138.630 113.880 138.690 ;
        RECT 116.780 138.630 117.100 138.890 ;
        RECT 117.240 138.630 117.560 138.890 ;
        RECT 118.160 138.630 118.480 138.890 ;
        RECT 120.000 138.830 120.320 138.890 ;
        RECT 124.140 138.830 124.460 138.890 ;
        RECT 125.980 138.830 126.300 138.890 ;
        RECT 120.000 138.690 126.300 138.830 ;
        RECT 120.000 138.630 120.320 138.690 ;
        RECT 124.140 138.630 124.460 138.690 ;
        RECT 125.980 138.630 126.300 138.690 ;
        RECT 130.120 138.630 130.440 138.890 ;
        RECT 134.260 138.630 134.580 138.890 ;
        RECT 135.180 138.630 135.500 138.890 ;
        RECT 137.020 138.630 137.340 138.890 ;
        RECT 137.480 138.630 137.800 138.890 ;
        RECT 138.860 138.830 139.180 138.890 ;
        RECT 143.000 138.830 143.320 138.890 ;
        RECT 138.860 138.690 143.320 138.830 ;
        RECT 138.860 138.630 139.180 138.690 ;
        RECT 143.000 138.630 143.320 138.690 ;
        RECT 99.315 138.350 107.810 138.490 ;
        RECT 99.315 138.305 99.605 138.350 ;
        RECT 81.910 138.010 83.980 138.150 ;
        RECT 81.910 137.870 82.050 138.010 ;
        RECT 82.295 137.965 82.585 138.010 ;
        RECT 83.660 137.950 83.980 138.010 ;
        RECT 86.895 138.150 87.185 138.195 ;
        RECT 88.720 138.150 89.040 138.210 ;
        RECT 86.895 138.010 89.040 138.150 ;
        RECT 92.950 138.150 93.090 138.290 ;
        RECT 95.175 138.150 95.465 138.195 ;
        RECT 92.950 138.010 95.465 138.150 ;
        RECT 86.895 137.965 87.185 138.010 ;
        RECT 88.720 137.950 89.040 138.010 ;
        RECT 95.175 137.965 95.465 138.010 ;
        RECT 99.775 137.965 100.065 138.195 ;
        RECT 100.680 138.150 101.000 138.210 ;
        RECT 100.310 138.010 101.000 138.150 ;
        RECT 81.820 137.610 82.140 137.870 ;
        RECT 85.515 137.810 85.805 137.855 ;
        RECT 87.340 137.810 87.660 137.870 ;
        RECT 85.515 137.670 87.660 137.810 ;
        RECT 85.515 137.625 85.805 137.670 ;
        RECT 87.340 137.610 87.660 137.670 ;
        RECT 98.380 137.810 98.700 137.870 ;
        RECT 99.850 137.810 99.990 137.965 ;
        RECT 98.380 137.670 99.990 137.810 ;
        RECT 98.380 137.610 98.700 137.670 ;
        RECT 82.280 137.470 82.600 137.530 ;
        RECT 77.770 137.330 82.600 137.470 ;
        RECT 82.280 137.270 82.600 137.330 ;
        RECT 96.095 137.470 96.385 137.515 ;
        RECT 100.310 137.470 100.450 138.010 ;
        RECT 100.680 137.950 101.000 138.010 ;
        RECT 103.440 138.150 103.760 138.210 ;
        RECT 107.670 138.195 107.810 138.350 ;
        RECT 108.130 138.350 110.200 138.490 ;
        RECT 108.130 138.195 108.270 138.350 ;
        RECT 109.880 138.290 110.200 138.350 ;
        RECT 112.655 138.305 112.945 138.535 ;
        RECT 114.020 138.490 114.340 138.550 ;
        RECT 115.415 138.490 115.705 138.535 ;
        RECT 114.020 138.350 115.705 138.490 ;
        RECT 114.020 138.290 114.340 138.350 ;
        RECT 115.415 138.305 115.705 138.350 ;
        RECT 116.870 138.195 117.010 138.630 ;
        RECT 117.330 138.490 117.470 138.630 ;
        RECT 118.250 138.490 118.390 138.630 ;
        RECT 128.295 138.490 128.585 138.535 ;
        RECT 130.210 138.490 130.350 138.630 ;
        RECT 117.330 138.350 117.930 138.490 ;
        RECT 118.250 138.350 120.690 138.490 ;
        RECT 107.135 138.150 107.425 138.195 ;
        RECT 103.440 138.010 107.425 138.150 ;
        RECT 103.440 137.950 103.760 138.010 ;
        RECT 107.135 137.965 107.425 138.010 ;
        RECT 107.595 137.965 107.885 138.195 ;
        RECT 108.055 137.965 108.345 138.195 ;
        RECT 108.975 137.965 109.265 138.195 ;
        RECT 113.575 138.150 113.865 138.195 ;
        RECT 116.795 138.150 117.085 138.195 ;
        RECT 113.575 138.010 117.085 138.150 ;
        RECT 113.575 137.965 113.865 138.010 ;
        RECT 116.795 137.965 117.085 138.010 ;
        RECT 107.670 137.810 107.810 137.965 ;
        RECT 109.050 137.810 109.190 137.965 ;
        RECT 117.240 137.950 117.560 138.210 ;
        RECT 117.790 138.195 117.930 138.350 ;
        RECT 117.715 137.965 118.005 138.195 ;
        RECT 118.160 138.150 118.480 138.210 ;
        RECT 118.635 138.150 118.925 138.195 ;
        RECT 118.160 138.010 118.925 138.150 ;
        RECT 118.160 137.950 118.480 138.010 ;
        RECT 118.635 137.965 118.925 138.010 ;
        RECT 119.080 138.150 119.400 138.210 ;
        RECT 120.550 138.195 120.690 138.350 ;
        RECT 128.295 138.350 130.350 138.490 ;
        RECT 128.295 138.305 128.585 138.350 ;
        RECT 119.555 138.150 119.845 138.195 ;
        RECT 119.080 138.010 119.845 138.150 ;
        RECT 119.080 137.950 119.400 138.010 ;
        RECT 119.555 137.965 119.845 138.010 ;
        RECT 120.475 137.965 120.765 138.195 ;
        RECT 122.760 138.150 123.080 138.210 ;
        RECT 122.760 138.010 128.050 138.150 ;
        RECT 122.760 137.950 123.080 138.010 ;
        RECT 118.250 137.810 118.390 137.950 ;
        RECT 107.670 137.670 108.270 137.810 ;
        RECT 109.050 137.670 118.390 137.810 ;
        RECT 96.095 137.330 100.450 137.470 ;
        RECT 100.695 137.470 100.985 137.515 ;
        RECT 103.440 137.470 103.760 137.530 ;
        RECT 108.130 137.470 108.270 137.670 ;
        RECT 120.000 137.610 120.320 137.870 ;
        RECT 120.935 137.625 121.225 137.855 ;
        RECT 121.855 137.810 122.145 137.855 ;
        RECT 127.360 137.810 127.680 137.870 ;
        RECT 121.855 137.670 127.680 137.810 ;
        RECT 127.910 137.810 128.050 138.010 ;
        RECT 128.740 137.950 129.060 138.210 ;
        RECT 130.210 138.195 130.350 138.350 ;
        RECT 134.350 138.195 134.490 138.630 ;
        RECT 135.270 138.490 135.410 138.630 ;
        RECT 134.810 138.350 135.410 138.490 ;
        RECT 134.810 138.195 134.950 138.350 ;
        RECT 137.110 138.195 137.250 138.630 ;
        RECT 139.870 138.350 141.850 138.490 ;
        RECT 130.095 137.965 130.385 138.195 ;
        RECT 131.055 138.150 131.345 138.195 ;
        RECT 131.055 138.010 131.455 138.150 ;
        RECT 131.055 137.965 131.345 138.010 ;
        RECT 133.355 137.965 133.645 138.195 ;
        RECT 134.275 137.965 134.565 138.195 ;
        RECT 134.735 137.965 135.025 138.195 ;
        RECT 135.195 138.150 135.485 138.195 ;
        RECT 135.195 138.010 136.790 138.150 ;
        RECT 135.195 137.965 135.485 138.010 ;
        RECT 131.130 137.810 131.270 137.965 ;
        RECT 132.420 137.810 132.740 137.870 ;
        RECT 127.910 137.670 132.740 137.810 ;
        RECT 121.855 137.625 122.145 137.670 ;
        RECT 112.640 137.470 112.960 137.530 ;
        RECT 100.695 137.330 103.760 137.470 ;
        RECT 96.095 137.285 96.385 137.330 ;
        RECT 100.695 137.285 100.985 137.330 ;
        RECT 103.440 137.270 103.760 137.330 ;
        RECT 103.990 137.330 107.810 137.470 ;
        RECT 108.130 137.330 112.960 137.470 ;
        RECT 77.220 136.930 77.540 137.190 ;
        RECT 79.980 136.930 80.300 137.190 ;
        RECT 97.475 137.130 97.765 137.175 ;
        RECT 97.920 137.130 98.240 137.190 ;
        RECT 97.475 136.990 98.240 137.130 ;
        RECT 97.475 136.945 97.765 136.990 ;
        RECT 97.920 136.930 98.240 136.990 ;
        RECT 102.060 137.130 102.380 137.190 ;
        RECT 103.990 137.130 104.130 137.330 ;
        RECT 102.060 136.990 104.130 137.130 ;
        RECT 105.755 137.130 106.045 137.175 ;
        RECT 107.120 137.130 107.440 137.190 ;
        RECT 105.755 136.990 107.440 137.130 ;
        RECT 107.670 137.130 107.810 137.330 ;
        RECT 112.640 137.270 112.960 137.330 ;
        RECT 114.495 137.470 114.785 137.515 ;
        RECT 121.010 137.470 121.150 137.625 ;
        RECT 127.360 137.610 127.680 137.670 ;
        RECT 132.420 137.610 132.740 137.670 ;
        RECT 133.430 137.810 133.570 137.965 ;
        RECT 135.640 137.810 135.960 137.870 ;
        RECT 133.430 137.670 135.960 137.810 ;
        RECT 136.650 137.810 136.790 138.010 ;
        RECT 137.035 137.965 137.325 138.195 ;
        RECT 137.940 137.950 138.260 138.210 ;
        RECT 139.870 138.150 140.010 138.350 ;
        RECT 141.710 138.210 141.850 138.350 ;
        RECT 150.450 138.350 152.430 138.490 ;
        RECT 138.490 138.010 140.010 138.150 ;
        RECT 138.490 137.810 138.630 138.010 ;
        RECT 140.240 137.950 140.560 138.210 ;
        RECT 141.620 137.950 141.940 138.210 ;
        RECT 150.450 138.195 150.590 138.350 ;
        RECT 152.290 138.210 152.430 138.350 ;
        RECT 150.375 137.965 150.665 138.195 ;
        RECT 151.755 137.965 152.045 138.195 ;
        RECT 136.650 137.670 138.630 137.810 ;
        RECT 114.495 137.330 121.150 137.470 ;
        RECT 125.520 137.470 125.840 137.530 ;
        RECT 126.455 137.470 126.745 137.515 ;
        RECT 125.520 137.330 126.745 137.470 ;
        RECT 114.495 137.285 114.785 137.330 ;
        RECT 125.520 137.270 125.840 137.330 ;
        RECT 126.455 137.285 126.745 137.330 ;
        RECT 126.900 137.470 127.220 137.530 ;
        RECT 129.675 137.470 129.965 137.515 ;
        RECT 133.430 137.470 133.570 137.670 ;
        RECT 135.640 137.610 135.960 137.670 ;
        RECT 138.860 137.610 139.180 137.870 ;
        RECT 139.335 137.625 139.625 137.855 ;
        RECT 139.795 137.810 140.085 137.855 ;
        RECT 141.160 137.810 141.480 137.870 ;
        RECT 139.795 137.670 141.480 137.810 ;
        RECT 139.795 137.625 140.085 137.670 ;
        RECT 139.410 137.470 139.550 137.625 ;
        RECT 141.160 137.610 141.480 137.670 ;
        RECT 143.000 137.810 143.320 137.870 ;
        RECT 144.840 137.810 145.160 137.870 ;
        RECT 143.000 137.670 145.160 137.810 ;
        RECT 143.000 137.610 143.320 137.670 ;
        RECT 144.840 137.610 145.160 137.670 ;
        RECT 148.980 137.810 149.300 137.870 ;
        RECT 149.915 137.810 150.205 137.855 ;
        RECT 148.980 137.670 150.205 137.810 ;
        RECT 151.830 137.810 151.970 137.965 ;
        RECT 152.200 137.950 152.520 138.210 ;
        RECT 153.120 137.810 153.440 137.870 ;
        RECT 151.830 137.670 153.440 137.810 ;
        RECT 148.980 137.610 149.300 137.670 ;
        RECT 149.915 137.625 150.205 137.670 ;
        RECT 153.120 137.610 153.440 137.670 ;
        RECT 126.900 137.330 133.570 137.470 ;
        RECT 138.030 137.330 139.550 137.470 ;
        RECT 140.700 137.470 141.020 137.530 ;
        RECT 148.535 137.470 148.825 137.515 ;
        RECT 140.700 137.330 148.825 137.470 ;
        RECT 126.900 137.270 127.220 137.330 ;
        RECT 129.675 137.285 129.965 137.330 ;
        RECT 138.030 137.190 138.170 137.330 ;
        RECT 140.700 137.270 141.020 137.330 ;
        RECT 148.535 137.285 148.825 137.330 ;
        RECT 120.000 137.130 120.320 137.190 ;
        RECT 107.670 136.990 120.320 137.130 ;
        RECT 102.060 136.930 102.380 136.990 ;
        RECT 105.755 136.945 106.045 136.990 ;
        RECT 107.120 136.930 107.440 136.990 ;
        RECT 120.000 136.930 120.320 136.990 ;
        RECT 123.220 137.130 123.540 137.190 ;
        RECT 125.995 137.130 126.285 137.175 ;
        RECT 123.220 136.990 126.285 137.130 ;
        RECT 123.220 136.930 123.540 136.990 ;
        RECT 125.995 136.945 126.285 136.990 ;
        RECT 129.200 137.130 129.520 137.190 ;
        RECT 130.595 137.130 130.885 137.175 ;
        RECT 129.200 136.990 130.885 137.130 ;
        RECT 129.200 136.930 129.520 136.990 ;
        RECT 130.595 136.945 130.885 136.990 ;
        RECT 136.575 137.130 136.865 137.175 ;
        RECT 137.480 137.130 137.800 137.190 ;
        RECT 136.575 136.990 137.800 137.130 ;
        RECT 136.575 136.945 136.865 136.990 ;
        RECT 137.480 136.930 137.800 136.990 ;
        RECT 137.940 136.930 138.260 137.190 ;
        RECT 141.160 136.930 141.480 137.190 ;
        RECT 151.740 137.130 152.060 137.190 ;
        RECT 152.215 137.130 152.505 137.175 ;
        RECT 151.740 136.990 152.505 137.130 ;
        RECT 151.740 136.930 152.060 136.990 ;
        RECT 152.215 136.945 152.505 136.990 ;
        RECT 154.055 137.130 154.345 137.175 ;
        RECT 154.055 136.990 156.570 137.130 ;
        RECT 154.055 136.945 154.345 136.990 ;
        RECT 70.710 136.310 156.270 136.790 ;
        RECT 78.600 135.910 78.920 136.170 ;
        RECT 79.520 135.910 79.840 136.170 ;
        RECT 79.980 135.910 80.300 136.170 ;
        RECT 91.940 135.910 92.260 136.170 ;
        RECT 102.060 136.110 102.380 136.170 ;
        RECT 94.330 135.970 97.230 136.110 ;
        RECT 78.690 135.770 78.830 135.910 ;
        RECT 76.850 135.630 78.830 135.770 ;
        RECT 76.850 135.475 76.990 135.630 ;
        RECT 76.775 135.245 77.065 135.475 ;
        RECT 79.610 135.430 79.750 135.910 ;
        RECT 78.690 135.290 79.750 135.430 ;
        RECT 78.690 135.135 78.830 135.290 ;
        RECT 76.315 134.905 76.605 135.135 ;
        RECT 78.615 134.905 78.905 135.135 ;
        RECT 79.535 135.090 79.825 135.135 ;
        RECT 80.070 135.090 80.210 135.910 ;
        RECT 87.815 135.430 88.105 135.475 ;
        RECT 89.180 135.430 89.500 135.490 ;
        RECT 92.030 135.430 92.170 135.910 ;
        RECT 86.510 135.290 89.500 135.430 ;
        RECT 86.510 135.135 86.650 135.290 ;
        RECT 87.815 135.245 88.105 135.290 ;
        RECT 89.180 135.230 89.500 135.290 ;
        RECT 91.110 135.290 92.170 135.430 ;
        RECT 79.535 134.950 80.210 135.090 ;
        RECT 79.535 134.905 79.825 134.950 ;
        RECT 86.435 134.905 86.725 135.135 ;
        RECT 87.355 135.090 87.645 135.135 ;
        RECT 88.735 135.090 89.025 135.135 ;
        RECT 90.100 135.090 90.420 135.150 ;
        RECT 91.110 135.135 91.250 135.290 ;
        RECT 94.330 135.150 94.470 135.970 ;
        RECT 96.540 135.570 96.860 135.830 ;
        RECT 96.630 135.430 96.770 135.570 ;
        RECT 95.250 135.290 96.770 135.430 ;
        RECT 87.355 134.950 90.420 135.090 ;
        RECT 87.355 134.905 87.645 134.950 ;
        RECT 88.735 134.905 89.025 134.950 ;
        RECT 76.390 134.750 76.530 134.905 ;
        RECT 90.100 134.890 90.420 134.950 ;
        RECT 91.035 134.905 91.325 135.135 ;
        RECT 91.495 134.905 91.785 135.135 ;
        RECT 81.820 134.750 82.140 134.810 ;
        RECT 76.390 134.610 82.140 134.750 ;
        RECT 81.820 134.550 82.140 134.610 ;
        RECT 88.260 134.750 88.580 134.810 ;
        RECT 91.570 134.750 91.710 134.905 ;
        RECT 94.240 134.890 94.560 135.150 ;
        RECT 95.250 135.135 95.390 135.290 ;
        RECT 95.175 134.905 95.465 135.135 ;
        RECT 96.540 134.890 96.860 135.150 ;
        RECT 97.090 135.135 97.230 135.970 ;
        RECT 100.310 135.970 102.380 136.110 ;
        RECT 97.015 134.905 97.305 135.135 ;
        RECT 97.460 134.890 97.780 135.150 ;
        RECT 97.920 135.135 98.240 135.150 ;
        RECT 97.920 134.905 98.355 135.135 ;
        RECT 98.855 135.090 99.145 135.135 ;
        RECT 99.300 135.090 99.620 135.150 ;
        RECT 98.855 134.950 99.620 135.090 ;
        RECT 98.855 134.905 99.145 134.950 ;
        RECT 97.920 134.890 98.240 134.905 ;
        RECT 99.300 134.890 99.620 134.950 ;
        RECT 99.760 134.890 100.080 135.150 ;
        RECT 100.310 135.135 100.450 135.970 ;
        RECT 102.060 135.910 102.380 135.970 ;
        RECT 102.980 135.910 103.300 136.170 ;
        RECT 103.915 136.110 104.205 136.155 ;
        RECT 104.360 136.110 104.680 136.170 ;
        RECT 103.915 135.970 104.680 136.110 ;
        RECT 103.915 135.925 104.205 135.970 ;
        RECT 104.360 135.910 104.680 135.970 ;
        RECT 107.120 135.910 107.440 136.170 ;
        RECT 113.100 135.910 113.420 136.170 ;
        RECT 114.020 136.110 114.340 136.170 ;
        RECT 118.160 136.110 118.480 136.170 ;
        RECT 126.900 136.110 127.220 136.170 ;
        RECT 140.700 136.110 141.020 136.170 ;
        RECT 114.020 135.970 117.470 136.110 ;
        RECT 114.020 135.910 114.340 135.970 ;
        RECT 100.680 135.770 101.000 135.830 ;
        RECT 100.680 135.630 101.370 135.770 ;
        RECT 100.680 135.570 101.000 135.630 ;
        RECT 101.230 135.475 101.370 135.630 ;
        RECT 101.195 135.245 101.485 135.475 ;
        RECT 103.070 135.430 103.210 135.910 ;
        RECT 104.450 135.430 104.590 135.910 ;
        RECT 106.215 135.430 106.505 135.475 ;
        RECT 107.210 135.430 107.350 135.910 ;
        RECT 103.070 135.290 104.130 135.430 ;
        RECT 104.450 135.290 105.970 135.430 ;
        RECT 100.235 134.905 100.525 135.135 ;
        RECT 100.695 134.905 100.985 135.135 ;
        RECT 102.995 135.090 103.285 135.135 ;
        RECT 103.440 135.090 103.760 135.150 ;
        RECT 102.995 134.950 103.760 135.090 ;
        RECT 102.995 134.905 103.285 134.950 ;
        RECT 88.260 134.610 91.710 134.750 ;
        RECT 94.715 134.750 95.005 134.795 ;
        RECT 94.715 134.610 99.990 134.750 ;
        RECT 88.260 134.550 88.580 134.610 ;
        RECT 94.715 134.565 95.005 134.610 ;
        RECT 78.140 134.210 78.460 134.470 ;
        RECT 86.880 134.210 87.200 134.470 ;
        RECT 89.180 134.410 89.500 134.470 ;
        RECT 89.655 134.410 89.945 134.455 ;
        RECT 89.180 134.270 89.945 134.410 ;
        RECT 89.180 134.210 89.500 134.270 ;
        RECT 89.655 134.225 89.945 134.270 ;
        RECT 90.115 134.410 90.405 134.455 ;
        RECT 91.940 134.410 92.260 134.470 ;
        RECT 90.115 134.270 92.260 134.410 ;
        RECT 90.115 134.225 90.405 134.270 ;
        RECT 91.940 134.210 92.260 134.270 ;
        RECT 95.635 134.410 95.925 134.455 ;
        RECT 98.840 134.410 99.160 134.470 ;
        RECT 95.635 134.270 99.160 134.410 ;
        RECT 99.850 134.410 99.990 134.610 ;
        RECT 100.770 134.410 100.910 134.905 ;
        RECT 103.440 134.890 103.760 134.950 ;
        RECT 99.850 134.270 100.910 134.410 ;
        RECT 102.075 134.410 102.365 134.455 ;
        RECT 102.980 134.410 103.300 134.470 ;
        RECT 102.075 134.270 103.300 134.410 ;
        RECT 103.990 134.410 104.130 135.290 ;
        RECT 104.360 135.090 104.680 135.150 ;
        RECT 105.830 135.090 105.970 135.290 ;
        RECT 106.215 135.290 107.350 135.430 ;
        RECT 107.595 135.430 107.885 135.475 ;
        RECT 113.190 135.430 113.330 135.910 ;
        RECT 107.595 135.290 108.270 135.430 ;
        RECT 113.190 135.290 116.550 135.430 ;
        RECT 106.215 135.245 106.505 135.290 ;
        RECT 107.595 135.245 107.885 135.290 ;
        RECT 108.130 135.150 108.270 135.290 ;
        RECT 106.675 135.090 106.965 135.135 ;
        RECT 104.360 134.950 105.510 135.090 ;
        RECT 105.830 134.950 106.965 135.090 ;
        RECT 104.360 134.890 104.680 134.950 ;
        RECT 105.370 134.750 105.510 134.950 ;
        RECT 106.675 134.905 106.965 134.950 ;
        RECT 107.120 134.890 107.440 135.150 ;
        RECT 108.040 135.090 108.360 135.150 ;
        RECT 116.410 135.135 116.550 135.290 ;
        RECT 116.780 135.230 117.100 135.490 ;
        RECT 117.330 135.475 117.470 135.970 ;
        RECT 118.160 135.970 127.220 136.110 ;
        RECT 118.160 135.910 118.480 135.970 ;
        RECT 126.900 135.910 127.220 135.970 ;
        RECT 128.340 135.970 141.020 136.110 ;
        RECT 117.255 135.245 117.545 135.475 ;
        RECT 128.340 135.430 128.480 135.970 ;
        RECT 140.700 135.910 141.020 135.970 ;
        RECT 148.520 135.910 148.840 136.170 ;
        RECT 148.980 136.110 149.300 136.170 ;
        RECT 152.215 136.110 152.505 136.155 ;
        RECT 148.980 135.970 152.505 136.110 ;
        RECT 148.980 135.910 149.300 135.970 ;
        RECT 152.215 135.925 152.505 135.970 ;
        RECT 132.420 135.770 132.740 135.830 ;
        RECT 136.560 135.770 136.880 135.830 ;
        RECT 132.420 135.630 136.880 135.770 ;
        RECT 132.420 135.570 132.740 135.630 ;
        RECT 136.560 135.570 136.880 135.630 ;
        RECT 137.480 135.570 137.800 135.830 ;
        RECT 143.000 135.770 143.320 135.830 ;
        RECT 139.410 135.630 143.320 135.770 ;
        RECT 130.580 135.430 130.900 135.490 ;
        RECT 127.910 135.290 128.480 135.430 ;
        RECT 129.290 135.290 130.900 135.430 ;
        RECT 115.875 135.090 116.165 135.135 ;
        RECT 108.040 134.950 116.165 135.090 ;
        RECT 108.040 134.890 108.360 134.950 ;
        RECT 115.875 134.905 116.165 134.950 ;
        RECT 116.335 134.905 116.625 135.135 ;
        RECT 123.220 134.890 123.540 135.150 ;
        RECT 126.900 134.890 127.220 135.150 ;
        RECT 127.910 135.135 128.050 135.290 ;
        RECT 127.835 134.905 128.125 135.135 ;
        RECT 128.280 134.890 128.600 135.150 ;
        RECT 129.290 135.135 129.430 135.290 ;
        RECT 130.580 135.230 130.900 135.290 ;
        RECT 132.880 135.430 133.200 135.490 ;
        RECT 135.655 135.430 135.945 135.475 ;
        RECT 132.880 135.290 135.945 135.430 ;
        RECT 132.880 135.230 133.200 135.290 ;
        RECT 135.655 135.245 135.945 135.290 ;
        RECT 137.020 135.230 137.340 135.490 ;
        RECT 137.570 135.430 137.710 135.570 ;
        RECT 137.955 135.430 138.245 135.475 ;
        RECT 139.410 135.430 139.550 135.630 ;
        RECT 143.000 135.570 143.320 135.630 ;
        RECT 145.775 135.430 146.065 135.475 ;
        RECT 148.610 135.430 148.750 135.910 ;
        RECT 137.570 135.290 138.245 135.430 ;
        RECT 137.955 135.245 138.245 135.290 ;
        RECT 138.490 135.290 139.550 135.430 ;
        RECT 139.870 135.290 148.750 135.430 ;
        RECT 129.215 134.905 129.505 135.135 ;
        RECT 129.675 134.905 129.965 135.135 ;
        RECT 133.815 134.905 134.105 135.135 ;
        RECT 134.720 135.090 135.040 135.150 ;
        RECT 136.575 135.090 136.865 135.135 ;
        RECT 134.720 134.950 136.865 135.090 ;
        RECT 123.310 134.750 123.450 134.890 ;
        RECT 129.750 134.750 129.890 134.905 ;
        RECT 133.890 134.750 134.030 134.905 ;
        RECT 134.720 134.890 135.040 134.950 ;
        RECT 136.575 134.905 136.865 134.950 ;
        RECT 137.495 135.090 137.785 135.135 ;
        RECT 138.490 135.090 138.630 135.290 ;
        RECT 139.870 135.090 140.010 135.290 ;
        RECT 145.775 135.245 146.065 135.290 ;
        RECT 152.200 135.230 152.520 135.490 ;
        RECT 153.135 135.430 153.425 135.475 ;
        RECT 156.430 135.430 156.570 136.990 ;
        RECT 153.135 135.290 156.570 135.430 ;
        RECT 153.135 135.245 153.425 135.290 ;
        RECT 141.620 135.090 141.940 135.150 ;
        RECT 137.495 134.950 138.630 135.090 ;
        RECT 138.950 134.950 140.010 135.090 ;
        RECT 140.330 134.950 141.940 135.090 ;
        RECT 137.495 134.905 137.785 134.950 ;
        RECT 138.950 134.750 139.090 134.950 ;
        RECT 105.370 134.610 116.320 134.750 ;
        RECT 123.310 134.610 129.890 134.750 ;
        RECT 133.430 134.610 139.090 134.750 ;
        RECT 139.795 134.750 140.085 134.795 ;
        RECT 140.330 134.750 140.470 134.950 ;
        RECT 141.620 134.890 141.940 134.950 ;
        RECT 144.380 134.890 144.700 135.150 ;
        RECT 148.520 135.090 148.840 135.150 ;
        RECT 149.915 135.090 150.205 135.135 ;
        RECT 148.520 134.950 150.205 135.090 ;
        RECT 148.520 134.890 148.840 134.950 ;
        RECT 149.915 134.905 150.205 134.950 ;
        RECT 151.755 135.090 152.045 135.135 ;
        RECT 152.290 135.090 152.430 135.230 ;
        RECT 151.755 134.950 152.430 135.090 ;
        RECT 151.755 134.905 152.045 134.950 ;
        RECT 153.580 134.890 153.900 135.150 ;
        RECT 154.515 134.905 154.805 135.135 ;
        RECT 139.795 134.610 140.470 134.750 ;
        RECT 105.295 134.410 105.585 134.455 ;
        RECT 108.040 134.410 108.360 134.470 ;
        RECT 103.990 134.270 108.360 134.410 ;
        RECT 95.635 134.225 95.925 134.270 ;
        RECT 98.840 134.210 99.160 134.270 ;
        RECT 102.075 134.225 102.365 134.270 ;
        RECT 102.980 134.210 103.300 134.270 ;
        RECT 105.295 134.225 105.585 134.270 ;
        RECT 108.040 134.210 108.360 134.270 ;
        RECT 108.500 134.210 108.820 134.470 ;
        RECT 114.940 134.210 115.260 134.470 ;
        RECT 116.180 134.410 116.320 134.610 ;
        RECT 133.430 134.410 133.570 134.610 ;
        RECT 139.795 134.565 140.085 134.610 ;
        RECT 140.715 134.565 141.005 134.795 ;
        RECT 144.470 134.750 144.610 134.890 ;
        RECT 152.660 134.750 152.980 134.810 ;
        RECT 144.470 134.610 152.980 134.750 ;
        RECT 116.180 134.270 133.570 134.410 ;
        RECT 133.800 134.410 134.120 134.470 ;
        RECT 134.720 134.410 135.040 134.470 ;
        RECT 133.800 134.270 135.040 134.410 ;
        RECT 133.800 134.210 134.120 134.270 ;
        RECT 134.720 134.210 135.040 134.270 ;
        RECT 138.860 134.210 139.180 134.470 ;
        RECT 139.320 134.410 139.640 134.470 ;
        RECT 140.790 134.410 140.930 134.565 ;
        RECT 152.660 134.550 152.980 134.610 ;
        RECT 153.135 134.750 153.425 134.795 ;
        RECT 154.040 134.750 154.360 134.810 ;
        RECT 154.590 134.750 154.730 134.905 ;
        RECT 153.135 134.610 154.730 134.750 ;
        RECT 153.135 134.565 153.425 134.610 ;
        RECT 154.040 134.550 154.360 134.610 ;
        RECT 142.540 134.410 142.860 134.470 ;
        RECT 139.320 134.270 142.860 134.410 ;
        RECT 139.320 134.210 139.640 134.270 ;
        RECT 142.540 134.210 142.860 134.270 ;
        RECT 143.460 134.410 143.780 134.470 ;
        RECT 145.760 134.410 146.080 134.470 ;
        RECT 143.460 134.270 146.080 134.410 ;
        RECT 143.460 134.210 143.780 134.270 ;
        RECT 145.760 134.210 146.080 134.270 ;
        RECT 150.835 134.410 151.125 134.455 ;
        RECT 151.740 134.410 152.060 134.470 ;
        RECT 150.835 134.270 152.060 134.410 ;
        RECT 150.835 134.225 151.125 134.270 ;
        RECT 151.740 134.210 152.060 134.270 ;
        RECT 154.500 134.210 154.820 134.470 ;
        RECT 70.710 133.590 156.270 134.070 ;
        RECT 84.135 133.390 84.425 133.435 ;
        RECT 85.040 133.390 85.360 133.450 ;
        RECT 90.100 133.390 90.420 133.450 ;
        RECT 84.135 133.250 90.420 133.390 ;
        RECT 84.135 133.205 84.425 133.250 ;
        RECT 85.040 133.190 85.360 133.250 ;
        RECT 90.100 133.190 90.420 133.250 ;
        RECT 97.000 133.190 97.320 133.450 ;
        RECT 111.260 133.390 111.580 133.450 ;
        RECT 98.010 133.250 111.580 133.390 ;
        RECT 83.675 133.050 83.965 133.095 ;
        RECT 85.960 133.050 86.280 133.110 ;
        RECT 83.675 132.910 86.280 133.050 ;
        RECT 83.675 132.865 83.965 132.910 ;
        RECT 85.960 132.850 86.280 132.910 ;
        RECT 98.010 132.770 98.150 133.250 ;
        RECT 111.260 133.190 111.580 133.250 ;
        RECT 123.695 133.390 123.985 133.435 ;
        RECT 124.140 133.390 124.460 133.450 ;
        RECT 123.695 133.250 124.460 133.390 ;
        RECT 123.695 133.205 123.985 133.250 ;
        RECT 124.140 133.190 124.460 133.250 ;
        RECT 141.620 133.390 141.940 133.450 ;
        RECT 148.980 133.390 149.300 133.450 ;
        RECT 149.535 133.390 149.825 133.435 ;
        RECT 153.580 133.390 153.900 133.450 ;
        RECT 141.620 133.250 148.750 133.390 ;
        RECT 141.620 133.190 141.940 133.250 ;
        RECT 103.440 133.050 103.760 133.110 ;
        RECT 105.295 133.050 105.585 133.095 ;
        RECT 103.440 132.910 105.585 133.050 ;
        RECT 103.440 132.850 103.760 132.910 ;
        RECT 105.295 132.865 105.585 132.910 ;
        RECT 106.200 133.050 106.520 133.110 ;
        RECT 108.960 133.050 109.280 133.110 ;
        RECT 106.200 132.910 109.280 133.050 ;
        RECT 106.200 132.850 106.520 132.910 ;
        RECT 108.960 132.850 109.280 132.910 ;
        RECT 109.420 132.850 109.740 133.110 ;
        RECT 123.235 133.050 123.525 133.095 ;
        RECT 129.660 133.050 129.980 133.110 ;
        RECT 131.500 133.050 131.820 133.110 ;
        RECT 137.940 133.050 138.260 133.110 ;
        RECT 143.000 133.050 143.320 133.110 ;
        RECT 113.650 132.910 124.830 133.050 ;
        RECT 73.095 132.710 73.385 132.755 ;
        RECT 76.760 132.710 77.080 132.770 ;
        RECT 73.095 132.570 77.080 132.710 ;
        RECT 73.095 132.525 73.385 132.570 ;
        RECT 76.760 132.510 77.080 132.570 ;
        RECT 82.740 132.710 83.060 132.770 ;
        RECT 83.215 132.710 83.505 132.755 ;
        RECT 82.740 132.570 83.505 132.710 ;
        RECT 82.740 132.510 83.060 132.570 ;
        RECT 83.215 132.525 83.505 132.570 ;
        RECT 85.055 132.710 85.345 132.755 ;
        RECT 86.420 132.710 86.740 132.770 ;
        RECT 85.055 132.570 86.740 132.710 ;
        RECT 85.055 132.525 85.345 132.570 ;
        RECT 86.420 132.510 86.740 132.570 ;
        RECT 86.880 132.710 87.200 132.770 ;
        RECT 88.275 132.710 88.565 132.755 ;
        RECT 86.880 132.570 88.565 132.710 ;
        RECT 86.880 132.510 87.200 132.570 ;
        RECT 88.275 132.525 88.565 132.570 ;
        RECT 89.180 132.510 89.500 132.770 ;
        RECT 97.920 132.510 98.240 132.770 ;
        RECT 98.840 132.510 99.160 132.770 ;
        RECT 100.695 132.710 100.985 132.755 ;
        RECT 104.360 132.710 104.680 132.770 ;
        RECT 100.695 132.570 104.680 132.710 ;
        RECT 100.695 132.525 100.985 132.570 ;
        RECT 104.360 132.510 104.680 132.570 ;
        RECT 73.555 132.370 73.845 132.415 ;
        RECT 85.500 132.370 85.820 132.430 ;
        RECT 73.555 132.230 85.820 132.370 ;
        RECT 73.555 132.185 73.845 132.230 ;
        RECT 85.500 132.170 85.820 132.230 ;
        RECT 99.315 132.370 99.605 132.415 ;
        RECT 102.060 132.370 102.380 132.430 ;
        RECT 109.510 132.370 109.650 132.850 ;
        RECT 113.100 132.510 113.420 132.770 ;
        RECT 113.650 132.755 113.790 132.910 ;
        RECT 123.235 132.865 123.525 132.910 ;
        RECT 113.575 132.525 113.865 132.755 ;
        RECT 114.480 132.510 114.800 132.770 ;
        RECT 114.955 132.710 115.245 132.755 ;
        RECT 120.920 132.710 121.240 132.770 ;
        RECT 124.140 132.710 124.460 132.770 ;
        RECT 124.690 132.755 124.830 132.910 ;
        RECT 129.660 132.910 130.350 133.050 ;
        RECT 129.660 132.850 129.980 132.910 ;
        RECT 130.210 132.755 130.350 132.910 ;
        RECT 131.130 132.910 140.010 133.050 ;
        RECT 114.955 132.570 116.320 132.710 ;
        RECT 114.955 132.525 115.245 132.570 ;
        RECT 116.180 132.370 116.320 132.570 ;
        RECT 120.920 132.570 124.460 132.710 ;
        RECT 120.920 132.510 121.240 132.570 ;
        RECT 124.140 132.510 124.460 132.570 ;
        RECT 124.615 132.525 124.905 132.755 ;
        RECT 130.090 132.525 130.380 132.755 ;
        RECT 123.220 132.370 123.540 132.430 ;
        RECT 99.315 132.230 102.380 132.370 ;
        RECT 99.315 132.185 99.605 132.230 ;
        RECT 102.060 132.170 102.380 132.230 ;
        RECT 102.610 132.230 109.190 132.370 ;
        RECT 109.510 132.230 113.330 132.370 ;
        RECT 116.180 132.230 123.540 132.370 ;
        RECT 74.935 132.030 75.225 132.075 ;
        RECT 76.760 132.030 77.080 132.090 ;
        RECT 74.935 131.890 77.080 132.030 ;
        RECT 74.935 131.845 75.225 131.890 ;
        RECT 76.760 131.830 77.080 131.890 ;
        RECT 84.120 132.030 84.440 132.090 ;
        RECT 89.640 132.030 89.960 132.090 ;
        RECT 96.540 132.030 96.860 132.090 ;
        RECT 99.775 132.030 100.065 132.075 ;
        RECT 84.120 131.890 100.065 132.030 ;
        RECT 84.120 131.830 84.440 131.890 ;
        RECT 89.640 131.830 89.960 131.890 ;
        RECT 96.540 131.830 96.860 131.890 ;
        RECT 99.775 131.845 100.065 131.890 ;
        RECT 84.580 131.490 84.900 131.750 ;
        RECT 88.260 131.490 88.580 131.750 ;
        RECT 95.620 131.690 95.940 131.750 ;
        RECT 102.610 131.690 102.750 132.230 ;
        RECT 102.980 132.030 103.300 132.090 ;
        RECT 108.040 132.030 108.360 132.090 ;
        RECT 102.980 131.890 108.360 132.030 ;
        RECT 109.050 132.030 109.190 132.230 ;
        RECT 113.190 132.090 113.330 132.230 ;
        RECT 123.220 132.170 123.540 132.230 ;
        RECT 109.050 131.890 112.870 132.030 ;
        RECT 102.980 131.830 103.300 131.890 ;
        RECT 108.040 131.830 108.360 131.890 ;
        RECT 95.620 131.550 102.750 131.690 ;
        RECT 95.620 131.490 95.940 131.550 ;
        RECT 104.360 131.490 104.680 131.750 ;
        RECT 112.180 131.490 112.500 131.750 ;
        RECT 112.730 131.690 112.870 131.890 ;
        RECT 113.100 131.830 113.420 132.090 ;
        RECT 120.920 132.030 121.240 132.090 ;
        RECT 116.180 131.890 121.240 132.030 ;
        RECT 124.690 132.030 124.830 132.525 ;
        RECT 130.580 132.510 130.900 132.770 ;
        RECT 131.130 132.370 131.270 132.910 ;
        RECT 131.500 132.850 131.820 132.910 ;
        RECT 137.940 132.850 138.260 132.910 ;
        RECT 131.975 132.700 132.265 132.755 ;
        RECT 129.750 132.230 131.270 132.370 ;
        RECT 131.590 132.560 132.265 132.700 ;
        RECT 128.280 132.030 128.600 132.090 ;
        RECT 129.215 132.030 129.505 132.075 ;
        RECT 124.690 131.890 129.505 132.030 ;
        RECT 116.180 131.690 116.320 131.890 ;
        RECT 120.920 131.830 121.240 131.890 ;
        RECT 128.280 131.830 128.600 131.890 ;
        RECT 129.215 131.845 129.505 131.890 ;
        RECT 112.730 131.550 116.320 131.690 ;
        RECT 116.780 131.690 117.100 131.750 ;
        RECT 125.535 131.690 125.825 131.735 ;
        RECT 129.750 131.690 129.890 132.230 ;
        RECT 130.120 132.030 130.440 132.090 ;
        RECT 131.590 132.030 131.730 132.560 ;
        RECT 131.975 132.525 132.265 132.560 ;
        RECT 139.320 132.510 139.640 132.770 ;
        RECT 139.870 132.710 140.010 132.910 ;
        RECT 141.710 132.910 143.320 133.050 ;
        RECT 140.210 132.710 140.500 132.755 ;
        RECT 139.870 132.570 140.500 132.710 ;
        RECT 140.210 132.525 140.500 132.570 ;
        RECT 140.700 132.510 141.020 132.770 ;
        RECT 141.710 132.755 141.850 132.910 ;
        RECT 143.000 132.850 143.320 132.910 ;
        RECT 143.920 133.050 144.240 133.110 ;
        RECT 148.610 133.095 148.750 133.250 ;
        RECT 148.980 133.250 149.825 133.390 ;
        RECT 148.980 133.190 149.300 133.250 ;
        RECT 149.535 133.205 149.825 133.250 ;
        RECT 149.990 133.250 153.900 133.390 ;
        RECT 148.535 133.050 148.825 133.095 ;
        RECT 149.990 133.050 150.130 133.250 ;
        RECT 153.580 133.190 153.900 133.250 ;
        RECT 143.920 132.910 146.450 133.050 ;
        RECT 143.920 132.850 144.240 132.910 ;
        RECT 141.635 132.525 141.925 132.755 ;
        RECT 142.540 132.510 142.860 132.770 ;
        RECT 143.475 132.525 143.765 132.755 ;
        RECT 144.395 132.525 144.685 132.755 ;
        RECT 139.795 132.370 140.085 132.415 ;
        RECT 142.095 132.370 142.385 132.415 ;
        RECT 139.795 132.230 142.385 132.370 ;
        RECT 139.795 132.185 140.085 132.230 ;
        RECT 142.095 132.185 142.385 132.230 ;
        RECT 130.120 131.890 131.730 132.030 ;
        RECT 131.960 132.030 132.280 132.090 ;
        RECT 132.895 132.030 133.185 132.075 ;
        RECT 131.960 131.890 133.185 132.030 ;
        RECT 143.550 132.030 143.690 132.525 ;
        RECT 144.470 132.370 144.610 132.525 ;
        RECT 144.840 132.510 145.160 132.770 ;
        RECT 145.760 132.510 146.080 132.770 ;
        RECT 146.310 132.755 146.450 132.910 ;
        RECT 148.535 132.910 150.130 133.050 ;
        RECT 153.135 133.050 153.425 133.095 ;
        RECT 155.420 133.050 155.740 133.110 ;
        RECT 153.135 132.910 155.740 133.050 ;
        RECT 148.535 132.865 148.825 132.910 ;
        RECT 153.135 132.865 153.425 132.910 ;
        RECT 154.590 132.755 154.730 132.910 ;
        RECT 155.420 132.850 155.740 132.910 ;
        RECT 155.880 132.850 156.200 133.110 ;
        RECT 146.235 132.525 146.525 132.755 ;
        RECT 152.215 132.710 152.505 132.755 ;
        RECT 153.595 132.710 153.885 132.755 ;
        RECT 152.215 132.570 153.885 132.710 ;
        RECT 152.215 132.525 152.505 132.570 ;
        RECT 153.595 132.525 153.885 132.570 ;
        RECT 154.515 132.525 154.805 132.755 ;
        RECT 145.315 132.370 145.605 132.415 ;
        RECT 144.470 132.230 145.605 132.370 ;
        RECT 153.670 132.370 153.810 132.525 ;
        RECT 155.970 132.370 156.110 132.850 ;
        RECT 153.670 132.230 156.110 132.370 ;
        RECT 145.315 132.185 145.605 132.230 ;
        RECT 145.760 132.030 146.080 132.090 ;
        RECT 155.420 132.030 155.740 132.090 ;
        RECT 143.550 131.890 145.070 132.030 ;
        RECT 130.120 131.830 130.440 131.890 ;
        RECT 131.960 131.830 132.280 131.890 ;
        RECT 132.895 131.845 133.185 131.890 ;
        RECT 116.780 131.550 129.890 131.690 ;
        RECT 131.515 131.690 131.805 131.735 ;
        RECT 137.940 131.690 138.260 131.750 ;
        RECT 131.515 131.550 138.260 131.690 ;
        RECT 116.780 131.490 117.100 131.550 ;
        RECT 125.535 131.505 125.825 131.550 ;
        RECT 131.515 131.505 131.805 131.550 ;
        RECT 137.940 131.490 138.260 131.550 ;
        RECT 138.415 131.690 138.705 131.735 ;
        RECT 139.320 131.690 139.640 131.750 ;
        RECT 138.415 131.550 139.640 131.690 ;
        RECT 138.415 131.505 138.705 131.550 ;
        RECT 139.320 131.490 139.640 131.550 ;
        RECT 140.700 131.690 141.020 131.750 ;
        RECT 141.620 131.690 141.940 131.750 ;
        RECT 140.700 131.550 141.940 131.690 ;
        RECT 140.700 131.490 141.020 131.550 ;
        RECT 141.620 131.490 141.940 131.550 ;
        RECT 144.380 131.490 144.700 131.750 ;
        RECT 144.930 131.690 145.070 131.890 ;
        RECT 145.760 131.890 155.740 132.030 ;
        RECT 145.760 131.830 146.080 131.890 ;
        RECT 155.420 131.830 155.740 131.890 ;
        RECT 145.300 131.690 145.620 131.750 ;
        RECT 144.930 131.550 145.620 131.690 ;
        RECT 145.300 131.490 145.620 131.550 ;
        RECT 147.140 131.490 147.460 131.750 ;
        RECT 148.060 131.690 148.380 131.750 ;
        RECT 149.455 131.690 149.745 131.735 ;
        RECT 149.900 131.690 150.220 131.750 ;
        RECT 148.060 131.550 150.220 131.690 ;
        RECT 148.060 131.490 148.380 131.550 ;
        RECT 149.455 131.505 149.745 131.550 ;
        RECT 149.900 131.490 150.220 131.550 ;
        RECT 150.360 131.490 150.680 131.750 ;
        RECT 151.295 131.690 151.585 131.735 ;
        RECT 152.200 131.690 152.520 131.750 ;
        RECT 151.295 131.550 152.520 131.690 ;
        RECT 151.295 131.505 151.585 131.550 ;
        RECT 152.200 131.490 152.520 131.550 ;
        RECT 70.710 130.870 156.270 131.350 ;
        RECT 76.760 130.470 77.080 130.730 ;
        RECT 84.580 130.670 84.900 130.730 ;
        RECT 85.055 130.670 85.345 130.715 ;
        RECT 84.580 130.530 85.345 130.670 ;
        RECT 84.580 130.470 84.900 130.530 ;
        RECT 85.055 130.485 85.345 130.530 ;
        RECT 85.590 130.530 91.250 130.670 ;
        RECT 75.395 129.990 75.685 130.035 ;
        RECT 76.850 129.990 76.990 130.470 ;
        RECT 85.590 130.390 85.730 130.530 ;
        RECT 78.140 130.130 78.460 130.390 ;
        RECT 85.500 130.130 85.820 130.390 ;
        RECT 85.975 130.330 86.265 130.375 ;
        RECT 90.560 130.330 90.880 130.390 ;
        RECT 85.975 130.190 90.880 130.330 ;
        RECT 85.975 130.145 86.265 130.190 ;
        RECT 90.560 130.130 90.880 130.190 ;
        RECT 75.395 129.850 76.990 129.990 ;
        RECT 75.395 129.805 75.685 129.850 ;
        RECT 74.935 129.650 75.225 129.695 ;
        RECT 77.220 129.650 77.540 129.710 ;
        RECT 74.935 129.510 77.540 129.650 ;
        RECT 74.935 129.465 75.225 129.510 ;
        RECT 77.220 129.450 77.540 129.510 ;
        RECT 77.680 129.450 78.000 129.710 ;
        RECT 78.230 129.650 78.370 130.130 ;
        RECT 89.180 129.990 89.500 130.050 ;
        RECT 79.610 129.850 85.350 129.990 ;
        RECT 79.610 129.710 79.750 129.850 ;
        RECT 78.615 129.650 78.905 129.695 ;
        RECT 78.230 129.510 78.905 129.650 ;
        RECT 78.615 129.465 78.905 129.510 ;
        RECT 79.075 129.650 79.365 129.695 ;
        RECT 79.520 129.650 79.840 129.710 ;
        RECT 79.075 129.510 79.840 129.650 ;
        RECT 79.075 129.465 79.365 129.510 ;
        RECT 79.520 129.450 79.840 129.510 ;
        RECT 80.455 129.465 80.745 129.695 ;
        RECT 81.360 129.650 81.680 129.710 ;
        RECT 81.835 129.650 82.125 129.695 ;
        RECT 81.360 129.510 82.125 129.650 ;
        RECT 80.530 129.310 80.670 129.465 ;
        RECT 81.360 129.450 81.680 129.510 ;
        RECT 81.835 129.465 82.125 129.510 ;
        RECT 82.755 129.465 83.045 129.695 ;
        RECT 85.210 129.650 85.350 129.850 ;
        RECT 86.510 129.850 89.500 129.990 ;
        RECT 85.500 129.650 85.820 129.710 ;
        RECT 86.510 129.695 86.650 129.850 ;
        RECT 89.180 129.790 89.500 129.850 ;
        RECT 89.640 129.790 89.960 130.050 ;
        RECT 90.100 129.790 90.420 130.050 ;
        RECT 91.110 129.990 91.250 130.530 ;
        RECT 98.380 130.470 98.700 130.730 ;
        RECT 121.380 130.670 121.700 130.730 ;
        RECT 121.855 130.670 122.145 130.715 ;
        RECT 128.280 130.670 128.600 130.730 ;
        RECT 99.390 130.530 111.490 130.670 ;
        RECT 91.480 130.330 91.800 130.390 ;
        RECT 94.255 130.330 94.545 130.375 ;
        RECT 91.480 130.190 94.545 130.330 ;
        RECT 91.480 130.130 91.800 130.190 ;
        RECT 94.255 130.145 94.545 130.190 ;
        RECT 94.700 130.130 95.020 130.390 ;
        RECT 97.460 129.990 97.780 130.050 ;
        RECT 99.390 129.990 99.530 130.530 ;
        RECT 111.350 130.390 111.490 130.530 ;
        RECT 115.950 130.530 128.600 130.670 ;
        RECT 100.220 130.130 100.540 130.390 ;
        RECT 105.740 130.330 106.060 130.390 ;
        RECT 109.420 130.330 109.740 130.390 ;
        RECT 100.770 130.190 109.740 130.330 ;
        RECT 91.110 129.850 91.710 129.990 ;
        RECT 82.830 129.310 82.970 129.465 ;
        RECT 85.210 129.450 85.820 129.650 ;
        RECT 86.435 129.465 86.725 129.695 ;
        RECT 86.880 129.450 87.200 129.710 ;
        RECT 87.340 129.650 87.660 129.710 ;
        RECT 87.815 129.650 88.105 129.695 ;
        RECT 87.340 129.510 88.105 129.650 ;
        RECT 87.340 129.450 87.660 129.510 ;
        RECT 87.815 129.465 88.105 129.510 ;
        RECT 88.260 129.450 88.580 129.710 ;
        RECT 90.190 129.650 90.330 129.790 ;
        RECT 91.570 129.695 91.710 129.850 ;
        RECT 93.870 129.850 99.530 129.990 ;
        RECT 91.035 129.650 91.325 129.695 ;
        RECT 88.810 129.510 89.970 129.650 ;
        RECT 90.190 129.510 91.325 129.650 ;
        RECT 76.850 129.170 80.670 129.310 ;
        RECT 80.990 129.170 82.970 129.310 ;
        RECT 76.850 129.015 76.990 129.170 ;
        RECT 76.775 128.970 77.065 129.015 ;
        RECT 77.220 128.970 77.540 129.030 ;
        RECT 76.775 128.830 77.540 128.970 ;
        RECT 76.775 128.785 77.065 128.830 ;
        RECT 77.220 128.770 77.540 128.830 ;
        RECT 78.615 128.970 78.905 129.015 ;
        RECT 79.535 128.970 79.825 129.015 ;
        RECT 79.980 128.970 80.300 129.030 ;
        RECT 80.990 128.970 81.130 129.170 ;
        RECT 84.120 129.110 84.440 129.370 ;
        RECT 85.210 129.340 85.575 129.450 ;
        RECT 85.285 129.295 85.575 129.340 ;
        RECT 78.615 128.830 81.130 128.970 ;
        RECT 81.375 128.970 81.665 129.015 ;
        RECT 81.820 128.970 82.140 129.030 ;
        RECT 81.375 128.830 82.140 128.970 ;
        RECT 78.615 128.785 78.905 128.830 ;
        RECT 79.535 128.785 79.825 128.830 ;
        RECT 79.980 128.770 80.300 128.830 ;
        RECT 81.375 128.785 81.665 128.830 ;
        RECT 81.820 128.770 82.140 128.830 ;
        RECT 82.740 128.770 83.060 129.030 ;
        RECT 84.580 128.970 84.900 129.030 ;
        RECT 88.810 128.970 88.950 129.510 ;
        RECT 89.830 129.310 89.970 129.510 ;
        RECT 91.035 129.465 91.325 129.510 ;
        RECT 91.495 129.465 91.785 129.695 ;
        RECT 92.860 129.450 93.180 129.710 ;
        RECT 93.870 129.695 94.010 129.850 ;
        RECT 97.460 129.790 97.780 129.850 ;
        RECT 93.795 129.465 94.085 129.695 ;
        RECT 95.175 129.650 95.465 129.695 ;
        RECT 97.920 129.650 98.240 129.710 ;
        RECT 99.390 129.695 99.530 129.850 ;
        RECT 100.770 129.695 100.910 130.190 ;
        RECT 105.740 130.130 106.060 130.190 ;
        RECT 109.420 130.130 109.740 130.190 ;
        RECT 111.260 130.130 111.580 130.390 ;
        RECT 113.560 130.130 113.880 130.390 ;
        RECT 101.600 129.990 101.920 130.050 ;
        RECT 102.535 129.990 102.825 130.035 ;
        RECT 101.600 129.850 102.825 129.990 ;
        RECT 101.600 129.790 101.920 129.850 ;
        RECT 102.535 129.805 102.825 129.850 ;
        RECT 103.455 129.990 103.745 130.035 ;
        RECT 104.360 129.990 104.680 130.050 ;
        RECT 103.455 129.850 104.680 129.990 ;
        RECT 103.455 129.805 103.745 129.850 ;
        RECT 104.360 129.790 104.680 129.850 ;
        RECT 104.835 129.990 105.125 130.035 ;
        RECT 108.960 129.990 109.280 130.050 ;
        RECT 104.835 129.850 109.280 129.990 ;
        RECT 104.835 129.805 105.125 129.850 ;
        RECT 108.960 129.790 109.280 129.850 ;
        RECT 112.640 129.990 112.960 130.050 ;
        RECT 115.950 130.035 116.090 130.530 ;
        RECT 121.380 130.470 121.700 130.530 ;
        RECT 121.855 130.485 122.145 130.530 ;
        RECT 128.280 130.470 128.600 130.530 ;
        RECT 138.860 130.670 139.180 130.730 ;
        RECT 142.080 130.670 142.400 130.730 ;
        RECT 138.860 130.530 142.400 130.670 ;
        RECT 138.860 130.470 139.180 130.530 ;
        RECT 142.080 130.470 142.400 130.530 ;
        RECT 145.300 130.670 145.620 130.730 ;
        RECT 145.300 130.530 149.670 130.670 ;
        RECT 145.300 130.470 145.620 130.530 ;
        RECT 120.475 130.330 120.765 130.375 ;
        RECT 123.695 130.330 123.985 130.375 ;
        RECT 130.120 130.330 130.440 130.390 ;
        RECT 117.330 130.190 120.765 130.330 ;
        RECT 112.640 129.850 114.710 129.990 ;
        RECT 112.640 129.790 112.960 129.850 ;
        RECT 95.175 129.510 98.240 129.650 ;
        RECT 95.175 129.465 95.465 129.510 ;
        RECT 97.920 129.450 98.240 129.510 ;
        RECT 99.315 129.465 99.605 129.695 ;
        RECT 99.775 129.465 100.065 129.695 ;
        RECT 100.695 129.465 100.985 129.695 ;
        RECT 102.075 129.465 102.365 129.695 ;
        RECT 99.850 129.310 99.990 129.465 ;
        RECT 89.830 129.170 99.990 129.310 ;
        RECT 102.150 129.310 102.290 129.465 ;
        RECT 102.980 129.450 103.300 129.710 ;
        RECT 106.200 129.650 106.520 129.710 ;
        RECT 107.120 129.650 107.440 129.710 ;
        RECT 106.200 129.510 107.440 129.650 ;
        RECT 106.200 129.450 106.520 129.510 ;
        RECT 107.120 129.450 107.440 129.510 ;
        RECT 108.040 129.450 108.360 129.710 ;
        RECT 109.895 129.650 110.185 129.695 ;
        RECT 111.275 129.650 111.565 129.695 ;
        RECT 109.895 129.510 111.565 129.650 ;
        RECT 109.895 129.465 110.185 129.510 ;
        RECT 111.275 129.465 111.565 129.510 ;
        RECT 112.180 129.450 112.500 129.710 ;
        RECT 113.100 129.450 113.420 129.710 ;
        RECT 114.570 129.695 114.710 129.850 ;
        RECT 115.875 129.805 116.165 130.035 ;
        RECT 117.330 129.710 117.470 130.190 ;
        RECT 120.475 130.145 120.765 130.190 ;
        RECT 121.470 130.190 130.440 130.330 ;
        RECT 114.495 129.465 114.785 129.695 ;
        RECT 115.415 129.465 115.705 129.695 ;
        RECT 103.900 129.310 104.220 129.370 ;
        RECT 102.150 129.170 104.220 129.310 ;
        RECT 108.130 129.310 108.270 129.450 ;
        RECT 115.490 129.310 115.630 129.465 ;
        RECT 116.320 129.450 116.640 129.710 ;
        RECT 116.780 129.450 117.100 129.710 ;
        RECT 117.240 129.450 117.560 129.710 ;
        RECT 121.470 129.695 121.610 130.190 ;
        RECT 123.695 130.145 123.985 130.190 ;
        RECT 130.120 130.130 130.440 130.190 ;
        RECT 130.595 130.330 130.885 130.375 ;
        RECT 133.340 130.330 133.660 130.390 ;
        RECT 138.415 130.330 138.705 130.375 ;
        RECT 130.595 130.190 133.660 130.330 ;
        RECT 130.595 130.145 130.885 130.190 ;
        RECT 133.340 130.130 133.660 130.190 ;
        RECT 135.730 130.190 138.705 130.330 ;
        RECT 123.220 129.790 123.540 130.050 ;
        RECT 127.820 129.790 128.140 130.050 ;
        RECT 129.215 129.990 129.505 130.035 ;
        RECT 130.210 129.990 130.350 130.130 ;
        RECT 129.215 129.850 130.350 129.990 ;
        RECT 131.040 129.990 131.360 130.050 ;
        RECT 134.720 129.990 135.040 130.050 ;
        RECT 131.040 129.850 133.110 129.990 ;
        RECT 129.215 129.805 129.505 129.850 ;
        RECT 131.040 129.790 131.360 129.850 ;
        RECT 117.715 129.650 118.005 129.695 ;
        RECT 120.015 129.650 120.305 129.695 ;
        RECT 121.395 129.650 121.685 129.695 ;
        RECT 117.715 129.510 119.770 129.650 ;
        RECT 117.715 129.465 118.005 129.510 ;
        RECT 118.160 129.310 118.480 129.370 ;
        RECT 119.630 129.310 119.770 129.510 ;
        RECT 120.015 129.510 121.685 129.650 ;
        RECT 120.015 129.465 120.305 129.510 ;
        RECT 121.395 129.465 121.685 129.510 ;
        RECT 122.775 129.650 123.065 129.695 ;
        RECT 123.310 129.650 123.450 129.790 ;
        RECT 124.615 129.650 124.905 129.695 ;
        RECT 122.775 129.510 124.905 129.650 ;
        RECT 122.775 129.465 123.065 129.510 ;
        RECT 124.615 129.465 124.905 129.510 ;
        RECT 129.660 129.450 129.980 129.710 ;
        RECT 130.120 129.650 130.440 129.710 ;
        RECT 132.970 129.695 133.110 129.850 ;
        RECT 133.430 129.850 135.040 129.990 ;
        RECT 133.430 129.695 133.570 129.850 ;
        RECT 134.720 129.790 135.040 129.850 ;
        RECT 132.435 129.650 132.725 129.695 ;
        RECT 130.120 129.510 132.725 129.650 ;
        RECT 130.120 129.450 130.440 129.510 ;
        RECT 132.435 129.465 132.725 129.510 ;
        RECT 132.895 129.465 133.185 129.695 ;
        RECT 133.355 129.465 133.645 129.695 ;
        RECT 134.275 129.650 134.565 129.695 ;
        RECT 135.730 129.650 135.870 130.190 ;
        RECT 138.415 130.145 138.705 130.190 ;
        RECT 141.175 130.330 141.465 130.375 ;
        RECT 141.175 130.190 148.750 130.330 ;
        RECT 141.175 130.145 141.465 130.190 ;
        RECT 136.100 129.790 136.420 130.050 ;
        RECT 136.575 129.805 136.865 130.035 ;
        RECT 134.275 129.510 135.870 129.650 ;
        RECT 134.275 129.465 134.565 129.510 ;
        RECT 122.300 129.310 122.620 129.370 ;
        RECT 108.130 129.170 115.630 129.310 ;
        RECT 115.950 129.170 119.310 129.310 ;
        RECT 119.630 129.170 122.620 129.310 ;
        RECT 103.900 129.110 104.220 129.170 ;
        RECT 84.580 128.830 88.950 128.970 ;
        RECT 89.195 128.970 89.485 129.015 ;
        RECT 90.575 128.970 90.865 129.015 ;
        RECT 89.195 128.830 90.865 128.970 ;
        RECT 84.580 128.770 84.900 128.830 ;
        RECT 89.195 128.785 89.485 128.830 ;
        RECT 90.575 128.785 90.865 128.830 ;
        RECT 92.400 128.770 92.720 129.030 ;
        RECT 104.375 128.970 104.665 129.015 ;
        RECT 110.340 128.970 110.660 129.030 ;
        RECT 104.375 128.830 110.660 128.970 ;
        RECT 104.375 128.785 104.665 128.830 ;
        RECT 110.340 128.770 110.660 128.830 ;
        RECT 110.800 128.770 111.120 129.030 ;
        RECT 111.260 128.970 111.580 129.030 ;
        RECT 115.950 128.970 116.090 129.170 ;
        RECT 118.160 129.110 118.480 129.170 ;
        RECT 111.260 128.830 116.090 128.970 ;
        RECT 111.260 128.770 111.580 128.830 ;
        RECT 118.620 128.770 118.940 129.030 ;
        RECT 119.170 129.015 119.310 129.170 ;
        RECT 122.300 129.110 122.620 129.170 ;
        RECT 128.740 129.310 129.060 129.370 ;
        RECT 133.800 129.310 134.120 129.370 ;
        RECT 136.650 129.310 136.790 129.805 ;
        RECT 137.480 129.790 137.800 130.050 ;
        RECT 143.460 129.790 143.780 130.050 ;
        RECT 146.220 129.790 146.540 130.050 ;
        RECT 137.020 129.450 137.340 129.710 ;
        RECT 139.795 129.465 140.085 129.695 ;
        RECT 140.255 129.650 140.545 129.695 ;
        RECT 140.700 129.650 141.020 129.710 ;
        RECT 140.255 129.510 141.020 129.650 ;
        RECT 140.255 129.465 140.545 129.510 ;
        RECT 128.740 129.170 131.730 129.310 ;
        RECT 128.740 129.110 129.060 129.170 ;
        RECT 119.095 128.785 119.385 129.015 ;
        RECT 121.380 128.970 121.700 129.030 ;
        RECT 122.760 128.970 123.080 129.030 ;
        RECT 121.380 128.830 123.080 128.970 ;
        RECT 121.380 128.770 121.700 128.830 ;
        RECT 122.760 128.770 123.080 128.830 ;
        RECT 131.040 128.770 131.360 129.030 ;
        RECT 131.590 128.970 131.730 129.170 ;
        RECT 133.800 129.170 136.790 129.310 ;
        RECT 139.870 129.310 140.010 129.465 ;
        RECT 140.700 129.450 141.020 129.510 ;
        RECT 141.175 129.650 141.465 129.695 ;
        RECT 142.540 129.650 142.860 129.710 ;
        RECT 141.175 129.510 142.860 129.650 ;
        RECT 141.175 129.465 141.465 129.510 ;
        RECT 142.540 129.450 142.860 129.510 ;
        RECT 143.000 129.450 143.320 129.710 ;
        RECT 144.395 129.650 144.685 129.695 ;
        RECT 144.840 129.650 145.160 129.710 ;
        RECT 144.395 129.510 145.160 129.650 ;
        RECT 146.310 129.650 146.450 129.790 ;
        RECT 148.610 129.695 148.750 130.190 ;
        RECT 149.530 129.695 149.670 130.530 ;
        RECT 150.360 130.470 150.680 130.730 ;
        RECT 152.675 130.670 152.965 130.715 ;
        RECT 153.595 130.670 153.885 130.715 ;
        RECT 152.675 130.530 153.885 130.670 ;
        RECT 152.675 130.485 152.965 130.530 ;
        RECT 153.595 130.485 153.885 130.530 ;
        RECT 147.155 129.650 147.445 129.695 ;
        RECT 146.310 129.510 147.445 129.650 ;
        RECT 144.395 129.465 144.685 129.510 ;
        RECT 144.840 129.450 145.160 129.510 ;
        RECT 147.155 129.465 147.445 129.510 ;
        RECT 148.535 129.465 148.825 129.695 ;
        RECT 149.455 129.465 149.745 129.695 ;
        RECT 150.450 129.650 150.590 130.470 ;
        RECT 150.820 130.130 151.140 130.390 ;
        RECT 150.910 129.990 151.050 130.130 ;
        RECT 150.910 129.850 154.270 129.990 ;
        RECT 150.835 129.650 151.125 129.695 ;
        RECT 150.450 129.510 151.125 129.650 ;
        RECT 150.835 129.465 151.125 129.510 ;
        RECT 151.295 129.465 151.585 129.695 ;
        RECT 139.870 129.170 146.910 129.310 ;
        RECT 133.800 129.110 134.120 129.170 ;
        RECT 139.335 128.970 139.625 129.015 ;
        RECT 131.590 128.830 139.625 128.970 ;
        RECT 139.335 128.785 139.625 128.830 ;
        RECT 142.095 128.970 142.385 129.015 ;
        RECT 145.760 128.970 146.080 129.030 ;
        RECT 142.095 128.830 146.080 128.970 ;
        RECT 142.095 128.785 142.385 128.830 ;
        RECT 145.760 128.770 146.080 128.830 ;
        RECT 146.220 128.770 146.540 129.030 ;
        RECT 146.770 128.970 146.910 129.170 ;
        RECT 147.600 129.110 147.920 129.370 ;
        RECT 148.060 129.110 148.380 129.370 ;
        RECT 148.610 129.310 148.750 129.465 ;
        RECT 151.370 129.310 151.510 129.465 ;
        RECT 153.120 129.450 153.440 129.710 ;
        RECT 153.595 129.465 153.885 129.695 ;
        RECT 154.130 129.650 154.270 129.850 ;
        RECT 154.500 129.695 154.820 129.710 ;
        RECT 154.485 129.650 154.820 129.695 ;
        RECT 154.130 129.510 154.820 129.650 ;
        RECT 154.485 129.465 154.820 129.510 ;
        RECT 148.610 129.170 151.510 129.310 ;
        RECT 149.915 128.970 150.205 129.015 ;
        RECT 146.770 128.830 150.205 128.970 ;
        RECT 149.915 128.785 150.205 128.830 ;
        RECT 150.360 128.970 150.680 129.030 ;
        RECT 153.670 128.970 153.810 129.465 ;
        RECT 154.500 129.450 154.820 129.465 ;
        RECT 150.360 128.830 153.810 128.970 ;
        RECT 150.360 128.770 150.680 128.830 ;
        RECT 70.710 128.150 156.270 128.630 ;
        RECT 74.000 127.750 74.320 128.010 ;
        RECT 76.760 127.750 77.080 128.010 ;
        RECT 78.140 127.750 78.460 128.010 ;
        RECT 79.995 127.950 80.285 127.995 ;
        RECT 81.360 127.950 81.680 128.010 ;
        RECT 79.995 127.810 81.680 127.950 ;
        RECT 79.995 127.765 80.285 127.810 ;
        RECT 81.360 127.750 81.680 127.810 ;
        RECT 82.755 127.950 83.045 127.995 ;
        RECT 84.580 127.950 84.900 128.010 ;
        RECT 82.755 127.810 84.900 127.950 ;
        RECT 82.755 127.765 83.045 127.810 ;
        RECT 84.580 127.750 84.900 127.810 ;
        RECT 85.500 127.950 85.820 128.010 ;
        RECT 86.435 127.950 86.725 127.995 ;
        RECT 85.500 127.810 86.725 127.950 ;
        RECT 85.500 127.750 85.820 127.810 ;
        RECT 86.435 127.765 86.725 127.810 ;
        RECT 91.940 127.750 92.260 128.010 ;
        RECT 97.000 127.750 97.320 128.010 ;
        RECT 102.520 127.750 102.840 128.010 ;
        RECT 102.980 127.750 103.300 128.010 ;
        RECT 106.200 127.750 106.520 128.010 ;
        RECT 107.120 127.750 107.440 128.010 ;
        RECT 108.500 127.950 108.820 128.010 ;
        RECT 107.670 127.810 108.820 127.950 ;
        RECT 74.090 127.270 74.230 127.750 ;
        RECT 74.475 127.270 74.765 127.315 ;
        RECT 74.090 127.130 74.765 127.270 ;
        RECT 74.475 127.085 74.765 127.130 ;
        RECT 76.315 127.270 76.605 127.315 ;
        RECT 76.850 127.270 76.990 127.750 ;
        RECT 77.680 127.410 78.000 127.670 ;
        RECT 78.230 127.610 78.370 127.750 ;
        RECT 79.075 127.610 79.365 127.655 ;
        RECT 80.915 127.610 81.205 127.655 ;
        RECT 81.915 127.610 82.205 127.655 ;
        RECT 78.230 127.470 79.365 127.610 ;
        RECT 79.075 127.425 79.365 127.470 ;
        RECT 80.070 127.470 81.205 127.610 ;
        RECT 76.315 127.130 76.990 127.270 ;
        RECT 77.770 127.270 77.910 127.410 ;
        RECT 78.155 127.270 78.445 127.315 ;
        RECT 77.770 127.130 78.445 127.270 ;
        RECT 76.315 127.085 76.605 127.130 ;
        RECT 78.155 127.085 78.445 127.130 ;
        RECT 80.070 126.590 80.210 127.470 ;
        RECT 80.915 127.425 81.205 127.470 ;
        RECT 81.450 127.470 82.205 127.610 ;
        RECT 80.440 127.270 80.760 127.330 ;
        RECT 81.450 127.270 81.590 127.470 ;
        RECT 81.915 127.425 82.205 127.470 ;
        RECT 86.880 127.610 87.200 127.670 ;
        RECT 92.030 127.610 92.170 127.750 ;
        RECT 86.880 127.470 92.170 127.610 ;
        RECT 86.880 127.410 87.200 127.470 ;
        RECT 80.440 127.130 81.590 127.270 ;
        RECT 82.740 127.270 83.060 127.330 ;
        RECT 84.135 127.270 84.425 127.315 ;
        RECT 82.740 127.130 84.425 127.270 ;
        RECT 80.440 127.070 80.760 127.130 ;
        RECT 82.740 127.070 83.060 127.130 ;
        RECT 84.135 127.085 84.425 127.130 ;
        RECT 84.595 127.270 84.885 127.315 ;
        RECT 86.420 127.270 86.740 127.330 ;
        RECT 84.595 127.130 86.740 127.270 ;
        RECT 84.595 127.085 84.885 127.130 ;
        RECT 86.420 127.070 86.740 127.130 ;
        RECT 87.800 127.070 88.120 127.330 ;
        RECT 88.260 127.070 88.580 127.330 ;
        RECT 88.735 127.260 89.025 127.315 ;
        RECT 89.180 127.260 89.500 127.330 ;
        RECT 89.830 127.315 89.970 127.470 ;
        RECT 92.400 127.410 92.720 127.670 ;
        RECT 97.090 127.610 97.230 127.750 ;
        RECT 97.090 127.470 100.450 127.610 ;
        RECT 88.735 127.120 89.500 127.260 ;
        RECT 88.735 127.085 89.025 127.120 ;
        RECT 89.180 127.070 89.500 127.120 ;
        RECT 89.655 127.120 89.970 127.315 ;
        RECT 89.655 127.085 89.945 127.120 ;
        RECT 91.940 127.070 92.260 127.330 ;
        RECT 92.490 127.270 92.630 127.410 ;
        RECT 92.490 127.130 95.390 127.270 ;
        RECT 85.040 126.730 85.360 126.990 ;
        RECT 85.515 126.930 85.805 126.975 ;
        RECT 85.960 126.930 86.280 126.990 ;
        RECT 85.515 126.790 86.280 126.930 ;
        RECT 87.890 126.930 88.030 127.070 ;
        RECT 91.495 126.930 91.785 126.975 ;
        RECT 87.890 126.790 91.785 126.930 ;
        RECT 85.515 126.745 85.805 126.790 ;
        RECT 85.960 126.730 86.280 126.790 ;
        RECT 91.495 126.745 91.785 126.790 ;
        RECT 93.795 126.745 94.085 126.975 ;
        RECT 95.250 126.930 95.390 127.130 ;
        RECT 95.620 127.070 95.940 127.330 ;
        RECT 97.460 127.270 97.780 127.330 ;
        RECT 97.935 127.270 98.225 127.315 ;
        RECT 97.460 127.130 98.225 127.270 ;
        RECT 97.460 127.070 97.780 127.130 ;
        RECT 97.935 127.085 98.225 127.130 ;
        RECT 99.315 127.270 99.605 127.315 ;
        RECT 99.760 127.270 100.080 127.330 ;
        RECT 100.310 127.315 100.450 127.470 ;
        RECT 102.610 127.315 102.750 127.750 ;
        RECT 106.290 127.610 106.430 127.750 ;
        RECT 103.990 127.470 106.430 127.610 ;
        RECT 99.315 127.130 100.080 127.270 ;
        RECT 99.315 127.085 99.605 127.130 ;
        RECT 99.760 127.070 100.080 127.130 ;
        RECT 100.235 127.085 100.525 127.315 ;
        RECT 102.535 127.085 102.825 127.315 ;
        RECT 102.995 127.270 103.285 127.315 ;
        RECT 103.440 127.270 103.760 127.330 ;
        RECT 103.990 127.315 104.130 127.470 ;
        RECT 102.995 127.130 103.760 127.270 ;
        RECT 102.995 127.085 103.285 127.130 ;
        RECT 98.395 126.930 98.685 126.975 ;
        RECT 95.250 126.790 98.685 126.930 ;
        RECT 98.395 126.745 98.685 126.790 ;
        RECT 98.855 126.930 99.145 126.975 ;
        RECT 101.140 126.930 101.460 126.990 ;
        RECT 98.855 126.790 101.460 126.930 ;
        RECT 102.610 126.930 102.750 127.085 ;
        RECT 103.440 127.070 103.760 127.130 ;
        RECT 103.915 127.085 104.205 127.315 ;
        RECT 105.295 127.270 105.585 127.315 ;
        RECT 105.740 127.270 106.060 127.330 ;
        RECT 105.295 127.130 106.060 127.270 ;
        RECT 105.295 127.085 105.585 127.130 ;
        RECT 105.740 127.070 106.060 127.130 ;
        RECT 106.215 127.270 106.505 127.315 ;
        RECT 107.210 127.270 107.350 127.750 ;
        RECT 107.670 127.315 107.810 127.810 ;
        RECT 108.500 127.750 108.820 127.810 ;
        RECT 116.780 127.750 117.100 128.010 ;
        RECT 118.160 127.950 118.480 128.010 ;
        RECT 130.120 127.950 130.440 128.010 ;
        RECT 118.160 127.810 119.080 127.950 ;
        RECT 118.160 127.750 118.480 127.810 ;
        RECT 108.040 127.610 108.360 127.670 ;
        RECT 110.340 127.610 110.660 127.670 ;
        RECT 112.640 127.610 112.960 127.670 ;
        RECT 116.870 127.610 117.010 127.750 ;
        RECT 118.940 127.610 119.080 127.810 ;
        RECT 120.550 127.810 130.440 127.950 ;
        RECT 108.040 127.470 108.730 127.610 ;
        RECT 108.040 127.410 108.360 127.470 ;
        RECT 108.590 127.315 108.730 127.470 ;
        RECT 110.340 127.470 112.960 127.610 ;
        RECT 110.340 127.410 110.660 127.470 ;
        RECT 112.640 127.410 112.960 127.470 ;
        RECT 113.190 127.470 117.470 127.610 ;
        RECT 118.940 127.470 119.770 127.610 ;
        RECT 113.190 127.315 113.330 127.470 ;
        RECT 106.215 127.130 107.350 127.270 ;
        RECT 106.215 127.085 106.505 127.130 ;
        RECT 107.595 127.085 107.885 127.315 ;
        RECT 108.515 127.085 108.805 127.315 ;
        RECT 109.050 127.130 112.870 127.270 ;
        RECT 104.375 126.930 104.665 126.975 ;
        RECT 102.610 126.790 104.665 126.930 ;
        RECT 98.855 126.745 99.145 126.790 ;
        RECT 84.120 126.590 84.440 126.650 ;
        RECT 80.070 126.450 84.440 126.590 ;
        RECT 85.130 126.590 85.270 126.730 ;
        RECT 87.355 126.590 87.645 126.635 ;
        RECT 85.130 126.450 87.645 126.590 ;
        RECT 93.870 126.590 94.010 126.745 ;
        RECT 101.140 126.730 101.460 126.790 ;
        RECT 104.375 126.745 104.665 126.790 ;
        RECT 106.660 126.730 106.980 126.990 ;
        RECT 107.135 126.745 107.425 126.975 ;
        RECT 93.870 126.450 99.990 126.590 ;
        RECT 84.120 126.390 84.440 126.450 ;
        RECT 87.355 126.405 87.645 126.450 ;
        RECT 99.850 126.310 99.990 126.450 ;
        RECT 73.540 126.050 73.860 126.310 ;
        RECT 75.395 126.250 75.685 126.295 ;
        RECT 76.760 126.250 77.080 126.310 ;
        RECT 75.395 126.110 77.080 126.250 ;
        RECT 75.395 126.065 75.685 126.110 ;
        RECT 76.760 126.050 77.080 126.110 ;
        RECT 81.820 126.050 82.140 126.310 ;
        RECT 85.960 126.250 86.280 126.310 ;
        RECT 89.195 126.250 89.485 126.295 ;
        RECT 85.960 126.110 89.485 126.250 ;
        RECT 85.960 126.050 86.280 126.110 ;
        RECT 89.195 126.065 89.485 126.110 ;
        RECT 94.700 126.050 95.020 126.310 ;
        RECT 97.000 126.050 97.320 126.310 ;
        RECT 99.760 126.050 100.080 126.310 ;
        RECT 101.140 126.050 101.460 126.310 ;
        RECT 101.600 126.050 101.920 126.310 ;
        RECT 102.060 126.250 102.380 126.310 ;
        RECT 107.210 126.250 107.350 126.745 ;
        RECT 109.050 126.250 109.190 127.130 ;
        RECT 109.435 126.930 109.725 126.975 ;
        RECT 110.340 126.930 110.660 126.990 ;
        RECT 109.435 126.790 110.660 126.930 ;
        RECT 112.730 126.930 112.870 127.130 ;
        RECT 113.115 127.085 113.405 127.315 ;
        RECT 114.020 127.070 114.340 127.330 ;
        RECT 116.335 127.085 116.625 127.315 ;
        RECT 114.480 126.930 114.800 126.990 ;
        RECT 112.730 126.790 114.800 126.930 ;
        RECT 116.410 126.930 116.550 127.085 ;
        RECT 116.780 127.070 117.100 127.330 ;
        RECT 117.330 127.315 117.470 127.470 ;
        RECT 117.255 127.085 117.545 127.315 ;
        RECT 118.160 127.070 118.480 127.330 ;
        RECT 119.630 127.315 119.770 127.470 ;
        RECT 119.555 127.085 119.845 127.315 ;
        RECT 120.550 127.270 120.690 127.810 ;
        RECT 130.120 127.750 130.440 127.810 ;
        RECT 130.580 127.950 130.900 128.010 ;
        RECT 131.055 127.950 131.345 127.995 ;
        RECT 130.580 127.810 131.345 127.950 ;
        RECT 130.580 127.750 130.900 127.810 ;
        RECT 131.055 127.765 131.345 127.810 ;
        RECT 135.180 127.950 135.500 128.010 ;
        RECT 143.015 127.950 143.305 127.995 ;
        RECT 144.380 127.950 144.700 128.010 ;
        RECT 135.180 127.810 140.930 127.950 ;
        RECT 135.180 127.750 135.500 127.810 ;
        RECT 121.380 127.610 121.700 127.670 ;
        RECT 125.060 127.610 125.380 127.670 ;
        RECT 121.380 127.470 123.910 127.610 ;
        RECT 121.380 127.410 121.700 127.470 ;
        RECT 120.090 127.130 120.690 127.270 ;
        RECT 120.935 127.270 121.225 127.315 ;
        RECT 120.935 127.130 123.450 127.270 ;
        RECT 120.090 126.930 120.230 127.130 ;
        RECT 120.935 127.085 121.225 127.130 ;
        RECT 123.310 126.990 123.450 127.130 ;
        RECT 116.410 126.790 120.230 126.930 ;
        RECT 109.435 126.745 109.725 126.790 ;
        RECT 110.340 126.730 110.660 126.790 ;
        RECT 114.480 126.730 114.800 126.790 ;
        RECT 120.460 126.730 120.780 126.990 ;
        RECT 122.760 126.730 123.080 126.990 ;
        RECT 123.220 126.730 123.540 126.990 ;
        RECT 123.770 126.930 123.910 127.470 ;
        RECT 124.230 127.470 125.380 127.610 ;
        RECT 124.230 127.315 124.370 127.470 ;
        RECT 125.060 127.410 125.380 127.470 ;
        RECT 127.375 127.610 127.665 127.655 ;
        RECT 127.375 127.470 130.850 127.610 ;
        RECT 127.375 127.425 127.665 127.470 ;
        RECT 124.155 127.085 124.445 127.315 ;
        RECT 129.675 127.270 129.965 127.315 ;
        RECT 124.690 127.130 129.965 127.270 ;
        RECT 124.690 126.930 124.830 127.130 ;
        RECT 129.675 127.085 129.965 127.130 ;
        RECT 123.770 126.790 124.830 126.930 ;
        RECT 128.280 126.730 128.600 126.990 ;
        RECT 128.740 126.730 129.060 126.990 ;
        RECT 112.180 126.390 112.500 126.650 ;
        RECT 112.640 126.590 112.960 126.650 ;
        RECT 118.160 126.590 118.480 126.650 ;
        RECT 118.635 126.590 118.925 126.635 ;
        RECT 112.640 126.450 117.930 126.590 ;
        RECT 112.640 126.390 112.960 126.450 ;
        RECT 102.060 126.110 109.190 126.250 ;
        RECT 109.880 126.250 110.200 126.310 ;
        RECT 114.955 126.250 115.245 126.295 ;
        RECT 109.880 126.110 115.245 126.250 ;
        RECT 117.790 126.250 117.930 126.450 ;
        RECT 118.160 126.450 118.925 126.590 ;
        RECT 118.160 126.390 118.480 126.450 ;
        RECT 118.635 126.405 118.925 126.450 ;
        RECT 120.015 126.590 120.305 126.635 ;
        RECT 128.830 126.590 128.970 126.730 ;
        RECT 120.015 126.450 128.970 126.590 ;
        RECT 130.710 126.590 130.850 127.470 ;
        RECT 133.800 127.410 134.120 127.670 ;
        RECT 134.260 127.610 134.580 127.670 ;
        RECT 134.260 127.470 135.870 127.610 ;
        RECT 134.260 127.410 134.580 127.470 ;
        RECT 131.500 127.070 131.820 127.330 ;
        RECT 131.975 127.270 132.265 127.315 ;
        RECT 132.420 127.270 132.740 127.330 ;
        RECT 131.975 127.130 132.740 127.270 ;
        RECT 131.975 127.085 132.265 127.130 ;
        RECT 132.420 127.070 132.740 127.130 ;
        RECT 132.880 127.070 133.200 127.330 ;
        RECT 134.720 127.070 135.040 127.330 ;
        RECT 135.730 127.315 135.870 127.470 ;
        RECT 135.655 127.085 135.945 127.315 ;
        RECT 137.480 127.070 137.800 127.330 ;
        RECT 138.400 127.070 138.720 127.330 ;
        RECT 139.780 127.070 140.100 127.330 ;
        RECT 140.790 127.315 140.930 127.810 ;
        RECT 143.015 127.810 144.700 127.950 ;
        RECT 143.015 127.765 143.305 127.810 ;
        RECT 144.380 127.750 144.700 127.810 ;
        RECT 145.300 127.950 145.620 128.010 ;
        RECT 146.695 127.950 146.985 127.995 ;
        RECT 145.300 127.810 146.985 127.950 ;
        RECT 145.300 127.750 145.620 127.810 ;
        RECT 146.695 127.765 146.985 127.810 ;
        RECT 148.060 127.950 148.380 128.010 ;
        RECT 148.060 127.810 152.430 127.950 ;
        RECT 148.060 127.750 148.380 127.810 ;
        RECT 152.290 127.655 152.430 127.810 ;
        RECT 148.995 127.610 149.285 127.655 ;
        RECT 143.090 127.470 149.285 127.610 ;
        RECT 140.715 127.085 141.005 127.315 ;
        RECT 141.620 127.270 141.940 127.330 ;
        RECT 142.095 127.270 142.385 127.315 ;
        RECT 141.620 127.130 142.385 127.270 ;
        RECT 141.620 127.070 141.940 127.130 ;
        RECT 142.095 127.085 142.385 127.130 ;
        RECT 131.590 126.930 131.730 127.070 ;
        RECT 133.355 126.930 133.645 126.975 ;
        RECT 136.115 126.930 136.405 126.975 ;
        RECT 138.875 126.930 139.165 126.975 ;
        RECT 131.590 126.790 139.165 126.930 ;
        RECT 133.355 126.745 133.645 126.790 ;
        RECT 136.115 126.745 136.405 126.790 ;
        RECT 138.875 126.745 139.165 126.790 ;
        RECT 139.335 126.745 139.625 126.975 ;
        RECT 143.090 126.930 143.230 127.470 ;
        RECT 148.995 127.425 149.285 127.470 ;
        RECT 152.215 127.610 152.505 127.655 ;
        RECT 154.040 127.610 154.360 127.670 ;
        RECT 152.215 127.470 154.360 127.610 ;
        RECT 152.215 127.425 152.505 127.470 ;
        RECT 154.040 127.410 154.360 127.470 ;
        RECT 154.960 127.410 155.280 127.670 ;
        RECT 143.460 127.270 143.780 127.330 ;
        RECT 144.855 127.270 145.145 127.315 ;
        RECT 143.460 127.130 145.145 127.270 ;
        RECT 143.460 127.070 143.780 127.130 ;
        RECT 144.855 127.085 145.145 127.130 ;
        RECT 146.680 127.070 147.000 127.330 ;
        RECT 147.600 127.270 147.920 127.330 ;
        RECT 153.120 127.270 153.440 127.330 ;
        RECT 155.050 127.270 155.190 127.410 ;
        RECT 147.600 127.130 155.190 127.270 ;
        RECT 147.600 127.070 147.920 127.130 ;
        RECT 153.120 127.070 153.440 127.130 ;
        RECT 141.250 126.790 143.230 126.930 ;
        RECT 144.395 126.930 144.685 126.975 ;
        RECT 146.770 126.930 146.910 127.070 ;
        RECT 151.295 126.930 151.585 126.975 ;
        RECT 144.395 126.790 145.070 126.930 ;
        RECT 146.770 126.790 151.585 126.930 ;
        RECT 136.575 126.590 136.865 126.635 ;
        RECT 130.710 126.450 136.865 126.590 ;
        RECT 120.015 126.405 120.305 126.450 ;
        RECT 136.575 126.405 136.865 126.450 ;
        RECT 138.400 126.590 138.720 126.650 ;
        RECT 139.410 126.590 139.550 126.745 ;
        RECT 138.400 126.450 139.550 126.590 ;
        RECT 138.400 126.390 138.720 126.450 ;
        RECT 123.235 126.250 123.525 126.295 ;
        RECT 117.790 126.110 123.525 126.250 ;
        RECT 102.060 126.050 102.380 126.110 ;
        RECT 109.880 126.050 110.200 126.110 ;
        RECT 114.955 126.065 115.245 126.110 ;
        RECT 123.235 126.065 123.525 126.110 ;
        RECT 125.075 126.250 125.365 126.295 ;
        RECT 125.520 126.250 125.840 126.310 ;
        RECT 125.075 126.110 125.840 126.250 ;
        RECT 125.075 126.065 125.365 126.110 ;
        RECT 125.520 126.050 125.840 126.110 ;
        RECT 125.980 126.050 126.300 126.310 ;
        RECT 127.360 126.250 127.680 126.310 ;
        RECT 128.755 126.250 129.045 126.295 ;
        RECT 127.360 126.110 129.045 126.250 ;
        RECT 127.360 126.050 127.680 126.110 ;
        RECT 128.755 126.065 129.045 126.110 ;
        RECT 130.595 126.250 130.885 126.295 ;
        RECT 141.250 126.250 141.390 126.790 ;
        RECT 144.395 126.745 144.685 126.790 ;
        RECT 144.930 126.650 145.070 126.790 ;
        RECT 151.295 126.745 151.585 126.790 ;
        RECT 141.635 126.590 141.925 126.635 ;
        RECT 143.920 126.590 144.240 126.650 ;
        RECT 141.635 126.450 144.240 126.590 ;
        RECT 141.635 126.405 141.925 126.450 ;
        RECT 143.920 126.390 144.240 126.450 ;
        RECT 144.840 126.390 145.160 126.650 ;
        RECT 145.850 126.450 149.670 126.590 ;
        RECT 130.595 126.110 141.390 126.250 ;
        RECT 142.540 126.250 142.860 126.310 ;
        RECT 145.850 126.250 145.990 126.450 ;
        RECT 149.530 126.295 149.670 126.450 ;
        RECT 142.540 126.110 145.990 126.250 ;
        RECT 130.595 126.065 130.885 126.110 ;
        RECT 142.540 126.050 142.860 126.110 ;
        RECT 149.455 126.065 149.745 126.295 ;
        RECT 70.710 125.430 156.270 125.910 ;
        RECT 80.440 125.030 80.760 125.290 ;
        RECT 97.000 125.030 97.320 125.290 ;
        RECT 112.180 125.030 112.500 125.290 ;
        RECT 114.480 125.030 114.800 125.290 ;
        RECT 117.255 125.230 117.545 125.275 ;
        RECT 117.700 125.230 118.020 125.290 ;
        RECT 117.255 125.090 118.020 125.230 ;
        RECT 117.255 125.045 117.545 125.090 ;
        RECT 117.700 125.030 118.020 125.090 ;
        RECT 120.475 125.045 120.765 125.275 ;
        RECT 123.235 125.230 123.525 125.275 ;
        RECT 123.680 125.230 124.000 125.290 ;
        RECT 123.235 125.090 124.000 125.230 ;
        RECT 123.235 125.045 123.525 125.090 ;
        RECT 78.140 124.890 78.460 124.950 ;
        RECT 81.375 124.890 81.665 124.935 ;
        RECT 78.140 124.750 81.665 124.890 ;
        RECT 78.140 124.690 78.460 124.750 ;
        RECT 81.375 124.705 81.665 124.750 ;
        RECT 79.980 124.550 80.300 124.610 ;
        RECT 97.090 124.550 97.230 125.030 ;
        RECT 108.500 124.550 108.820 124.610 ;
        RECT 112.270 124.550 112.410 125.030 ;
        RECT 79.980 124.410 80.670 124.550 ;
        RECT 79.980 124.350 80.300 124.410 ;
        RECT 73.540 124.010 73.860 124.270 ;
        RECT 75.855 124.210 76.145 124.255 ;
        RECT 76.760 124.210 77.080 124.270 ;
        RECT 75.855 124.070 77.080 124.210 ;
        RECT 75.855 124.025 76.145 124.070 ;
        RECT 76.760 124.010 77.080 124.070 ;
        RECT 77.220 124.210 77.540 124.270 ;
        RECT 79.075 124.210 79.365 124.255 ;
        RECT 77.220 124.070 79.365 124.210 ;
        RECT 77.220 124.010 77.540 124.070 ;
        RECT 79.075 124.025 79.365 124.070 ;
        RECT 79.520 124.010 79.840 124.270 ;
        RECT 80.530 124.255 80.670 124.410 ;
        RECT 82.370 124.410 97.230 124.550 ;
        RECT 98.010 124.410 108.820 124.550 ;
        RECT 82.370 124.255 82.510 124.410 ;
        RECT 80.455 124.025 80.745 124.255 ;
        RECT 82.295 124.025 82.585 124.255 ;
        RECT 85.515 124.025 85.805 124.255 ;
        RECT 87.355 124.210 87.645 124.255 ;
        RECT 88.720 124.210 89.040 124.270 ;
        RECT 87.355 124.070 89.040 124.210 ;
        RECT 87.355 124.025 87.645 124.070 ;
        RECT 79.610 123.870 79.750 124.010 ;
        RECT 79.995 123.870 80.285 123.915 ;
        RECT 79.610 123.730 80.285 123.870 ;
        RECT 85.590 123.870 85.730 124.025 ;
        RECT 88.720 124.010 89.040 124.070 ;
        RECT 91.035 124.210 91.325 124.255 ;
        RECT 94.240 124.210 94.560 124.270 ;
        RECT 91.035 124.070 94.560 124.210 ;
        RECT 91.035 124.025 91.325 124.070 ;
        RECT 94.240 124.010 94.560 124.070 ;
        RECT 94.700 124.010 95.020 124.270 ;
        RECT 98.010 123.870 98.150 124.410 ;
        RECT 108.500 124.350 108.820 124.410 ;
        RECT 109.050 124.410 112.410 124.550 ;
        RECT 98.380 124.010 98.700 124.270 ;
        RECT 101.140 124.010 101.460 124.270 ;
        RECT 101.600 124.210 101.920 124.270 ;
        RECT 109.050 124.255 109.190 124.410 ;
        RECT 102.075 124.210 102.365 124.255 ;
        RECT 101.600 124.070 102.365 124.210 ;
        RECT 101.600 124.010 101.920 124.070 ;
        RECT 102.075 124.025 102.365 124.070 ;
        RECT 104.375 124.025 104.665 124.255 ;
        RECT 108.975 124.025 109.265 124.255 ;
        RECT 85.590 123.730 98.150 123.870 ;
        RECT 101.230 123.870 101.370 124.010 ;
        RECT 104.450 123.870 104.590 124.025 ;
        RECT 110.340 124.010 110.660 124.270 ;
        RECT 101.230 123.730 104.590 123.870 ;
        RECT 108.500 123.870 108.820 123.930 ;
        RECT 114.570 123.870 114.710 125.030 ;
        RECT 114.940 124.890 115.260 124.950 ;
        RECT 120.550 124.890 120.690 125.045 ;
        RECT 123.680 125.030 124.000 125.090 ;
        RECT 124.140 125.230 124.460 125.290 ;
        RECT 125.995 125.230 126.285 125.275 ;
        RECT 124.140 125.090 126.285 125.230 ;
        RECT 124.140 125.030 124.460 125.090 ;
        RECT 125.995 125.045 126.285 125.090 ;
        RECT 131.515 125.230 131.805 125.275 ;
        RECT 131.960 125.230 132.280 125.290 ;
        RECT 133.800 125.230 134.120 125.290 ;
        RECT 138.860 125.230 139.180 125.290 ;
        RECT 131.515 125.090 132.280 125.230 ;
        RECT 131.515 125.045 131.805 125.090 ;
        RECT 131.960 125.030 132.280 125.090 ;
        RECT 132.510 125.090 134.120 125.230 ;
        RECT 132.510 124.890 132.650 125.090 ;
        RECT 133.800 125.030 134.120 125.090 ;
        RECT 137.570 125.090 139.180 125.230 ;
        RECT 114.940 124.750 120.690 124.890 ;
        RECT 129.980 124.750 132.650 124.890 ;
        RECT 133.355 124.890 133.645 124.935 ;
        RECT 137.570 124.890 137.710 125.090 ;
        RECT 138.860 125.030 139.180 125.090 ;
        RECT 139.320 125.230 139.640 125.290 ;
        RECT 139.795 125.230 140.085 125.275 ;
        RECT 139.320 125.090 140.085 125.230 ;
        RECT 139.320 125.030 139.640 125.090 ;
        RECT 139.795 125.045 140.085 125.090 ;
        RECT 141.160 125.230 141.480 125.290 ;
        RECT 142.555 125.230 142.845 125.275 ;
        RECT 141.160 125.090 142.845 125.230 ;
        RECT 141.160 125.030 141.480 125.090 ;
        RECT 142.555 125.045 142.845 125.090 ;
        RECT 143.000 125.230 143.320 125.290 ;
        RECT 144.395 125.230 144.685 125.275 ;
        RECT 143.000 125.090 144.685 125.230 ;
        RECT 143.000 125.030 143.320 125.090 ;
        RECT 144.395 125.045 144.685 125.090 ;
        RECT 149.455 125.045 149.745 125.275 ;
        RECT 133.355 124.750 137.710 124.890 ;
        RECT 137.940 124.890 138.260 124.950 ;
        RECT 149.530 124.890 149.670 125.045 ;
        RECT 153.120 125.030 153.440 125.290 ;
        RECT 137.940 124.750 149.670 124.890 ;
        RECT 114.940 124.690 115.260 124.750 ;
        RECT 129.980 124.550 130.120 124.750 ;
        RECT 133.355 124.705 133.645 124.750 ;
        RECT 137.940 124.690 138.260 124.750 ;
        RECT 115.950 124.410 130.120 124.550 ;
        RECT 131.500 124.550 131.820 124.610 ;
        RECT 133.815 124.550 134.105 124.595 ;
        RECT 131.500 124.410 134.105 124.550 ;
        RECT 115.950 124.255 116.090 124.410 ;
        RECT 131.500 124.350 131.820 124.410 ;
        RECT 133.815 124.365 134.105 124.410 ;
        RECT 134.720 124.550 135.040 124.610 ;
        RECT 146.695 124.550 146.985 124.595 ;
        RECT 134.720 124.410 146.985 124.550 ;
        RECT 134.720 124.350 135.040 124.410 ;
        RECT 146.695 124.365 146.985 124.410 ;
        RECT 151.295 124.550 151.585 124.595 ;
        RECT 153.580 124.550 153.900 124.610 ;
        RECT 151.295 124.410 153.900 124.550 ;
        RECT 151.295 124.365 151.585 124.410 ;
        RECT 153.580 124.350 153.900 124.410 ;
        RECT 115.875 124.025 116.165 124.255 ;
        RECT 116.795 124.210 117.085 124.255 ;
        RECT 117.240 124.210 117.560 124.270 ;
        RECT 116.795 124.070 117.560 124.210 ;
        RECT 116.795 124.025 117.085 124.070 ;
        RECT 116.870 123.870 117.010 124.025 ;
        RECT 117.240 124.010 117.560 124.070 ;
        RECT 118.175 124.210 118.465 124.255 ;
        RECT 118.175 124.070 122.070 124.210 ;
        RECT 118.175 124.025 118.465 124.070 ;
        RECT 108.500 123.730 111.030 123.870 ;
        RECT 114.570 123.730 117.010 123.870 ;
        RECT 119.095 123.870 119.385 123.915 ;
        RECT 120.015 123.870 120.305 123.915 ;
        RECT 119.095 123.730 120.305 123.870 ;
        RECT 121.930 123.870 122.070 124.070 ;
        RECT 122.760 124.010 123.080 124.270 ;
        RECT 124.155 124.210 124.445 124.255 ;
        RECT 123.310 124.070 124.445 124.210 ;
        RECT 123.310 123.930 123.450 124.070 ;
        RECT 124.155 124.025 124.445 124.070 ;
        RECT 126.900 124.010 127.220 124.270 ;
        RECT 127.835 124.025 128.125 124.255 ;
        RECT 123.220 123.870 123.540 123.930 ;
        RECT 121.930 123.730 123.540 123.870 ;
        RECT 79.995 123.685 80.285 123.730 ;
        RECT 108.500 123.670 108.820 123.730 ;
        RECT 70.780 123.530 71.100 123.590 ;
        RECT 72.635 123.530 72.925 123.575 ;
        RECT 70.780 123.390 72.925 123.530 ;
        RECT 70.780 123.330 71.100 123.390 ;
        RECT 72.635 123.345 72.925 123.390 ;
        RECT 74.460 123.330 74.780 123.590 ;
        RECT 81.820 123.530 82.140 123.590 ;
        RECT 84.595 123.530 84.885 123.575 ;
        RECT 81.820 123.390 84.885 123.530 ;
        RECT 81.820 123.330 82.140 123.390 ;
        RECT 84.595 123.345 84.885 123.390 ;
        RECT 86.420 123.330 86.740 123.590 ;
        RECT 89.180 123.530 89.500 123.590 ;
        RECT 90.115 123.530 90.405 123.575 ;
        RECT 89.180 123.390 90.405 123.530 ;
        RECT 89.180 123.330 89.500 123.390 ;
        RECT 90.115 123.345 90.405 123.390 ;
        RECT 93.780 123.330 94.100 123.590 ;
        RECT 97.460 123.330 97.780 123.590 ;
        RECT 101.140 123.330 101.460 123.590 ;
        RECT 103.900 123.530 104.220 123.590 ;
        RECT 105.295 123.530 105.585 123.575 ;
        RECT 103.900 123.390 105.585 123.530 ;
        RECT 103.900 123.330 104.220 123.390 ;
        RECT 105.295 123.345 105.585 123.390 ;
        RECT 108.055 123.530 108.345 123.575 ;
        RECT 109.880 123.530 110.200 123.590 ;
        RECT 110.890 123.575 111.030 123.730 ;
        RECT 119.095 123.685 119.385 123.730 ;
        RECT 120.015 123.685 120.305 123.730 ;
        RECT 123.220 123.670 123.540 123.730 ;
        RECT 123.680 123.870 124.000 123.930 ;
        RECT 127.910 123.870 128.050 124.025 ;
        RECT 130.120 124.010 130.440 124.270 ;
        RECT 132.435 124.210 132.725 124.255 ;
        RECT 134.260 124.210 134.580 124.270 ;
        RECT 136.115 124.210 136.405 124.255 ;
        RECT 132.435 124.070 133.570 124.210 ;
        RECT 132.435 124.025 132.725 124.070 ;
        RECT 129.660 123.870 129.980 123.930 ;
        RECT 133.430 123.870 133.570 124.070 ;
        RECT 134.260 124.070 136.405 124.210 ;
        RECT 134.260 124.010 134.580 124.070 ;
        RECT 136.115 124.025 136.405 124.070 ;
        RECT 137.480 124.010 137.800 124.270 ;
        RECT 138.400 124.210 138.720 124.270 ;
        RECT 139.335 124.210 139.625 124.255 ;
        RECT 138.400 124.070 139.625 124.210 ;
        RECT 138.400 124.010 138.720 124.070 ;
        RECT 139.335 124.025 139.625 124.070 ;
        RECT 139.780 124.210 140.100 124.270 ;
        RECT 140.715 124.210 141.005 124.255 ;
        RECT 142.095 124.210 142.385 124.255 ;
        RECT 139.780 124.070 141.005 124.210 ;
        RECT 137.570 123.870 137.710 124.010 ;
        RECT 123.680 123.730 125.750 123.870 ;
        RECT 127.910 123.730 129.430 123.870 ;
        RECT 123.680 123.670 124.000 123.730 ;
        RECT 108.055 123.390 110.200 123.530 ;
        RECT 108.055 123.345 108.345 123.390 ;
        RECT 109.880 123.330 110.200 123.390 ;
        RECT 110.815 123.345 111.105 123.575 ;
        RECT 115.415 123.530 115.705 123.575 ;
        RECT 118.620 123.530 118.940 123.590 ;
        RECT 115.415 123.390 118.940 123.530 ;
        RECT 115.415 123.345 115.705 123.390 ;
        RECT 118.620 123.330 118.940 123.390 ;
        RECT 125.060 123.330 125.380 123.590 ;
        RECT 125.610 123.530 125.750 123.730 ;
        RECT 128.755 123.530 129.045 123.575 ;
        RECT 125.610 123.390 129.045 123.530 ;
        RECT 129.290 123.530 129.430 123.730 ;
        RECT 129.660 123.730 133.110 123.870 ;
        RECT 133.430 123.730 137.710 123.870 ;
        RECT 139.410 123.870 139.550 124.025 ;
        RECT 139.780 124.010 140.100 124.070 ;
        RECT 140.715 124.025 141.005 124.070 ;
        RECT 141.250 124.070 142.385 124.210 ;
        RECT 141.250 123.870 141.390 124.070 ;
        RECT 142.095 124.025 142.385 124.070 ;
        RECT 143.460 124.010 143.780 124.270 ;
        RECT 143.920 124.210 144.240 124.270 ;
        RECT 143.920 124.070 145.530 124.210 ;
        RECT 143.920 124.010 144.240 124.070 ;
        RECT 145.390 123.915 145.530 124.070 ;
        RECT 152.200 124.010 152.520 124.270 ;
        RECT 139.410 123.730 141.390 123.870 ;
        RECT 129.660 123.670 129.980 123.730 ;
        RECT 132.420 123.530 132.740 123.590 ;
        RECT 129.290 123.390 132.740 123.530 ;
        RECT 132.970 123.530 133.110 123.730 ;
        RECT 141.635 123.685 141.925 123.915 ;
        RECT 145.315 123.685 145.605 123.915 ;
        RECT 136.575 123.530 136.865 123.575 ;
        RECT 132.970 123.390 136.865 123.530 ;
        RECT 141.710 123.530 141.850 123.685 ;
        RECT 148.980 123.670 149.300 123.930 ;
        RECT 148.520 123.530 148.840 123.590 ;
        RECT 141.710 123.390 148.840 123.530 ;
        RECT 128.755 123.345 129.045 123.390 ;
        RECT 132.420 123.330 132.740 123.390 ;
        RECT 136.575 123.345 136.865 123.390 ;
        RECT 148.520 123.330 148.840 123.390 ;
        RECT 70.710 122.710 156.270 123.190 ;
        RECT 94.240 122.310 94.560 122.570 ;
        RECT 98.380 122.510 98.700 122.570 ;
        RECT 131.960 122.510 132.280 122.570 ;
        RECT 98.380 122.370 132.280 122.510 ;
        RECT 98.380 122.310 98.700 122.370 ;
        RECT 131.960 122.310 132.280 122.370 ;
        RECT 132.420 122.510 132.740 122.570 ;
        RECT 139.780 122.510 140.100 122.570 ;
        RECT 132.420 122.370 140.100 122.510 ;
        RECT 132.420 122.310 132.740 122.370 ;
        RECT 139.780 122.310 140.100 122.370 ;
        RECT 141.620 122.310 141.940 122.570 ;
        RECT 148.980 122.310 149.300 122.570 ;
        RECT 94.330 121.830 94.470 122.310 ;
        RECT 99.760 122.170 100.080 122.230 ;
        RECT 116.320 122.170 116.640 122.230 ;
        RECT 99.760 122.030 116.640 122.170 ;
        RECT 99.760 121.970 100.080 122.030 ;
        RECT 116.320 121.970 116.640 122.030 ;
        RECT 125.060 122.170 125.380 122.230 ;
        RECT 141.710 122.170 141.850 122.310 ;
        RECT 125.060 122.030 141.850 122.170 ;
        RECT 125.060 121.970 125.380 122.030 ;
        RECT 130.580 121.830 130.900 121.890 ;
        RECT 94.330 121.690 130.900 121.830 ;
        RECT 130.580 121.630 130.900 121.690 ;
        RECT 107.120 121.490 107.440 121.550 ;
        RECT 127.820 121.490 128.140 121.550 ;
        RECT 138.400 121.490 138.720 121.550 ;
        RECT 107.120 121.350 138.720 121.490 ;
        RECT 107.120 121.290 107.440 121.350 ;
        RECT 127.820 121.290 128.140 121.350 ;
        RECT 138.400 121.290 138.720 121.350 ;
        RECT 88.720 121.150 89.040 121.210 ;
        RECT 118.160 121.150 118.480 121.210 ;
        RECT 88.720 121.010 118.480 121.150 ;
        RECT 88.720 120.950 89.040 121.010 ;
        RECT 118.160 120.950 118.480 121.010 ;
        RECT 125.520 121.150 125.840 121.210 ;
        RECT 149.070 121.150 149.210 122.310 ;
        RECT 125.520 121.010 149.210 121.150 ;
        RECT 125.520 120.950 125.840 121.010 ;
        RECT 51.580 101.330 52.580 105.830 ;
        RECT 55.580 101.330 56.580 105.830 ;
        RECT 59.580 101.330 60.580 105.830 ;
        RECT 63.580 101.330 64.580 105.830 ;
        RECT 67.580 101.330 68.580 105.830 ;
        RECT 71.580 101.330 72.580 105.830 ;
        RECT 75.580 101.330 76.580 105.830 ;
        RECT 51.810 100.865 52.400 101.330 ;
        RECT 55.810 100.865 56.400 101.330 ;
        RECT 59.810 100.865 60.400 101.330 ;
        RECT 63.810 100.865 64.400 101.330 ;
        RECT 67.810 100.865 68.400 101.330 ;
        RECT 71.810 100.865 72.400 101.330 ;
        RECT 75.810 100.865 76.400 101.330 ;
        RECT 77.580 80.110 78.580 105.830 ;
        RECT 79.580 101.330 80.580 105.830 ;
        RECT 79.810 100.865 80.400 101.330 ;
        RECT 77.580 80.080 78.600 80.110 ;
        RECT 50.900 79.080 81.410 80.080 ;
        RECT 77.600 79.050 78.600 79.080 ;
        RECT 51.810 60.650 52.400 61.075 ;
        RECT 55.810 60.650 56.400 61.075 ;
        RECT 59.810 60.650 60.400 61.075 ;
        RECT 63.810 60.650 64.400 61.075 ;
        RECT 67.810 60.650 68.400 61.075 ;
        RECT 71.810 60.650 72.400 61.075 ;
        RECT 75.810 60.650 76.400 61.075 ;
        RECT 79.810 60.650 80.400 61.075 ;
        RECT 51.580 57.530 52.580 60.650 ;
        RECT 50.000 56.530 52.580 57.530 ;
        RECT 51.580 53.430 52.580 56.530 ;
        RECT 55.580 54.430 56.580 60.650 ;
        RECT 59.580 54.430 60.580 60.650 ;
        RECT 63.580 54.430 64.580 60.650 ;
        RECT 67.580 54.430 68.580 60.650 ;
        RECT 71.580 54.430 72.580 60.650 ;
        RECT 75.580 54.430 76.580 60.650 ;
        RECT 79.580 54.430 80.580 60.650 ;
        RECT 53.630 53.430 56.610 54.430 ;
        RECT 57.630 53.430 60.610 54.430 ;
        RECT 61.630 53.430 64.610 54.430 ;
        RECT 65.630 53.430 68.610 54.430 ;
        RECT 69.630 53.430 72.610 54.430 ;
        RECT 73.630 53.430 76.610 54.430 ;
        RECT 77.630 53.430 80.610 54.430 ;
        RECT 51.810 52.865 52.400 53.430 ;
        RECT 51.810 32.940 52.400 33.425 ;
        RECT 53.630 32.940 54.630 53.430 ;
        RECT 55.810 52.865 56.400 53.430 ;
        RECT 55.810 32.940 56.400 33.425 ;
        RECT 57.630 32.940 58.630 53.430 ;
        RECT 59.810 52.865 60.400 53.430 ;
        RECT 59.810 32.940 60.400 33.425 ;
        RECT 61.630 32.940 62.630 53.430 ;
        RECT 63.810 52.865 64.400 53.430 ;
        RECT 63.810 32.940 64.400 33.425 ;
        RECT 65.630 32.940 66.630 53.430 ;
        RECT 67.810 52.865 68.400 53.430 ;
        RECT 67.810 32.940 68.400 33.425 ;
        RECT 69.630 32.940 70.630 53.430 ;
        RECT 71.810 52.865 72.400 53.430 ;
        RECT 71.810 32.940 72.400 33.425 ;
        RECT 73.630 32.940 74.630 53.430 ;
        RECT 75.810 52.865 76.400 53.430 ;
        RECT 75.810 32.940 76.400 33.425 ;
        RECT 77.630 32.940 78.630 53.430 ;
        RECT 79.810 52.865 80.400 53.430 ;
        RECT 51.490 31.940 54.630 32.940 ;
        RECT 55.490 31.940 58.630 32.940 ;
        RECT 59.490 31.940 62.630 32.940 ;
        RECT 63.490 31.940 66.630 32.940 ;
        RECT 67.490 31.940 70.630 32.940 ;
        RECT 71.490 31.940 74.630 32.940 ;
        RECT 75.490 31.940 78.630 32.940 ;
        RECT 79.810 32.930 80.400 33.425 ;
        RECT 81.930 32.930 82.930 105.830 ;
        RECT 88.580 101.330 89.580 105.830 ;
        RECT 92.580 101.330 93.580 105.830 ;
        RECT 96.580 101.330 97.580 105.830 ;
        RECT 100.580 101.330 101.580 105.830 ;
        RECT 104.580 101.330 105.580 105.830 ;
        RECT 108.580 101.330 109.580 105.830 ;
        RECT 112.580 101.330 113.580 105.830 ;
        RECT 88.810 100.865 89.400 101.330 ;
        RECT 92.810 100.865 93.400 101.330 ;
        RECT 96.810 100.865 97.400 101.330 ;
        RECT 100.810 100.865 101.400 101.330 ;
        RECT 104.810 100.865 105.400 101.330 ;
        RECT 108.810 100.865 109.400 101.330 ;
        RECT 112.810 100.865 113.400 101.330 ;
        RECT 114.580 80.110 115.580 105.830 ;
        RECT 116.580 101.330 117.580 105.830 ;
        RECT 116.810 100.865 117.400 101.330 ;
        RECT 114.580 80.080 115.600 80.110 ;
        RECT 87.900 79.080 118.410 80.080 ;
        RECT 114.600 79.050 115.600 79.080 ;
        RECT 88.810 60.650 89.400 61.075 ;
        RECT 92.810 60.650 93.400 61.075 ;
        RECT 96.810 60.650 97.400 61.075 ;
        RECT 100.810 60.650 101.400 61.075 ;
        RECT 104.810 60.650 105.400 61.075 ;
        RECT 108.810 60.650 109.400 61.075 ;
        RECT 112.810 60.650 113.400 61.075 ;
        RECT 116.810 60.650 117.400 61.075 ;
        RECT 88.580 57.530 89.580 60.650 ;
        RECT 87.000 56.530 89.580 57.530 ;
        RECT 88.580 53.430 89.580 56.530 ;
        RECT 92.580 54.430 93.580 60.650 ;
        RECT 96.580 54.430 97.580 60.650 ;
        RECT 100.580 54.430 101.580 60.650 ;
        RECT 104.580 54.430 105.580 60.650 ;
        RECT 108.580 54.430 109.580 60.650 ;
        RECT 112.580 54.430 113.580 60.650 ;
        RECT 116.580 54.430 117.580 60.650 ;
        RECT 90.630 53.430 93.610 54.430 ;
        RECT 94.630 53.430 97.610 54.430 ;
        RECT 98.630 53.430 101.610 54.430 ;
        RECT 102.630 53.430 105.610 54.430 ;
        RECT 106.630 53.430 109.610 54.430 ;
        RECT 110.630 53.430 113.610 54.430 ;
        RECT 114.630 53.430 117.610 54.430 ;
        RECT 88.810 52.865 89.400 53.430 ;
        RECT 88.810 32.940 89.400 33.425 ;
        RECT 90.630 32.940 91.630 53.430 ;
        RECT 92.810 52.865 93.400 53.430 ;
        RECT 92.810 32.940 93.400 33.425 ;
        RECT 94.630 32.940 95.630 53.430 ;
        RECT 96.810 52.865 97.400 53.430 ;
        RECT 96.810 32.940 97.400 33.425 ;
        RECT 98.630 32.940 99.630 53.430 ;
        RECT 100.810 52.865 101.400 53.430 ;
        RECT 100.810 32.940 101.400 33.425 ;
        RECT 102.630 32.940 103.630 53.430 ;
        RECT 104.810 52.865 105.400 53.430 ;
        RECT 104.810 32.940 105.400 33.425 ;
        RECT 106.630 32.940 107.630 53.430 ;
        RECT 108.810 52.865 109.400 53.430 ;
        RECT 108.810 32.940 109.400 33.425 ;
        RECT 110.630 32.940 111.630 53.430 ;
        RECT 112.810 52.865 113.400 53.430 ;
        RECT 112.810 32.940 113.400 33.425 ;
        RECT 114.630 32.940 115.630 53.430 ;
        RECT 116.810 52.865 117.400 53.430 ;
        RECT 51.810 31.320 52.400 31.940 ;
        RECT 55.810 31.320 56.400 31.940 ;
        RECT 59.810 31.320 60.400 31.940 ;
        RECT 63.810 31.320 64.400 31.940 ;
        RECT 67.810 31.320 68.400 31.940 ;
        RECT 71.810 31.320 72.400 31.940 ;
        RECT 75.810 31.320 76.400 31.940 ;
        RECT 79.520 31.930 82.930 32.930 ;
        RECT 88.490 31.940 91.630 32.940 ;
        RECT 92.490 31.940 95.630 32.940 ;
        RECT 96.490 31.940 99.630 32.940 ;
        RECT 100.490 31.940 103.630 32.940 ;
        RECT 104.490 31.940 107.630 32.940 ;
        RECT 108.490 31.940 111.630 32.940 ;
        RECT 112.490 31.940 115.630 32.940 ;
        RECT 116.810 32.930 117.400 33.425 ;
        RECT 118.930 32.930 119.930 105.830 ;
        RECT 125.580 101.330 126.580 105.830 ;
        RECT 129.580 101.330 130.580 105.830 ;
        RECT 133.580 101.330 134.580 105.830 ;
        RECT 137.580 101.330 138.580 105.830 ;
        RECT 141.580 101.330 142.580 105.830 ;
        RECT 145.580 101.330 146.580 105.830 ;
        RECT 149.580 101.330 150.580 105.830 ;
        RECT 125.810 100.865 126.400 101.330 ;
        RECT 129.810 100.865 130.400 101.330 ;
        RECT 133.810 100.865 134.400 101.330 ;
        RECT 137.810 100.865 138.400 101.330 ;
        RECT 141.810 100.865 142.400 101.330 ;
        RECT 145.810 100.865 146.400 101.330 ;
        RECT 149.810 100.865 150.400 101.330 ;
        RECT 151.580 80.110 152.580 105.830 ;
        RECT 153.580 101.330 154.580 105.830 ;
        RECT 153.810 100.865 154.400 101.330 ;
        RECT 151.580 80.080 152.600 80.110 ;
        RECT 124.900 79.080 155.410 80.080 ;
        RECT 151.600 79.050 152.600 79.080 ;
        RECT 125.810 60.650 126.400 61.075 ;
        RECT 129.810 60.650 130.400 61.075 ;
        RECT 133.810 60.650 134.400 61.075 ;
        RECT 137.810 60.650 138.400 61.075 ;
        RECT 141.810 60.650 142.400 61.075 ;
        RECT 145.810 60.650 146.400 61.075 ;
        RECT 149.810 60.650 150.400 61.075 ;
        RECT 153.810 60.650 154.400 61.075 ;
        RECT 125.580 57.530 126.580 60.650 ;
        RECT 124.000 56.530 126.580 57.530 ;
        RECT 125.580 53.430 126.580 56.530 ;
        RECT 129.580 54.430 130.580 60.650 ;
        RECT 133.580 54.430 134.580 60.650 ;
        RECT 137.580 54.430 138.580 60.650 ;
        RECT 141.580 54.430 142.580 60.650 ;
        RECT 145.580 54.430 146.580 60.650 ;
        RECT 149.580 54.430 150.580 60.650 ;
        RECT 153.580 54.430 154.580 60.650 ;
        RECT 127.630 53.430 130.610 54.430 ;
        RECT 131.630 53.430 134.610 54.430 ;
        RECT 135.630 53.430 138.610 54.430 ;
        RECT 139.630 53.430 142.610 54.430 ;
        RECT 143.630 53.430 146.610 54.430 ;
        RECT 147.630 53.430 150.610 54.430 ;
        RECT 151.630 53.430 154.610 54.430 ;
        RECT 125.810 52.865 126.400 53.430 ;
        RECT 125.810 32.940 126.400 33.425 ;
        RECT 127.630 32.940 128.630 53.430 ;
        RECT 129.810 52.865 130.400 53.430 ;
        RECT 129.810 32.940 130.400 33.425 ;
        RECT 131.630 32.940 132.630 53.430 ;
        RECT 133.810 52.865 134.400 53.430 ;
        RECT 133.810 32.940 134.400 33.425 ;
        RECT 135.630 32.940 136.630 53.430 ;
        RECT 137.810 52.865 138.400 53.430 ;
        RECT 137.810 32.940 138.400 33.425 ;
        RECT 139.630 32.940 140.630 53.430 ;
        RECT 141.810 52.865 142.400 53.430 ;
        RECT 141.810 32.940 142.400 33.425 ;
        RECT 143.630 32.940 144.630 53.430 ;
        RECT 145.810 52.865 146.400 53.430 ;
        RECT 145.810 32.940 146.400 33.425 ;
        RECT 147.630 32.940 148.630 53.430 ;
        RECT 149.810 52.865 150.400 53.430 ;
        RECT 149.810 32.940 150.400 33.425 ;
        RECT 151.630 32.940 152.630 53.430 ;
        RECT 153.810 52.865 154.400 53.430 ;
        RECT 79.810 31.320 80.400 31.930 ;
        RECT 88.810 31.320 89.400 31.940 ;
        RECT 92.810 31.320 93.400 31.940 ;
        RECT 96.810 31.320 97.400 31.940 ;
        RECT 100.810 31.320 101.400 31.940 ;
        RECT 104.810 31.320 105.400 31.940 ;
        RECT 108.810 31.320 109.400 31.940 ;
        RECT 112.810 31.320 113.400 31.940 ;
        RECT 116.520 31.930 119.930 32.930 ;
        RECT 125.490 31.940 128.630 32.940 ;
        RECT 129.490 31.940 132.630 32.940 ;
        RECT 133.490 31.940 136.630 32.940 ;
        RECT 137.490 31.940 140.630 32.940 ;
        RECT 141.490 31.940 144.630 32.940 ;
        RECT 145.490 31.940 148.630 32.940 ;
        RECT 149.490 31.940 152.630 32.940 ;
        RECT 153.810 32.930 154.400 33.425 ;
        RECT 155.930 32.930 156.930 105.830 ;
        RECT 116.810 31.320 117.400 31.930 ;
        RECT 125.810 31.320 126.400 31.940 ;
        RECT 129.810 31.320 130.400 31.940 ;
        RECT 133.810 31.320 134.400 31.940 ;
        RECT 137.810 31.320 138.400 31.940 ;
        RECT 141.810 31.320 142.400 31.940 ;
        RECT 145.810 31.320 146.400 31.940 ;
        RECT 149.810 31.320 150.400 31.940 ;
        RECT 153.520 31.930 156.930 32.930 ;
        RECT 153.810 31.320 154.400 31.930 ;
        RECT 50.980 30.030 80.920 31.030 ;
        RECT 87.980 30.030 117.920 31.030 ;
        RECT 124.980 30.030 154.920 31.030 ;
        RECT 32.020 26.310 35.120 26.345 ;
        RECT 32.015 26.080 35.120 26.310 ;
        RECT 32.020 26.045 35.120 26.080 ;
        RECT 31.825 22.595 32.055 25.875 ;
        RECT 32.265 22.845 32.495 25.875 ;
        RECT 34.820 24.345 35.120 26.045 ;
        RECT 36.020 24.345 36.320 24.375 ;
        RECT 34.720 24.045 36.320 24.345 ;
        RECT 36.020 24.015 36.320 24.045 ;
        RECT 34.640 22.845 34.870 23.895 ;
        RECT 35.080 23.745 35.310 23.895 ;
        RECT 36.470 23.745 37.470 28.095 ;
        RECT 29.320 21.595 32.070 22.595 ;
        RECT 32.265 21.595 34.870 22.845 ;
        RECT 35.070 22.745 37.470 23.745 ;
        RECT 31.825 17.875 32.055 21.595 ;
        RECT 32.265 17.875 32.495 21.595 ;
        RECT 33.470 18.345 33.770 21.595 ;
        RECT 34.640 19.895 34.870 21.595 ;
        RECT 35.080 19.895 35.310 22.745 ;
        RECT 36.020 21.995 36.320 22.025 ;
        RECT 36.470 21.995 37.470 22.345 ;
        RECT 36.020 21.695 37.470 21.995 ;
        RECT 36.020 21.665 36.320 21.695 ;
        RECT 36.470 21.345 37.470 21.695 ;
        RECT 36.020 19.745 36.320 19.775 ;
        RECT 34.720 19.445 36.320 19.745 ;
        RECT 34.320 18.345 34.620 18.375 ;
        RECT 33.470 18.045 34.620 18.345 ;
        RECT 34.320 18.015 34.620 18.045 ;
        RECT 34.820 17.695 35.120 19.445 ;
        RECT 36.020 19.415 36.320 19.445 ;
        RECT 36.470 18.345 37.470 18.695 ;
        RECT 35.340 18.045 37.470 18.345 ;
        RECT 36.470 17.695 37.470 18.045 ;
        RECT 31.970 17.395 35.120 17.695 ;
      LAYER via ;
        RECT 131.990 208.330 132.250 208.590 ;
        RECT 138.430 208.330 138.690 208.590 ;
        RECT 104.390 207.990 104.650 208.250 ;
        RECT 126.930 207.990 127.190 208.250 ;
        RECT 142.110 207.990 142.370 208.250 ;
        RECT 82.770 207.650 83.030 207.910 ;
        RECT 103.930 207.650 104.190 207.910 ;
        RECT 125.090 207.650 125.350 207.910 ;
        RECT 132.910 207.650 133.170 207.910 ;
        RECT 136.130 207.650 136.390 207.910 ;
        RECT 140.730 207.650 140.990 207.910 ;
        RECT 74.780 207.140 75.040 207.400 ;
        RECT 75.100 207.140 75.360 207.400 ;
        RECT 75.420 207.140 75.680 207.400 ;
        RECT 75.740 207.140 76.000 207.400 ;
        RECT 76.060 207.140 76.320 207.400 ;
        RECT 76.380 207.140 76.640 207.400 ;
        RECT 104.780 207.140 105.040 207.400 ;
        RECT 105.100 207.140 105.360 207.400 ;
        RECT 105.420 207.140 105.680 207.400 ;
        RECT 105.740 207.140 106.000 207.400 ;
        RECT 106.060 207.140 106.320 207.400 ;
        RECT 106.380 207.140 106.640 207.400 ;
        RECT 134.780 207.140 135.040 207.400 ;
        RECT 135.100 207.140 135.360 207.400 ;
        RECT 135.420 207.140 135.680 207.400 ;
        RECT 135.740 207.140 136.000 207.400 ;
        RECT 136.060 207.140 136.320 207.400 ;
        RECT 136.380 207.140 136.640 207.400 ;
        RECT 74.030 206.630 74.290 206.890 ;
        RECT 78.170 206.630 78.430 206.890 ;
        RECT 82.310 206.630 82.570 206.890 ;
        RECT 86.450 206.630 86.710 206.890 ;
        RECT 90.590 206.630 90.850 206.890 ;
        RECT 94.730 206.630 94.990 206.890 ;
        RECT 98.870 206.630 99.130 206.890 ;
        RECT 101.630 206.290 101.890 206.550 ;
        RECT 103.010 206.630 103.270 206.890 ;
        RECT 107.150 206.630 107.410 206.890 ;
        RECT 111.290 206.630 111.550 206.890 ;
        RECT 123.710 206.630 123.970 206.890 ;
        RECT 81.850 205.610 82.110 205.870 ;
        RECT 82.770 205.950 83.030 206.210 ;
        RECT 83.230 205.950 83.490 206.210 ;
        RECT 76.330 204.930 76.590 205.190 ;
        RECT 104.390 205.950 104.650 206.210 ;
        RECT 132.910 206.290 133.170 206.550 ;
        RECT 89.210 205.610 89.470 205.870 ;
        RECT 92.430 205.610 92.690 205.870 ;
        RECT 102.090 205.610 102.350 205.870 ;
        RECT 103.470 205.610 103.730 205.870 ;
        RECT 100.250 205.270 100.510 205.530 ;
        RECT 100.710 205.270 100.970 205.530 ;
        RECT 126.010 205.950 126.270 206.210 ;
        RECT 86.910 204.930 87.170 205.190 ;
        RECT 89.210 204.930 89.470 205.190 ;
        RECT 95.190 204.930 95.450 205.190 ;
        RECT 99.790 204.930 100.050 205.190 ;
        RECT 107.610 205.610 107.870 205.870 ;
        RECT 113.130 205.610 113.390 205.870 ;
        RECT 115.430 205.610 115.690 205.870 ;
        RECT 119.570 205.610 119.830 205.870 ;
        RECT 121.870 205.610 122.130 205.870 ;
        RECT 125.090 205.610 125.350 205.870 ;
        RECT 127.850 205.610 128.110 205.870 ;
        RECT 110.830 204.930 111.090 205.190 ;
        RECT 114.510 204.930 114.770 205.190 ;
        RECT 114.970 204.930 115.230 205.190 ;
        RECT 118.190 204.930 118.450 205.190 ;
        RECT 118.650 204.930 118.910 205.190 ;
        RECT 123.250 204.930 123.510 205.190 ;
        RECT 131.530 205.270 131.790 205.530 ;
        RECT 135.210 205.610 135.470 205.870 ;
        RECT 144.410 206.630 144.670 206.890 ;
        RECT 149.010 206.630 149.270 206.890 ;
        RECT 137.050 206.290 137.310 206.550 ;
        RECT 148.550 205.950 148.810 206.210 ;
        RECT 138.430 205.610 138.690 205.870 ;
        RECT 139.810 205.610 140.070 205.870 ;
        RECT 144.870 205.610 145.130 205.870 ;
        RECT 128.310 204.930 128.570 205.190 ;
        RECT 143.490 205.270 143.750 205.530 ;
        RECT 147.170 204.930 147.430 205.190 ;
        RECT 89.780 204.420 90.040 204.680 ;
        RECT 90.100 204.420 90.360 204.680 ;
        RECT 90.420 204.420 90.680 204.680 ;
        RECT 90.740 204.420 91.000 204.680 ;
        RECT 91.060 204.420 91.320 204.680 ;
        RECT 91.380 204.420 91.640 204.680 ;
        RECT 119.780 204.420 120.040 204.680 ;
        RECT 120.100 204.420 120.360 204.680 ;
        RECT 120.420 204.420 120.680 204.680 ;
        RECT 120.740 204.420 121.000 204.680 ;
        RECT 121.060 204.420 121.320 204.680 ;
        RECT 121.380 204.420 121.640 204.680 ;
        RECT 149.780 204.420 150.040 204.680 ;
        RECT 150.100 204.420 150.360 204.680 ;
        RECT 150.420 204.420 150.680 204.680 ;
        RECT 150.740 204.420 151.000 204.680 ;
        RECT 151.060 204.420 151.320 204.680 ;
        RECT 151.380 204.420 151.640 204.680 ;
        RECT 76.330 203.910 76.590 204.170 ;
        RECT 86.910 203.910 87.170 204.170 ;
        RECT 95.650 203.910 95.910 204.170 ;
        RECT 99.790 203.910 100.050 204.170 ;
        RECT 100.710 203.910 100.970 204.170 ;
        RECT 114.510 203.910 114.770 204.170 ;
        RECT 118.650 203.910 118.910 204.170 ;
        RECT 131.990 203.910 132.250 204.170 ;
        RECT 136.590 203.910 136.850 204.170 ;
        RECT 140.270 203.910 140.530 204.170 ;
        RECT 81.850 203.230 82.110 203.490 ;
        RECT 82.770 203.230 83.030 203.490 ;
        RECT 83.230 203.230 83.490 203.490 ;
        RECT 84.150 203.230 84.410 203.490 ;
        RECT 72.190 202.890 72.450 203.150 ;
        RECT 89.210 202.890 89.470 203.150 ;
        RECT 97.490 203.230 97.750 203.490 ;
        RECT 97.950 203.230 98.210 203.490 ;
        RECT 99.330 203.230 99.590 203.490 ;
        RECT 114.050 203.570 114.310 203.830 ;
        RECT 98.870 202.890 99.130 203.150 ;
        RECT 81.850 202.210 82.110 202.470 ;
        RECT 99.790 202.550 100.050 202.810 ;
        RECT 89.210 202.210 89.470 202.470 ;
        RECT 91.050 202.210 91.310 202.470 ;
        RECT 94.730 202.210 94.990 202.470 ;
        RECT 103.010 202.890 103.270 203.150 ;
        RECT 104.850 202.550 105.110 202.810 ;
        RECT 103.010 202.210 103.270 202.470 ;
        RECT 115.890 203.230 116.150 203.490 ;
        RECT 118.190 203.230 118.450 203.490 ;
        RECT 123.250 203.230 123.510 203.490 ;
        RECT 133.830 203.230 134.090 203.490 ;
        RECT 134.750 203.230 135.010 203.490 ;
        RECT 139.810 203.570 140.070 203.830 ;
        RECT 110.830 202.210 111.090 202.470 ;
        RECT 114.050 202.210 114.310 202.470 ;
        RECT 116.350 202.210 116.610 202.470 ;
        RECT 125.550 202.550 125.810 202.810 ;
        RECT 135.210 202.890 135.470 203.150 ;
        RECT 140.730 203.230 140.990 203.490 ;
        RECT 149.010 203.910 149.270 204.170 ;
        RECT 148.090 203.230 148.350 203.490 ;
        RECT 142.110 202.890 142.370 203.150 ;
        RECT 147.170 202.890 147.430 203.150 ;
        RECT 130.610 202.210 130.870 202.470 ;
        RECT 133.370 202.210 133.630 202.470 ;
        RECT 138.890 202.210 139.150 202.470 ;
        RECT 143.030 202.550 143.290 202.810 ;
        RECT 144.410 202.210 144.670 202.470 ;
        RECT 145.790 202.210 146.050 202.470 ;
        RECT 148.550 202.210 148.810 202.470 ;
        RECT 74.780 201.700 75.040 201.960 ;
        RECT 75.100 201.700 75.360 201.960 ;
        RECT 75.420 201.700 75.680 201.960 ;
        RECT 75.740 201.700 76.000 201.960 ;
        RECT 76.060 201.700 76.320 201.960 ;
        RECT 76.380 201.700 76.640 201.960 ;
        RECT 104.780 201.700 105.040 201.960 ;
        RECT 105.100 201.700 105.360 201.960 ;
        RECT 105.420 201.700 105.680 201.960 ;
        RECT 105.740 201.700 106.000 201.960 ;
        RECT 106.060 201.700 106.320 201.960 ;
        RECT 106.380 201.700 106.640 201.960 ;
        RECT 134.780 201.700 135.040 201.960 ;
        RECT 135.100 201.700 135.360 201.960 ;
        RECT 135.420 201.700 135.680 201.960 ;
        RECT 135.740 201.700 136.000 201.960 ;
        RECT 136.060 201.700 136.320 201.960 ;
        RECT 136.380 201.700 136.640 201.960 ;
        RECT 101.630 201.190 101.890 201.450 ;
        RECT 102.090 201.190 102.350 201.450 ;
        RECT 103.930 201.190 104.190 201.450 ;
        RECT 104.390 201.190 104.650 201.450 ;
        RECT 84.150 200.850 84.410 201.110 ;
        RECT 72.190 200.170 72.450 200.430 ;
        RECT 81.850 200.510 82.110 200.770 ;
        RECT 83.230 200.170 83.490 200.430 ;
        RECT 100.250 200.510 100.510 200.770 ;
        RECT 115.890 201.190 116.150 201.450 ;
        RECT 121.870 201.190 122.130 201.450 ;
        RECT 125.550 201.190 125.810 201.450 ;
        RECT 123.710 200.850 123.970 201.110 ;
        RECT 129.690 201.190 129.950 201.450 ;
        RECT 134.290 201.190 134.550 201.450 ;
        RECT 131.070 200.850 131.330 201.110 ;
        RECT 133.370 200.850 133.630 201.110 ;
        RECT 94.730 200.170 94.990 200.430 ;
        RECT 75.410 199.830 75.670 200.090 ;
        RECT 80.930 199.490 81.190 199.750 ;
        RECT 84.150 199.490 84.410 199.750 ;
        RECT 91.050 199.830 91.310 200.090 ;
        RECT 95.650 199.830 95.910 200.090 ;
        RECT 96.110 199.830 96.370 200.090 ;
        RECT 107.150 200.170 107.410 200.430 ;
        RECT 107.610 200.170 107.870 200.430 ;
        RECT 125.090 200.510 125.350 200.770 ;
        RECT 126.010 200.510 126.270 200.770 ;
        RECT 129.230 200.510 129.490 200.770 ;
        RECT 108.990 200.170 109.250 200.430 ;
        RECT 112.210 199.830 112.470 200.090 ;
        RECT 114.970 200.170 115.230 200.430 ;
        RECT 122.790 200.170 123.050 200.430 ;
        RECT 131.530 200.170 131.790 200.430 ;
        RECT 114.510 199.830 114.770 200.090 ;
        RECT 116.350 199.830 116.610 200.090 ;
        RECT 126.470 199.830 126.730 200.090 ;
        RECT 131.990 199.830 132.250 200.090 ;
        RECT 137.050 200.510 137.310 200.770 ;
        RECT 140.270 200.850 140.530 201.110 ;
        RECT 143.030 200.510 143.290 200.770 ;
        RECT 134.290 200.170 134.550 200.430 ;
        RECT 144.410 200.170 144.670 200.430 ;
        RECT 145.790 200.170 146.050 200.430 ;
        RECT 142.110 199.830 142.370 200.090 ;
        RECT 143.950 199.830 144.210 200.090 ;
        RECT 146.710 199.830 146.970 200.090 ;
        RECT 96.570 199.490 96.830 199.750 ;
        RECT 98.870 199.490 99.130 199.750 ;
        RECT 105.310 199.490 105.570 199.750 ;
        RECT 110.370 199.490 110.630 199.750 ;
        RECT 112.670 199.490 112.930 199.750 ;
        RECT 121.870 199.490 122.130 199.750 ;
        RECT 128.770 199.490 129.030 199.750 ;
        RECT 132.450 199.490 132.710 199.750 ;
        RECT 133.370 199.490 133.630 199.750 ;
        RECT 137.510 199.490 137.770 199.750 ;
        RECT 139.350 199.490 139.610 199.750 ;
        RECT 145.330 199.490 145.590 199.750 ;
        RECT 145.790 199.490 146.050 199.750 ;
        RECT 153.150 199.490 153.410 199.750 ;
        RECT 89.780 198.980 90.040 199.240 ;
        RECT 90.100 198.980 90.360 199.240 ;
        RECT 90.420 198.980 90.680 199.240 ;
        RECT 90.740 198.980 91.000 199.240 ;
        RECT 91.060 198.980 91.320 199.240 ;
        RECT 91.380 198.980 91.640 199.240 ;
        RECT 119.780 198.980 120.040 199.240 ;
        RECT 120.100 198.980 120.360 199.240 ;
        RECT 120.420 198.980 120.680 199.240 ;
        RECT 120.740 198.980 121.000 199.240 ;
        RECT 121.060 198.980 121.320 199.240 ;
        RECT 121.380 198.980 121.640 199.240 ;
        RECT 149.780 198.980 150.040 199.240 ;
        RECT 150.100 198.980 150.360 199.240 ;
        RECT 150.420 198.980 150.680 199.240 ;
        RECT 150.740 198.980 151.000 199.240 ;
        RECT 151.060 198.980 151.320 199.240 ;
        RECT 151.380 198.980 151.640 199.240 ;
        RECT 75.410 198.470 75.670 198.730 ;
        RECT 78.170 198.470 78.430 198.730 ;
        RECT 80.930 198.470 81.190 198.730 ;
        RECT 78.170 197.790 78.430 198.050 ;
        RECT 81.850 198.130 82.110 198.390 ;
        RECT 83.230 198.130 83.490 198.390 ;
        RECT 81.390 197.110 81.650 197.370 ;
        RECT 84.150 198.470 84.410 198.730 ;
        RECT 87.830 198.470 88.090 198.730 ;
        RECT 92.430 198.470 92.690 198.730 ;
        RECT 91.050 198.130 91.310 198.390 ;
        RECT 92.890 198.130 93.150 198.390 ;
        RECT 88.290 197.790 88.550 198.050 ;
        RECT 88.750 197.790 89.010 198.050 ;
        RECT 89.210 197.790 89.470 198.050 ;
        RECT 94.270 198.130 94.530 198.390 ;
        RECT 97.030 198.470 97.290 198.730 ;
        RECT 99.330 198.470 99.590 198.730 ;
        RECT 99.790 198.470 100.050 198.730 ;
        RECT 87.370 197.450 87.630 197.710 ;
        RECT 94.730 197.790 94.990 198.050 ;
        RECT 96.570 197.790 96.830 198.050 ;
        RECT 100.250 198.130 100.510 198.390 ;
        RECT 86.910 197.110 87.170 197.370 ;
        RECT 99.330 197.790 99.590 198.050 ;
        RECT 105.310 198.130 105.570 198.390 ;
        RECT 107.610 198.470 107.870 198.730 ;
        RECT 114.510 198.470 114.770 198.730 ;
        RECT 122.790 198.470 123.050 198.730 ;
        RECT 101.170 197.450 101.430 197.710 ;
        RECT 103.930 197.450 104.190 197.710 ;
        RECT 104.390 197.450 104.650 197.710 ;
        RECT 111.750 197.790 112.010 198.050 ;
        RECT 113.590 197.450 113.850 197.710 ;
        RECT 118.190 197.790 118.450 198.050 ;
        RECT 119.110 197.790 119.370 198.050 ;
        RECT 133.370 198.470 133.630 198.730 ;
        RECT 133.830 198.470 134.090 198.730 ;
        RECT 143.030 198.470 143.290 198.730 ;
        RECT 145.790 198.470 146.050 198.730 ;
        RECT 146.710 198.470 146.970 198.730 ;
        RECT 148.550 198.470 148.810 198.730 ;
        RECT 153.150 198.470 153.410 198.730 ;
        RECT 127.850 198.130 128.110 198.390 ;
        RECT 128.770 198.130 129.030 198.390 ;
        RECT 125.550 197.790 125.810 198.050 ;
        RECT 129.690 197.790 129.950 198.050 ;
        RECT 124.630 197.450 124.890 197.710 ;
        RECT 131.530 197.790 131.790 198.050 ;
        RECT 117.730 197.110 117.990 197.370 ;
        RECT 123.710 197.110 123.970 197.370 ;
        RECT 126.010 197.110 126.270 197.370 ;
        RECT 133.370 197.790 133.630 198.050 ;
        RECT 137.510 197.790 137.770 198.050 ;
        RECT 139.350 197.790 139.610 198.050 ;
        RECT 143.950 197.790 144.210 198.050 ;
        RECT 132.910 197.450 133.170 197.710 ;
        RECT 140.730 197.450 140.990 197.710 ;
        RECT 148.090 197.450 148.350 197.710 ;
        RECT 131.990 197.110 132.250 197.370 ;
        RECT 134.290 197.110 134.550 197.370 ;
        RECT 135.210 197.110 135.470 197.370 ;
        RECT 137.510 197.110 137.770 197.370 ;
        RECT 138.890 197.110 139.150 197.370 ;
        RECT 145.330 197.110 145.590 197.370 ;
        RECT 82.310 196.770 82.570 197.030 ;
        RECT 85.530 196.770 85.790 197.030 ;
        RECT 88.750 196.770 89.010 197.030 ;
        RECT 89.210 196.770 89.470 197.030 ;
        RECT 91.970 196.770 92.230 197.030 ;
        RECT 92.890 196.770 93.150 197.030 ;
        RECT 93.810 196.770 94.070 197.030 ;
        RECT 96.110 196.770 96.370 197.030 ;
        RECT 107.610 196.770 107.870 197.030 ;
        RECT 110.830 196.770 111.090 197.030 ;
        RECT 112.210 196.770 112.470 197.030 ;
        RECT 118.650 196.770 118.910 197.030 ;
        RECT 131.530 196.770 131.790 197.030 ;
        RECT 132.910 196.770 133.170 197.030 ;
        RECT 139.350 196.770 139.610 197.030 ;
        RECT 143.490 196.770 143.750 197.030 ;
        RECT 147.630 196.770 147.890 197.030 ;
        RECT 152.230 196.770 152.490 197.030 ;
        RECT 74.780 196.260 75.040 196.520 ;
        RECT 75.100 196.260 75.360 196.520 ;
        RECT 75.420 196.260 75.680 196.520 ;
        RECT 75.740 196.260 76.000 196.520 ;
        RECT 76.060 196.260 76.320 196.520 ;
        RECT 76.380 196.260 76.640 196.520 ;
        RECT 104.780 196.260 105.040 196.520 ;
        RECT 105.100 196.260 105.360 196.520 ;
        RECT 105.420 196.260 105.680 196.520 ;
        RECT 105.740 196.260 106.000 196.520 ;
        RECT 106.060 196.260 106.320 196.520 ;
        RECT 106.380 196.260 106.640 196.520 ;
        RECT 134.780 196.260 135.040 196.520 ;
        RECT 135.100 196.260 135.360 196.520 ;
        RECT 135.420 196.260 135.680 196.520 ;
        RECT 135.740 196.260 136.000 196.520 ;
        RECT 136.060 196.260 136.320 196.520 ;
        RECT 136.380 196.260 136.640 196.520 ;
        RECT 81.390 195.750 81.650 196.010 ;
        RECT 82.770 195.750 83.030 196.010 ;
        RECT 85.530 195.750 85.790 196.010 ;
        RECT 72.190 194.730 72.450 194.990 ;
        RECT 74.950 194.390 75.210 194.650 ;
        RECT 78.170 194.050 78.430 194.310 ;
        RECT 83.690 195.410 83.950 195.670 ;
        RECT 85.530 195.070 85.790 195.330 ;
        RECT 93.810 195.750 94.070 196.010 ;
        RECT 97.950 195.750 98.210 196.010 ;
        RECT 100.710 195.750 100.970 196.010 ;
        RECT 106.230 195.750 106.490 196.010 ;
        RECT 89.210 195.410 89.470 195.670 ;
        RECT 85.070 194.730 85.330 194.990 ;
        RECT 87.830 194.730 88.090 194.990 ;
        RECT 88.750 194.730 89.010 194.990 ;
        RECT 92.430 195.070 92.690 195.330 ;
        RECT 95.650 195.070 95.910 195.330 ;
        RECT 98.410 195.070 98.670 195.330 ;
        RECT 98.870 195.070 99.130 195.330 ;
        RECT 101.170 195.410 101.430 195.670 ;
        RECT 104.850 195.070 105.110 195.330 ;
        RECT 86.910 194.390 87.170 194.650 ;
        RECT 94.270 194.730 94.530 194.990 ;
        RECT 97.030 194.730 97.290 194.990 ;
        RECT 99.330 194.730 99.590 194.990 ;
        RECT 100.710 194.730 100.970 194.990 ;
        RECT 101.630 194.730 101.890 194.990 ;
        RECT 102.550 194.730 102.810 194.990 ;
        RECT 108.070 195.410 108.330 195.670 ;
        RECT 106.690 194.730 106.950 194.990 ;
        RECT 110.830 195.750 111.090 196.010 ;
        RECT 111.750 195.750 112.010 196.010 ;
        RECT 109.910 195.410 110.170 195.670 ;
        RECT 135.210 195.750 135.470 196.010 ;
        RECT 137.510 195.750 137.770 196.010 ;
        RECT 143.030 195.750 143.290 196.010 ;
        RECT 144.870 195.750 145.130 196.010 ;
        RECT 126.930 195.410 127.190 195.670 ;
        RECT 132.450 195.410 132.710 195.670 ;
        RECT 118.190 195.070 118.450 195.330 ;
        RECT 110.830 194.730 111.090 194.990 ;
        RECT 112.210 194.730 112.470 194.990 ;
        RECT 115.890 194.730 116.150 194.990 ;
        RECT 140.730 195.410 140.990 195.670 ;
        RECT 141.650 195.410 141.910 195.670 ;
        RECT 134.290 195.070 134.550 195.330 ;
        RECT 138.890 195.070 139.150 195.330 ;
        RECT 139.810 195.070 140.070 195.330 ;
        RECT 99.790 194.390 100.050 194.650 ;
        RECT 108.990 194.390 109.250 194.650 ;
        RECT 86.450 194.050 86.710 194.310 ;
        RECT 91.050 194.050 91.310 194.310 ;
        RECT 92.890 194.050 93.150 194.310 ;
        RECT 94.270 194.050 94.530 194.310 ;
        RECT 94.730 194.050 94.990 194.310 ;
        RECT 97.950 194.050 98.210 194.310 ;
        RECT 100.710 194.050 100.970 194.310 ;
        RECT 103.470 194.050 103.730 194.310 ;
        RECT 104.850 194.050 105.110 194.310 ;
        RECT 117.270 194.050 117.530 194.310 ;
        RECT 127.390 194.730 127.650 194.990 ;
        RECT 129.230 194.730 129.490 194.990 ;
        RECT 125.090 194.050 125.350 194.310 ;
        RECT 129.690 194.390 129.950 194.650 ;
        RECT 131.070 194.390 131.330 194.650 ;
        RECT 132.450 194.730 132.710 194.990 ;
        RECT 135.210 194.390 135.470 194.650 ;
        RECT 137.970 194.730 138.230 194.990 ;
        RECT 140.730 194.730 140.990 194.990 ;
        RECT 137.510 194.390 137.770 194.650 ;
        RECT 126.470 194.050 126.730 194.310 ;
        RECT 133.370 194.050 133.630 194.310 ;
        RECT 138.430 194.050 138.690 194.310 ;
        RECT 153.150 194.050 153.410 194.310 ;
        RECT 89.780 193.540 90.040 193.800 ;
        RECT 90.100 193.540 90.360 193.800 ;
        RECT 90.420 193.540 90.680 193.800 ;
        RECT 90.740 193.540 91.000 193.800 ;
        RECT 91.060 193.540 91.320 193.800 ;
        RECT 91.380 193.540 91.640 193.800 ;
        RECT 119.780 193.540 120.040 193.800 ;
        RECT 120.100 193.540 120.360 193.800 ;
        RECT 120.420 193.540 120.680 193.800 ;
        RECT 120.740 193.540 121.000 193.800 ;
        RECT 121.060 193.540 121.320 193.800 ;
        RECT 121.380 193.540 121.640 193.800 ;
        RECT 149.780 193.540 150.040 193.800 ;
        RECT 150.100 193.540 150.360 193.800 ;
        RECT 150.420 193.540 150.680 193.800 ;
        RECT 150.740 193.540 151.000 193.800 ;
        RECT 151.060 193.540 151.320 193.800 ;
        RECT 151.380 193.540 151.640 193.800 ;
        RECT 74.950 193.030 75.210 193.290 ;
        RECT 82.310 193.030 82.570 193.290 ;
        RECT 85.530 193.030 85.790 193.290 ;
        RECT 78.170 192.350 78.430 192.610 ;
        RECT 80.470 192.350 80.730 192.610 ;
        RECT 81.390 192.350 81.650 192.610 ;
        RECT 76.790 192.010 77.050 192.270 ;
        RECT 80.930 192.010 81.190 192.270 ;
        RECT 82.770 192.350 83.030 192.610 ;
        RECT 86.910 192.350 87.170 192.610 ;
        RECT 93.350 193.030 93.610 193.290 ;
        RECT 94.270 193.030 94.530 193.290 ;
        RECT 90.590 192.690 90.850 192.950 ;
        RECT 95.650 192.690 95.910 192.950 ;
        RECT 96.110 192.690 96.370 192.950 ;
        RECT 99.330 192.690 99.590 192.950 ;
        RECT 91.050 192.350 91.310 192.610 ;
        RECT 93.350 192.350 93.610 192.610 ;
        RECT 92.430 192.010 92.690 192.270 ;
        RECT 97.030 192.350 97.290 192.610 ;
        RECT 104.850 193.030 105.110 193.290 ;
        RECT 106.230 193.030 106.490 193.290 ;
        RECT 107.610 192.690 107.870 192.950 ;
        RECT 110.830 193.030 111.090 193.290 ;
        RECT 111.750 193.030 112.010 193.290 ;
        RECT 114.050 193.030 114.310 193.290 ;
        RECT 128.770 193.030 129.030 193.290 ;
        RECT 129.690 193.030 129.950 193.290 ;
        RECT 99.790 192.010 100.050 192.270 ;
        RECT 102.090 192.010 102.350 192.270 ;
        RECT 109.450 192.350 109.710 192.610 ;
        RECT 109.910 192.350 110.170 192.610 ;
        RECT 113.590 192.350 113.850 192.610 ;
        RECT 111.290 192.010 111.550 192.270 ;
        RECT 112.210 192.010 112.470 192.270 ;
        RECT 115.430 192.350 115.690 192.610 ;
        RECT 117.730 192.350 117.990 192.610 ;
        RECT 120.950 192.350 121.210 192.610 ;
        RECT 127.390 192.690 127.650 192.950 ;
        RECT 124.630 192.350 124.890 192.610 ;
        RECT 129.690 192.350 129.950 192.610 ;
        RECT 122.330 192.010 122.590 192.270 ;
        RECT 116.810 191.670 117.070 191.930 ;
        RECT 117.270 191.670 117.530 191.930 ;
        RECT 126.010 192.010 126.270 192.270 ;
        RECT 77.250 191.330 77.510 191.590 ;
        RECT 82.770 191.330 83.030 191.590 ;
        RECT 95.650 191.330 95.910 191.590 ;
        RECT 97.030 191.330 97.290 191.590 ;
        RECT 107.150 191.330 107.410 191.590 ;
        RECT 130.610 192.010 130.870 192.270 ;
        RECT 137.050 192.350 137.310 192.610 ;
        RECT 137.510 192.350 137.770 192.610 ;
        RECT 137.970 192.350 138.230 192.610 ;
        RECT 132.450 192.010 132.710 192.270 ;
        RECT 139.810 192.350 140.070 192.610 ;
        RECT 120.950 191.330 121.210 191.590 ;
        RECT 123.250 191.330 123.510 191.590 ;
        RECT 123.710 191.330 123.970 191.590 ;
        RECT 125.550 191.330 125.810 191.590 ;
        RECT 126.470 191.330 126.730 191.590 ;
        RECT 126.930 191.330 127.190 191.590 ;
        RECT 137.970 191.670 138.230 191.930 ;
        RECT 147.630 192.350 147.890 192.610 ;
        RECT 146.710 191.670 146.970 191.930 ;
        RECT 148.090 191.670 148.350 191.930 ;
        RECT 130.150 191.330 130.410 191.590 ;
        RECT 131.530 191.330 131.790 191.590 ;
        RECT 74.780 190.820 75.040 191.080 ;
        RECT 75.100 190.820 75.360 191.080 ;
        RECT 75.420 190.820 75.680 191.080 ;
        RECT 75.740 190.820 76.000 191.080 ;
        RECT 76.060 190.820 76.320 191.080 ;
        RECT 76.380 190.820 76.640 191.080 ;
        RECT 104.780 190.820 105.040 191.080 ;
        RECT 105.100 190.820 105.360 191.080 ;
        RECT 105.420 190.820 105.680 191.080 ;
        RECT 105.740 190.820 106.000 191.080 ;
        RECT 106.060 190.820 106.320 191.080 ;
        RECT 106.380 190.820 106.640 191.080 ;
        RECT 134.780 190.820 135.040 191.080 ;
        RECT 135.100 190.820 135.360 191.080 ;
        RECT 135.420 190.820 135.680 191.080 ;
        RECT 135.740 190.820 136.000 191.080 ;
        RECT 136.060 190.820 136.320 191.080 ;
        RECT 136.380 190.820 136.640 191.080 ;
        RECT 85.070 190.310 85.330 190.570 ;
        RECT 92.890 190.310 93.150 190.570 ;
        RECT 94.730 190.310 94.990 190.570 ;
        RECT 77.250 189.970 77.510 190.230 ;
        RECT 80.470 189.630 80.730 189.890 ;
        RECT 85.990 189.630 86.250 189.890 ;
        RECT 89.670 189.630 89.930 189.890 ;
        RECT 80.930 189.290 81.190 189.550 ;
        RECT 86.450 189.290 86.710 189.550 ;
        RECT 87.370 189.290 87.630 189.550 ;
        RECT 87.830 189.290 88.090 189.550 ;
        RECT 88.290 189.290 88.550 189.550 ;
        RECT 89.210 189.290 89.470 189.550 ;
        RECT 91.970 189.290 92.230 189.550 ;
        RECT 94.270 189.290 94.530 189.550 ;
        RECT 97.030 190.310 97.290 190.570 ;
        RECT 101.170 190.310 101.430 190.570 ;
        RECT 102.090 190.310 102.350 190.570 ;
        RECT 103.930 190.310 104.190 190.570 ;
        RECT 100.250 189.970 100.510 190.230 ;
        RECT 108.070 190.310 108.330 190.570 ;
        RECT 98.410 189.630 98.670 189.890 ;
        RECT 99.330 189.290 99.590 189.550 ;
        RECT 104.390 189.630 104.650 189.890 ;
        RECT 108.990 189.630 109.250 189.890 ;
        RECT 109.450 189.630 109.710 189.890 ;
        RECT 111.750 189.630 112.010 189.890 ;
        RECT 89.210 188.610 89.470 188.870 ;
        RECT 97.950 188.610 98.210 188.870 ;
        RECT 99.790 188.950 100.050 189.210 ;
        RECT 104.850 189.290 105.110 189.550 ;
        RECT 106.690 189.290 106.950 189.550 ;
        RECT 107.610 189.290 107.870 189.550 ;
        RECT 114.050 190.310 114.310 190.570 ;
        RECT 120.950 190.310 121.210 190.570 ;
        RECT 126.930 190.310 127.190 190.570 ;
        RECT 122.790 189.970 123.050 190.230 ;
        RECT 124.170 189.970 124.430 190.230 ;
        RECT 128.770 189.970 129.030 190.230 ;
        RECT 129.230 189.970 129.490 190.230 ;
        RECT 115.430 189.290 115.690 189.550 ;
        RECT 115.890 189.290 116.150 189.550 ;
        RECT 113.590 188.950 113.850 189.210 ;
        RECT 116.350 188.950 116.610 189.210 ;
        RECT 118.190 188.950 118.450 189.210 ;
        RECT 128.310 189.630 128.570 189.890 ;
        RECT 109.910 188.610 110.170 188.870 ;
        RECT 111.750 188.610 112.010 188.870 ;
        RECT 117.270 188.610 117.530 188.870 ;
        RECT 119.110 188.610 119.370 188.870 ;
        RECT 123.250 188.950 123.510 189.210 ;
        RECT 124.630 188.950 124.890 189.210 ;
        RECT 126.010 188.950 126.270 189.210 ;
        RECT 127.390 189.290 127.650 189.550 ;
        RECT 136.590 190.310 136.850 190.570 ;
        RECT 138.430 190.310 138.690 190.570 ;
        RECT 137.970 189.970 138.230 190.230 ;
        RECT 137.510 189.630 137.770 189.890 ;
        RECT 130.610 189.290 130.870 189.550 ;
        RECT 131.070 189.290 131.330 189.550 ;
        RECT 139.810 189.290 140.070 189.550 ;
        RECT 120.950 188.610 121.210 188.870 ;
        RECT 130.150 188.610 130.410 188.870 ;
        RECT 137.050 188.610 137.310 188.870 ;
        RECT 138.430 188.950 138.690 189.210 ;
        RECT 146.710 189.290 146.970 189.550 ;
        RECT 147.630 189.970 147.890 190.230 ;
        RECT 153.610 189.970 153.870 190.230 ;
        RECT 149.010 189.630 149.270 189.890 ;
        RECT 149.930 189.630 150.190 189.890 ;
        RECT 151.770 189.290 152.030 189.550 ;
        RECT 152.230 189.290 152.490 189.550 ;
        RECT 141.650 188.950 141.910 189.210 ;
        RECT 153.150 188.950 153.410 189.210 ;
        RECT 154.990 188.610 155.250 188.870 ;
        RECT 89.780 188.100 90.040 188.360 ;
        RECT 90.100 188.100 90.360 188.360 ;
        RECT 90.420 188.100 90.680 188.360 ;
        RECT 90.740 188.100 91.000 188.360 ;
        RECT 91.060 188.100 91.320 188.360 ;
        RECT 91.380 188.100 91.640 188.360 ;
        RECT 119.780 188.100 120.040 188.360 ;
        RECT 120.100 188.100 120.360 188.360 ;
        RECT 120.420 188.100 120.680 188.360 ;
        RECT 120.740 188.100 121.000 188.360 ;
        RECT 121.060 188.100 121.320 188.360 ;
        RECT 121.380 188.100 121.640 188.360 ;
        RECT 149.780 188.100 150.040 188.360 ;
        RECT 150.100 188.100 150.360 188.360 ;
        RECT 150.420 188.100 150.680 188.360 ;
        RECT 150.740 188.100 151.000 188.360 ;
        RECT 151.060 188.100 151.320 188.360 ;
        RECT 151.380 188.100 151.640 188.360 ;
        RECT 78.630 187.590 78.890 187.850 ;
        RECT 80.930 187.250 81.190 187.510 ;
        RECT 85.530 187.590 85.790 187.850 ;
        RECT 85.990 187.590 86.250 187.850 ;
        RECT 87.830 187.590 88.090 187.850 ;
        RECT 89.670 187.590 89.930 187.850 ;
        RECT 74.030 186.910 74.290 187.170 ;
        RECT 72.190 186.570 72.450 186.830 ;
        RECT 79.550 185.890 79.810 186.150 ;
        RECT 80.010 185.890 80.270 186.150 ;
        RECT 80.470 185.890 80.730 186.150 ;
        RECT 84.150 185.890 84.410 186.150 ;
        RECT 99.790 187.250 100.050 187.510 ;
        RECT 102.550 187.590 102.810 187.850 ;
        RECT 106.230 187.590 106.490 187.850 ;
        RECT 113.590 187.590 113.850 187.850 ;
        RECT 118.190 187.590 118.450 187.850 ;
        RECT 122.330 187.590 122.590 187.850 ;
        RECT 128.310 187.590 128.570 187.850 ;
        RECT 102.090 187.250 102.350 187.510 ;
        RECT 104.850 187.250 105.110 187.510 ;
        RECT 107.610 187.250 107.870 187.510 ;
        RECT 89.670 186.910 89.930 187.170 ;
        RECT 91.050 186.910 91.310 187.170 ;
        RECT 92.430 186.910 92.690 187.170 ;
        RECT 94.730 186.570 94.990 186.830 ;
        RECT 96.110 186.910 96.370 187.170 ;
        RECT 98.410 186.910 98.670 187.170 ;
        RECT 102.550 186.910 102.810 187.170 ;
        RECT 109.910 187.250 110.170 187.510 ;
        RECT 115.890 187.250 116.150 187.510 ;
        RECT 110.830 186.910 111.090 187.170 ;
        RECT 111.290 186.910 111.550 187.170 ;
        RECT 114.970 186.910 115.230 187.170 ;
        RECT 107.150 186.570 107.410 186.830 ;
        RECT 116.810 186.570 117.070 186.830 ;
        RECT 92.890 186.230 93.150 186.490 ;
        RECT 96.570 186.230 96.830 186.490 ;
        RECT 116.350 186.230 116.610 186.490 ;
        RECT 119.110 187.250 119.370 187.510 ;
        RECT 131.070 187.250 131.330 187.510 ;
        RECT 131.990 187.590 132.250 187.850 ;
        RECT 132.450 187.590 132.710 187.850 ;
        RECT 133.370 187.590 133.630 187.850 ;
        RECT 134.750 187.250 135.010 187.510 ;
        RECT 146.710 187.590 146.970 187.850 ;
        RECT 137.970 187.250 138.230 187.510 ;
        RECT 153.610 187.590 153.870 187.850 ;
        RECT 120.950 186.910 121.210 187.170 ;
        RECT 124.630 186.910 124.890 187.170 ;
        RECT 125.550 186.910 125.810 187.170 ;
        RECT 128.770 186.910 129.030 187.170 ;
        RECT 137.050 186.910 137.310 187.170 ;
        RECT 142.570 186.910 142.830 187.170 ;
        RECT 145.790 186.910 146.050 187.170 ;
        RECT 147.630 186.910 147.890 187.170 ;
        RECT 148.090 186.910 148.350 187.170 ;
        RECT 149.930 186.910 150.190 187.170 ;
        RECT 119.110 186.230 119.370 186.490 ;
        RECT 119.570 186.230 119.830 186.490 ;
        RECT 93.810 185.890 94.070 186.150 ;
        RECT 107.610 185.890 107.870 186.150 ;
        RECT 117.270 185.890 117.530 186.150 ;
        RECT 120.950 185.890 121.210 186.150 ;
        RECT 121.410 185.890 121.670 186.150 ;
        RECT 125.090 186.570 125.350 186.830 ;
        RECT 140.730 186.570 140.990 186.830 ;
        RECT 151.770 186.910 152.030 187.170 ;
        RECT 141.650 186.230 141.910 186.490 ;
        RECT 144.410 186.230 144.670 186.490 ;
        RECT 133.830 185.890 134.090 186.150 ;
        RECT 144.870 185.890 145.130 186.150 ;
        RECT 146.710 185.890 146.970 186.150 ;
        RECT 153.610 185.890 153.870 186.150 ;
        RECT 74.780 185.380 75.040 185.640 ;
        RECT 75.100 185.380 75.360 185.640 ;
        RECT 75.420 185.380 75.680 185.640 ;
        RECT 75.740 185.380 76.000 185.640 ;
        RECT 76.060 185.380 76.320 185.640 ;
        RECT 76.380 185.380 76.640 185.640 ;
        RECT 104.780 185.380 105.040 185.640 ;
        RECT 105.100 185.380 105.360 185.640 ;
        RECT 105.420 185.380 105.680 185.640 ;
        RECT 105.740 185.380 106.000 185.640 ;
        RECT 106.060 185.380 106.320 185.640 ;
        RECT 106.380 185.380 106.640 185.640 ;
        RECT 134.780 185.380 135.040 185.640 ;
        RECT 135.100 185.380 135.360 185.640 ;
        RECT 135.420 185.380 135.680 185.640 ;
        RECT 135.740 185.380 136.000 185.640 ;
        RECT 136.060 185.380 136.320 185.640 ;
        RECT 136.380 185.380 136.640 185.640 ;
        RECT 74.030 184.870 74.290 185.130 ;
        RECT 76.790 184.870 77.050 185.130 ;
        RECT 82.310 184.870 82.570 185.130 ;
        RECT 76.330 184.530 76.590 184.790 ;
        RECT 94.730 184.870 94.990 185.130 ;
        RECT 97.490 184.870 97.750 185.130 ;
        RECT 103.010 184.870 103.270 185.130 ;
        RECT 109.910 184.870 110.170 185.130 ;
        RECT 115.430 184.870 115.690 185.130 ;
        RECT 116.350 184.870 116.610 185.130 ;
        RECT 91.050 184.530 91.310 184.790 ;
        RECT 76.790 183.850 77.050 184.110 ;
        RECT 93.810 184.190 94.070 184.450 ;
        RECT 100.710 184.190 100.970 184.450 ;
        RECT 101.170 184.190 101.430 184.450 ;
        RECT 126.930 184.530 127.190 184.790 ;
        RECT 116.810 184.190 117.070 184.450 ;
        RECT 125.090 184.190 125.350 184.450 ;
        RECT 77.710 183.850 77.970 184.110 ;
        RECT 80.010 183.850 80.270 184.110 ;
        RECT 93.350 183.850 93.610 184.110 ;
        RECT 80.930 183.510 81.190 183.770 ;
        RECT 81.850 183.170 82.110 183.430 ;
        RECT 82.770 183.170 83.030 183.430 ;
        RECT 83.230 183.170 83.490 183.430 ;
        RECT 85.530 183.510 85.790 183.770 ;
        RECT 85.990 183.510 86.250 183.770 ;
        RECT 88.750 183.510 89.010 183.770 ;
        RECT 92.430 183.170 92.690 183.430 ;
        RECT 99.330 183.850 99.590 184.110 ;
        RECT 98.870 183.510 99.130 183.770 ;
        RECT 103.470 183.850 103.730 184.110 ;
        RECT 109.910 183.850 110.170 184.110 ;
        RECT 115.890 183.850 116.150 184.110 ;
        RECT 101.630 183.510 101.890 183.770 ;
        RECT 102.090 183.510 102.350 183.770 ;
        RECT 109.450 183.510 109.710 183.770 ;
        RECT 103.010 183.170 103.270 183.430 ;
        RECT 107.150 183.170 107.410 183.430 ;
        RECT 114.970 183.510 115.230 183.770 ;
        RECT 121.410 183.850 121.670 184.110 ;
        RECT 127.850 184.190 128.110 184.450 ;
        RECT 128.770 184.190 129.030 184.450 ;
        RECT 130.610 184.190 130.870 184.450 ;
        RECT 117.730 183.510 117.990 183.770 ;
        RECT 111.290 183.170 111.550 183.430 ;
        RECT 113.590 183.170 113.850 183.430 ;
        RECT 115.430 183.170 115.690 183.430 ;
        RECT 119.570 183.510 119.830 183.770 ;
        RECT 122.330 183.510 122.590 183.770 ;
        RECT 131.990 184.190 132.250 184.450 ;
        RECT 134.290 184.870 134.550 185.130 ;
        RECT 140.730 184.870 140.990 185.130 ;
        RECT 152.230 184.870 152.490 185.130 ;
        RECT 154.070 184.870 154.330 185.130 ;
        RECT 131.070 183.850 131.330 184.110 ;
        RECT 136.590 183.850 136.850 184.110 ;
        RECT 137.970 183.850 138.230 184.110 ;
        RECT 139.350 183.850 139.610 184.110 ;
        RECT 142.570 183.850 142.830 184.110 ;
        RECT 143.950 183.850 144.210 184.110 ;
        RECT 153.610 183.850 153.870 184.110 ;
        RECT 133.370 183.510 133.630 183.770 ;
        RECT 138.890 183.510 139.150 183.770 ;
        RECT 144.410 183.510 144.670 183.770 ;
        RECT 145.330 183.510 145.590 183.770 ;
        RECT 149.930 183.510 150.190 183.770 ;
        RECT 126.930 183.170 127.190 183.430 ;
        RECT 131.070 183.170 131.330 183.430 ;
        RECT 131.990 183.170 132.250 183.430 ;
        RECT 136.130 183.170 136.390 183.430 ;
        RECT 142.110 183.170 142.370 183.430 ;
        RECT 147.630 183.170 147.890 183.430 ;
        RECT 89.780 182.660 90.040 182.920 ;
        RECT 90.100 182.660 90.360 182.920 ;
        RECT 90.420 182.660 90.680 182.920 ;
        RECT 90.740 182.660 91.000 182.920 ;
        RECT 91.060 182.660 91.320 182.920 ;
        RECT 91.380 182.660 91.640 182.920 ;
        RECT 119.780 182.660 120.040 182.920 ;
        RECT 120.100 182.660 120.360 182.920 ;
        RECT 120.420 182.660 120.680 182.920 ;
        RECT 120.740 182.660 121.000 182.920 ;
        RECT 121.060 182.660 121.320 182.920 ;
        RECT 121.380 182.660 121.640 182.920 ;
        RECT 149.780 182.660 150.040 182.920 ;
        RECT 150.100 182.660 150.360 182.920 ;
        RECT 150.420 182.660 150.680 182.920 ;
        RECT 150.740 182.660 151.000 182.920 ;
        RECT 151.060 182.660 151.320 182.920 ;
        RECT 151.380 182.660 151.640 182.920 ;
        RECT 82.770 182.150 83.030 182.410 ;
        RECT 85.530 182.150 85.790 182.410 ;
        RECT 88.750 182.150 89.010 182.410 ;
        RECT 102.090 182.150 102.350 182.410 ;
        RECT 107.610 182.150 107.870 182.410 ;
        RECT 109.910 182.150 110.170 182.410 ;
        RECT 130.610 182.150 130.870 182.410 ;
        RECT 134.290 182.150 134.550 182.410 ;
        RECT 73.570 181.470 73.830 181.730 ;
        RECT 82.770 181.470 83.030 181.730 ;
        RECT 96.570 181.810 96.830 182.070 ;
        RECT 72.190 181.130 72.450 181.390 ;
        RECT 79.090 181.130 79.350 181.390 ;
        RECT 89.210 181.130 89.470 181.390 ;
        RECT 98.870 181.470 99.130 181.730 ;
        RECT 100.250 181.810 100.510 182.070 ;
        RECT 101.630 181.470 101.890 181.730 ;
        RECT 104.390 181.470 104.650 181.730 ;
        RECT 109.450 181.810 109.710 182.070 ;
        RECT 124.170 181.810 124.430 182.070 ;
        RECT 78.630 180.450 78.890 180.710 ;
        RECT 85.070 180.450 85.330 180.710 ;
        RECT 92.890 180.790 93.150 181.050 ;
        RECT 101.170 181.130 101.430 181.390 ;
        RECT 103.470 180.790 103.730 181.050 ;
        RECT 107.150 181.130 107.410 181.390 ;
        RECT 109.450 181.130 109.710 181.390 ;
        RECT 114.510 181.470 114.770 181.730 ;
        RECT 122.790 181.470 123.050 181.730 ;
        RECT 126.470 181.470 126.730 181.730 ;
        RECT 108.530 180.790 108.790 181.050 ;
        RECT 110.830 180.790 111.090 181.050 ;
        RECT 112.670 180.790 112.930 181.050 ;
        RECT 114.970 180.790 115.230 181.050 ;
        RECT 92.430 180.450 92.690 180.710 ;
        RECT 100.710 180.450 100.970 180.710 ;
        RECT 103.930 180.450 104.190 180.710 ;
        RECT 106.690 180.450 106.950 180.710 ;
        RECT 107.610 180.450 107.870 180.710 ;
        RECT 110.370 180.450 110.630 180.710 ;
        RECT 124.630 180.450 124.890 180.710 ;
        RECT 130.610 180.450 130.870 180.710 ;
        RECT 131.990 180.450 132.250 180.710 ;
        RECT 136.130 181.810 136.390 182.070 ;
        RECT 140.730 181.810 140.990 182.070 ;
        RECT 145.330 182.150 145.590 182.410 ;
        RECT 152.690 182.150 152.950 182.410 ;
        RECT 154.070 182.150 154.330 182.410 ;
        RECT 137.050 181.470 137.310 181.730 ;
        RECT 137.510 181.470 137.770 181.730 ;
        RECT 139.350 180.790 139.610 181.050 ;
        RECT 142.570 180.450 142.830 180.710 ;
        RECT 143.950 180.450 144.210 180.710 ;
        RECT 153.150 181.130 153.410 181.390 ;
        RECT 154.990 181.130 155.250 181.390 ;
        RECT 149.010 180.450 149.270 180.710 ;
        RECT 152.690 180.450 152.950 180.710 ;
        RECT 74.780 179.940 75.040 180.200 ;
        RECT 75.100 179.940 75.360 180.200 ;
        RECT 75.420 179.940 75.680 180.200 ;
        RECT 75.740 179.940 76.000 180.200 ;
        RECT 76.060 179.940 76.320 180.200 ;
        RECT 76.380 179.940 76.640 180.200 ;
        RECT 104.780 179.940 105.040 180.200 ;
        RECT 105.100 179.940 105.360 180.200 ;
        RECT 105.420 179.940 105.680 180.200 ;
        RECT 105.740 179.940 106.000 180.200 ;
        RECT 106.060 179.940 106.320 180.200 ;
        RECT 106.380 179.940 106.640 180.200 ;
        RECT 134.780 179.940 135.040 180.200 ;
        RECT 135.100 179.940 135.360 180.200 ;
        RECT 135.420 179.940 135.680 180.200 ;
        RECT 135.740 179.940 136.000 180.200 ;
        RECT 136.060 179.940 136.320 180.200 ;
        RECT 136.380 179.940 136.640 180.200 ;
        RECT 73.570 179.430 73.830 179.690 ;
        RECT 76.790 179.430 77.050 179.690 ;
        RECT 81.390 179.430 81.650 179.690 ;
        RECT 83.690 179.430 83.950 179.690 ;
        RECT 104.390 179.430 104.650 179.690 ;
        RECT 107.150 179.430 107.410 179.690 ;
        RECT 80.930 179.090 81.190 179.350 ;
        RECT 84.610 179.090 84.870 179.350 ;
        RECT 78.170 178.410 78.430 178.670 ;
        RECT 80.010 178.410 80.270 178.670 ;
        RECT 98.870 179.090 99.130 179.350 ;
        RECT 114.970 179.430 115.230 179.690 ;
        RECT 126.470 179.430 126.730 179.690 ;
        RECT 133.370 179.430 133.630 179.690 ;
        RECT 85.990 178.750 86.250 179.010 ;
        RECT 97.490 178.750 97.750 179.010 ;
        RECT 99.790 178.750 100.050 179.010 ;
        RECT 101.170 178.750 101.430 179.010 ;
        RECT 114.510 179.090 114.770 179.350 ;
        RECT 87.830 178.410 88.090 178.670 ;
        RECT 89.670 178.410 89.930 178.670 ;
        RECT 91.970 178.410 92.230 178.670 ;
        RECT 77.710 177.730 77.970 177.990 ;
        RECT 85.070 178.070 85.330 178.330 ;
        RECT 100.250 178.410 100.510 178.670 ;
        RECT 103.010 178.410 103.270 178.670 ;
        RECT 106.230 178.410 106.490 178.670 ;
        RECT 106.690 178.410 106.950 178.670 ;
        RECT 108.070 178.410 108.330 178.670 ;
        RECT 98.870 178.070 99.130 178.330 ;
        RECT 88.750 177.730 89.010 177.990 ;
        RECT 92.890 177.730 93.150 177.990 ;
        RECT 94.730 177.730 94.990 177.990 ;
        RECT 104.850 177.730 105.110 177.990 ;
        RECT 113.130 178.410 113.390 178.670 ;
        RECT 113.590 178.070 113.850 178.330 ;
        RECT 114.970 178.410 115.230 178.670 ;
        RECT 115.430 178.410 115.690 178.670 ;
        RECT 115.890 178.070 116.150 178.330 ;
        RECT 117.730 178.410 117.990 178.670 ;
        RECT 119.110 178.750 119.370 179.010 ;
        RECT 124.170 178.410 124.430 178.670 ;
        RECT 133.830 179.090 134.090 179.350 ;
        RECT 145.790 179.430 146.050 179.690 ;
        RECT 142.110 179.090 142.370 179.350 ;
        RECT 126.470 178.410 126.730 178.670 ;
        RECT 131.990 178.750 132.250 179.010 ;
        RECT 128.310 178.070 128.570 178.330 ;
        RECT 116.350 177.730 116.610 177.990 ;
        RECT 118.650 177.730 118.910 177.990 ;
        RECT 123.250 177.730 123.510 177.990 ;
        RECT 125.550 177.730 125.810 177.990 ;
        RECT 133.370 178.410 133.630 178.670 ;
        RECT 137.050 178.750 137.310 179.010 ;
        RECT 129.690 177.730 129.950 177.990 ;
        RECT 131.530 177.730 131.790 177.990 ;
        RECT 136.590 177.730 136.850 177.990 ;
        RECT 141.650 178.410 141.910 178.670 ;
        RECT 142.570 178.410 142.830 178.670 ;
        RECT 139.810 177.730 140.070 177.990 ;
        RECT 143.490 178.070 143.750 178.330 ;
        RECT 148.550 178.070 148.810 178.330 ;
        RECT 89.780 177.220 90.040 177.480 ;
        RECT 90.100 177.220 90.360 177.480 ;
        RECT 90.420 177.220 90.680 177.480 ;
        RECT 90.740 177.220 91.000 177.480 ;
        RECT 91.060 177.220 91.320 177.480 ;
        RECT 91.380 177.220 91.640 177.480 ;
        RECT 119.780 177.220 120.040 177.480 ;
        RECT 120.100 177.220 120.360 177.480 ;
        RECT 120.420 177.220 120.680 177.480 ;
        RECT 120.740 177.220 121.000 177.480 ;
        RECT 121.060 177.220 121.320 177.480 ;
        RECT 121.380 177.220 121.640 177.480 ;
        RECT 149.780 177.220 150.040 177.480 ;
        RECT 150.100 177.220 150.360 177.480 ;
        RECT 150.420 177.220 150.680 177.480 ;
        RECT 150.740 177.220 151.000 177.480 ;
        RECT 151.060 177.220 151.320 177.480 ;
        RECT 151.380 177.220 151.640 177.480 ;
        RECT 76.790 176.710 77.050 176.970 ;
        RECT 80.010 176.710 80.270 176.970 ;
        RECT 89.670 176.710 89.930 176.970 ;
        RECT 72.190 176.370 72.450 176.630 ;
        RECT 77.710 176.030 77.970 176.290 ;
        RECT 88.290 176.370 88.550 176.630 ;
        RECT 88.750 176.370 89.010 176.630 ;
        RECT 91.970 176.710 92.230 176.970 ;
        RECT 102.550 176.710 102.810 176.970 ;
        RECT 107.610 176.710 107.870 176.970 ;
        RECT 108.070 176.710 108.330 176.970 ;
        RECT 109.910 176.710 110.170 176.970 ;
        RECT 110.830 176.710 111.090 176.970 ;
        RECT 113.130 176.710 113.390 176.970 ;
        RECT 115.890 176.710 116.150 176.970 ;
        RECT 119.110 176.710 119.370 176.970 ;
        RECT 124.170 176.710 124.430 176.970 ;
        RECT 126.470 176.710 126.730 176.970 ;
        RECT 129.690 176.710 129.950 176.970 ;
        RECT 132.450 176.710 132.710 176.970 ;
        RECT 133.370 176.710 133.630 176.970 ;
        RECT 137.510 176.710 137.770 176.970 ;
        RECT 148.550 176.710 148.810 176.970 ;
        RECT 149.010 176.710 149.270 176.970 ;
        RECT 152.690 176.710 152.950 176.970 ;
        RECT 79.550 175.690 79.810 175.950 ;
        RECT 79.550 175.010 79.810 175.270 ;
        RECT 85.990 176.030 86.250 176.290 ;
        RECT 88.750 175.690 89.010 175.950 ;
        RECT 91.970 176.030 92.230 176.290 ;
        RECT 92.890 176.030 93.150 176.290 ;
        RECT 93.350 176.030 93.610 176.290 ;
        RECT 93.810 175.350 94.070 175.610 ;
        RECT 97.030 176.030 97.290 176.290 ;
        RECT 96.570 175.690 96.830 175.950 ;
        RECT 99.790 175.690 100.050 175.950 ;
        RECT 101.170 176.030 101.430 176.290 ;
        RECT 101.630 176.030 101.890 176.290 ;
        RECT 102.090 176.030 102.350 176.290 ;
        RECT 104.850 176.030 105.110 176.290 ;
        RECT 108.070 176.030 108.330 176.290 ;
        RECT 114.050 176.030 114.310 176.290 ;
        RECT 124.630 176.370 124.890 176.630 ;
        RECT 141.650 176.370 141.910 176.630 ;
        RECT 126.010 176.030 126.270 176.290 ;
        RECT 131.530 176.030 131.790 176.290 ;
        RECT 138.430 176.030 138.690 176.290 ;
        RECT 142.570 176.030 142.830 176.290 ;
        RECT 143.490 176.030 143.750 176.290 ;
        RECT 108.530 175.690 108.790 175.950 ;
        RECT 84.610 175.010 84.870 175.270 ;
        RECT 86.450 175.010 86.710 175.270 ;
        RECT 94.730 175.010 94.990 175.270 ;
        RECT 95.650 175.010 95.910 175.270 ;
        RECT 100.250 175.010 100.510 175.270 ;
        RECT 101.630 175.010 101.890 175.270 ;
        RECT 110.830 175.350 111.090 175.610 ;
        RECT 114.510 175.690 114.770 175.950 ;
        RECT 117.730 175.690 117.990 175.950 ;
        RECT 123.250 175.690 123.510 175.950 ;
        RECT 129.230 175.690 129.490 175.950 ;
        RECT 140.730 175.690 140.990 175.950 ;
        RECT 143.030 175.690 143.290 175.950 ;
        RECT 136.130 175.350 136.390 175.610 ;
        RECT 139.350 175.350 139.610 175.610 ;
        RECT 115.890 175.010 116.150 175.270 ;
        RECT 118.650 175.010 118.910 175.270 ;
        RECT 123.710 175.010 123.970 175.270 ;
        RECT 128.310 175.010 128.570 175.270 ;
        RECT 140.730 175.010 140.990 175.270 ;
        RECT 149.470 176.030 149.730 176.290 ;
        RECT 150.850 176.030 151.110 176.290 ;
        RECT 155.450 175.350 155.710 175.610 ;
        RECT 147.170 175.010 147.430 175.270 ;
        RECT 74.780 174.500 75.040 174.760 ;
        RECT 75.100 174.500 75.360 174.760 ;
        RECT 75.420 174.500 75.680 174.760 ;
        RECT 75.740 174.500 76.000 174.760 ;
        RECT 76.060 174.500 76.320 174.760 ;
        RECT 76.380 174.500 76.640 174.760 ;
        RECT 104.780 174.500 105.040 174.760 ;
        RECT 105.100 174.500 105.360 174.760 ;
        RECT 105.420 174.500 105.680 174.760 ;
        RECT 105.740 174.500 106.000 174.760 ;
        RECT 106.060 174.500 106.320 174.760 ;
        RECT 106.380 174.500 106.640 174.760 ;
        RECT 134.780 174.500 135.040 174.760 ;
        RECT 135.100 174.500 135.360 174.760 ;
        RECT 135.420 174.500 135.680 174.760 ;
        RECT 135.740 174.500 136.000 174.760 ;
        RECT 136.060 174.500 136.320 174.760 ;
        RECT 136.380 174.500 136.640 174.760 ;
        RECT 89.210 173.990 89.470 174.250 ;
        RECT 97.030 173.990 97.290 174.250 ;
        RECT 102.550 173.990 102.810 174.250 ;
        RECT 103.010 173.990 103.270 174.250 ;
        RECT 89.670 173.650 89.930 173.910 ;
        RECT 100.250 173.650 100.510 173.910 ;
        RECT 100.710 173.650 100.970 173.910 ;
        RECT 108.070 173.990 108.330 174.250 ;
        RECT 114.970 173.990 115.230 174.250 ;
        RECT 115.890 173.990 116.150 174.250 ;
        RECT 131.990 173.990 132.250 174.250 ;
        RECT 133.830 173.990 134.090 174.250 ;
        RECT 137.510 173.990 137.770 174.250 ;
        RECT 142.110 173.990 142.370 174.250 ;
        RECT 149.470 173.990 149.730 174.250 ;
        RECT 88.290 173.310 88.550 173.570 ;
        RECT 94.270 173.310 94.530 173.570 ;
        RECT 76.790 172.970 77.050 173.230 ;
        RECT 79.550 172.970 79.810 173.230 ;
        RECT 91.050 172.970 91.310 173.230 ;
        RECT 93.350 172.970 93.610 173.230 ;
        RECT 99.790 173.310 100.050 173.570 ;
        RECT 94.270 172.630 94.530 172.890 ;
        RECT 75.870 172.290 76.130 172.550 ;
        RECT 89.210 172.290 89.470 172.550 ;
        RECT 94.730 172.290 94.990 172.550 ;
        RECT 99.790 172.630 100.050 172.890 ;
        RECT 100.250 172.630 100.510 172.890 ;
        RECT 102.090 172.970 102.350 173.230 ;
        RECT 103.470 173.310 103.730 173.570 ;
        RECT 107.610 173.650 107.870 173.910 ;
        RECT 110.830 173.650 111.090 173.910 ;
        RECT 113.130 173.650 113.390 173.910 ;
        RECT 124.170 173.650 124.430 173.910 ;
        RECT 124.630 173.650 124.890 173.910 ;
        RECT 105.310 172.970 105.570 173.230 ;
        RECT 108.530 173.310 108.790 173.570 ;
        RECT 101.630 172.630 101.890 172.890 ;
        RECT 104.850 172.630 105.110 172.890 ;
        RECT 96.570 172.290 96.830 172.550 ;
        RECT 99.330 172.290 99.590 172.550 ;
        RECT 103.470 172.290 103.730 172.550 ;
        RECT 106.230 172.290 106.490 172.550 ;
        RECT 122.330 172.970 122.590 173.230 ;
        RECT 131.530 173.310 131.790 173.570 ;
        RECT 126.470 172.970 126.730 173.230 ;
        RECT 137.970 173.310 138.230 173.570 ;
        RECT 143.950 173.650 144.210 173.910 ;
        RECT 147.170 173.650 147.430 173.910 ;
        RECT 144.410 173.310 144.670 173.570 ;
        RECT 145.790 173.310 146.050 173.570 ;
        RECT 149.010 173.310 149.270 173.570 ;
        RECT 113.130 172.630 113.390 172.890 ;
        RECT 134.750 172.970 135.010 173.230 ;
        RECT 137.050 172.970 137.310 173.230 ;
        RECT 138.430 172.970 138.690 173.230 ;
        RECT 110.370 172.290 110.630 172.550 ;
        RECT 110.830 172.290 111.090 172.550 ;
        RECT 119.110 172.290 119.370 172.550 ;
        RECT 139.810 172.630 140.070 172.890 ;
        RECT 147.170 172.970 147.430 173.230 ;
        RECT 135.670 172.290 135.930 172.550 ;
        RECT 143.490 172.630 143.750 172.890 ;
        RECT 149.010 172.290 149.270 172.550 ;
        RECT 152.690 172.290 152.950 172.550 ;
        RECT 89.780 171.780 90.040 172.040 ;
        RECT 90.100 171.780 90.360 172.040 ;
        RECT 90.420 171.780 90.680 172.040 ;
        RECT 90.740 171.780 91.000 172.040 ;
        RECT 91.060 171.780 91.320 172.040 ;
        RECT 91.380 171.780 91.640 172.040 ;
        RECT 119.780 171.780 120.040 172.040 ;
        RECT 120.100 171.780 120.360 172.040 ;
        RECT 120.420 171.780 120.680 172.040 ;
        RECT 120.740 171.780 121.000 172.040 ;
        RECT 121.060 171.780 121.320 172.040 ;
        RECT 121.380 171.780 121.640 172.040 ;
        RECT 149.780 171.780 150.040 172.040 ;
        RECT 150.100 171.780 150.360 172.040 ;
        RECT 150.420 171.780 150.680 172.040 ;
        RECT 150.740 171.780 151.000 172.040 ;
        RECT 151.060 171.780 151.320 172.040 ;
        RECT 151.380 171.780 151.640 172.040 ;
        RECT 87.830 171.270 88.090 171.530 ;
        RECT 88.750 171.270 89.010 171.530 ;
        RECT 91.510 171.270 91.770 171.530 ;
        RECT 92.890 171.270 93.150 171.530 ;
        RECT 93.350 171.270 93.610 171.530 ;
        RECT 94.730 171.270 94.990 171.530 ;
        RECT 97.490 171.270 97.750 171.530 ;
        RECT 99.790 171.270 100.050 171.530 ;
        RECT 113.590 171.270 113.850 171.530 ;
        RECT 120.030 171.270 120.290 171.530 ;
        RECT 124.630 171.270 124.890 171.530 ;
        RECT 129.690 171.270 129.950 171.530 ;
        RECT 130.610 171.270 130.870 171.530 ;
        RECT 131.990 171.270 132.250 171.530 ;
        RECT 137.050 171.270 137.310 171.530 ;
        RECT 143.950 171.270 144.210 171.530 ;
        RECT 144.410 171.270 144.670 171.530 ;
        RECT 75.870 170.590 76.130 170.850 ;
        RECT 87.370 170.590 87.630 170.850 ;
        RECT 88.290 170.590 88.550 170.850 ;
        RECT 91.970 170.590 92.230 170.850 ;
        RECT 93.350 170.590 93.610 170.850 ;
        RECT 72.190 170.250 72.450 170.510 ;
        RECT 89.670 170.250 89.930 170.510 ;
        RECT 94.270 170.590 94.530 170.850 ;
        RECT 96.570 170.590 96.830 170.850 ;
        RECT 105.310 170.930 105.570 171.190 ;
        RECT 102.090 170.590 102.350 170.850 ;
        RECT 103.930 170.590 104.190 170.850 ;
        RECT 89.210 169.910 89.470 170.170 ;
        RECT 98.410 170.250 98.670 170.510 ;
        RECT 99.330 170.250 99.590 170.510 ;
        RECT 108.530 170.250 108.790 170.510 ;
        RECT 93.810 169.910 94.070 170.170 ;
        RECT 110.830 170.250 111.090 170.510 ;
        RECT 81.390 169.570 81.650 169.830 ;
        RECT 88.750 169.570 89.010 169.830 ;
        RECT 91.970 169.570 92.230 169.830 ;
        RECT 114.050 170.590 114.310 170.850 ;
        RECT 121.870 170.930 122.130 171.190 ;
        RECT 126.010 170.930 126.270 171.190 ;
        RECT 155.910 171.270 156.170 171.530 ;
        RECT 116.810 170.590 117.070 170.850 ;
        RECT 117.730 170.590 117.990 170.850 ;
        RECT 119.570 170.590 119.830 170.850 ;
        RECT 120.030 170.590 120.290 170.850 ;
        RECT 121.410 170.590 121.670 170.850 ;
        RECT 122.790 170.590 123.050 170.850 ;
        RECT 113.590 170.250 113.850 170.510 ;
        RECT 135.670 170.590 135.930 170.850 ;
        RECT 140.270 170.590 140.530 170.850 ;
        RECT 144.410 170.590 144.670 170.850 ;
        RECT 146.710 170.590 146.970 170.850 ;
        RECT 137.510 170.250 137.770 170.510 ;
        RECT 141.650 170.250 141.910 170.510 ;
        RECT 143.490 170.250 143.750 170.510 ;
        RECT 151.770 170.590 152.030 170.850 ;
        RECT 103.470 169.570 103.730 169.830 ;
        RECT 107.610 169.570 107.870 169.830 ;
        RECT 116.350 169.570 116.610 169.830 ;
        RECT 117.730 169.570 117.990 169.830 ;
        RECT 118.190 169.570 118.450 169.830 ;
        RECT 120.030 169.570 120.290 169.830 ;
        RECT 121.870 169.570 122.130 169.830 ;
        RECT 129.690 169.910 129.950 170.170 ;
        RECT 148.090 170.250 148.350 170.510 ;
        RECT 153.150 170.590 153.410 170.850 ;
        RECT 130.150 169.570 130.410 169.830 ;
        RECT 145.330 169.570 145.590 169.830 ;
        RECT 153.610 169.570 153.870 169.830 ;
        RECT 74.780 169.060 75.040 169.320 ;
        RECT 75.100 169.060 75.360 169.320 ;
        RECT 75.420 169.060 75.680 169.320 ;
        RECT 75.740 169.060 76.000 169.320 ;
        RECT 76.060 169.060 76.320 169.320 ;
        RECT 76.380 169.060 76.640 169.320 ;
        RECT 104.780 169.060 105.040 169.320 ;
        RECT 105.100 169.060 105.360 169.320 ;
        RECT 105.420 169.060 105.680 169.320 ;
        RECT 105.740 169.060 106.000 169.320 ;
        RECT 106.060 169.060 106.320 169.320 ;
        RECT 106.380 169.060 106.640 169.320 ;
        RECT 134.780 169.060 135.040 169.320 ;
        RECT 135.100 169.060 135.360 169.320 ;
        RECT 135.420 169.060 135.680 169.320 ;
        RECT 135.740 169.060 136.000 169.320 ;
        RECT 136.060 169.060 136.320 169.320 ;
        RECT 136.380 169.060 136.640 169.320 ;
        RECT 88.750 168.550 89.010 168.810 ;
        RECT 94.270 168.550 94.530 168.810 ;
        RECT 97.030 168.550 97.290 168.810 ;
        RECT 116.810 168.550 117.070 168.810 ;
        RECT 126.010 168.550 126.270 168.810 ;
        RECT 129.690 168.550 129.950 168.810 ;
        RECT 87.370 168.210 87.630 168.470 ;
        RECT 96.570 168.210 96.830 168.470 ;
        RECT 101.170 168.210 101.430 168.470 ;
        RECT 102.090 168.210 102.350 168.470 ;
        RECT 103.930 168.210 104.190 168.470 ;
        RECT 113.590 168.210 113.850 168.470 ;
        RECT 119.110 168.210 119.370 168.470 ;
        RECT 120.030 168.210 120.290 168.470 ;
        RECT 137.510 168.550 137.770 168.810 ;
        RECT 77.710 167.870 77.970 168.130 ;
        RECT 79.090 167.870 79.350 168.130 ;
        RECT 85.530 167.870 85.790 168.130 ;
        RECT 93.810 167.870 94.070 168.130 ;
        RECT 114.510 167.870 114.770 168.130 ;
        RECT 117.730 167.870 117.990 168.130 ;
        RECT 139.350 168.210 139.610 168.470 ;
        RECT 153.150 168.210 153.410 168.470 ;
        RECT 72.190 167.530 72.450 167.790 ;
        RECT 77.250 167.190 77.510 167.450 ;
        RECT 86.910 167.530 87.170 167.790 ;
        RECT 88.290 167.530 88.550 167.790 ;
        RECT 88.750 167.530 89.010 167.790 ;
        RECT 90.590 167.530 90.850 167.790 ;
        RECT 87.370 167.190 87.630 167.450 ;
        RECT 91.050 167.190 91.310 167.450 ;
        RECT 94.270 167.530 94.530 167.790 ;
        RECT 98.870 167.530 99.130 167.790 ;
        RECT 99.790 167.530 100.050 167.790 ;
        RECT 100.250 167.530 100.510 167.790 ;
        RECT 101.170 167.530 101.430 167.790 ;
        RECT 113.130 167.530 113.390 167.790 ;
        RECT 116.810 167.530 117.070 167.790 ;
        RECT 118.650 167.530 118.910 167.790 ;
        RECT 119.570 167.530 119.830 167.790 ;
        RECT 123.250 167.530 123.510 167.790 ;
        RECT 126.470 167.530 126.730 167.790 ;
        RECT 129.230 167.530 129.490 167.790 ;
        RECT 134.290 167.870 134.550 168.130 ;
        RECT 101.630 167.190 101.890 167.450 ;
        RECT 92.430 166.850 92.690 167.110 ;
        RECT 98.870 166.850 99.130 167.110 ;
        RECT 99.330 166.850 99.590 167.110 ;
        RECT 101.170 166.850 101.430 167.110 ;
        RECT 102.550 166.850 102.810 167.110 ;
        RECT 104.390 166.850 104.650 167.110 ;
        RECT 114.510 166.850 114.770 167.110 ;
        RECT 119.110 166.850 119.370 167.110 ;
        RECT 131.990 167.530 132.250 167.790 ;
        RECT 154.990 167.870 155.250 168.130 ;
        RECT 139.350 167.530 139.610 167.790 ;
        RECT 139.810 167.530 140.070 167.790 ;
        RECT 140.270 167.530 140.530 167.790 ;
        RECT 142.570 167.530 142.830 167.790 ;
        RECT 149.010 167.530 149.270 167.790 ;
        RECT 123.250 166.850 123.510 167.110 ;
        RECT 123.710 166.850 123.970 167.110 ;
        RECT 129.690 166.850 129.950 167.110 ;
        RECT 130.150 166.850 130.410 167.110 ;
        RECT 131.070 167.190 131.330 167.450 ;
        RECT 131.990 166.850 132.250 167.110 ;
        RECT 137.970 166.850 138.230 167.110 ;
        RECT 139.810 166.850 140.070 167.110 ;
        RECT 140.730 166.850 140.990 167.110 ;
        RECT 152.230 166.850 152.490 167.110 ;
        RECT 89.780 166.340 90.040 166.600 ;
        RECT 90.100 166.340 90.360 166.600 ;
        RECT 90.420 166.340 90.680 166.600 ;
        RECT 90.740 166.340 91.000 166.600 ;
        RECT 91.060 166.340 91.320 166.600 ;
        RECT 91.380 166.340 91.640 166.600 ;
        RECT 119.780 166.340 120.040 166.600 ;
        RECT 120.100 166.340 120.360 166.600 ;
        RECT 120.420 166.340 120.680 166.600 ;
        RECT 120.740 166.340 121.000 166.600 ;
        RECT 121.060 166.340 121.320 166.600 ;
        RECT 121.380 166.340 121.640 166.600 ;
        RECT 149.780 166.340 150.040 166.600 ;
        RECT 150.100 166.340 150.360 166.600 ;
        RECT 150.420 166.340 150.680 166.600 ;
        RECT 150.740 166.340 151.000 166.600 ;
        RECT 151.060 166.340 151.320 166.600 ;
        RECT 151.380 166.340 151.640 166.600 ;
        RECT 88.750 165.830 89.010 166.090 ;
        RECT 92.430 165.830 92.690 166.090 ;
        RECT 98.870 165.830 99.130 166.090 ;
        RECT 100.250 165.830 100.510 166.090 ;
        RECT 117.730 165.830 117.990 166.090 ;
        RECT 118.650 165.830 118.910 166.090 ;
        RECT 72.190 165.150 72.450 165.410 ;
        RECT 80.930 165.150 81.190 165.410 ;
        RECT 86.910 165.150 87.170 165.410 ;
        RECT 95.650 165.150 95.910 165.410 ;
        RECT 104.390 165.490 104.650 165.750 ;
        RECT 112.670 165.490 112.930 165.750 ;
        RECT 113.590 165.490 113.850 165.750 ;
        RECT 123.250 165.830 123.510 166.090 ;
        RECT 137.050 165.830 137.310 166.090 ;
        RECT 91.970 164.810 92.230 165.070 ;
        RECT 93.810 164.810 94.070 165.070 ;
        RECT 99.790 165.150 100.050 165.410 ;
        RECT 101.630 165.150 101.890 165.410 ;
        RECT 102.090 165.150 102.350 165.410 ;
        RECT 102.550 165.150 102.810 165.410 ;
        RECT 99.330 164.470 99.590 164.730 ;
        RECT 101.170 164.810 101.430 165.070 ;
        RECT 104.390 164.810 104.650 165.070 ;
        RECT 98.410 164.130 98.670 164.390 ;
        RECT 100.250 164.130 100.510 164.390 ;
        RECT 103.470 164.470 103.730 164.730 ;
        RECT 107.150 165.150 107.410 165.410 ;
        RECT 114.510 165.150 114.770 165.410 ;
        RECT 110.370 164.470 110.630 164.730 ;
        RECT 116.810 164.810 117.070 165.070 ;
        RECT 118.190 165.150 118.450 165.410 ;
        RECT 120.030 165.150 120.290 165.410 ;
        RECT 120.490 165.150 120.750 165.410 ;
        RECT 121.870 165.150 122.130 165.410 ;
        RECT 124.630 165.490 124.890 165.750 ;
        RECT 126.470 165.490 126.730 165.750 ;
        RECT 128.310 165.150 128.570 165.410 ;
        RECT 130.150 165.490 130.410 165.750 ;
        RECT 131.530 165.150 131.790 165.410 ;
        RECT 131.990 165.270 132.250 165.530 ;
        RECT 133.830 165.490 134.090 165.750 ;
        RECT 137.510 165.490 137.770 165.750 ;
        RECT 137.050 165.150 137.310 165.410 ;
        RECT 139.350 165.830 139.610 166.090 ;
        RECT 151.770 165.830 152.030 166.090 ;
        RECT 153.150 165.830 153.410 166.090 ;
        RECT 140.730 165.150 140.990 165.410 ;
        RECT 131.990 164.810 132.250 165.070 ;
        RECT 129.230 164.470 129.490 164.730 ;
        RECT 116.350 164.130 116.610 164.390 ;
        RECT 131.070 164.130 131.330 164.390 ;
        RECT 140.270 164.470 140.530 164.730 ;
        RECT 146.710 165.150 146.970 165.410 ;
        RECT 152.230 165.150 152.490 165.410 ;
        RECT 148.090 164.810 148.350 165.070 ;
        RECT 153.610 164.810 153.870 165.070 ;
        RECT 143.950 164.130 144.210 164.390 ;
        RECT 153.610 164.130 153.870 164.390 ;
        RECT 154.990 164.130 155.250 164.390 ;
        RECT 74.780 163.620 75.040 163.880 ;
        RECT 75.100 163.620 75.360 163.880 ;
        RECT 75.420 163.620 75.680 163.880 ;
        RECT 75.740 163.620 76.000 163.880 ;
        RECT 76.060 163.620 76.320 163.880 ;
        RECT 76.380 163.620 76.640 163.880 ;
        RECT 104.780 163.620 105.040 163.880 ;
        RECT 105.100 163.620 105.360 163.880 ;
        RECT 105.420 163.620 105.680 163.880 ;
        RECT 105.740 163.620 106.000 163.880 ;
        RECT 106.060 163.620 106.320 163.880 ;
        RECT 106.380 163.620 106.640 163.880 ;
        RECT 134.780 163.620 135.040 163.880 ;
        RECT 135.100 163.620 135.360 163.880 ;
        RECT 135.420 163.620 135.680 163.880 ;
        RECT 135.740 163.620 136.000 163.880 ;
        RECT 136.060 163.620 136.320 163.880 ;
        RECT 136.380 163.620 136.640 163.880 ;
        RECT 83.690 163.110 83.950 163.370 ;
        RECT 95.650 163.110 95.910 163.370 ;
        RECT 96.570 163.110 96.830 163.370 ;
        RECT 98.410 163.110 98.670 163.370 ;
        RECT 102.090 163.110 102.350 163.370 ;
        RECT 102.550 163.110 102.810 163.370 ;
        RECT 107.150 163.110 107.410 163.370 ;
        RECT 114.510 163.110 114.770 163.370 ;
        RECT 116.810 163.110 117.070 163.370 ;
        RECT 129.690 163.110 129.950 163.370 ;
        RECT 133.830 163.110 134.090 163.370 ;
        RECT 152.230 163.110 152.490 163.370 ;
        RECT 72.190 162.430 72.450 162.690 ;
        RECT 87.830 162.430 88.090 162.690 ;
        RECT 97.490 162.770 97.750 163.030 ;
        RECT 87.370 162.090 87.630 162.350 ;
        RECT 86.910 161.750 87.170 162.010 ;
        RECT 96.110 162.090 96.370 162.350 ;
        RECT 97.490 162.090 97.750 162.350 ;
        RECT 100.710 161.750 100.970 162.010 ;
        RECT 101.630 162.430 101.890 162.690 ;
        RECT 103.010 162.090 103.270 162.350 ;
        RECT 104.850 162.430 105.110 162.690 ;
        RECT 121.870 162.770 122.130 163.030 ;
        RECT 125.090 162.770 125.350 163.030 ;
        RECT 105.310 162.090 105.570 162.350 ;
        RECT 93.810 161.410 94.070 161.670 ;
        RECT 104.850 161.750 105.110 162.010 ;
        RECT 107.150 162.090 107.410 162.350 ;
        RECT 108.530 162.090 108.790 162.350 ;
        RECT 113.590 162.090 113.850 162.350 ;
        RECT 116.350 162.430 116.610 162.690 ;
        RECT 119.570 162.430 119.830 162.690 ;
        RECT 108.070 161.750 108.330 162.010 ;
        RECT 117.730 162.090 117.990 162.350 ;
        RECT 118.190 162.090 118.450 162.350 ;
        RECT 129.230 162.430 129.490 162.690 ;
        RECT 137.050 162.430 137.310 162.690 ;
        RECT 142.570 162.430 142.830 162.690 ;
        RECT 126.470 162.090 126.730 162.350 ;
        RECT 119.110 161.750 119.370 162.010 ;
        RECT 122.790 161.410 123.050 161.670 ;
        RECT 123.250 161.410 123.510 161.670 ;
        RECT 125.090 161.750 125.350 162.010 ;
        RECT 127.390 161.750 127.650 162.010 ;
        RECT 138.890 162.090 139.150 162.350 ;
        RECT 151.770 161.750 152.030 162.010 ;
        RECT 128.770 161.410 129.030 161.670 ;
        RECT 135.670 161.410 135.930 161.670 ;
        RECT 136.130 161.410 136.390 161.670 ;
        RECT 137.050 161.410 137.310 161.670 ;
        RECT 138.890 161.410 139.150 161.670 ;
        RECT 139.350 161.410 139.610 161.670 ;
        RECT 139.810 161.410 140.070 161.670 ;
        RECT 89.780 160.900 90.040 161.160 ;
        RECT 90.100 160.900 90.360 161.160 ;
        RECT 90.420 160.900 90.680 161.160 ;
        RECT 90.740 160.900 91.000 161.160 ;
        RECT 91.060 160.900 91.320 161.160 ;
        RECT 91.380 160.900 91.640 161.160 ;
        RECT 119.780 160.900 120.040 161.160 ;
        RECT 120.100 160.900 120.360 161.160 ;
        RECT 120.420 160.900 120.680 161.160 ;
        RECT 120.740 160.900 121.000 161.160 ;
        RECT 121.060 160.900 121.320 161.160 ;
        RECT 121.380 160.900 121.640 161.160 ;
        RECT 149.780 160.900 150.040 161.160 ;
        RECT 150.100 160.900 150.360 161.160 ;
        RECT 150.420 160.900 150.680 161.160 ;
        RECT 150.740 160.900 151.000 161.160 ;
        RECT 151.060 160.900 151.320 161.160 ;
        RECT 151.380 160.900 151.640 161.160 ;
        RECT 79.090 160.390 79.350 160.650 ;
        RECT 81.390 160.390 81.650 160.650 ;
        RECT 84.150 160.390 84.410 160.650 ;
        RECT 89.210 160.390 89.470 160.650 ;
        RECT 103.010 160.390 103.270 160.650 ;
        RECT 118.650 160.390 118.910 160.650 ;
        RECT 77.710 159.710 77.970 159.970 ;
        RECT 79.090 159.710 79.350 159.970 ;
        RECT 79.550 159.710 79.810 159.970 ;
        RECT 80.930 159.710 81.190 159.970 ;
        RECT 77.250 159.370 77.510 159.630 ;
        RECT 83.690 159.710 83.950 159.970 ;
        RECT 88.290 159.710 88.550 159.970 ;
        RECT 93.810 160.050 94.070 160.310 ;
        RECT 97.490 160.050 97.750 160.310 ;
        RECT 89.670 159.710 89.930 159.970 ;
        RECT 92.430 159.710 92.690 159.970 ;
        RECT 94.270 159.710 94.530 159.970 ;
        RECT 95.650 159.710 95.910 159.970 ;
        RECT 108.530 160.050 108.790 160.310 ;
        RECT 109.450 160.050 109.710 160.310 ;
        RECT 114.050 160.050 114.310 160.310 ;
        RECT 137.050 160.390 137.310 160.650 ;
        RECT 108.070 159.710 108.330 159.970 ;
        RECT 77.710 159.030 77.970 159.290 ;
        RECT 85.530 159.030 85.790 159.290 ;
        RECT 87.830 159.030 88.090 159.290 ;
        RECT 98.410 159.370 98.670 159.630 ;
        RECT 124.170 159.710 124.430 159.970 ;
        RECT 76.790 158.690 77.050 158.950 ;
        RECT 80.930 158.690 81.190 158.950 ;
        RECT 92.890 158.690 93.150 158.950 ;
        RECT 103.470 159.030 103.730 159.290 ;
        RECT 125.550 159.370 125.810 159.630 ;
        RECT 128.770 159.710 129.030 159.970 ;
        RECT 130.610 159.710 130.870 159.970 ;
        RECT 133.830 159.710 134.090 159.970 ;
        RECT 135.670 159.710 135.930 159.970 ;
        RECT 136.130 159.710 136.390 159.970 ;
        RECT 137.050 159.710 137.310 159.970 ;
        RECT 138.890 159.710 139.150 159.970 ;
        RECT 121.870 159.030 122.130 159.290 ;
        RECT 94.270 158.690 94.530 158.950 ;
        RECT 95.190 158.690 95.450 158.950 ;
        RECT 100.710 158.690 100.970 158.950 ;
        RECT 110.370 158.690 110.630 158.950 ;
        RECT 118.190 158.690 118.450 158.950 ;
        RECT 120.030 158.690 120.290 158.950 ;
        RECT 121.410 158.690 121.670 158.950 ;
        RECT 126.470 159.030 126.730 159.290 ;
        RECT 126.010 158.690 126.270 158.950 ;
        RECT 135.670 159.030 135.930 159.290 ;
        RECT 140.730 159.710 140.990 159.970 ;
        RECT 143.950 160.390 144.210 160.650 ;
        RECT 151.770 160.390 152.030 160.650 ;
        RECT 141.650 159.710 141.910 159.970 ;
        RECT 142.570 159.710 142.830 159.970 ;
        RECT 143.950 159.710 144.210 159.970 ;
        RECT 146.710 160.050 146.970 160.310 ;
        RECT 141.190 159.030 141.450 159.290 ;
        RECT 129.690 158.690 129.950 158.950 ;
        RECT 137.050 158.690 137.310 158.950 ;
        RECT 142.570 158.690 142.830 158.950 ;
        RECT 143.030 158.690 143.290 158.950 ;
        RECT 74.780 158.180 75.040 158.440 ;
        RECT 75.100 158.180 75.360 158.440 ;
        RECT 75.420 158.180 75.680 158.440 ;
        RECT 75.740 158.180 76.000 158.440 ;
        RECT 76.060 158.180 76.320 158.440 ;
        RECT 76.380 158.180 76.640 158.440 ;
        RECT 104.780 158.180 105.040 158.440 ;
        RECT 105.100 158.180 105.360 158.440 ;
        RECT 105.420 158.180 105.680 158.440 ;
        RECT 105.740 158.180 106.000 158.440 ;
        RECT 106.060 158.180 106.320 158.440 ;
        RECT 106.380 158.180 106.640 158.440 ;
        RECT 134.780 158.180 135.040 158.440 ;
        RECT 135.100 158.180 135.360 158.440 ;
        RECT 135.420 158.180 135.680 158.440 ;
        RECT 135.740 158.180 136.000 158.440 ;
        RECT 136.060 158.180 136.320 158.440 ;
        RECT 136.380 158.180 136.640 158.440 ;
        RECT 77.250 157.670 77.510 157.930 ;
        RECT 77.710 157.670 77.970 157.930 ;
        RECT 80.930 157.670 81.190 157.930 ;
        RECT 89.210 157.670 89.470 157.930 ;
        RECT 88.750 157.330 89.010 157.590 ;
        RECT 92.890 157.670 93.150 157.930 ;
        RECT 95.190 157.670 95.450 157.930 ;
        RECT 97.030 157.670 97.290 157.930 ;
        RECT 97.490 157.670 97.750 157.930 ;
        RECT 100.250 157.670 100.510 157.930 ;
        RECT 115.430 157.670 115.690 157.930 ;
        RECT 116.350 157.670 116.610 157.930 ;
        RECT 94.270 157.330 94.530 157.590 ;
        RECT 107.610 157.330 107.870 157.590 ;
        RECT 93.810 156.990 94.070 157.250 ;
        RECT 79.550 156.650 79.810 156.910 ;
        RECT 76.790 155.970 77.050 156.230 ;
        RECT 78.170 155.970 78.430 156.230 ;
        RECT 79.090 155.970 79.350 156.230 ;
        RECT 80.470 156.650 80.730 156.910 ;
        RECT 81.390 156.650 81.650 156.910 ;
        RECT 84.150 156.310 84.410 156.570 ;
        RECT 87.830 156.650 88.090 156.910 ;
        RECT 87.370 156.310 87.630 156.570 ;
        RECT 89.670 156.310 89.930 156.570 ;
        RECT 92.430 156.650 92.690 156.910 ;
        RECT 95.650 156.650 95.910 156.910 ;
        RECT 97.950 156.990 98.210 157.250 ;
        RECT 100.710 156.990 100.970 157.250 ;
        RECT 102.090 156.650 102.350 156.910 ;
        RECT 108.530 156.650 108.790 156.910 ;
        RECT 116.810 157.330 117.070 157.590 ;
        RECT 118.650 157.670 118.910 157.930 ;
        RECT 120.030 157.670 120.290 157.930 ;
        RECT 121.410 157.670 121.670 157.930 ;
        RECT 126.010 157.670 126.270 157.930 ;
        RECT 126.470 157.670 126.730 157.930 ;
        RECT 128.770 157.670 129.030 157.930 ;
        RECT 129.690 157.670 129.950 157.930 ;
        RECT 130.150 157.670 130.410 157.930 ;
        RECT 132.450 157.670 132.710 157.930 ;
        RECT 137.050 157.670 137.310 157.930 ;
        RECT 141.650 157.670 141.910 157.930 ;
        RECT 119.570 157.330 119.830 157.590 ;
        RECT 92.430 155.970 92.690 156.230 ;
        RECT 93.810 155.970 94.070 156.230 ;
        RECT 99.790 155.970 100.050 156.230 ;
        RECT 103.470 155.970 103.730 156.230 ;
        RECT 110.830 155.970 111.090 156.230 ;
        RECT 113.590 156.650 113.850 156.910 ;
        RECT 114.050 156.650 114.310 156.910 ;
        RECT 115.430 156.650 115.690 156.910 ;
        RECT 123.250 156.990 123.510 157.250 ;
        RECT 145.790 157.330 146.050 157.590 ;
        RECT 146.710 157.330 146.970 157.590 ;
        RECT 127.850 156.990 128.110 157.250 ;
        RECT 139.810 156.990 140.070 157.250 ;
        RECT 142.570 156.990 142.830 157.250 ;
        RECT 143.030 156.990 143.290 157.250 ;
        RECT 120.490 156.650 120.750 156.910 ;
        RECT 126.010 156.650 126.270 156.910 ;
        RECT 129.690 156.650 129.950 156.910 ;
        RECT 132.450 156.650 132.710 156.910 ;
        RECT 139.350 156.650 139.610 156.910 ;
        RECT 144.870 156.650 145.130 156.910 ;
        RECT 145.790 156.650 146.050 156.910 ;
        RECT 146.250 156.650 146.510 156.910 ;
        RECT 149.010 156.650 149.270 156.910 ;
        RECT 154.070 156.650 154.330 156.910 ;
        RECT 113.130 155.970 113.390 156.230 ;
        RECT 113.590 155.970 113.850 156.230 ;
        RECT 114.510 155.970 114.770 156.230 ;
        RECT 118.650 155.970 118.910 156.230 ;
        RECT 123.250 155.970 123.510 156.230 ;
        RECT 133.830 155.970 134.090 156.230 ;
        RECT 142.570 155.970 142.830 156.230 ;
        RECT 143.030 155.970 143.290 156.230 ;
        RECT 89.780 155.460 90.040 155.720 ;
        RECT 90.100 155.460 90.360 155.720 ;
        RECT 90.420 155.460 90.680 155.720 ;
        RECT 90.740 155.460 91.000 155.720 ;
        RECT 91.060 155.460 91.320 155.720 ;
        RECT 91.380 155.460 91.640 155.720 ;
        RECT 119.780 155.460 120.040 155.720 ;
        RECT 120.100 155.460 120.360 155.720 ;
        RECT 120.420 155.460 120.680 155.720 ;
        RECT 120.740 155.460 121.000 155.720 ;
        RECT 121.060 155.460 121.320 155.720 ;
        RECT 121.380 155.460 121.640 155.720 ;
        RECT 149.780 155.460 150.040 155.720 ;
        RECT 150.100 155.460 150.360 155.720 ;
        RECT 150.420 155.460 150.680 155.720 ;
        RECT 150.740 155.460 151.000 155.720 ;
        RECT 151.060 155.460 151.320 155.720 ;
        RECT 151.380 155.460 151.640 155.720 ;
        RECT 87.370 154.950 87.630 155.210 ;
        RECT 89.670 154.950 89.930 155.210 ;
        RECT 97.950 154.950 98.210 155.210 ;
        RECT 85.530 154.610 85.790 154.870 ;
        RECT 77.250 154.270 77.510 154.530 ;
        RECT 72.190 153.930 72.450 154.190 ;
        RECT 80.470 154.270 80.730 154.530 ;
        RECT 87.370 154.270 87.630 154.530 ;
        RECT 88.750 154.610 89.010 154.870 ;
        RECT 89.670 154.270 89.930 154.530 ;
        RECT 94.270 154.610 94.530 154.870 ;
        RECT 103.010 154.610 103.270 154.870 ;
        RECT 103.930 154.610 104.190 154.870 ;
        RECT 108.530 154.610 108.790 154.870 ;
        RECT 104.390 154.270 104.650 154.530 ;
        RECT 113.130 154.950 113.390 155.210 ;
        RECT 122.790 154.950 123.050 155.210 ;
        RECT 143.950 154.950 144.210 155.210 ;
        RECT 144.870 154.950 145.130 155.210 ;
        RECT 110.830 154.610 111.090 154.870 ;
        RECT 115.430 154.610 115.690 154.870 ;
        RECT 88.290 153.590 88.550 153.850 ;
        RECT 103.010 153.930 103.270 154.190 ;
        RECT 103.470 153.930 103.730 154.190 ;
        RECT 105.310 153.930 105.570 154.190 ;
        RECT 106.690 153.930 106.950 154.190 ;
        RECT 91.970 153.590 92.230 153.850 ;
        RECT 107.610 153.930 107.870 154.190 ;
        RECT 85.990 153.250 86.250 153.510 ;
        RECT 89.210 153.250 89.470 153.510 ;
        RECT 89.670 153.250 89.930 153.510 ;
        RECT 100.710 153.250 100.970 153.510 ;
        RECT 107.610 153.250 107.870 153.510 ;
        RECT 113.590 154.270 113.850 154.530 ;
        RECT 118.190 154.270 118.450 154.530 ;
        RECT 118.650 154.270 118.910 154.530 ;
        RECT 122.790 154.270 123.050 154.530 ;
        RECT 127.390 154.610 127.650 154.870 ;
        RECT 134.290 154.610 134.550 154.870 ;
        RECT 138.430 154.610 138.690 154.870 ;
        RECT 139.810 154.610 140.070 154.870 ;
        RECT 141.190 154.610 141.450 154.870 ;
        RECT 149.010 154.610 149.270 154.870 ;
        RECT 150.390 154.610 150.650 154.870 ;
        RECT 124.630 154.270 124.890 154.530 ;
        RECT 110.830 153.930 111.090 154.190 ;
        RECT 114.050 153.930 114.310 154.190 ;
        RECT 115.430 153.930 115.690 154.190 ;
        RECT 119.570 153.930 119.830 154.190 ;
        RECT 120.030 153.930 120.290 154.190 ;
        RECT 120.490 153.930 120.750 154.190 ;
        RECT 123.250 153.930 123.510 154.190 ;
        RECT 125.090 153.930 125.350 154.190 ;
        RECT 116.810 153.590 117.070 153.850 ;
        RECT 110.370 153.250 110.630 153.510 ;
        RECT 147.630 154.270 147.890 154.530 ;
        RECT 148.550 154.270 148.810 154.530 ;
        RECT 126.470 153.590 126.730 153.850 ;
        RECT 142.570 153.930 142.830 154.190 ;
        RECT 139.810 153.590 140.070 153.850 ;
        RECT 142.110 153.590 142.370 153.850 ;
        RECT 128.770 153.250 129.030 153.510 ;
        RECT 130.610 153.250 130.870 153.510 ;
        RECT 133.370 153.250 133.630 153.510 ;
        RECT 74.780 152.740 75.040 153.000 ;
        RECT 75.100 152.740 75.360 153.000 ;
        RECT 75.420 152.740 75.680 153.000 ;
        RECT 75.740 152.740 76.000 153.000 ;
        RECT 76.060 152.740 76.320 153.000 ;
        RECT 76.380 152.740 76.640 153.000 ;
        RECT 104.780 152.740 105.040 153.000 ;
        RECT 105.100 152.740 105.360 153.000 ;
        RECT 105.420 152.740 105.680 153.000 ;
        RECT 105.740 152.740 106.000 153.000 ;
        RECT 106.060 152.740 106.320 153.000 ;
        RECT 106.380 152.740 106.640 153.000 ;
        RECT 134.780 152.740 135.040 153.000 ;
        RECT 135.100 152.740 135.360 153.000 ;
        RECT 135.420 152.740 135.680 153.000 ;
        RECT 135.740 152.740 136.000 153.000 ;
        RECT 136.060 152.740 136.320 153.000 ;
        RECT 136.380 152.740 136.640 153.000 ;
        RECT 86.450 152.230 86.710 152.490 ;
        RECT 100.250 152.230 100.510 152.490 ;
        RECT 103.010 152.230 103.270 152.490 ;
        RECT 110.830 152.230 111.090 152.490 ;
        RECT 97.030 151.890 97.290 152.150 ;
        RECT 99.330 151.890 99.590 152.150 ;
        RECT 80.930 151.210 81.190 151.470 ;
        RECT 102.090 151.550 102.350 151.810 ;
        RECT 103.470 151.550 103.730 151.810 ;
        RECT 79.090 150.870 79.350 151.130 ;
        RECT 103.930 151.210 104.190 151.470 ;
        RECT 104.850 151.210 105.110 151.470 ;
        RECT 78.170 150.530 78.430 150.790 ;
        RECT 103.010 150.870 103.270 151.130 ;
        RECT 80.470 150.530 80.730 150.790 ;
        RECT 96.570 150.530 96.830 150.790 ;
        RECT 98.870 150.530 99.130 150.790 ;
        RECT 103.930 150.530 104.190 150.790 ;
        RECT 108.530 151.210 108.790 151.470 ;
        RECT 113.590 152.230 113.850 152.490 ;
        RECT 114.970 152.230 115.230 152.490 ;
        RECT 116.810 152.230 117.070 152.490 ;
        RECT 123.250 152.230 123.510 152.490 ;
        RECT 124.170 152.230 124.430 152.490 ;
        RECT 112.670 151.890 112.930 152.150 ;
        RECT 124.630 151.890 124.890 152.150 ;
        RECT 129.230 152.230 129.490 152.490 ;
        RECT 145.790 152.230 146.050 152.490 ;
        RECT 147.170 152.230 147.430 152.490 ;
        RECT 149.010 152.230 149.270 152.490 ;
        RECT 111.290 151.210 111.550 151.470 ;
        RECT 125.090 151.550 125.350 151.810 ;
        RECT 117.730 151.210 117.990 151.470 ;
        RECT 119.570 151.210 119.830 151.470 ;
        RECT 122.790 151.210 123.050 151.470 ;
        RECT 126.930 151.210 127.190 151.470 ;
        RECT 108.070 150.530 108.330 150.790 ;
        RECT 126.470 150.530 126.730 150.790 ;
        RECT 129.230 151.210 129.490 151.470 ;
        RECT 131.990 151.210 132.250 151.470 ;
        RECT 137.050 151.550 137.310 151.810 ;
        RECT 128.770 150.870 129.030 151.130 ;
        RECT 129.230 150.530 129.490 150.790 ;
        RECT 138.890 151.210 139.150 151.470 ;
        RECT 140.730 151.210 140.990 151.470 ;
        RECT 142.110 151.550 142.370 151.810 ;
        RECT 143.950 150.870 144.210 151.130 ;
        RECT 145.790 151.210 146.050 151.470 ;
        RECT 148.550 151.210 148.810 151.470 ;
        RECT 150.850 151.210 151.110 151.470 ;
        RECT 154.070 151.210 154.330 151.470 ;
        RECT 142.110 150.530 142.370 150.790 ;
        RECT 145.790 150.530 146.050 150.790 ;
        RECT 148.550 150.530 148.810 150.790 ;
        RECT 152.230 150.530 152.490 150.790 ;
        RECT 89.780 150.020 90.040 150.280 ;
        RECT 90.100 150.020 90.360 150.280 ;
        RECT 90.420 150.020 90.680 150.280 ;
        RECT 90.740 150.020 91.000 150.280 ;
        RECT 91.060 150.020 91.320 150.280 ;
        RECT 91.380 150.020 91.640 150.280 ;
        RECT 119.780 150.020 120.040 150.280 ;
        RECT 120.100 150.020 120.360 150.280 ;
        RECT 120.420 150.020 120.680 150.280 ;
        RECT 120.740 150.020 121.000 150.280 ;
        RECT 121.060 150.020 121.320 150.280 ;
        RECT 121.380 150.020 121.640 150.280 ;
        RECT 149.780 150.020 150.040 150.280 ;
        RECT 150.100 150.020 150.360 150.280 ;
        RECT 150.420 150.020 150.680 150.280 ;
        RECT 150.740 150.020 151.000 150.280 ;
        RECT 151.060 150.020 151.320 150.280 ;
        RECT 151.380 150.020 151.640 150.280 ;
        RECT 77.250 149.510 77.510 149.770 ;
        RECT 84.610 149.510 84.870 149.770 ;
        RECT 87.830 149.510 88.090 149.770 ;
        RECT 72.190 148.490 72.450 148.750 ;
        RECT 80.010 148.490 80.270 148.750 ;
        RECT 83.230 148.830 83.490 149.090 ;
        RECT 85.990 148.830 86.250 149.090 ;
        RECT 87.830 148.830 88.090 149.090 ;
        RECT 85.530 148.490 85.790 148.750 ;
        RECT 86.450 148.490 86.710 148.750 ;
        RECT 96.110 149.170 96.370 149.430 ;
        RECT 103.470 149.510 103.730 149.770 ;
        RECT 104.390 149.510 104.650 149.770 ;
        RECT 104.850 149.510 105.110 149.770 ;
        RECT 109.910 149.510 110.170 149.770 ;
        RECT 145.790 149.510 146.050 149.770 ;
        RECT 148.090 149.510 148.350 149.770 ;
        RECT 148.550 149.510 148.810 149.770 ;
        RECT 149.010 149.510 149.270 149.770 ;
        RECT 85.990 148.150 86.250 148.410 ;
        RECT 92.430 148.490 92.690 148.750 ;
        RECT 95.650 148.490 95.910 148.750 ;
        RECT 94.270 148.150 94.530 148.410 ;
        RECT 99.790 148.830 100.050 149.090 ;
        RECT 100.710 148.830 100.970 149.090 ;
        RECT 103.010 148.830 103.270 149.090 ;
        RECT 98.870 148.490 99.130 148.750 ;
        RECT 102.090 148.490 102.350 148.750 ;
        RECT 115.890 148.830 116.150 149.090 ;
        RECT 104.390 148.490 104.650 148.750 ;
        RECT 110.830 148.490 111.090 148.750 ;
        RECT 124.630 148.830 124.890 149.090 ;
        RECT 129.230 148.830 129.490 149.090 ;
        RECT 131.990 148.830 132.250 149.090 ;
        RECT 134.290 148.830 134.550 149.090 ;
        RECT 136.130 148.830 136.390 149.090 ;
        RECT 137.050 148.830 137.310 149.090 ;
        RECT 111.290 148.150 111.550 148.410 ;
        RECT 112.670 148.150 112.930 148.410 ;
        RECT 114.970 148.150 115.230 148.410 ;
        RECT 119.110 148.150 119.370 148.410 ;
        RECT 126.930 148.150 127.190 148.410 ;
        RECT 132.450 148.150 132.710 148.410 ;
        RECT 135.670 148.150 135.930 148.410 ;
        RECT 140.730 148.830 140.990 149.090 ;
        RECT 143.950 149.170 144.210 149.430 ;
        RECT 146.710 148.830 146.970 149.090 ;
        RECT 149.930 148.830 150.190 149.090 ;
        RECT 153.610 148.830 153.870 149.090 ;
        RECT 151.770 148.150 152.030 148.410 ;
        RECT 79.090 147.810 79.350 148.070 ;
        RECT 84.150 147.810 84.410 148.070 ;
        RECT 98.870 147.810 99.130 148.070 ;
        RECT 100.250 147.810 100.510 148.070 ;
        RECT 114.050 147.810 114.310 148.070 ;
        RECT 115.430 147.810 115.690 148.070 ;
        RECT 118.190 147.810 118.450 148.070 ;
        RECT 121.870 147.810 122.130 148.070 ;
        RECT 124.170 147.810 124.430 148.070 ;
        RECT 126.470 147.810 126.730 148.070 ;
        RECT 127.850 147.810 128.110 148.070 ;
        RECT 130.610 147.810 130.870 148.070 ;
        RECT 134.290 147.810 134.550 148.070 ;
        RECT 138.430 147.810 138.690 148.070 ;
        RECT 138.890 147.810 139.150 148.070 ;
        RECT 143.950 147.810 144.210 148.070 ;
        RECT 152.690 147.810 152.950 148.070 ;
        RECT 74.780 147.300 75.040 147.560 ;
        RECT 75.100 147.300 75.360 147.560 ;
        RECT 75.420 147.300 75.680 147.560 ;
        RECT 75.740 147.300 76.000 147.560 ;
        RECT 76.060 147.300 76.320 147.560 ;
        RECT 76.380 147.300 76.640 147.560 ;
        RECT 104.780 147.300 105.040 147.560 ;
        RECT 105.100 147.300 105.360 147.560 ;
        RECT 105.420 147.300 105.680 147.560 ;
        RECT 105.740 147.300 106.000 147.560 ;
        RECT 106.060 147.300 106.320 147.560 ;
        RECT 106.380 147.300 106.640 147.560 ;
        RECT 134.780 147.300 135.040 147.560 ;
        RECT 135.100 147.300 135.360 147.560 ;
        RECT 135.420 147.300 135.680 147.560 ;
        RECT 135.740 147.300 136.000 147.560 ;
        RECT 136.060 147.300 136.320 147.560 ;
        RECT 136.380 147.300 136.640 147.560 ;
        RECT 102.090 146.790 102.350 147.050 ;
        RECT 108.530 146.790 108.790 147.050 ;
        RECT 110.830 146.790 111.090 147.050 ;
        RECT 78.170 146.110 78.430 146.370 ;
        RECT 80.010 145.770 80.270 146.030 ;
        RECT 80.930 145.770 81.190 146.030 ;
        RECT 75.410 145.430 75.670 145.690 ;
        RECT 78.630 145.430 78.890 145.690 ;
        RECT 84.610 146.110 84.870 146.370 ;
        RECT 100.710 146.450 100.970 146.710 ;
        RECT 116.810 146.790 117.070 147.050 ;
        RECT 93.810 146.110 94.070 146.370 ;
        RECT 97.030 146.110 97.290 146.370 ;
        RECT 97.950 146.110 98.210 146.370 ;
        RECT 99.330 146.110 99.590 146.370 ;
        RECT 99.790 146.110 100.050 146.370 ;
        RECT 111.750 146.450 112.010 146.710 ;
        RECT 114.970 146.450 115.230 146.710 ;
        RECT 116.350 146.450 116.610 146.710 ;
        RECT 108.070 146.110 108.330 146.370 ;
        RECT 85.990 145.770 86.250 146.030 ;
        RECT 85.530 145.430 85.790 145.690 ;
        RECT 87.370 145.770 87.630 146.030 ;
        RECT 87.830 145.430 88.090 145.690 ;
        RECT 77.250 145.090 77.510 145.350 ;
        RECT 80.930 145.090 81.190 145.350 ;
        RECT 81.390 145.090 81.650 145.350 ;
        RECT 82.770 145.090 83.030 145.350 ;
        RECT 87.370 145.090 87.630 145.350 ;
        RECT 92.430 145.770 92.690 146.030 ;
        RECT 95.650 145.770 95.910 146.030 ;
        RECT 96.570 145.770 96.830 146.030 ;
        RECT 104.850 145.770 105.110 146.030 ;
        RECT 105.770 145.770 106.030 146.030 ;
        RECT 109.910 145.770 110.170 146.030 ;
        RECT 110.370 145.770 110.630 146.030 ;
        RECT 111.290 145.770 111.550 146.030 ;
        RECT 113.130 145.770 113.390 146.030 ;
        RECT 121.870 146.110 122.130 146.370 ;
        RECT 125.550 146.110 125.810 146.370 ;
        RECT 115.890 145.770 116.150 146.030 ;
        RECT 116.810 145.770 117.070 146.030 ;
        RECT 117.270 145.770 117.530 146.030 ;
        RECT 118.190 145.770 118.450 146.030 ;
        RECT 118.650 145.770 118.910 146.030 ;
        RECT 97.950 145.430 98.210 145.690 ;
        RECT 88.750 145.090 89.010 145.350 ;
        RECT 108.530 145.430 108.790 145.690 ;
        RECT 124.170 145.770 124.430 146.030 ;
        RECT 102.550 145.090 102.810 145.350 ;
        RECT 104.390 145.090 104.650 145.350 ;
        RECT 110.370 145.090 110.630 145.350 ;
        RECT 116.350 145.090 116.610 145.350 ;
        RECT 118.190 145.090 118.450 145.350 ;
        RECT 118.650 145.090 118.910 145.350 ;
        RECT 121.870 145.090 122.130 145.350 ;
        RECT 127.390 145.770 127.650 146.030 ;
        RECT 128.770 146.110 129.030 146.370 ;
        RECT 131.990 146.790 132.250 147.050 ;
        RECT 132.450 146.450 132.710 146.710 ;
        RECT 146.710 146.450 146.970 146.710 ;
        RECT 128.770 145.430 129.030 145.690 ;
        RECT 131.070 145.430 131.330 145.690 ;
        RECT 132.450 145.770 132.710 146.030 ;
        RECT 134.750 145.770 135.010 146.030 ;
        RECT 136.590 145.770 136.850 146.030 ;
        RECT 138.430 146.110 138.690 146.370 ;
        RECT 140.730 146.110 140.990 146.370 ;
        RECT 139.350 145.770 139.610 146.030 ;
        RECT 89.780 144.580 90.040 144.840 ;
        RECT 90.100 144.580 90.360 144.840 ;
        RECT 90.420 144.580 90.680 144.840 ;
        RECT 90.740 144.580 91.000 144.840 ;
        RECT 91.060 144.580 91.320 144.840 ;
        RECT 91.380 144.580 91.640 144.840 ;
        RECT 119.780 144.580 120.040 144.840 ;
        RECT 120.100 144.580 120.360 144.840 ;
        RECT 120.420 144.580 120.680 144.840 ;
        RECT 120.740 144.580 121.000 144.840 ;
        RECT 121.060 144.580 121.320 144.840 ;
        RECT 121.380 144.580 121.640 144.840 ;
        RECT 149.780 144.580 150.040 144.840 ;
        RECT 150.100 144.580 150.360 144.840 ;
        RECT 150.420 144.580 150.680 144.840 ;
        RECT 150.740 144.580 151.000 144.840 ;
        RECT 151.060 144.580 151.320 144.840 ;
        RECT 151.380 144.580 151.640 144.840 ;
        RECT 75.410 144.070 75.670 144.330 ;
        RECT 77.250 144.070 77.510 144.330 ;
        RECT 81.390 144.070 81.650 144.330 ;
        RECT 83.230 144.070 83.490 144.330 ;
        RECT 76.790 143.390 77.050 143.650 ;
        RECT 84.610 143.390 84.870 143.650 ;
        RECT 92.430 143.390 92.690 143.650 ;
        RECT 92.890 143.390 93.150 143.650 ;
        RECT 97.030 144.070 97.290 144.330 ;
        RECT 84.150 143.050 84.410 143.310 ;
        RECT 85.530 143.050 85.790 143.310 ;
        RECT 95.190 143.390 95.450 143.650 ;
        RECT 97.950 143.390 98.210 143.650 ;
        RECT 104.390 144.070 104.650 144.330 ;
        RECT 110.370 144.070 110.630 144.330 ;
        RECT 111.290 144.070 111.550 144.330 ;
        RECT 100.710 143.390 100.970 143.650 ;
        RECT 103.930 143.390 104.190 143.650 ;
        RECT 104.390 143.390 104.650 143.650 ;
        RECT 105.770 143.390 106.030 143.650 ;
        RECT 74.030 142.370 74.290 142.630 ;
        RECT 76.330 142.370 76.590 142.630 ;
        RECT 91.510 142.710 91.770 142.970 ;
        RECT 97.030 143.050 97.290 143.310 ;
        RECT 98.410 143.050 98.670 143.310 ;
        RECT 103.010 143.050 103.270 143.310 ;
        RECT 108.070 143.390 108.330 143.650 ;
        RECT 115.430 143.730 115.690 143.990 ;
        RECT 110.370 143.390 110.630 143.650 ;
        RECT 101.170 142.710 101.430 142.970 ;
        RECT 108.530 143.050 108.790 143.310 ;
        RECT 113.130 143.050 113.390 143.310 ;
        RECT 114.970 143.050 115.230 143.310 ;
        RECT 115.890 143.390 116.150 143.650 ;
        RECT 116.350 143.390 116.610 143.650 ;
        RECT 123.250 144.070 123.510 144.330 ;
        RECT 124.630 144.070 124.890 144.330 ;
        RECT 127.390 144.070 127.650 144.330 ;
        RECT 128.310 144.070 128.570 144.330 ;
        RECT 128.770 144.070 129.030 144.330 ;
        RECT 126.470 143.730 126.730 143.990 ;
        RECT 126.930 143.730 127.190 143.990 ;
        RECT 125.550 143.390 125.810 143.650 ;
        RECT 140.270 143.730 140.530 143.990 ;
        RECT 133.830 143.390 134.090 143.650 ;
        RECT 146.250 143.730 146.510 143.990 ;
        RECT 85.530 142.370 85.790 142.630 ;
        RECT 99.330 142.370 99.590 142.630 ;
        RECT 102.550 142.370 102.810 142.630 ;
        RECT 116.350 142.710 116.610 142.970 ;
        RECT 117.270 142.710 117.530 142.970 ;
        RECT 121.870 143.050 122.130 143.310 ;
        RECT 129.230 143.050 129.490 143.310 ;
        RECT 131.530 143.050 131.790 143.310 ;
        RECT 137.510 143.050 137.770 143.310 ;
        RECT 137.970 143.050 138.230 143.310 ;
        RECT 143.490 143.390 143.750 143.650 ;
        RECT 151.770 143.390 152.030 143.650 ;
        RECT 152.230 143.050 152.490 143.310 ;
        RECT 153.150 143.050 153.410 143.310 ;
        RECT 138.890 142.370 139.150 142.630 ;
        RECT 140.270 142.370 140.530 142.630 ;
        RECT 141.190 142.370 141.450 142.630 ;
        RECT 149.010 142.370 149.270 142.630 ;
        RECT 74.780 141.860 75.040 142.120 ;
        RECT 75.100 141.860 75.360 142.120 ;
        RECT 75.420 141.860 75.680 142.120 ;
        RECT 75.740 141.860 76.000 142.120 ;
        RECT 76.060 141.860 76.320 142.120 ;
        RECT 76.380 141.860 76.640 142.120 ;
        RECT 104.780 141.860 105.040 142.120 ;
        RECT 105.100 141.860 105.360 142.120 ;
        RECT 105.420 141.860 105.680 142.120 ;
        RECT 105.740 141.860 106.000 142.120 ;
        RECT 106.060 141.860 106.320 142.120 ;
        RECT 106.380 141.860 106.640 142.120 ;
        RECT 134.780 141.860 135.040 142.120 ;
        RECT 135.100 141.860 135.360 142.120 ;
        RECT 135.420 141.860 135.680 142.120 ;
        RECT 135.740 141.860 136.000 142.120 ;
        RECT 136.060 141.860 136.320 142.120 ;
        RECT 136.380 141.860 136.640 142.120 ;
        RECT 88.750 141.350 89.010 141.610 ;
        RECT 95.190 141.350 95.450 141.610 ;
        RECT 91.510 141.010 91.770 141.270 ;
        RECT 93.810 141.010 94.070 141.270 ;
        RECT 72.190 140.330 72.450 140.590 ;
        RECT 79.550 140.330 79.810 140.590 ;
        RECT 74.030 139.990 74.290 140.250 ;
        RECT 85.530 140.330 85.790 140.590 ;
        RECT 87.370 140.330 87.630 140.590 ;
        RECT 96.110 140.330 96.370 140.590 ;
        RECT 100.710 141.010 100.970 141.270 ;
        RECT 103.930 141.350 104.190 141.610 ;
        RECT 124.170 141.350 124.430 141.610 ;
        RECT 102.090 140.670 102.350 140.930 ;
        RECT 97.950 140.330 98.210 140.590 ;
        RECT 95.650 139.990 95.910 140.250 ;
        RECT 99.330 140.330 99.590 140.590 ;
        RECT 102.550 140.330 102.810 140.590 ;
        RECT 108.070 141.010 108.330 141.270 ;
        RECT 110.370 141.010 110.630 141.270 ;
        RECT 123.250 141.010 123.510 141.270 ;
        RECT 108.530 140.670 108.790 140.930 ;
        RECT 122.790 140.670 123.050 140.930 ;
        RECT 106.690 140.330 106.950 140.590 ;
        RECT 113.130 140.330 113.390 140.590 ;
        RECT 116.810 140.330 117.070 140.590 ;
        RECT 117.270 140.330 117.530 140.590 ;
        RECT 118.190 140.330 118.450 140.590 ;
        RECT 129.230 140.670 129.490 140.930 ;
        RECT 131.990 140.670 132.250 140.930 ;
        RECT 137.970 141.350 138.230 141.610 ;
        RECT 139.810 141.350 140.070 141.610 ;
        RECT 140.730 141.350 140.990 141.610 ;
        RECT 143.490 141.350 143.750 141.610 ;
        RECT 146.250 141.350 146.510 141.610 ;
        RECT 125.550 140.330 125.810 140.590 ;
        RECT 114.050 139.990 114.310 140.250 ;
        RECT 116.350 139.990 116.610 140.250 ;
        RECT 133.830 140.330 134.090 140.590 ;
        RECT 142.110 140.670 142.370 140.930 ;
        RECT 137.050 140.330 137.310 140.590 ;
        RECT 135.210 139.990 135.470 140.250 ;
        RECT 138.430 140.330 138.690 140.590 ;
        RECT 143.950 140.670 144.210 140.930 ;
        RECT 151.770 141.010 152.030 141.270 ;
        RECT 76.790 139.650 77.050 139.910 ;
        RECT 79.550 139.650 79.810 139.910 ;
        RECT 81.390 139.650 81.650 139.910 ;
        RECT 85.070 139.650 85.330 139.910 ;
        RECT 92.430 139.650 92.690 139.910 ;
        RECT 94.730 139.650 94.990 139.910 ;
        RECT 96.570 139.650 96.830 139.910 ;
        RECT 99.790 139.650 100.050 139.910 ;
        RECT 103.930 139.650 104.190 139.910 ;
        RECT 118.190 139.650 118.450 139.910 ;
        RECT 134.750 139.650 135.010 139.910 ;
        RECT 135.670 139.650 135.930 139.910 ;
        RECT 148.550 140.330 148.810 140.590 ;
        RECT 151.770 140.330 152.030 140.590 ;
        RECT 152.690 140.330 152.950 140.590 ;
        RECT 154.530 140.330 154.790 140.590 ;
        RECT 152.230 139.990 152.490 140.250 ;
        RECT 139.350 139.650 139.610 139.910 ;
        RECT 140.730 139.650 140.990 139.910 ;
        RECT 142.110 139.650 142.370 139.910 ;
        RECT 89.780 139.140 90.040 139.400 ;
        RECT 90.100 139.140 90.360 139.400 ;
        RECT 90.420 139.140 90.680 139.400 ;
        RECT 90.740 139.140 91.000 139.400 ;
        RECT 91.060 139.140 91.320 139.400 ;
        RECT 91.380 139.140 91.640 139.400 ;
        RECT 119.780 139.140 120.040 139.400 ;
        RECT 120.100 139.140 120.360 139.400 ;
        RECT 120.420 139.140 120.680 139.400 ;
        RECT 120.740 139.140 121.000 139.400 ;
        RECT 121.060 139.140 121.320 139.400 ;
        RECT 121.380 139.140 121.640 139.400 ;
        RECT 149.780 139.140 150.040 139.400 ;
        RECT 150.100 139.140 150.360 139.400 ;
        RECT 150.420 139.140 150.680 139.400 ;
        RECT 150.740 139.140 151.000 139.400 ;
        RECT 151.060 139.140 151.320 139.400 ;
        RECT 151.380 139.140 151.640 139.400 ;
        RECT 79.550 138.630 79.810 138.890 ;
        RECT 82.310 138.630 82.570 138.890 ;
        RECT 95.190 138.630 95.450 138.890 ;
        RECT 97.950 138.630 98.210 138.890 ;
        RECT 108.530 138.630 108.790 138.890 ;
        RECT 78.630 137.950 78.890 138.210 ;
        RECT 80.010 137.950 80.270 138.210 ;
        RECT 81.390 138.290 81.650 138.550 ;
        RECT 83.690 137.950 83.950 138.210 ;
        RECT 92.890 138.290 93.150 138.550 ;
        RECT 94.270 138.290 94.530 138.550 ;
        RECT 97.490 138.290 97.750 138.550 ;
        RECT 88.750 137.950 89.010 138.210 ;
        RECT 81.850 137.610 82.110 137.870 ;
        RECT 87.370 137.610 87.630 137.870 ;
        RECT 98.410 137.610 98.670 137.870 ;
        RECT 82.310 137.270 82.570 137.530 ;
        RECT 100.710 137.950 100.970 138.210 ;
        RECT 103.470 137.950 103.730 138.210 ;
        RECT 109.910 138.290 110.170 138.550 ;
        RECT 113.590 138.630 113.850 138.890 ;
        RECT 116.810 138.630 117.070 138.890 ;
        RECT 117.270 138.630 117.530 138.890 ;
        RECT 118.190 138.630 118.450 138.890 ;
        RECT 120.030 138.630 120.290 138.890 ;
        RECT 124.170 138.630 124.430 138.890 ;
        RECT 126.010 138.630 126.270 138.890 ;
        RECT 130.150 138.630 130.410 138.890 ;
        RECT 134.290 138.630 134.550 138.890 ;
        RECT 135.210 138.630 135.470 138.890 ;
        RECT 137.050 138.630 137.310 138.890 ;
        RECT 137.510 138.630 137.770 138.890 ;
        RECT 138.890 138.630 139.150 138.890 ;
        RECT 143.030 138.630 143.290 138.890 ;
        RECT 114.050 138.290 114.310 138.550 ;
        RECT 117.270 137.950 117.530 138.210 ;
        RECT 118.190 137.950 118.450 138.210 ;
        RECT 119.110 137.950 119.370 138.210 ;
        RECT 122.790 137.950 123.050 138.210 ;
        RECT 103.470 137.270 103.730 137.530 ;
        RECT 120.030 137.610 120.290 137.870 ;
        RECT 77.250 136.930 77.510 137.190 ;
        RECT 80.010 136.930 80.270 137.190 ;
        RECT 97.950 136.930 98.210 137.190 ;
        RECT 102.090 136.930 102.350 137.190 ;
        RECT 107.150 136.930 107.410 137.190 ;
        RECT 112.670 137.270 112.930 137.530 ;
        RECT 127.390 137.610 127.650 137.870 ;
        RECT 128.770 137.950 129.030 138.210 ;
        RECT 132.450 137.610 132.710 137.870 ;
        RECT 125.550 137.270 125.810 137.530 ;
        RECT 126.930 137.270 127.190 137.530 ;
        RECT 135.670 137.610 135.930 137.870 ;
        RECT 137.970 137.950 138.230 138.210 ;
        RECT 140.270 137.950 140.530 138.210 ;
        RECT 141.650 137.950 141.910 138.210 ;
        RECT 138.890 137.610 139.150 137.870 ;
        RECT 141.190 137.610 141.450 137.870 ;
        RECT 143.030 137.610 143.290 137.870 ;
        RECT 144.870 137.610 145.130 137.870 ;
        RECT 149.010 137.610 149.270 137.870 ;
        RECT 152.230 137.950 152.490 138.210 ;
        RECT 153.150 137.610 153.410 137.870 ;
        RECT 140.730 137.270 140.990 137.530 ;
        RECT 120.030 136.930 120.290 137.190 ;
        RECT 123.250 136.930 123.510 137.190 ;
        RECT 129.230 136.930 129.490 137.190 ;
        RECT 137.510 136.930 137.770 137.190 ;
        RECT 137.970 136.930 138.230 137.190 ;
        RECT 141.190 136.930 141.450 137.190 ;
        RECT 151.770 136.930 152.030 137.190 ;
        RECT 74.780 136.420 75.040 136.680 ;
        RECT 75.100 136.420 75.360 136.680 ;
        RECT 75.420 136.420 75.680 136.680 ;
        RECT 75.740 136.420 76.000 136.680 ;
        RECT 76.060 136.420 76.320 136.680 ;
        RECT 76.380 136.420 76.640 136.680 ;
        RECT 104.780 136.420 105.040 136.680 ;
        RECT 105.100 136.420 105.360 136.680 ;
        RECT 105.420 136.420 105.680 136.680 ;
        RECT 105.740 136.420 106.000 136.680 ;
        RECT 106.060 136.420 106.320 136.680 ;
        RECT 106.380 136.420 106.640 136.680 ;
        RECT 134.780 136.420 135.040 136.680 ;
        RECT 135.100 136.420 135.360 136.680 ;
        RECT 135.420 136.420 135.680 136.680 ;
        RECT 135.740 136.420 136.000 136.680 ;
        RECT 136.060 136.420 136.320 136.680 ;
        RECT 136.380 136.420 136.640 136.680 ;
        RECT 78.630 135.910 78.890 136.170 ;
        RECT 79.550 135.910 79.810 136.170 ;
        RECT 80.010 135.910 80.270 136.170 ;
        RECT 91.970 135.910 92.230 136.170 ;
        RECT 89.210 135.230 89.470 135.490 ;
        RECT 90.130 134.890 90.390 135.150 ;
        RECT 96.570 135.570 96.830 135.830 ;
        RECT 81.850 134.550 82.110 134.810 ;
        RECT 88.290 134.550 88.550 134.810 ;
        RECT 94.270 134.890 94.530 135.150 ;
        RECT 96.570 134.890 96.830 135.150 ;
        RECT 97.490 134.890 97.750 135.150 ;
        RECT 97.950 134.890 98.210 135.150 ;
        RECT 99.330 134.890 99.590 135.150 ;
        RECT 99.790 134.890 100.050 135.150 ;
        RECT 102.090 135.910 102.350 136.170 ;
        RECT 103.010 135.910 103.270 136.170 ;
        RECT 104.390 135.910 104.650 136.170 ;
        RECT 107.150 135.910 107.410 136.170 ;
        RECT 113.130 135.910 113.390 136.170 ;
        RECT 114.050 135.910 114.310 136.170 ;
        RECT 100.710 135.570 100.970 135.830 ;
        RECT 78.170 134.210 78.430 134.470 ;
        RECT 86.910 134.210 87.170 134.470 ;
        RECT 89.210 134.210 89.470 134.470 ;
        RECT 91.970 134.210 92.230 134.470 ;
        RECT 98.870 134.210 99.130 134.470 ;
        RECT 103.470 134.890 103.730 135.150 ;
        RECT 103.010 134.210 103.270 134.470 ;
        RECT 104.390 134.890 104.650 135.150 ;
        RECT 107.150 134.890 107.410 135.150 ;
        RECT 108.070 134.890 108.330 135.150 ;
        RECT 116.810 135.230 117.070 135.490 ;
        RECT 118.190 135.910 118.450 136.170 ;
        RECT 126.930 135.910 127.190 136.170 ;
        RECT 140.730 135.910 140.990 136.170 ;
        RECT 148.550 135.910 148.810 136.170 ;
        RECT 149.010 135.910 149.270 136.170 ;
        RECT 132.450 135.570 132.710 135.830 ;
        RECT 136.590 135.570 136.850 135.830 ;
        RECT 137.510 135.570 137.770 135.830 ;
        RECT 123.250 134.890 123.510 135.150 ;
        RECT 126.930 134.890 127.190 135.150 ;
        RECT 128.310 134.890 128.570 135.150 ;
        RECT 130.610 135.230 130.870 135.490 ;
        RECT 132.910 135.230 133.170 135.490 ;
        RECT 137.050 135.230 137.310 135.490 ;
        RECT 143.030 135.570 143.290 135.830 ;
        RECT 134.750 134.890 135.010 135.150 ;
        RECT 152.230 135.230 152.490 135.490 ;
        RECT 141.650 134.890 141.910 135.150 ;
        RECT 144.410 134.890 144.670 135.150 ;
        RECT 148.550 134.890 148.810 135.150 ;
        RECT 153.610 134.890 153.870 135.150 ;
        RECT 108.070 134.210 108.330 134.470 ;
        RECT 108.530 134.210 108.790 134.470 ;
        RECT 114.970 134.210 115.230 134.470 ;
        RECT 133.830 134.210 134.090 134.470 ;
        RECT 134.750 134.210 135.010 134.470 ;
        RECT 138.890 134.210 139.150 134.470 ;
        RECT 139.350 134.210 139.610 134.470 ;
        RECT 152.690 134.550 152.950 134.810 ;
        RECT 154.070 134.550 154.330 134.810 ;
        RECT 142.570 134.210 142.830 134.470 ;
        RECT 143.490 134.210 143.750 134.470 ;
        RECT 145.790 134.210 146.050 134.470 ;
        RECT 151.770 134.210 152.030 134.470 ;
        RECT 154.530 134.210 154.790 134.470 ;
        RECT 89.780 133.700 90.040 133.960 ;
        RECT 90.100 133.700 90.360 133.960 ;
        RECT 90.420 133.700 90.680 133.960 ;
        RECT 90.740 133.700 91.000 133.960 ;
        RECT 91.060 133.700 91.320 133.960 ;
        RECT 91.380 133.700 91.640 133.960 ;
        RECT 119.780 133.700 120.040 133.960 ;
        RECT 120.100 133.700 120.360 133.960 ;
        RECT 120.420 133.700 120.680 133.960 ;
        RECT 120.740 133.700 121.000 133.960 ;
        RECT 121.060 133.700 121.320 133.960 ;
        RECT 121.380 133.700 121.640 133.960 ;
        RECT 149.780 133.700 150.040 133.960 ;
        RECT 150.100 133.700 150.360 133.960 ;
        RECT 150.420 133.700 150.680 133.960 ;
        RECT 150.740 133.700 151.000 133.960 ;
        RECT 151.060 133.700 151.320 133.960 ;
        RECT 151.380 133.700 151.640 133.960 ;
        RECT 85.070 133.190 85.330 133.450 ;
        RECT 90.130 133.190 90.390 133.450 ;
        RECT 97.030 133.190 97.290 133.450 ;
        RECT 85.990 132.850 86.250 133.110 ;
        RECT 111.290 133.190 111.550 133.450 ;
        RECT 124.170 133.190 124.430 133.450 ;
        RECT 141.650 133.190 141.910 133.450 ;
        RECT 103.470 132.850 103.730 133.110 ;
        RECT 106.230 132.850 106.490 133.110 ;
        RECT 108.990 132.850 109.250 133.110 ;
        RECT 109.450 132.850 109.710 133.110 ;
        RECT 76.790 132.510 77.050 132.770 ;
        RECT 82.770 132.510 83.030 132.770 ;
        RECT 86.450 132.510 86.710 132.770 ;
        RECT 86.910 132.510 87.170 132.770 ;
        RECT 89.210 132.510 89.470 132.770 ;
        RECT 97.950 132.510 98.210 132.770 ;
        RECT 98.870 132.510 99.130 132.770 ;
        RECT 104.390 132.510 104.650 132.770 ;
        RECT 85.530 132.170 85.790 132.430 ;
        RECT 102.090 132.170 102.350 132.430 ;
        RECT 113.130 132.510 113.390 132.770 ;
        RECT 114.510 132.510 114.770 132.770 ;
        RECT 120.950 132.510 121.210 132.770 ;
        RECT 124.170 132.510 124.430 132.770 ;
        RECT 129.690 132.850 129.950 133.110 ;
        RECT 76.790 131.830 77.050 132.090 ;
        RECT 84.150 131.830 84.410 132.090 ;
        RECT 89.670 131.830 89.930 132.090 ;
        RECT 96.570 131.830 96.830 132.090 ;
        RECT 84.610 131.490 84.870 131.750 ;
        RECT 88.290 131.490 88.550 131.750 ;
        RECT 95.650 131.490 95.910 131.750 ;
        RECT 103.010 131.830 103.270 132.090 ;
        RECT 108.070 131.830 108.330 132.090 ;
        RECT 123.250 132.170 123.510 132.430 ;
        RECT 104.390 131.490 104.650 131.750 ;
        RECT 112.210 131.490 112.470 131.750 ;
        RECT 113.130 131.830 113.390 132.090 ;
        RECT 120.950 131.830 121.210 132.090 ;
        RECT 130.610 132.510 130.870 132.770 ;
        RECT 131.530 132.850 131.790 133.110 ;
        RECT 137.970 132.850 138.230 133.110 ;
        RECT 128.310 131.830 128.570 132.090 ;
        RECT 116.810 131.490 117.070 131.750 ;
        RECT 130.150 131.830 130.410 132.090 ;
        RECT 139.350 132.510 139.610 132.770 ;
        RECT 140.730 132.510 140.990 132.770 ;
        RECT 143.030 132.850 143.290 133.110 ;
        RECT 143.950 132.850 144.210 133.110 ;
        RECT 149.010 133.190 149.270 133.450 ;
        RECT 153.610 133.190 153.870 133.450 ;
        RECT 142.570 132.510 142.830 132.770 ;
        RECT 131.990 131.830 132.250 132.090 ;
        RECT 144.870 132.510 145.130 132.770 ;
        RECT 145.790 132.510 146.050 132.770 ;
        RECT 155.450 132.850 155.710 133.110 ;
        RECT 155.910 132.850 156.170 133.110 ;
        RECT 137.970 131.490 138.230 131.750 ;
        RECT 139.350 131.490 139.610 131.750 ;
        RECT 140.730 131.490 140.990 131.750 ;
        RECT 141.650 131.490 141.910 131.750 ;
        RECT 144.410 131.490 144.670 131.750 ;
        RECT 145.790 131.830 146.050 132.090 ;
        RECT 155.450 131.830 155.710 132.090 ;
        RECT 145.330 131.490 145.590 131.750 ;
        RECT 147.170 131.490 147.430 131.750 ;
        RECT 148.090 131.490 148.350 131.750 ;
        RECT 149.930 131.490 150.190 131.750 ;
        RECT 150.390 131.490 150.650 131.750 ;
        RECT 152.230 131.490 152.490 131.750 ;
        RECT 74.780 130.980 75.040 131.240 ;
        RECT 75.100 130.980 75.360 131.240 ;
        RECT 75.420 130.980 75.680 131.240 ;
        RECT 75.740 130.980 76.000 131.240 ;
        RECT 76.060 130.980 76.320 131.240 ;
        RECT 76.380 130.980 76.640 131.240 ;
        RECT 104.780 130.980 105.040 131.240 ;
        RECT 105.100 130.980 105.360 131.240 ;
        RECT 105.420 130.980 105.680 131.240 ;
        RECT 105.740 130.980 106.000 131.240 ;
        RECT 106.060 130.980 106.320 131.240 ;
        RECT 106.380 130.980 106.640 131.240 ;
        RECT 134.780 130.980 135.040 131.240 ;
        RECT 135.100 130.980 135.360 131.240 ;
        RECT 135.420 130.980 135.680 131.240 ;
        RECT 135.740 130.980 136.000 131.240 ;
        RECT 136.060 130.980 136.320 131.240 ;
        RECT 136.380 130.980 136.640 131.240 ;
        RECT 76.790 130.470 77.050 130.730 ;
        RECT 84.610 130.470 84.870 130.730 ;
        RECT 78.170 130.130 78.430 130.390 ;
        RECT 85.530 130.130 85.790 130.390 ;
        RECT 90.590 130.130 90.850 130.390 ;
        RECT 77.250 129.450 77.510 129.710 ;
        RECT 77.710 129.450 77.970 129.710 ;
        RECT 79.550 129.450 79.810 129.710 ;
        RECT 81.390 129.450 81.650 129.710 ;
        RECT 85.530 129.450 85.790 129.710 ;
        RECT 89.210 129.790 89.470 130.050 ;
        RECT 89.670 129.790 89.930 130.050 ;
        RECT 90.130 129.790 90.390 130.050 ;
        RECT 98.410 130.470 98.670 130.730 ;
        RECT 91.510 130.130 91.770 130.390 ;
        RECT 94.730 130.130 94.990 130.390 ;
        RECT 86.910 129.450 87.170 129.710 ;
        RECT 87.370 129.450 87.630 129.710 ;
        RECT 88.290 129.450 88.550 129.710 ;
        RECT 77.250 128.770 77.510 129.030 ;
        RECT 80.010 128.770 80.270 129.030 ;
        RECT 84.150 129.110 84.410 129.370 ;
        RECT 81.850 128.770 82.110 129.030 ;
        RECT 82.770 128.770 83.030 129.030 ;
        RECT 84.610 128.770 84.870 129.030 ;
        RECT 92.890 129.450 93.150 129.710 ;
        RECT 97.490 129.790 97.750 130.050 ;
        RECT 100.250 130.130 100.510 130.390 ;
        RECT 97.950 129.450 98.210 129.710 ;
        RECT 105.770 130.130 106.030 130.390 ;
        RECT 109.450 130.130 109.710 130.390 ;
        RECT 111.290 130.130 111.550 130.390 ;
        RECT 113.590 130.130 113.850 130.390 ;
        RECT 101.630 129.790 101.890 130.050 ;
        RECT 104.390 129.790 104.650 130.050 ;
        RECT 108.990 129.790 109.250 130.050 ;
        RECT 112.670 129.790 112.930 130.050 ;
        RECT 121.410 130.470 121.670 130.730 ;
        RECT 128.310 130.470 128.570 130.730 ;
        RECT 138.890 130.470 139.150 130.730 ;
        RECT 142.110 130.470 142.370 130.730 ;
        RECT 145.330 130.470 145.590 130.730 ;
        RECT 103.010 129.450 103.270 129.710 ;
        RECT 106.230 129.450 106.490 129.710 ;
        RECT 107.150 129.450 107.410 129.710 ;
        RECT 108.070 129.450 108.330 129.710 ;
        RECT 112.210 129.450 112.470 129.710 ;
        RECT 113.130 129.450 113.390 129.710 ;
        RECT 103.930 129.110 104.190 129.370 ;
        RECT 116.350 129.450 116.610 129.710 ;
        RECT 116.810 129.450 117.070 129.710 ;
        RECT 117.270 129.450 117.530 129.710 ;
        RECT 130.150 130.130 130.410 130.390 ;
        RECT 133.370 130.130 133.630 130.390 ;
        RECT 123.250 129.790 123.510 130.050 ;
        RECT 127.850 129.790 128.110 130.050 ;
        RECT 131.070 129.790 131.330 130.050 ;
        RECT 92.430 128.770 92.690 129.030 ;
        RECT 110.370 128.770 110.630 129.030 ;
        RECT 110.830 128.770 111.090 129.030 ;
        RECT 111.290 128.770 111.550 129.030 ;
        RECT 118.190 129.110 118.450 129.370 ;
        RECT 129.690 129.450 129.950 129.710 ;
        RECT 130.150 129.450 130.410 129.710 ;
        RECT 134.750 129.790 135.010 130.050 ;
        RECT 136.130 129.790 136.390 130.050 ;
        RECT 118.650 128.770 118.910 129.030 ;
        RECT 122.330 129.110 122.590 129.370 ;
        RECT 128.770 129.110 129.030 129.370 ;
        RECT 121.410 128.770 121.670 129.030 ;
        RECT 122.790 128.770 123.050 129.030 ;
        RECT 131.070 128.770 131.330 129.030 ;
        RECT 133.830 129.110 134.090 129.370 ;
        RECT 137.510 129.790 137.770 130.050 ;
        RECT 143.490 129.790 143.750 130.050 ;
        RECT 146.250 129.790 146.510 130.050 ;
        RECT 137.050 129.450 137.310 129.710 ;
        RECT 140.730 129.450 140.990 129.710 ;
        RECT 142.570 129.450 142.830 129.710 ;
        RECT 143.030 129.450 143.290 129.710 ;
        RECT 144.870 129.450 145.130 129.710 ;
        RECT 150.390 130.470 150.650 130.730 ;
        RECT 150.850 130.130 151.110 130.390 ;
        RECT 145.790 128.770 146.050 129.030 ;
        RECT 146.250 128.770 146.510 129.030 ;
        RECT 147.630 129.110 147.890 129.370 ;
        RECT 148.090 129.110 148.350 129.370 ;
        RECT 153.150 129.450 153.410 129.710 ;
        RECT 150.390 128.770 150.650 129.030 ;
        RECT 154.530 129.450 154.790 129.710 ;
        RECT 89.780 128.260 90.040 128.520 ;
        RECT 90.100 128.260 90.360 128.520 ;
        RECT 90.420 128.260 90.680 128.520 ;
        RECT 90.740 128.260 91.000 128.520 ;
        RECT 91.060 128.260 91.320 128.520 ;
        RECT 91.380 128.260 91.640 128.520 ;
        RECT 119.780 128.260 120.040 128.520 ;
        RECT 120.100 128.260 120.360 128.520 ;
        RECT 120.420 128.260 120.680 128.520 ;
        RECT 120.740 128.260 121.000 128.520 ;
        RECT 121.060 128.260 121.320 128.520 ;
        RECT 121.380 128.260 121.640 128.520 ;
        RECT 149.780 128.260 150.040 128.520 ;
        RECT 150.100 128.260 150.360 128.520 ;
        RECT 150.420 128.260 150.680 128.520 ;
        RECT 150.740 128.260 151.000 128.520 ;
        RECT 151.060 128.260 151.320 128.520 ;
        RECT 151.380 128.260 151.640 128.520 ;
        RECT 74.030 127.750 74.290 128.010 ;
        RECT 76.790 127.750 77.050 128.010 ;
        RECT 78.170 127.750 78.430 128.010 ;
        RECT 81.390 127.750 81.650 128.010 ;
        RECT 84.610 127.750 84.870 128.010 ;
        RECT 85.530 127.750 85.790 128.010 ;
        RECT 91.970 127.750 92.230 128.010 ;
        RECT 97.030 127.750 97.290 128.010 ;
        RECT 102.550 127.750 102.810 128.010 ;
        RECT 103.010 127.750 103.270 128.010 ;
        RECT 106.230 127.750 106.490 128.010 ;
        RECT 107.150 127.750 107.410 128.010 ;
        RECT 77.710 127.410 77.970 127.670 ;
        RECT 80.470 127.070 80.730 127.330 ;
        RECT 86.910 127.410 87.170 127.670 ;
        RECT 82.770 127.070 83.030 127.330 ;
        RECT 86.450 127.070 86.710 127.330 ;
        RECT 87.830 127.070 88.090 127.330 ;
        RECT 88.290 127.070 88.550 127.330 ;
        RECT 89.210 127.070 89.470 127.330 ;
        RECT 92.430 127.410 92.690 127.670 ;
        RECT 91.970 127.070 92.230 127.330 ;
        RECT 85.070 126.730 85.330 126.990 ;
        RECT 85.990 126.730 86.250 126.990 ;
        RECT 95.650 127.070 95.910 127.330 ;
        RECT 97.490 127.070 97.750 127.330 ;
        RECT 99.790 127.070 100.050 127.330 ;
        RECT 84.150 126.390 84.410 126.650 ;
        RECT 101.170 126.730 101.430 126.990 ;
        RECT 103.470 127.070 103.730 127.330 ;
        RECT 105.770 127.070 106.030 127.330 ;
        RECT 108.530 127.750 108.790 128.010 ;
        RECT 116.810 127.750 117.070 128.010 ;
        RECT 118.190 127.750 118.450 128.010 ;
        RECT 108.070 127.410 108.330 127.670 ;
        RECT 110.370 127.410 110.630 127.670 ;
        RECT 112.670 127.410 112.930 127.670 ;
        RECT 106.690 126.730 106.950 126.990 ;
        RECT 73.570 126.050 73.830 126.310 ;
        RECT 76.790 126.050 77.050 126.310 ;
        RECT 81.850 126.050 82.110 126.310 ;
        RECT 85.990 126.050 86.250 126.310 ;
        RECT 94.730 126.050 94.990 126.310 ;
        RECT 97.030 126.050 97.290 126.310 ;
        RECT 99.790 126.050 100.050 126.310 ;
        RECT 101.170 126.050 101.430 126.310 ;
        RECT 101.630 126.050 101.890 126.310 ;
        RECT 102.090 126.050 102.350 126.310 ;
        RECT 110.370 126.730 110.630 126.990 ;
        RECT 114.050 127.070 114.310 127.330 ;
        RECT 114.510 126.730 114.770 126.990 ;
        RECT 116.810 127.070 117.070 127.330 ;
        RECT 118.190 127.070 118.450 127.330 ;
        RECT 130.150 127.750 130.410 128.010 ;
        RECT 130.610 127.750 130.870 128.010 ;
        RECT 135.210 127.750 135.470 128.010 ;
        RECT 121.410 127.410 121.670 127.670 ;
        RECT 120.490 126.730 120.750 126.990 ;
        RECT 122.790 126.730 123.050 126.990 ;
        RECT 123.250 126.730 123.510 126.990 ;
        RECT 125.090 127.410 125.350 127.670 ;
        RECT 128.310 126.730 128.570 126.990 ;
        RECT 128.770 126.730 129.030 126.990 ;
        RECT 112.210 126.390 112.470 126.650 ;
        RECT 112.670 126.390 112.930 126.650 ;
        RECT 109.910 126.050 110.170 126.310 ;
        RECT 118.190 126.390 118.450 126.650 ;
        RECT 133.830 127.410 134.090 127.670 ;
        RECT 134.290 127.410 134.550 127.670 ;
        RECT 131.530 127.070 131.790 127.330 ;
        RECT 132.450 127.070 132.710 127.330 ;
        RECT 132.910 127.070 133.170 127.330 ;
        RECT 134.750 127.070 135.010 127.330 ;
        RECT 137.510 127.070 137.770 127.330 ;
        RECT 138.430 127.070 138.690 127.330 ;
        RECT 139.810 127.070 140.070 127.330 ;
        RECT 144.410 127.750 144.670 128.010 ;
        RECT 145.330 127.750 145.590 128.010 ;
        RECT 148.090 127.750 148.350 128.010 ;
        RECT 141.650 127.070 141.910 127.330 ;
        RECT 154.070 127.410 154.330 127.670 ;
        RECT 154.990 127.410 155.250 127.670 ;
        RECT 143.490 127.070 143.750 127.330 ;
        RECT 146.710 127.070 146.970 127.330 ;
        RECT 147.630 127.070 147.890 127.330 ;
        RECT 153.150 127.070 153.410 127.330 ;
        RECT 138.430 126.390 138.690 126.650 ;
        RECT 125.550 126.050 125.810 126.310 ;
        RECT 126.010 126.050 126.270 126.310 ;
        RECT 127.390 126.050 127.650 126.310 ;
        RECT 143.950 126.390 144.210 126.650 ;
        RECT 144.870 126.390 145.130 126.650 ;
        RECT 142.570 126.050 142.830 126.310 ;
        RECT 74.780 125.540 75.040 125.800 ;
        RECT 75.100 125.540 75.360 125.800 ;
        RECT 75.420 125.540 75.680 125.800 ;
        RECT 75.740 125.540 76.000 125.800 ;
        RECT 76.060 125.540 76.320 125.800 ;
        RECT 76.380 125.540 76.640 125.800 ;
        RECT 104.780 125.540 105.040 125.800 ;
        RECT 105.100 125.540 105.360 125.800 ;
        RECT 105.420 125.540 105.680 125.800 ;
        RECT 105.740 125.540 106.000 125.800 ;
        RECT 106.060 125.540 106.320 125.800 ;
        RECT 106.380 125.540 106.640 125.800 ;
        RECT 134.780 125.540 135.040 125.800 ;
        RECT 135.100 125.540 135.360 125.800 ;
        RECT 135.420 125.540 135.680 125.800 ;
        RECT 135.740 125.540 136.000 125.800 ;
        RECT 136.060 125.540 136.320 125.800 ;
        RECT 136.380 125.540 136.640 125.800 ;
        RECT 80.470 125.030 80.730 125.290 ;
        RECT 97.030 125.030 97.290 125.290 ;
        RECT 112.210 125.030 112.470 125.290 ;
        RECT 114.510 125.030 114.770 125.290 ;
        RECT 117.730 125.030 117.990 125.290 ;
        RECT 78.170 124.690 78.430 124.950 ;
        RECT 80.010 124.350 80.270 124.610 ;
        RECT 73.570 124.010 73.830 124.270 ;
        RECT 76.790 124.010 77.050 124.270 ;
        RECT 77.250 124.010 77.510 124.270 ;
        RECT 79.550 124.010 79.810 124.270 ;
        RECT 88.750 124.010 89.010 124.270 ;
        RECT 94.270 124.010 94.530 124.270 ;
        RECT 94.730 124.010 94.990 124.270 ;
        RECT 108.530 124.350 108.790 124.610 ;
        RECT 98.410 124.010 98.670 124.270 ;
        RECT 101.170 124.010 101.430 124.270 ;
        RECT 101.630 124.010 101.890 124.270 ;
        RECT 110.370 124.010 110.630 124.270 ;
        RECT 108.530 123.670 108.790 123.930 ;
        RECT 114.970 124.690 115.230 124.950 ;
        RECT 123.710 125.030 123.970 125.290 ;
        RECT 124.170 125.030 124.430 125.290 ;
        RECT 131.990 125.030 132.250 125.290 ;
        RECT 133.830 125.030 134.090 125.290 ;
        RECT 138.890 125.030 139.150 125.290 ;
        RECT 139.350 125.030 139.610 125.290 ;
        RECT 141.190 125.030 141.450 125.290 ;
        RECT 143.030 125.030 143.290 125.290 ;
        RECT 137.970 124.690 138.230 124.950 ;
        RECT 153.150 125.030 153.410 125.290 ;
        RECT 131.530 124.350 131.790 124.610 ;
        RECT 134.750 124.350 135.010 124.610 ;
        RECT 153.610 124.350 153.870 124.610 ;
        RECT 117.270 124.010 117.530 124.270 ;
        RECT 122.790 124.010 123.050 124.270 ;
        RECT 126.930 124.010 127.190 124.270 ;
        RECT 70.810 123.330 71.070 123.590 ;
        RECT 74.490 123.330 74.750 123.590 ;
        RECT 81.850 123.330 82.110 123.590 ;
        RECT 86.450 123.330 86.710 123.590 ;
        RECT 89.210 123.330 89.470 123.590 ;
        RECT 93.810 123.330 94.070 123.590 ;
        RECT 97.490 123.330 97.750 123.590 ;
        RECT 101.170 123.330 101.430 123.590 ;
        RECT 103.930 123.330 104.190 123.590 ;
        RECT 109.910 123.330 110.170 123.590 ;
        RECT 123.250 123.670 123.510 123.930 ;
        RECT 123.710 123.670 123.970 123.930 ;
        RECT 130.150 124.010 130.410 124.270 ;
        RECT 118.650 123.330 118.910 123.590 ;
        RECT 125.090 123.330 125.350 123.590 ;
        RECT 129.690 123.670 129.950 123.930 ;
        RECT 134.290 124.010 134.550 124.270 ;
        RECT 137.510 124.010 137.770 124.270 ;
        RECT 138.430 124.010 138.690 124.270 ;
        RECT 139.810 124.010 140.070 124.270 ;
        RECT 143.490 124.010 143.750 124.270 ;
        RECT 143.950 124.010 144.210 124.270 ;
        RECT 152.230 124.010 152.490 124.270 ;
        RECT 132.450 123.330 132.710 123.590 ;
        RECT 149.010 123.670 149.270 123.930 ;
        RECT 148.550 123.330 148.810 123.590 ;
        RECT 89.780 122.820 90.040 123.080 ;
        RECT 90.100 122.820 90.360 123.080 ;
        RECT 90.420 122.820 90.680 123.080 ;
        RECT 90.740 122.820 91.000 123.080 ;
        RECT 91.060 122.820 91.320 123.080 ;
        RECT 91.380 122.820 91.640 123.080 ;
        RECT 119.780 122.820 120.040 123.080 ;
        RECT 120.100 122.820 120.360 123.080 ;
        RECT 120.420 122.820 120.680 123.080 ;
        RECT 120.740 122.820 121.000 123.080 ;
        RECT 121.060 122.820 121.320 123.080 ;
        RECT 121.380 122.820 121.640 123.080 ;
        RECT 149.780 122.820 150.040 123.080 ;
        RECT 150.100 122.820 150.360 123.080 ;
        RECT 150.420 122.820 150.680 123.080 ;
        RECT 150.740 122.820 151.000 123.080 ;
        RECT 151.060 122.820 151.320 123.080 ;
        RECT 151.380 122.820 151.640 123.080 ;
        RECT 94.270 122.310 94.530 122.570 ;
        RECT 98.410 122.310 98.670 122.570 ;
        RECT 131.990 122.310 132.250 122.570 ;
        RECT 132.450 122.310 132.710 122.570 ;
        RECT 139.810 122.310 140.070 122.570 ;
        RECT 141.650 122.310 141.910 122.570 ;
        RECT 149.010 122.310 149.270 122.570 ;
        RECT 99.790 121.970 100.050 122.230 ;
        RECT 116.350 121.970 116.610 122.230 ;
        RECT 125.090 121.970 125.350 122.230 ;
        RECT 130.610 121.630 130.870 121.890 ;
        RECT 107.150 121.290 107.410 121.550 ;
        RECT 127.850 121.290 128.110 121.550 ;
        RECT 138.430 121.290 138.690 121.550 ;
        RECT 88.750 120.950 89.010 121.210 ;
        RECT 118.190 120.950 118.450 121.210 ;
        RECT 125.550 120.950 125.810 121.210 ;
        RECT 77.600 79.080 78.600 80.080 ;
        RECT 114.600 79.080 115.600 80.080 ;
        RECT 151.600 79.080 152.600 80.080 ;
        RECT 77.600 30.030 78.600 31.030 ;
        RECT 114.600 30.030 115.600 31.030 ;
        RECT 151.600 30.030 152.600 31.030 ;
        RECT 36.020 24.045 36.320 24.345 ;
        RECT 36.020 19.445 36.320 19.745 ;
        RECT 34.320 18.045 34.620 18.345 ;
        RECT 35.370 18.045 35.670 18.345 ;
      LAYER met2 ;
        RECT 121.990 216.885 122.410 216.910 ;
        RECT 121.970 216.515 122.430 216.885 ;
        RECT 118.290 215.390 118.715 215.415 ;
        RECT 113.800 215.275 114.200 215.300 ;
        RECT 113.780 214.925 114.220 215.275 ;
        RECT 118.270 215.015 118.735 215.390 ;
        RECT 110.265 214.660 110.735 214.680 ;
        RECT 107.040 214.140 110.760 214.660 ;
        RECT 74.020 209.455 74.300 211.455 ;
        RECT 78.160 209.455 78.440 211.455 ;
        RECT 82.300 209.455 82.580 211.455 ;
        RECT 86.440 209.455 86.720 211.455 ;
        RECT 90.580 209.455 90.860 211.455 ;
        RECT 94.720 209.455 95.000 211.455 ;
        RECT 98.860 209.455 99.140 211.455 ;
        RECT 103.000 209.455 103.280 211.455 ;
        RECT 107.040 209.740 107.560 214.140 ;
        RECT 110.265 214.120 110.735 214.140 ;
        RECT 113.800 213.900 114.200 214.925 ;
        RECT 118.290 213.915 118.715 215.015 ;
        RECT 111.200 213.500 114.200 213.900 ;
        RECT 111.200 209.800 111.600 213.500 ;
        RECT 115.390 213.490 118.715 213.915 ;
        RECT 121.990 213.910 122.410 216.515 ;
        RECT 126.520 214.605 126.880 214.625 ;
        RECT 135.965 214.615 136.440 214.640 ;
        RECT 119.490 213.490 122.410 213.910 ;
        RECT 123.595 214.195 126.905 214.605 ;
        RECT 127.805 214.575 128.200 214.600 ;
        RECT 127.785 214.230 128.220 214.575 ;
        RECT 131.910 214.570 132.295 214.595 ;
        RECT 131.890 214.235 132.315 214.570 ;
        RECT 107.140 209.455 107.420 209.740 ;
        RECT 111.280 209.455 111.560 209.800 ;
        RECT 115.390 209.790 115.815 213.490 ;
        RECT 119.490 209.790 119.910 213.490 ;
        RECT 115.420 209.455 115.700 209.790 ;
        RECT 119.560 209.455 119.840 209.790 ;
        RECT 123.595 209.695 124.005 214.195 ;
        RECT 126.520 214.175 126.880 214.195 ;
        RECT 127.805 209.705 128.200 214.230 ;
        RECT 131.910 209.710 132.295 214.235 ;
        RECT 135.945 214.190 136.460 214.615 ;
        RECT 144.270 214.605 144.730 214.630 ;
        RECT 140.205 214.575 140.600 214.600 ;
        RECT 140.185 214.230 140.620 214.575 ;
        RECT 135.965 209.765 136.440 214.190 ;
        RECT 123.700 209.455 123.980 209.695 ;
        RECT 127.840 209.455 128.120 209.705 ;
        RECT 131.980 209.455 132.260 209.710 ;
        RECT 136.120 209.455 136.400 209.765 ;
        RECT 140.205 209.705 140.600 214.230 ;
        RECT 144.250 214.195 144.750 214.605 ;
        RECT 148.485 214.590 148.915 214.615 ;
        RECT 152.570 214.605 153.030 214.630 ;
        RECT 148.465 214.210 148.935 214.590 ;
        RECT 140.260 209.455 140.540 209.705 ;
        RECT 144.270 209.670 144.730 214.195 ;
        RECT 148.485 209.685 148.915 214.210 ;
        RECT 152.550 214.195 153.050 214.605 ;
        RECT 152.570 209.770 153.030 214.195 ;
        RECT 144.400 209.455 144.680 209.670 ;
        RECT 148.540 209.455 148.820 209.685 ;
        RECT 152.680 209.455 152.960 209.770 ;
        RECT 74.090 206.920 74.230 209.455 ;
        RECT 74.770 207.085 76.650 207.455 ;
        RECT 78.230 206.920 78.370 209.455 ;
        RECT 82.370 206.920 82.510 209.455 ;
        RECT 82.770 207.620 83.030 207.940 ;
        RECT 74.030 206.600 74.290 206.920 ;
        RECT 78.170 206.600 78.430 206.920 ;
        RECT 82.310 206.600 82.570 206.920 ;
        RECT 82.830 206.240 82.970 207.620 ;
        RECT 86.510 206.920 86.650 209.455 ;
        RECT 90.650 206.920 90.790 209.455 ;
        RECT 94.790 206.920 94.930 209.455 ;
        RECT 98.930 206.920 99.070 209.455 ;
        RECT 103.070 206.920 103.210 209.455 ;
        RECT 104.390 207.960 104.650 208.280 ;
        RECT 103.930 207.620 104.190 207.940 ;
        RECT 86.450 206.600 86.710 206.920 ;
        RECT 90.590 206.600 90.850 206.920 ;
        RECT 94.730 206.600 94.990 206.920 ;
        RECT 98.870 206.600 99.130 206.920 ;
        RECT 103.010 206.600 103.270 206.920 ;
        RECT 101.630 206.260 101.890 206.580 ;
        RECT 82.770 205.920 83.030 206.240 ;
        RECT 83.230 205.920 83.490 206.240 ;
        RECT 81.850 205.580 82.110 205.900 ;
        RECT 76.330 204.900 76.590 205.220 ;
        RECT 76.390 204.200 76.530 204.900 ;
        RECT 76.330 203.880 76.590 204.200 ;
        RECT 81.910 203.520 82.050 205.580 ;
        RECT 83.290 203.520 83.430 205.920 ;
        RECT 89.210 205.580 89.470 205.900 ;
        RECT 92.430 205.580 92.690 205.900 ;
        RECT 89.270 205.220 89.410 205.580 ;
        RECT 86.910 204.900 87.170 205.220 ;
        RECT 89.210 204.900 89.470 205.220 ;
        RECT 86.970 204.200 87.110 204.900 ;
        RECT 89.770 204.365 91.650 204.735 ;
        RECT 86.910 203.880 87.170 204.200 ;
        RECT 92.490 203.715 92.630 205.580 ;
        RECT 100.250 205.240 100.510 205.560 ;
        RECT 100.710 205.240 100.970 205.560 ;
        RECT 95.190 204.900 95.450 205.220 ;
        RECT 99.790 204.900 100.050 205.220 ;
        RECT 81.850 203.200 82.110 203.520 ;
        RECT 82.770 203.200 83.030 203.520 ;
        RECT 83.230 203.200 83.490 203.520 ;
        RECT 84.150 203.200 84.410 203.520 ;
        RECT 92.420 203.345 92.700 203.715 ;
        RECT 72.190 202.860 72.450 203.180 ;
        RECT 72.250 200.460 72.390 202.860 ;
        RECT 81.850 202.180 82.110 202.500 ;
        RECT 74.770 201.645 76.650 202.015 ;
        RECT 81.910 200.800 82.050 202.180 ;
        RECT 81.850 200.480 82.110 200.800 ;
        RECT 72.190 200.140 72.450 200.460 ;
        RECT 72.250 195.020 72.390 200.140 ;
        RECT 75.410 199.800 75.670 200.120 ;
        RECT 75.470 198.760 75.610 199.800 ;
        RECT 80.930 199.460 81.190 199.780 ;
        RECT 75.410 198.440 75.670 198.760 ;
        RECT 78.160 198.585 78.440 198.955 ;
        RECT 80.990 198.760 81.130 199.460 ;
        RECT 78.170 198.440 78.430 198.585 ;
        RECT 80.930 198.440 81.190 198.760 ;
        RECT 78.230 198.080 78.370 198.440 ;
        RECT 81.850 198.100 82.110 198.420 ;
        RECT 78.170 197.760 78.430 198.080 ;
        RECT 81.390 197.080 81.650 197.400 ;
        RECT 74.770 196.205 76.650 196.575 ;
        RECT 81.450 196.040 81.590 197.080 ;
        RECT 81.390 195.720 81.650 196.040 ;
        RECT 72.190 194.700 72.450 195.020 ;
        RECT 72.250 186.860 72.390 194.700 ;
        RECT 74.950 194.360 75.210 194.680 ;
        RECT 81.380 194.505 81.660 194.875 ;
        RECT 75.010 193.320 75.150 194.360 ;
        RECT 78.170 194.020 78.430 194.340 ;
        RECT 74.950 193.000 75.210 193.320 ;
        RECT 78.230 192.640 78.370 194.020 ;
        RECT 81.450 192.640 81.590 194.505 ;
        RECT 78.170 192.320 78.430 192.640 ;
        RECT 80.470 192.320 80.730 192.640 ;
        RECT 81.390 192.320 81.650 192.640 ;
        RECT 76.790 191.980 77.050 192.300 ;
        RECT 74.770 190.765 76.650 191.135 ;
        RECT 74.030 186.880 74.290 187.200 ;
        RECT 72.190 186.540 72.450 186.860 ;
        RECT 72.250 181.420 72.390 186.540 ;
        RECT 74.090 185.160 74.230 186.880 ;
        RECT 74.770 185.325 76.650 185.695 ;
        RECT 76.850 185.160 76.990 191.980 ;
        RECT 77.250 191.300 77.510 191.620 ;
        RECT 77.310 190.260 77.450 191.300 ;
        RECT 77.250 189.940 77.510 190.260 ;
        RECT 74.030 184.840 74.290 185.160 ;
        RECT 76.790 184.840 77.050 185.160 ;
        RECT 76.330 184.560 76.590 184.820 ;
        RECT 77.310 184.560 77.450 189.940 ;
        RECT 80.530 189.920 80.670 192.320 ;
        RECT 80.930 192.040 81.190 192.300 ;
        RECT 81.380 192.040 81.660 192.155 ;
        RECT 80.930 191.980 81.660 192.040 ;
        RECT 80.990 191.900 81.660 191.980 ;
        RECT 80.470 189.600 80.730 189.920 ;
        RECT 78.630 187.560 78.890 187.880 ;
        RECT 76.330 184.500 77.450 184.560 ;
        RECT 76.390 184.420 77.450 184.500 ;
        RECT 76.790 183.820 77.050 184.140 ;
        RECT 77.710 183.820 77.970 184.140 ;
        RECT 73.570 181.440 73.830 181.760 ;
        RECT 72.190 181.100 72.450 181.420 ;
        RECT 72.250 176.660 72.390 181.100 ;
        RECT 73.630 179.720 73.770 181.440 ;
        RECT 74.770 179.885 76.650 180.255 ;
        RECT 76.850 179.720 76.990 183.820 ;
        RECT 73.570 179.400 73.830 179.720 ;
        RECT 76.790 179.400 77.050 179.720 ;
        RECT 77.770 178.020 77.910 183.820 ;
        RECT 78.690 180.740 78.830 187.560 ;
        RECT 80.530 186.180 80.670 189.600 ;
        RECT 80.990 189.580 81.130 191.900 ;
        RECT 81.380 191.785 81.660 191.900 ;
        RECT 80.930 189.260 81.190 189.580 ;
        RECT 80.990 187.540 81.130 189.260 ;
        RECT 80.930 187.220 81.190 187.540 ;
        RECT 79.550 185.860 79.810 186.180 ;
        RECT 80.010 185.860 80.270 186.180 ;
        RECT 80.470 185.860 80.730 186.180 ;
        RECT 79.090 181.100 79.350 181.420 ;
        RECT 78.630 180.420 78.890 180.740 ;
        RECT 78.170 178.380 78.430 178.700 ;
        RECT 77.710 177.700 77.970 178.020 ;
        RECT 76.790 176.680 77.050 177.000 ;
        RECT 72.190 176.340 72.450 176.660 ;
        RECT 74.770 174.445 76.650 174.815 ;
        RECT 76.850 173.260 76.990 176.680 ;
        RECT 77.770 176.320 77.910 177.700 ;
        RECT 77.710 176.000 77.970 176.320 ;
        RECT 76.790 172.940 77.050 173.260 ;
        RECT 75.870 172.260 76.130 172.580 ;
        RECT 75.930 170.880 76.070 172.260 ;
        RECT 75.870 170.560 76.130 170.880 ;
        RECT 72.190 170.220 72.450 170.540 ;
        RECT 72.250 167.820 72.390 170.220 ;
        RECT 74.770 169.005 76.650 169.375 ;
        RECT 77.710 167.840 77.970 168.160 ;
        RECT 72.190 167.500 72.450 167.820 ;
        RECT 72.250 165.440 72.390 167.500 ;
        RECT 77.250 167.160 77.510 167.480 ;
        RECT 72.190 165.120 72.450 165.440 ;
        RECT 72.250 162.720 72.390 165.120 ;
        RECT 77.310 164.955 77.450 167.160 ;
        RECT 77.240 164.585 77.520 164.955 ;
        RECT 74.770 163.565 76.650 163.935 ;
        RECT 72.190 162.400 72.450 162.720 ;
        RECT 72.250 154.220 72.390 162.400 ;
        RECT 77.770 160.000 77.910 167.840 ;
        RECT 77.710 159.680 77.970 160.000 ;
        RECT 77.250 159.340 77.510 159.660 ;
        RECT 76.790 158.660 77.050 158.980 ;
        RECT 74.770 158.125 76.650 158.495 ;
        RECT 76.850 156.680 76.990 158.660 ;
        RECT 77.310 157.960 77.450 159.340 ;
        RECT 77.710 159.000 77.970 159.320 ;
        RECT 77.770 157.960 77.910 159.000 ;
        RECT 77.250 157.640 77.510 157.960 ;
        RECT 77.710 157.640 77.970 157.960 ;
        RECT 76.850 156.540 77.910 156.680 ;
        RECT 76.790 155.940 77.050 156.260 ;
        RECT 72.190 153.900 72.450 154.220 ;
        RECT 72.250 148.780 72.390 153.900 ;
        RECT 74.770 152.685 76.650 153.055 ;
        RECT 72.190 148.460 72.450 148.780 ;
        RECT 72.250 140.620 72.390 148.460 ;
        RECT 74.770 147.245 76.650 147.615 ;
        RECT 75.410 145.400 75.670 145.720 ;
        RECT 75.470 144.360 75.610 145.400 ;
        RECT 76.850 145.120 76.990 155.940 ;
        RECT 77.250 154.240 77.510 154.560 ;
        RECT 77.310 149.800 77.450 154.240 ;
        RECT 77.250 149.480 77.510 149.800 ;
        RECT 76.390 144.980 76.990 145.120 ;
        RECT 77.250 145.060 77.510 145.380 ;
        RECT 75.410 144.040 75.670 144.360 ;
        RECT 76.390 142.660 76.530 144.980 ;
        RECT 77.310 144.360 77.450 145.060 ;
        RECT 77.250 144.040 77.510 144.360 ;
        RECT 76.790 143.360 77.050 143.680 ;
        RECT 74.030 142.340 74.290 142.660 ;
        RECT 76.330 142.340 76.590 142.660 ;
        RECT 72.190 140.300 72.450 140.620 ;
        RECT 74.090 140.280 74.230 142.340 ;
        RECT 74.770 141.805 76.650 142.175 ;
        RECT 74.030 139.960 74.290 140.280 ;
        RECT 76.850 139.940 76.990 143.360 ;
        RECT 76.790 139.620 77.050 139.940 ;
        RECT 74.770 136.365 76.650 136.735 ;
        RECT 74.480 132.880 74.760 132.995 ;
        RECT 74.090 132.740 74.760 132.880 ;
        RECT 76.850 132.800 76.990 139.620 ;
        RECT 77.250 136.900 77.510 137.220 ;
        RECT 74.090 128.040 74.230 132.740 ;
        RECT 74.480 132.625 74.760 132.740 ;
        RECT 76.790 132.480 77.050 132.800 ;
        RECT 76.790 131.800 77.050 132.120 ;
        RECT 74.770 130.925 76.650 131.295 ;
        RECT 76.850 130.760 76.990 131.800 ;
        RECT 76.790 130.440 77.050 130.760 ;
        RECT 77.310 129.740 77.450 136.900 ;
        RECT 77.770 129.740 77.910 156.540 ;
        RECT 78.230 156.260 78.370 178.380 ;
        RECT 78.690 160.080 78.830 180.420 ;
        RECT 79.150 175.890 79.290 181.100 ;
        RECT 79.610 176.400 79.750 185.860 ;
        RECT 80.070 184.140 80.210 185.860 ;
        RECT 80.010 183.820 80.270 184.140 ;
        RECT 80.930 183.480 81.190 183.800 ;
        RECT 81.380 183.625 81.660 183.995 ;
        RECT 80.990 179.380 81.130 183.480 ;
        RECT 81.450 179.720 81.590 183.625 ;
        RECT 81.910 183.460 82.050 198.100 ;
        RECT 82.830 197.480 82.970 203.200 ;
        RECT 83.290 200.880 83.430 203.200 ;
        RECT 84.210 201.140 84.350 203.200 ;
        RECT 89.210 202.860 89.470 203.180 ;
        RECT 89.270 202.500 89.410 202.860 ;
        RECT 89.210 202.180 89.470 202.500 ;
        RECT 91.050 202.180 91.310 202.500 ;
        RECT 94.730 202.180 94.990 202.500 ;
        RECT 83.290 200.740 83.890 200.880 ;
        RECT 84.150 200.820 84.410 201.140 ;
        RECT 83.230 200.140 83.490 200.460 ;
        RECT 83.290 198.420 83.430 200.140 ;
        RECT 83.230 198.100 83.490 198.420 ;
        RECT 82.830 197.340 83.430 197.480 ;
        RECT 82.310 196.740 82.570 197.060 ;
        RECT 82.370 193.320 82.510 196.740 ;
        RECT 82.770 195.720 83.030 196.040 ;
        RECT 82.310 193.000 82.570 193.320 ;
        RECT 82.830 192.640 82.970 195.720 ;
        RECT 83.290 194.930 83.430 197.340 ;
        RECT 83.750 195.700 83.890 200.740 ;
        RECT 84.150 199.690 84.410 199.780 ;
        RECT 84.150 199.550 84.810 199.690 ;
        RECT 84.150 199.460 84.410 199.550 ;
        RECT 84.140 198.585 84.420 198.955 ;
        RECT 84.150 198.440 84.410 198.585 ;
        RECT 83.690 195.380 83.950 195.700 ;
        RECT 83.290 194.790 83.890 194.930 ;
        RECT 82.770 192.320 83.030 192.640 ;
        RECT 82.770 191.300 83.030 191.620 ;
        RECT 82.310 184.840 82.570 185.160 ;
        RECT 82.370 184.675 82.510 184.840 ;
        RECT 82.300 184.305 82.580 184.675 ;
        RECT 82.830 184.050 82.970 191.300 ;
        RECT 82.370 183.910 82.970 184.050 ;
        RECT 81.850 183.140 82.110 183.460 ;
        RECT 81.390 179.400 81.650 179.720 ;
        RECT 80.930 179.060 81.190 179.380 ;
        RECT 80.010 178.380 80.270 178.700 ;
        RECT 80.070 177.000 80.210 178.380 ;
        RECT 80.010 176.680 80.270 177.000 ;
        RECT 79.610 176.260 80.210 176.400 ;
        RECT 79.550 175.890 79.810 175.980 ;
        RECT 79.150 175.750 79.810 175.890 ;
        RECT 79.550 175.660 79.810 175.750 ;
        RECT 79.550 174.980 79.810 175.300 ;
        RECT 79.610 173.260 79.750 174.980 ;
        RECT 79.550 172.940 79.810 173.260 ;
        RECT 79.090 167.840 79.350 168.160 ;
        RECT 79.150 160.680 79.290 167.840 ;
        RECT 79.090 160.360 79.350 160.680 ;
        RECT 78.690 160.000 79.290 160.080 ;
        RECT 78.690 159.940 79.350 160.000 ;
        RECT 79.090 159.680 79.350 159.940 ;
        RECT 79.550 159.680 79.810 160.000 ;
        RECT 78.620 159.145 78.900 159.515 ;
        RECT 78.170 155.940 78.430 156.260 ;
        RECT 78.170 150.500 78.430 150.820 ;
        RECT 78.230 146.400 78.370 150.500 ;
        RECT 78.170 146.080 78.430 146.400 ;
        RECT 78.690 145.720 78.830 159.145 ;
        RECT 79.150 156.260 79.290 159.680 ;
        RECT 79.610 156.940 79.750 159.680 ;
        RECT 79.550 156.620 79.810 156.940 ;
        RECT 79.090 155.940 79.350 156.260 ;
        RECT 80.070 154.800 80.210 176.260 ;
        RECT 81.390 169.540 81.650 169.860 ;
        RECT 80.920 165.265 81.200 165.635 ;
        RECT 80.930 165.120 81.190 165.265 ;
        RECT 81.450 160.680 81.590 169.540 ;
        RECT 81.390 160.360 81.650 160.680 ;
        RECT 80.930 159.680 81.190 160.000 ;
        RECT 80.990 159.400 81.130 159.680 ;
        RECT 80.530 159.260 81.130 159.400 ;
        RECT 80.530 157.360 80.670 159.260 ;
        RECT 80.930 158.660 81.190 158.980 ;
        RECT 80.990 157.960 81.130 158.660 ;
        RECT 80.930 157.640 81.190 157.960 ;
        RECT 80.530 157.220 81.130 157.360 ;
        RECT 80.470 156.620 80.730 156.940 ;
        RECT 79.610 154.660 80.210 154.800 ;
        RECT 79.090 150.840 79.350 151.160 ;
        RECT 79.150 148.100 79.290 150.840 ;
        RECT 79.090 147.780 79.350 148.100 ;
        RECT 78.630 145.400 78.890 145.720 ;
        RECT 79.610 140.620 79.750 154.660 ;
        RECT 80.530 154.560 80.670 156.620 ;
        RECT 80.470 154.240 80.730 154.560 ;
        RECT 80.990 151.500 81.130 157.220 ;
        RECT 81.450 156.940 81.590 160.360 ;
        RECT 81.390 156.620 81.650 156.940 ;
        RECT 82.370 156.795 82.510 183.910 ;
        RECT 82.770 183.140 83.030 183.460 ;
        RECT 83.230 183.140 83.490 183.460 ;
        RECT 82.830 182.440 82.970 183.140 ;
        RECT 82.770 182.120 83.030 182.440 ;
        RECT 83.290 181.840 83.430 183.140 ;
        RECT 82.830 181.760 83.430 181.840 ;
        RECT 82.770 181.700 83.430 181.760 ;
        RECT 82.770 181.440 83.030 181.700 ;
        RECT 83.750 179.720 83.890 194.790 ;
        RECT 84.150 185.860 84.410 186.180 ;
        RECT 83.690 179.400 83.950 179.720 ;
        RECT 83.690 163.080 83.950 163.400 ;
        RECT 83.750 160.000 83.890 163.080 ;
        RECT 84.210 160.680 84.350 185.860 ;
        RECT 84.670 179.380 84.810 199.550 ;
        RECT 87.830 198.440 88.090 198.760 ;
        RECT 87.370 197.420 87.630 197.740 ;
        RECT 86.910 197.080 87.170 197.400 ;
        RECT 85.530 196.740 85.790 197.060 ;
        RECT 85.590 196.040 85.730 196.740 ;
        RECT 85.530 195.720 85.790 196.040 ;
        RECT 85.590 195.360 85.730 195.720 ;
        RECT 85.530 195.040 85.790 195.360 ;
        RECT 85.070 194.700 85.330 195.020 ;
        RECT 85.130 190.600 85.270 194.700 ;
        RECT 85.590 193.320 85.730 195.040 ;
        RECT 86.970 194.680 87.110 197.080 ;
        RECT 86.910 194.360 87.170 194.680 ;
        RECT 86.450 194.020 86.710 194.340 ;
        RECT 85.530 193.000 85.790 193.320 ;
        RECT 85.070 190.280 85.330 190.600 ;
        RECT 85.520 189.745 85.800 190.115 ;
        RECT 85.590 187.880 85.730 189.745 ;
        RECT 85.990 189.600 86.250 189.920 ;
        RECT 86.050 187.880 86.190 189.600 ;
        RECT 86.510 189.580 86.650 194.020 ;
        RECT 86.970 192.640 87.110 194.360 ;
        RECT 86.910 192.320 87.170 192.640 ;
        RECT 87.430 189.580 87.570 197.420 ;
        RECT 87.890 195.020 88.030 198.440 ;
        RECT 89.270 198.080 89.410 202.180 ;
        RECT 91.110 200.120 91.250 202.180 ;
        RECT 94.790 200.460 94.930 202.180 ;
        RECT 94.730 200.140 94.990 200.460 ;
        RECT 91.050 199.800 91.310 200.120 ;
        RECT 89.770 198.925 91.650 199.295 ;
        RECT 92.430 198.440 92.690 198.760 ;
        RECT 93.410 198.700 94.930 198.840 ;
        RECT 91.050 198.100 91.310 198.420 ;
        RECT 88.290 197.760 88.550 198.080 ;
        RECT 88.750 197.760 89.010 198.080 ;
        RECT 89.210 197.760 89.470 198.080 ;
        RECT 88.350 196.970 88.490 197.760 ;
        RECT 88.810 197.480 88.950 197.760 ;
        RECT 88.810 197.340 89.410 197.480 ;
        RECT 89.270 197.060 89.410 197.340 ;
        RECT 88.750 196.970 89.010 197.060 ;
        RECT 88.350 196.830 89.010 196.970 ;
        RECT 88.750 196.740 89.010 196.830 ;
        RECT 89.210 196.740 89.470 197.060 ;
        RECT 88.810 195.020 88.950 196.740 ;
        RECT 89.270 195.700 89.410 196.740 ;
        RECT 89.210 195.380 89.470 195.700 ;
        RECT 87.830 194.700 88.090 195.020 ;
        RECT 88.750 194.700 89.010 195.020 ;
        RECT 87.890 192.720 88.030 194.700 ;
        RECT 89.270 194.250 89.410 195.380 ;
        RECT 91.110 194.340 91.250 198.100 ;
        RECT 91.970 196.740 92.230 197.060 ;
        RECT 88.810 194.110 89.410 194.250 ;
        RECT 88.280 192.720 88.560 192.835 ;
        RECT 87.890 192.580 88.560 192.720 ;
        RECT 88.280 192.465 88.560 192.580 ;
        RECT 86.450 189.260 86.710 189.580 ;
        RECT 87.370 189.260 87.630 189.580 ;
        RECT 87.830 189.260 88.090 189.580 ;
        RECT 88.290 189.260 88.550 189.580 ;
        RECT 88.810 189.490 88.950 194.110 ;
        RECT 91.050 194.020 91.310 194.340 ;
        RECT 89.770 193.485 91.650 193.855 ;
        RECT 90.590 192.835 90.850 192.980 ;
        RECT 90.580 192.465 90.860 192.835 ;
        RECT 91.050 192.320 91.310 192.640 ;
        RECT 91.110 190.795 91.250 192.320 ;
        RECT 91.040 190.425 91.320 190.795 ;
        RECT 89.660 189.745 89.940 190.115 ;
        RECT 89.670 189.600 89.930 189.745 ;
        RECT 92.030 189.580 92.170 196.740 ;
        RECT 92.490 195.360 92.630 198.440 ;
        RECT 92.890 198.330 93.150 198.420 ;
        RECT 93.410 198.330 93.550 198.700 ;
        RECT 92.890 198.190 93.550 198.330 ;
        RECT 92.890 198.100 93.150 198.190 ;
        RECT 94.270 198.100 94.530 198.420 ;
        RECT 92.890 196.740 93.150 197.060 ;
        RECT 93.810 196.740 94.070 197.060 ;
        RECT 92.430 195.040 92.690 195.360 ;
        RECT 92.490 194.875 92.630 195.040 ;
        RECT 92.420 194.505 92.700 194.875 ;
        RECT 92.950 194.340 93.090 196.740 ;
        RECT 93.870 196.040 94.010 196.740 ;
        RECT 93.810 195.720 94.070 196.040 ;
        RECT 93.340 195.185 93.620 195.555 ;
        RECT 92.890 194.020 93.150 194.340 ;
        RECT 92.950 192.550 93.090 194.020 ;
        RECT 93.410 193.320 93.550 195.185 ;
        RECT 93.350 193.000 93.610 193.320 ;
        RECT 93.350 192.550 93.610 192.640 ;
        RECT 92.950 192.410 93.610 192.550 ;
        RECT 93.350 192.320 93.610 192.410 ;
        RECT 92.430 191.980 92.690 192.300 ;
        RECT 89.210 189.490 89.470 189.580 ;
        RECT 88.810 189.350 89.470 189.490 ;
        RECT 87.890 187.880 88.030 189.260 ;
        RECT 85.530 187.560 85.790 187.880 ;
        RECT 85.990 187.560 86.250 187.880 ;
        RECT 87.830 187.560 88.090 187.880 ;
        RECT 88.350 187.395 88.490 189.260 ;
        RECT 88.280 187.025 88.560 187.395 ;
        RECT 88.810 186.770 88.950 189.350 ;
        RECT 89.210 189.260 89.470 189.350 ;
        RECT 91.970 189.260 92.230 189.580 ;
        RECT 89.210 188.580 89.470 188.900 ;
        RECT 89.270 187.790 89.410 188.580 ;
        RECT 89.770 188.045 91.650 188.415 ;
        RECT 89.670 187.790 89.930 187.880 ;
        RECT 89.270 187.650 89.930 187.790 ;
        RECT 89.670 187.560 89.930 187.650 ;
        RECT 86.970 186.630 88.950 186.770 ;
        RECT 89.270 187.200 89.870 187.280 ;
        RECT 92.490 187.200 92.630 191.980 ;
        RECT 92.890 190.280 93.150 190.600 ;
        RECT 89.270 187.140 89.930 187.200 ;
        RECT 85.530 183.480 85.790 183.800 ;
        RECT 85.990 183.480 86.250 183.800 ;
        RECT 85.590 182.440 85.730 183.480 ;
        RECT 85.530 182.120 85.790 182.440 ;
        RECT 85.070 180.420 85.330 180.740 ;
        RECT 84.610 179.060 84.870 179.380 ;
        RECT 85.130 178.360 85.270 180.420 ;
        RECT 86.050 179.040 86.190 183.480 ;
        RECT 85.990 178.720 86.250 179.040 ;
        RECT 85.070 178.040 85.330 178.360 ;
        RECT 86.050 176.320 86.190 178.720 ;
        RECT 85.990 176.000 86.250 176.320 ;
        RECT 84.610 175.210 84.870 175.300 ;
        RECT 84.610 175.070 85.270 175.210 ;
        RECT 84.610 174.980 84.870 175.070 ;
        RECT 84.150 160.360 84.410 160.680 ;
        RECT 83.690 159.680 83.950 160.000 ;
        RECT 82.300 156.425 82.580 156.795 ;
        RECT 80.930 151.180 81.190 151.500 ;
        RECT 80.470 150.500 80.730 150.820 ;
        RECT 80.010 148.460 80.270 148.780 ;
        RECT 80.070 146.060 80.210 148.460 ;
        RECT 80.010 145.740 80.270 146.060 ;
        RECT 80.530 145.290 80.670 150.500 ;
        RECT 83.230 148.800 83.490 149.120 ;
        RECT 80.930 145.800 81.190 146.060 ;
        RECT 81.680 145.830 82.970 145.970 ;
        RECT 81.680 145.800 81.820 145.830 ;
        RECT 80.930 145.740 81.820 145.800 ;
        RECT 80.990 145.660 81.820 145.740 ;
        RECT 82.830 145.380 82.970 145.830 ;
        RECT 80.930 145.290 81.190 145.380 ;
        RECT 80.530 145.235 81.190 145.290 ;
        RECT 80.530 145.150 81.200 145.235 ;
        RECT 80.920 144.865 81.200 145.150 ;
        RECT 81.390 145.060 81.650 145.380 ;
        RECT 82.770 145.060 83.030 145.380 ;
        RECT 81.450 144.360 81.590 145.060 ;
        RECT 83.290 144.360 83.430 148.800 ;
        RECT 81.390 144.040 81.650 144.360 ;
        RECT 83.230 144.040 83.490 144.360 ;
        RECT 79.550 140.530 79.810 140.620 ;
        RECT 79.550 140.390 80.210 140.530 ;
        RECT 79.550 140.300 79.810 140.390 ;
        RECT 79.550 139.620 79.810 139.940 ;
        RECT 79.610 138.920 79.750 139.620 ;
        RECT 79.550 138.600 79.810 138.920 ;
        RECT 78.630 137.920 78.890 138.240 ;
        RECT 78.690 136.200 78.830 137.920 ;
        RECT 79.610 136.200 79.750 138.600 ;
        RECT 80.070 138.240 80.210 140.390 ;
        RECT 81.390 139.620 81.650 139.940 ;
        RECT 81.450 138.580 81.590 139.620 ;
        RECT 82.310 138.600 82.570 138.920 ;
        RECT 81.390 138.260 81.650 138.580 ;
        RECT 80.010 137.920 80.270 138.240 ;
        RECT 81.850 137.580 82.110 137.900 ;
        RECT 80.010 136.900 80.270 137.220 ;
        RECT 80.070 136.200 80.210 136.900 ;
        RECT 78.630 135.880 78.890 136.200 ;
        RECT 79.550 135.880 79.810 136.200 ;
        RECT 80.010 135.880 80.270 136.200 ;
        RECT 81.910 134.840 82.050 137.580 ;
        RECT 82.370 137.560 82.510 138.600 ;
        RECT 83.750 138.240 83.890 159.680 ;
        RECT 84.210 156.600 84.350 160.360 ;
        RECT 84.150 156.280 84.410 156.600 ;
        RECT 84.610 149.480 84.870 149.800 ;
        RECT 84.150 147.780 84.410 148.100 ;
        RECT 84.210 143.340 84.350 147.780 ;
        RECT 84.670 146.400 84.810 149.480 ;
        RECT 84.610 146.080 84.870 146.400 ;
        RECT 84.670 143.680 84.810 146.080 ;
        RECT 84.610 143.360 84.870 143.680 ;
        RECT 84.150 143.020 84.410 143.340 ;
        RECT 85.130 139.940 85.270 175.070 ;
        RECT 86.450 174.980 86.710 175.300 ;
        RECT 86.510 169.715 86.650 174.980 ;
        RECT 86.970 170.395 87.110 186.630 ;
        RECT 88.750 183.480 89.010 183.800 ;
        RECT 88.810 182.440 88.950 183.480 ;
        RECT 88.750 182.120 89.010 182.440 ;
        RECT 89.270 181.420 89.410 187.140 ;
        RECT 89.670 186.880 89.930 187.140 ;
        RECT 91.050 186.880 91.310 187.200 ;
        RECT 92.430 186.880 92.690 187.200 ;
        RECT 91.110 184.820 91.250 186.880 ;
        RECT 92.950 186.520 93.090 190.280 ;
        RECT 92.890 186.200 93.150 186.520 ;
        RECT 93.870 186.180 94.010 195.720 ;
        RECT 94.330 195.020 94.470 198.100 ;
        RECT 94.790 198.080 94.930 198.700 ;
        RECT 94.730 197.760 94.990 198.080 ;
        RECT 94.270 194.700 94.530 195.020 ;
        RECT 94.270 194.020 94.530 194.340 ;
        RECT 94.730 194.020 94.990 194.340 ;
        RECT 94.330 193.320 94.470 194.020 ;
        RECT 94.270 193.000 94.530 193.320 ;
        RECT 94.790 190.600 94.930 194.020 ;
        RECT 94.730 190.280 94.990 190.600 ;
        RECT 94.270 189.435 94.530 189.580 ;
        RECT 94.260 189.065 94.540 189.435 ;
        RECT 94.730 186.540 94.990 186.860 ;
        RECT 93.810 185.860 94.070 186.180 ;
        RECT 91.050 184.500 91.310 184.820 ;
        RECT 93.870 184.480 94.010 185.860 ;
        RECT 94.790 185.160 94.930 186.540 ;
        RECT 94.730 184.840 94.990 185.160 ;
        RECT 93.810 184.160 94.070 184.480 ;
        RECT 93.350 183.820 93.610 184.140 ;
        RECT 94.790 183.880 94.930 184.840 ;
        RECT 92.430 183.140 92.690 183.460 ;
        RECT 89.770 182.605 91.650 182.975 ;
        RECT 89.210 181.100 89.470 181.420 ;
        RECT 89.270 178.950 89.410 181.100 ;
        RECT 92.490 180.740 92.630 183.140 ;
        RECT 93.410 182.400 93.550 183.820 ;
        RECT 92.950 182.260 93.550 182.400 ;
        RECT 93.870 183.740 94.930 183.880 ;
        RECT 93.870 182.400 94.010 183.740 ;
        RECT 95.250 183.200 95.390 204.900 ;
        RECT 99.850 204.200 99.990 204.900 ;
        RECT 95.650 203.880 95.910 204.200 ;
        RECT 99.790 203.880 100.050 204.200 ;
        RECT 95.710 200.120 95.850 203.880 ;
        RECT 100.310 203.600 100.450 205.240 ;
        RECT 100.770 204.200 100.910 205.240 ;
        RECT 100.710 203.880 100.970 204.200 ;
        RECT 97.490 203.200 97.750 203.520 ;
        RECT 97.950 203.200 98.210 203.520 ;
        RECT 99.330 203.200 99.590 203.520 ;
        RECT 100.310 203.460 100.910 203.600 ;
        RECT 95.650 199.800 95.910 200.120 ;
        RECT 96.110 199.800 96.370 200.120 ;
        RECT 95.710 195.360 95.850 199.800 ;
        RECT 96.170 197.060 96.310 199.800 ;
        RECT 96.570 199.460 96.830 199.780 ;
        RECT 96.630 198.080 96.770 199.460 ;
        RECT 97.030 198.440 97.290 198.760 ;
        RECT 96.570 197.760 96.830 198.080 ;
        RECT 96.110 196.740 96.370 197.060 ;
        RECT 95.650 195.040 95.910 195.360 ;
        RECT 96.170 192.980 96.310 196.740 ;
        RECT 97.090 195.020 97.230 198.440 ;
        RECT 97.030 194.700 97.290 195.020 ;
        RECT 95.650 192.660 95.910 192.980 ;
        RECT 96.110 192.660 96.370 192.980 ;
        RECT 95.710 192.040 95.850 192.660 ;
        RECT 97.090 192.640 97.230 194.700 ;
        RECT 97.030 192.320 97.290 192.640 ;
        RECT 95.710 191.900 96.310 192.040 ;
        RECT 95.650 191.300 95.910 191.620 ;
        RECT 94.790 183.060 95.390 183.200 ;
        RECT 93.870 182.260 94.470 182.400 ;
        RECT 92.950 181.080 93.090 182.260 ;
        RECT 92.890 180.760 93.150 181.080 ;
        RECT 92.430 180.420 92.690 180.740 ;
        RECT 88.810 178.810 89.410 178.950 ;
        RECT 87.830 178.380 88.090 178.700 ;
        RECT 87.360 174.785 87.640 175.155 ;
        RECT 87.430 170.880 87.570 174.785 ;
        RECT 87.890 171.560 88.030 178.380 ;
        RECT 88.810 178.020 88.950 178.810 ;
        RECT 89.670 178.610 89.930 178.700 ;
        RECT 89.270 178.470 89.930 178.610 ;
        RECT 88.750 177.700 89.010 178.020 ;
        RECT 88.810 176.660 88.950 177.700 ;
        RECT 88.290 176.340 88.550 176.660 ;
        RECT 88.750 176.340 89.010 176.660 ;
        RECT 88.350 174.475 88.490 176.340 ;
        RECT 88.750 175.660 89.010 175.980 ;
        RECT 88.280 174.105 88.560 174.475 ;
        RECT 88.290 173.280 88.550 173.600 ;
        RECT 87.830 171.240 88.090 171.560 ;
        RECT 88.350 170.880 88.490 173.280 ;
        RECT 88.810 171.560 88.950 175.660 ;
        RECT 89.270 174.280 89.410 178.470 ;
        RECT 89.670 178.380 89.930 178.470 ;
        RECT 91.970 178.380 92.230 178.700 ;
        RECT 89.770 177.165 91.650 177.535 ;
        RECT 92.030 177.000 92.170 178.380 ;
        RECT 92.890 177.930 93.150 178.020 ;
        RECT 92.490 177.790 93.150 177.930 ;
        RECT 89.670 176.680 89.930 177.000 ;
        RECT 91.970 176.680 92.230 177.000 ;
        RECT 89.210 173.960 89.470 174.280 ;
        RECT 89.730 173.940 89.870 176.680 ;
        RECT 91.970 176.000 92.230 176.320 ;
        RECT 89.670 173.620 89.930 173.940 ;
        RECT 91.050 173.115 91.310 173.260 ;
        RECT 91.040 172.745 91.320 173.115 ;
        RECT 89.210 172.260 89.470 172.580 ;
        RECT 88.750 171.240 89.010 171.560 ;
        RECT 87.370 170.560 87.630 170.880 ;
        RECT 88.290 170.560 88.550 170.880 ;
        RECT 86.900 170.025 87.180 170.395 ;
        RECT 88.810 169.860 88.950 171.240 ;
        RECT 89.270 170.200 89.410 172.260 ;
        RECT 89.770 171.725 91.650 172.095 ;
        RECT 91.510 171.240 91.770 171.560 ;
        RECT 89.660 170.705 89.940 171.075 ;
        RECT 89.730 170.540 89.870 170.705 ;
        RECT 89.670 170.220 89.930 170.540 ;
        RECT 89.210 169.880 89.470 170.200 ;
        RECT 86.440 169.345 86.720 169.715 ;
        RECT 88.750 169.540 89.010 169.860 ;
        RECT 88.810 168.840 88.950 169.540 ;
        RECT 88.750 168.520 89.010 168.840 ;
        RECT 85.520 167.985 85.800 168.355 ;
        RECT 87.370 168.240 87.630 168.500 ;
        RECT 89.730 168.240 89.870 170.220 ;
        RECT 91.040 170.025 91.320 170.395 ;
        RECT 91.570 170.280 91.710 171.240 ;
        RECT 92.030 170.880 92.170 176.000 ;
        RECT 92.490 170.960 92.630 177.790 ;
        RECT 92.890 177.700 93.150 177.790 ;
        RECT 92.890 176.000 93.150 176.320 ;
        RECT 93.350 176.000 93.610 176.320 ;
        RECT 92.950 171.560 93.090 176.000 ;
        RECT 93.410 175.835 93.550 176.000 ;
        RECT 93.340 175.465 93.620 175.835 ;
        RECT 94.330 175.720 94.470 182.260 ;
        RECT 94.790 178.020 94.930 183.060 ;
        RECT 95.710 182.400 95.850 191.300 ;
        RECT 96.170 187.200 96.310 191.900 ;
        RECT 97.030 191.300 97.290 191.620 ;
        RECT 97.090 190.600 97.230 191.300 ;
        RECT 97.030 190.280 97.290 190.600 ;
        RECT 96.110 186.880 96.370 187.200 ;
        RECT 96.570 186.200 96.830 186.520 ;
        RECT 95.710 182.260 96.310 182.400 ;
        RECT 96.170 179.630 96.310 182.260 ;
        RECT 96.630 182.100 96.770 186.200 ;
        RECT 97.550 185.160 97.690 203.200 ;
        RECT 98.010 196.040 98.150 203.200 ;
        RECT 98.870 202.860 99.130 203.180 ;
        RECT 98.930 199.780 99.070 202.860 ;
        RECT 98.870 199.460 99.130 199.780 ;
        RECT 97.950 195.720 98.210 196.040 ;
        RECT 98.930 195.360 99.070 199.460 ;
        RECT 99.390 198.760 99.530 203.200 ;
        RECT 99.790 202.520 100.050 202.840 ;
        RECT 100.240 202.665 100.520 203.035 ;
        RECT 99.850 198.760 99.990 202.520 ;
        RECT 100.310 200.800 100.450 202.665 ;
        RECT 100.250 200.480 100.510 200.800 ;
        RECT 99.330 198.440 99.590 198.760 ;
        RECT 99.790 198.440 100.050 198.760 ;
        RECT 100.250 198.100 100.510 198.420 ;
        RECT 99.330 197.760 99.590 198.080 ;
        RECT 99.390 195.555 99.530 197.760 ;
        RECT 98.410 195.040 98.670 195.360 ;
        RECT 98.870 195.040 99.130 195.360 ;
        RECT 99.320 195.185 99.600 195.555 ;
        RECT 97.950 194.020 98.210 194.340 ;
        RECT 98.010 188.900 98.150 194.020 ;
        RECT 98.470 189.920 98.610 195.040 ;
        RECT 99.330 194.760 99.590 195.020 ;
        RECT 98.930 194.700 99.590 194.760 ;
        RECT 98.930 194.620 99.530 194.700 ;
        RECT 98.930 190.115 99.070 194.620 ;
        RECT 99.780 194.505 100.060 194.875 ;
        RECT 99.790 194.360 100.050 194.505 ;
        RECT 99.330 192.660 99.590 192.980 ;
        RECT 98.410 189.600 98.670 189.920 ;
        RECT 98.860 189.745 99.140 190.115 ;
        RECT 97.950 188.755 98.210 188.900 ;
        RECT 97.940 188.385 98.220 188.755 ;
        RECT 98.930 187.960 99.070 189.745 ;
        RECT 99.390 189.580 99.530 192.660 ;
        RECT 99.790 191.980 100.050 192.300 ;
        RECT 99.330 189.260 99.590 189.580 ;
        RECT 99.850 189.240 99.990 191.980 ;
        RECT 100.310 190.260 100.450 198.100 ;
        RECT 100.770 197.595 100.910 203.460 ;
        RECT 101.690 201.480 101.830 206.260 ;
        RECT 102.090 205.580 102.350 205.900 ;
        RECT 103.470 205.580 103.730 205.900 ;
        RECT 102.150 201.480 102.290 205.580 ;
        RECT 103.010 202.920 103.270 203.180 ;
        RECT 102.610 202.860 103.270 202.920 ;
        RECT 102.610 202.780 103.210 202.860 ;
        RECT 101.630 201.160 101.890 201.480 ;
        RECT 102.090 201.160 102.350 201.480 ;
        RECT 100.700 197.225 100.980 197.595 ;
        RECT 101.170 197.420 101.430 197.740 ;
        RECT 100.710 195.720 100.970 196.040 ;
        RECT 100.770 195.020 100.910 195.720 ;
        RECT 101.230 195.700 101.370 197.420 ;
        RECT 101.170 195.380 101.430 195.700 ;
        RECT 100.710 194.700 100.970 195.020 ;
        RECT 100.710 194.020 100.970 194.340 ;
        RECT 100.250 189.940 100.510 190.260 ;
        RECT 99.790 188.920 100.050 189.240 ;
        RECT 99.780 187.960 100.060 188.075 ;
        RECT 98.930 187.820 100.060 187.960 ;
        RECT 99.780 187.705 100.060 187.820 ;
        RECT 98.400 187.025 98.680 187.395 ;
        RECT 99.790 187.220 100.050 187.540 ;
        RECT 98.410 186.880 98.670 187.025 ;
        RECT 97.490 184.840 97.750 185.160 ;
        RECT 99.330 183.820 99.590 184.140 ;
        RECT 99.850 183.995 99.990 187.220 ;
        RECT 98.870 183.480 99.130 183.800 ;
        RECT 96.570 181.780 96.830 182.100 ;
        RECT 98.930 181.760 99.070 183.480 ;
        RECT 99.390 182.635 99.530 183.820 ;
        RECT 99.780 183.625 100.060 183.995 ;
        RECT 99.320 182.265 99.600 182.635 ;
        RECT 100.310 182.100 100.450 189.940 ;
        RECT 100.770 184.480 100.910 194.020 ;
        RECT 101.230 190.600 101.370 195.380 ;
        RECT 102.610 195.020 102.750 202.780 ;
        RECT 103.010 202.180 103.270 202.500 ;
        RECT 101.630 194.700 101.890 195.020 ;
        RECT 102.550 194.700 102.810 195.020 ;
        RECT 101.170 190.280 101.430 190.600 ;
        RECT 100.710 184.160 100.970 184.480 ;
        RECT 101.170 184.160 101.430 184.480 ;
        RECT 100.250 181.780 100.510 182.100 ;
        RECT 101.230 181.840 101.370 184.160 ;
        RECT 101.690 183.800 101.830 194.700 ;
        RECT 102.090 192.210 102.350 192.300 ;
        RECT 102.090 192.070 102.750 192.210 ;
        RECT 102.090 191.980 102.350 192.070 ;
        RECT 102.090 190.280 102.350 190.600 ;
        RECT 102.150 187.540 102.290 190.280 ;
        RECT 102.610 187.880 102.750 192.070 ;
        RECT 102.550 187.560 102.810 187.880 ;
        RECT 102.090 187.220 102.350 187.540 ;
        RECT 102.550 186.880 102.810 187.200 ;
        RECT 102.610 186.715 102.750 186.880 ;
        RECT 102.540 186.345 102.820 186.715 ;
        RECT 103.070 185.160 103.210 202.180 ;
        RECT 103.530 196.915 103.670 205.580 ;
        RECT 103.990 201.480 104.130 207.620 ;
        RECT 104.450 206.830 104.590 207.960 ;
        RECT 104.770 207.085 106.650 207.455 ;
        RECT 107.210 206.920 107.350 209.455 ;
        RECT 111.350 206.920 111.490 209.455 ;
        RECT 104.450 206.690 105.050 206.830 ;
        RECT 104.390 205.920 104.650 206.240 ;
        RECT 104.450 201.480 104.590 205.920 ;
        RECT 104.910 203.035 105.050 206.690 ;
        RECT 107.150 206.600 107.410 206.920 ;
        RECT 111.290 206.600 111.550 206.920 ;
        RECT 115.490 205.900 115.630 209.455 ;
        RECT 119.630 205.900 119.770 209.455 ;
        RECT 123.770 206.920 123.910 209.455 ;
        RECT 126.930 207.960 127.190 208.280 ;
        RECT 125.090 207.620 125.350 207.940 ;
        RECT 123.710 206.600 123.970 206.920 ;
        RECT 125.150 205.900 125.290 207.620 ;
        RECT 126.010 205.920 126.270 206.240 ;
        RECT 107.610 205.580 107.870 205.900 ;
        RECT 113.130 205.580 113.390 205.900 ;
        RECT 115.430 205.580 115.690 205.900 ;
        RECT 119.570 205.580 119.830 205.900 ;
        RECT 121.870 205.580 122.130 205.900 ;
        RECT 125.090 205.580 125.350 205.900 ;
        RECT 104.840 202.665 105.120 203.035 ;
        RECT 104.850 202.520 105.110 202.665 ;
        RECT 104.770 201.645 106.650 202.015 ;
        RECT 103.930 201.160 104.190 201.480 ;
        RECT 104.390 201.160 104.650 201.480 ;
        RECT 107.670 200.880 107.810 205.580 ;
        RECT 110.830 204.900 111.090 205.220 ;
        RECT 110.890 202.500 111.030 204.900 ;
        RECT 113.190 203.715 113.330 205.580 ;
        RECT 114.510 204.900 114.770 205.220 ;
        RECT 114.970 204.900 115.230 205.220 ;
        RECT 118.190 204.900 118.450 205.220 ;
        RECT 118.650 204.900 118.910 205.220 ;
        RECT 114.570 204.200 114.710 204.900 ;
        RECT 114.510 203.880 114.770 204.200 ;
        RECT 113.120 203.345 113.400 203.715 ;
        RECT 114.050 203.600 114.310 203.860 ;
        RECT 115.030 203.600 115.170 204.900 ;
        RECT 114.050 203.540 115.170 203.600 ;
        RECT 114.110 203.460 115.170 203.540 ;
        RECT 118.250 203.520 118.390 204.900 ;
        RECT 118.710 204.200 118.850 204.900 ;
        RECT 119.770 204.365 121.650 204.735 ;
        RECT 118.650 203.880 118.910 204.200 ;
        RECT 110.830 202.180 111.090 202.500 ;
        RECT 114.050 202.180 114.310 202.500 ;
        RECT 107.670 200.740 108.730 200.880 ;
        RECT 107.150 200.140 107.410 200.460 ;
        RECT 107.610 200.140 107.870 200.460 ;
        RECT 105.310 199.460 105.570 199.780 ;
        RECT 105.370 198.420 105.510 199.460 ;
        RECT 105.310 198.100 105.570 198.420 ;
        RECT 103.930 197.420 104.190 197.740 ;
        RECT 104.390 197.420 104.650 197.740 ;
        RECT 103.460 196.545 103.740 196.915 ;
        RECT 103.460 195.440 103.740 195.555 ;
        RECT 103.990 195.440 104.130 197.420 ;
        RECT 103.460 195.300 104.130 195.440 ;
        RECT 103.460 195.185 103.740 195.300 ;
        RECT 103.470 194.020 103.730 194.340 ;
        RECT 103.010 185.070 103.270 185.160 ;
        RECT 102.610 184.930 103.270 185.070 ;
        RECT 101.630 183.480 101.890 183.800 ;
        RECT 102.090 183.480 102.350 183.800 ;
        RECT 102.150 182.440 102.290 183.480 ;
        RECT 102.090 182.120 102.350 182.440 ;
        RECT 98.870 181.440 99.130 181.760 ;
        RECT 96.170 179.490 98.150 179.630 ;
        RECT 97.490 178.720 97.750 179.040 ;
        RECT 94.730 177.700 94.990 178.020 ;
        RECT 97.020 176.145 97.300 176.515 ;
        RECT 97.030 176.000 97.290 176.145 ;
        RECT 93.810 175.320 94.070 175.640 ;
        RECT 94.330 175.580 95.390 175.720 ;
        RECT 96.570 175.660 96.830 175.980 ;
        RECT 93.350 172.940 93.610 173.260 ;
        RECT 93.410 171.560 93.550 172.940 ;
        RECT 92.890 171.240 93.150 171.560 ;
        RECT 93.350 171.240 93.610 171.560 ;
        RECT 91.970 170.560 92.230 170.880 ;
        RECT 92.490 170.820 93.090 170.960 ;
        RECT 91.570 170.140 92.630 170.280 ;
        RECT 90.580 169.345 90.860 169.715 ;
        RECT 87.370 168.180 89.870 168.240 ;
        RECT 87.430 168.100 89.870 168.180 ;
        RECT 85.530 167.840 85.790 167.985 ;
        RECT 86.910 167.500 87.170 167.820 ;
        RECT 86.970 165.440 87.110 167.500 ;
        RECT 87.370 167.160 87.630 167.480 ;
        RECT 86.910 165.120 87.170 165.440 ;
        RECT 87.430 162.380 87.570 167.160 ;
        RECT 87.890 162.720 88.030 168.100 ;
        RECT 90.650 167.820 90.790 169.345 ;
        RECT 88.290 167.500 88.550 167.820 ;
        RECT 88.750 167.500 89.010 167.820 ;
        RECT 90.590 167.500 90.850 167.820 ;
        RECT 87.830 162.400 88.090 162.720 ;
        RECT 87.370 162.060 87.630 162.380 ;
        RECT 86.910 161.720 87.170 162.040 ;
        RECT 85.530 159.000 85.790 159.320 ;
        RECT 85.590 154.900 85.730 159.000 ;
        RECT 85.530 154.580 85.790 154.900 ;
        RECT 85.990 153.220 86.250 153.540 ;
        RECT 86.050 149.120 86.190 153.220 ;
        RECT 86.450 152.200 86.710 152.520 ;
        RECT 85.990 148.800 86.250 149.120 ;
        RECT 86.510 148.780 86.650 152.200 ;
        RECT 85.530 148.460 85.790 148.780 ;
        RECT 86.450 148.460 86.710 148.780 ;
        RECT 85.590 145.720 85.730 148.460 ;
        RECT 85.990 148.120 86.250 148.440 ;
        RECT 86.050 146.060 86.190 148.120 ;
        RECT 85.990 145.740 86.250 146.060 ;
        RECT 85.530 145.400 85.790 145.720 ;
        RECT 85.590 143.340 85.730 145.400 ;
        RECT 85.530 143.020 85.790 143.340 ;
        RECT 85.530 142.340 85.790 142.660 ;
        RECT 85.590 140.620 85.730 142.340 ;
        RECT 85.530 140.300 85.790 140.620 ;
        RECT 85.070 139.620 85.330 139.940 ;
        RECT 86.970 138.490 87.110 161.720 ;
        RECT 88.350 160.000 88.490 167.500 ;
        RECT 88.810 166.120 88.950 167.500 ;
        RECT 91.110 167.480 91.250 170.025 ;
        RECT 91.970 169.540 92.230 169.860 ;
        RECT 91.050 167.160 91.310 167.480 ;
        RECT 89.770 166.285 91.650 166.655 ;
        RECT 88.750 166.030 89.010 166.120 ;
        RECT 88.750 165.890 89.410 166.030 ;
        RECT 88.750 165.800 89.010 165.890 ;
        RECT 89.270 160.680 89.410 165.890 ;
        RECT 92.030 165.100 92.170 169.540 ;
        RECT 92.490 167.560 92.630 170.140 ;
        RECT 92.950 168.240 93.090 170.820 ;
        RECT 93.350 170.790 93.610 170.880 ;
        RECT 93.870 170.790 94.010 175.320 ;
        RECT 94.730 174.980 94.990 175.300 ;
        RECT 94.260 173.425 94.540 173.795 ;
        RECT 94.270 173.280 94.530 173.425 ;
        RECT 94.270 172.600 94.530 172.920 ;
        RECT 94.330 170.880 94.470 172.600 ;
        RECT 94.790 172.580 94.930 174.980 ;
        RECT 94.730 172.260 94.990 172.580 ;
        RECT 94.790 171.560 94.930 172.260 ;
        RECT 94.730 171.240 94.990 171.560 ;
        RECT 93.350 170.650 94.010 170.790 ;
        RECT 93.350 170.560 93.610 170.650 ;
        RECT 94.270 170.560 94.530 170.880 ;
        RECT 93.810 169.880 94.070 170.200 ;
        RECT 92.950 168.100 93.550 168.240 ;
        RECT 93.870 168.160 94.010 169.880 ;
        RECT 94.330 168.840 94.470 170.560 ;
        RECT 95.250 170.280 95.390 175.580 ;
        RECT 95.650 175.155 95.910 175.300 ;
        RECT 95.640 174.785 95.920 175.155 ;
        RECT 96.630 173.680 96.770 175.660 ;
        RECT 97.030 173.960 97.290 174.280 ;
        RECT 94.790 170.140 95.390 170.280 ;
        RECT 95.710 173.540 96.770 173.680 ;
        RECT 94.270 168.520 94.530 168.840 ;
        RECT 92.490 167.420 93.090 167.560 ;
        RECT 92.430 166.820 92.690 167.140 ;
        RECT 92.490 166.120 92.630 166.820 ;
        RECT 92.430 165.800 92.690 166.120 ;
        RECT 91.970 164.780 92.230 165.100 ;
        RECT 89.770 160.845 91.650 161.215 ;
        RECT 89.210 160.360 89.470 160.680 ;
        RECT 88.290 159.680 88.550 160.000 ;
        RECT 89.670 159.680 89.930 160.000 ;
        RECT 92.430 159.910 92.690 160.000 ;
        RECT 92.950 159.910 93.090 167.420 ;
        RECT 92.430 159.770 93.090 159.910 ;
        RECT 92.430 159.680 92.690 159.770 ;
        RECT 87.830 159.000 88.090 159.320 ;
        RECT 87.890 156.940 88.030 159.000 ;
        RECT 89.210 157.640 89.470 157.960 ;
        RECT 88.750 157.300 89.010 157.620 ;
        RECT 87.830 156.620 88.090 156.940 ;
        RECT 87.370 156.280 87.630 156.600 ;
        RECT 87.430 155.240 87.570 156.280 ;
        RECT 87.370 154.920 87.630 155.240 ;
        RECT 87.430 154.560 87.570 154.920 ;
        RECT 88.810 154.900 88.950 157.300 ;
        RECT 88.750 154.580 89.010 154.900 ;
        RECT 87.370 154.240 87.630 154.560 ;
        RECT 88.290 153.560 88.550 153.880 ;
        RECT 87.830 149.480 88.090 149.800 ;
        RECT 87.890 149.120 88.030 149.480 ;
        RECT 87.830 148.800 88.090 149.120 ;
        RECT 87.370 145.740 87.630 146.060 ;
        RECT 87.430 145.380 87.570 145.740 ;
        RECT 87.890 145.720 88.030 148.800 ;
        RECT 87.830 145.400 88.090 145.720 ;
        RECT 87.370 145.060 87.630 145.380 ;
        RECT 87.430 140.620 87.570 145.060 ;
        RECT 87.370 140.300 87.630 140.620 ;
        RECT 85.590 138.350 87.110 138.490 ;
        RECT 83.690 137.920 83.950 138.240 ;
        RECT 82.310 137.240 82.570 137.560 ;
        RECT 81.850 134.520 82.110 134.840 ;
        RECT 78.170 134.180 78.430 134.500 ;
        RECT 78.230 130.420 78.370 134.180 ;
        RECT 85.070 133.160 85.330 133.480 ;
        RECT 82.770 132.480 83.030 132.800 ;
        RECT 78.170 130.100 78.430 130.420 ;
        RECT 76.780 129.225 77.060 129.595 ;
        RECT 77.250 129.420 77.510 129.740 ;
        RECT 77.710 129.420 77.970 129.740 ;
        RECT 76.850 128.040 76.990 129.225 ;
        RECT 77.250 128.740 77.510 129.060 ;
        RECT 74.030 127.720 74.290 128.040 ;
        RECT 76.790 127.720 77.050 128.040 ;
        RECT 73.570 126.020 73.830 126.340 ;
        RECT 76.790 126.020 77.050 126.340 ;
        RECT 73.630 124.300 73.770 126.020 ;
        RECT 74.770 125.485 76.650 125.855 ;
        RECT 76.850 124.300 76.990 126.020 ;
        RECT 77.310 124.300 77.450 128.740 ;
        RECT 77.770 127.700 77.910 129.420 ;
        RECT 78.230 128.040 78.370 130.100 ;
        RECT 79.550 129.420 79.810 129.740 ;
        RECT 81.390 129.420 81.650 129.740 ;
        RECT 78.170 127.720 78.430 128.040 ;
        RECT 77.710 127.380 77.970 127.700 ;
        RECT 78.170 124.660 78.430 124.980 ;
        RECT 73.570 123.980 73.830 124.300 ;
        RECT 76.790 123.980 77.050 124.300 ;
        RECT 77.250 123.980 77.510 124.300 ;
        RECT 70.810 123.300 71.070 123.620 ;
        RECT 74.490 123.300 74.750 123.620 ;
        RECT 70.870 122.230 71.010 123.300 ;
        RECT 74.550 122.230 74.690 123.300 ;
        RECT 78.230 122.230 78.370 124.660 ;
        RECT 79.610 124.300 79.750 129.420 ;
        RECT 80.010 128.740 80.270 129.060 ;
        RECT 80.070 124.640 80.210 128.740 ;
        RECT 81.450 128.040 81.590 129.420 ;
        RECT 82.830 129.060 82.970 132.480 ;
        RECT 84.150 131.800 84.410 132.120 ;
        RECT 84.210 129.400 84.350 131.800 ;
        RECT 84.610 131.460 84.870 131.780 ;
        RECT 84.670 130.760 84.810 131.460 ;
        RECT 84.610 130.440 84.870 130.760 ;
        RECT 84.150 129.080 84.410 129.400 ;
        RECT 81.850 128.740 82.110 129.060 ;
        RECT 82.770 128.740 83.030 129.060 ;
        RECT 81.390 127.720 81.650 128.040 ;
        RECT 80.470 127.040 80.730 127.360 ;
        RECT 80.530 125.320 80.670 127.040 ;
        RECT 81.910 126.340 82.050 128.740 ;
        RECT 82.830 127.360 82.970 128.740 ;
        RECT 82.770 127.040 83.030 127.360 ;
        RECT 84.210 126.680 84.350 129.080 ;
        RECT 84.610 128.740 84.870 129.060 ;
        RECT 84.670 128.040 84.810 128.740 ;
        RECT 84.610 127.720 84.870 128.040 ;
        RECT 85.130 127.020 85.270 133.160 ;
        RECT 85.590 132.995 85.730 138.350 ;
        RECT 87.430 137.900 87.570 140.300 ;
        RECT 87.370 137.580 87.630 137.900 ;
        RECT 88.350 134.920 88.490 153.560 ;
        RECT 89.270 153.540 89.410 157.640 ;
        RECT 89.730 156.600 89.870 159.680 ;
        RECT 92.490 156.940 92.630 159.680 ;
        RECT 92.950 158.980 93.090 159.770 ;
        RECT 92.890 158.660 93.150 158.980 ;
        RECT 92.890 157.640 93.150 157.960 ;
        RECT 92.430 156.620 92.690 156.940 ;
        RECT 89.670 156.280 89.930 156.600 ;
        RECT 92.430 155.940 92.690 156.260 ;
        RECT 89.770 155.405 91.650 155.775 ;
        RECT 89.670 154.920 89.930 155.240 ;
        RECT 89.730 154.560 89.870 154.920 ;
        RECT 89.670 154.240 89.930 154.560 ;
        RECT 91.970 153.560 92.230 153.880 ;
        RECT 89.210 153.220 89.470 153.540 ;
        RECT 89.670 153.220 89.930 153.540 ;
        RECT 89.730 150.730 89.870 153.220 ;
        RECT 89.270 150.590 89.870 150.730 ;
        RECT 88.750 145.235 89.010 145.380 ;
        RECT 88.740 144.865 89.020 145.235 ;
        RECT 88.750 141.320 89.010 141.640 ;
        RECT 88.810 138.240 88.950 141.320 ;
        RECT 88.750 137.920 89.010 138.240 ;
        RECT 89.270 135.520 89.410 150.590 ;
        RECT 89.770 149.965 91.650 150.335 ;
        RECT 89.770 144.525 91.650 144.895 ;
        RECT 91.510 142.680 91.770 143.000 ;
        RECT 91.570 141.300 91.710 142.680 ;
        RECT 91.510 140.980 91.770 141.300 ;
        RECT 89.770 139.085 91.650 139.455 ;
        RECT 90.120 136.705 90.400 137.075 ;
        RECT 89.210 135.200 89.470 135.520 ;
        RECT 90.190 135.180 90.330 136.705 ;
        RECT 92.030 136.200 92.170 153.560 ;
        RECT 92.490 148.780 92.630 155.940 ;
        RECT 92.430 148.460 92.690 148.780 ;
        RECT 92.430 145.740 92.690 146.060 ;
        RECT 92.950 145.915 93.090 157.640 ;
        RECT 92.490 143.680 92.630 145.740 ;
        RECT 92.880 145.545 93.160 145.915 ;
        RECT 92.950 143.680 93.090 145.545 ;
        RECT 92.430 143.360 92.690 143.680 ;
        RECT 92.890 143.360 93.150 143.680 ;
        RECT 92.490 143.195 92.630 143.360 ;
        RECT 92.420 142.825 92.700 143.195 ;
        RECT 92.420 140.105 92.700 140.475 ;
        RECT 92.490 139.940 92.630 140.105 ;
        RECT 92.430 139.620 92.690 139.940 ;
        RECT 92.950 138.580 93.090 143.360 ;
        RECT 92.890 138.260 93.150 138.580 ;
        RECT 91.970 135.880 92.230 136.200 ;
        RECT 86.510 134.840 88.490 134.920 ;
        RECT 90.130 134.860 90.390 135.180 ;
        RECT 86.510 134.780 88.550 134.840 ;
        RECT 85.520 132.625 85.800 132.995 ;
        RECT 85.990 132.820 86.250 133.140 ;
        RECT 85.590 132.460 85.730 132.625 ;
        RECT 85.530 132.140 85.790 132.460 ;
        RECT 85.530 130.330 85.790 130.420 ;
        RECT 86.050 130.330 86.190 132.820 ;
        RECT 86.510 132.800 86.650 134.780 ;
        RECT 88.290 134.520 88.550 134.780 ;
        RECT 86.910 134.180 87.170 134.500 ;
        RECT 89.210 134.180 89.470 134.500 ;
        RECT 91.970 134.180 92.230 134.500 ;
        RECT 86.970 132.800 87.110 134.180 ;
        RECT 89.270 132.800 89.410 134.180 ;
        RECT 89.770 133.645 91.650 134.015 ;
        RECT 90.130 133.160 90.390 133.480 ;
        RECT 86.450 132.480 86.710 132.800 ;
        RECT 86.910 132.480 87.170 132.800 ;
        RECT 89.210 132.480 89.470 132.800 ;
        RECT 85.530 130.190 86.190 130.330 ;
        RECT 85.530 130.100 85.790 130.190 ;
        RECT 85.530 129.420 85.790 129.740 ;
        RECT 85.590 128.040 85.730 129.420 ;
        RECT 85.530 127.720 85.790 128.040 ;
        RECT 86.050 127.020 86.190 130.190 ;
        RECT 86.510 127.360 86.650 132.480 ;
        RECT 88.290 131.460 88.550 131.780 ;
        RECT 88.350 129.740 88.490 131.460 ;
        RECT 89.270 130.080 89.410 132.480 ;
        RECT 89.670 131.800 89.930 132.120 ;
        RECT 89.730 130.080 89.870 131.800 ;
        RECT 90.190 130.080 90.330 133.160 ;
        RECT 90.590 130.330 90.850 130.420 ;
        RECT 91.510 130.330 91.770 130.420 ;
        RECT 90.590 130.190 91.770 130.330 ;
        RECT 90.590 130.100 90.850 130.190 ;
        RECT 91.510 130.100 91.770 130.190 ;
        RECT 89.210 129.760 89.470 130.080 ;
        RECT 89.670 129.760 89.930 130.080 ;
        RECT 90.130 129.760 90.390 130.080 ;
        RECT 86.910 129.420 87.170 129.740 ;
        RECT 87.370 129.420 87.630 129.740 ;
        RECT 88.290 129.650 88.550 129.740 ;
        RECT 87.890 129.510 88.550 129.650 ;
        RECT 86.970 127.700 87.110 129.420 ;
        RECT 86.910 127.380 87.170 127.700 ;
        RECT 86.450 127.040 86.710 127.360 ;
        RECT 85.070 126.700 85.330 127.020 ;
        RECT 85.990 126.700 86.250 127.020 ;
        RECT 87.430 126.760 87.570 129.420 ;
        RECT 87.890 127.360 88.030 129.510 ;
        RECT 88.290 129.420 88.550 129.510 ;
        RECT 87.830 127.040 88.090 127.360 ;
        RECT 88.280 127.185 88.560 127.555 ;
        RECT 89.270 127.360 89.410 129.760 ;
        RECT 89.770 128.205 91.650 128.575 ;
        RECT 92.030 128.040 92.170 134.180 ;
        RECT 93.410 134.100 93.550 168.100 ;
        RECT 93.810 167.840 94.070 168.160 ;
        RECT 94.270 167.500 94.530 167.820 ;
        RECT 93.810 164.780 94.070 165.100 ;
        RECT 93.870 161.700 94.010 164.780 ;
        RECT 93.810 161.380 94.070 161.700 ;
        RECT 93.870 160.340 94.010 161.380 ;
        RECT 93.810 160.020 94.070 160.340 ;
        RECT 93.870 157.280 94.010 160.020 ;
        RECT 94.330 160.000 94.470 167.500 ;
        RECT 94.270 159.680 94.530 160.000 ;
        RECT 94.270 158.660 94.530 158.980 ;
        RECT 94.330 157.620 94.470 158.660 ;
        RECT 94.270 157.300 94.530 157.620 ;
        RECT 93.810 156.960 94.070 157.280 ;
        RECT 93.810 155.940 94.070 156.260 ;
        RECT 93.870 146.400 94.010 155.940 ;
        RECT 94.270 154.580 94.530 154.900 ;
        RECT 94.330 148.440 94.470 154.580 ;
        RECT 94.270 148.120 94.530 148.440 ;
        RECT 94.790 147.840 94.930 170.140 ;
        RECT 95.710 165.440 95.850 173.540 ;
        RECT 96.570 172.260 96.830 172.580 ;
        RECT 96.630 170.880 96.770 172.260 ;
        RECT 96.570 170.560 96.830 170.880 ;
        RECT 97.090 168.840 97.230 173.960 ;
        RECT 97.550 171.560 97.690 178.720 ;
        RECT 97.490 171.240 97.750 171.560 ;
        RECT 97.030 168.520 97.290 168.840 ;
        RECT 96.570 168.180 96.830 168.500 ;
        RECT 95.650 165.120 95.910 165.440 ;
        RECT 96.630 163.400 96.770 168.180 ;
        RECT 95.650 163.080 95.910 163.400 ;
        RECT 96.570 163.080 96.830 163.400 ;
        RECT 95.710 160.000 95.850 163.080 ;
        RECT 97.490 162.800 97.750 163.060 ;
        RECT 97.090 162.740 97.750 162.800 ;
        RECT 97.090 162.660 97.690 162.740 ;
        RECT 96.110 162.060 96.370 162.380 ;
        RECT 95.650 159.680 95.910 160.000 ;
        RECT 95.190 158.660 95.450 158.980 ;
        RECT 95.250 157.960 95.390 158.660 ;
        RECT 95.190 157.640 95.450 157.960 ;
        RECT 95.710 156.940 95.850 159.680 ;
        RECT 95.650 156.620 95.910 156.940 ;
        RECT 96.170 156.000 96.310 162.060 ;
        RECT 97.090 157.960 97.230 162.660 ;
        RECT 97.490 162.235 97.750 162.380 ;
        RECT 97.480 161.865 97.760 162.235 ;
        RECT 97.490 160.020 97.750 160.340 ;
        RECT 98.010 160.080 98.150 179.490 ;
        RECT 98.930 179.380 99.070 181.440 ;
        RECT 98.870 179.060 99.130 179.380 ;
        RECT 99.790 178.720 100.050 179.040 ;
        RECT 98.870 178.040 99.130 178.360 ;
        RECT 98.400 177.505 98.680 177.875 ;
        RECT 98.470 170.540 98.610 177.505 ;
        RECT 98.930 172.435 99.070 178.040 ;
        RECT 99.850 175.980 99.990 178.720 ;
        RECT 100.310 178.700 100.450 181.780 ;
        RECT 101.230 181.760 101.830 181.840 ;
        RECT 101.230 181.700 101.890 181.760 ;
        RECT 101.630 181.440 101.890 181.700 ;
        RECT 101.170 181.100 101.430 181.420 ;
        RECT 100.710 180.420 100.970 180.740 ;
        RECT 100.250 178.380 100.510 178.700 ;
        RECT 99.790 175.660 100.050 175.980 ;
        RECT 100.250 174.980 100.510 175.300 ;
        RECT 100.310 173.940 100.450 174.980 ;
        RECT 100.770 173.940 100.910 180.420 ;
        RECT 101.230 179.040 101.370 181.100 ;
        RECT 102.610 179.235 102.750 184.930 ;
        RECT 103.010 184.840 103.270 184.930 ;
        RECT 103.530 184.140 103.670 194.020 ;
        RECT 104.450 193.400 104.590 197.420 ;
        RECT 104.770 196.205 106.650 196.575 ;
        RECT 106.230 195.950 106.490 196.040 ;
        RECT 107.210 195.950 107.350 200.140 ;
        RECT 107.670 198.760 107.810 200.140 ;
        RECT 107.610 198.440 107.870 198.760 ;
        RECT 107.610 196.740 107.870 197.060 ;
        RECT 106.230 195.810 107.350 195.950 ;
        RECT 106.230 195.720 106.490 195.810 ;
        RECT 107.670 195.610 107.810 196.740 ;
        RECT 107.210 195.470 107.810 195.610 ;
        RECT 104.850 195.270 105.110 195.360 ;
        RECT 104.850 195.130 106.430 195.270 ;
        RECT 104.850 195.040 105.110 195.130 ;
        RECT 104.850 194.020 105.110 194.340 ;
        RECT 103.990 193.260 104.590 193.400 ;
        RECT 104.910 193.320 105.050 194.020 ;
        RECT 106.290 193.320 106.430 195.130 ;
        RECT 106.690 194.875 106.950 195.020 ;
        RECT 106.680 194.505 106.960 194.875 ;
        RECT 103.990 190.600 104.130 193.260 ;
        RECT 104.850 193.000 105.110 193.320 ;
        RECT 106.230 193.000 106.490 193.320 ;
        RECT 104.380 191.785 104.660 192.155 ;
        RECT 103.930 190.280 104.190 190.600 ;
        RECT 104.450 189.920 104.590 191.785 ;
        RECT 107.210 191.620 107.350 195.470 ;
        RECT 108.070 195.380 108.330 195.700 ;
        RECT 107.610 192.660 107.870 192.980 ;
        RECT 107.150 191.300 107.410 191.620 ;
        RECT 104.770 190.765 106.650 191.135 ;
        RECT 107.140 190.510 107.420 190.795 ;
        RECT 105.370 190.425 107.420 190.510 ;
        RECT 105.370 190.370 107.350 190.425 ;
        RECT 105.370 190.115 105.510 190.370 ;
        RECT 104.390 189.600 104.650 189.920 ;
        RECT 105.300 189.745 105.580 190.115 ;
        RECT 106.220 189.745 106.500 190.115 ;
        RECT 104.850 189.260 105.110 189.580 ;
        RECT 104.910 187.540 105.050 189.260 ;
        RECT 106.290 187.880 106.430 189.745 ;
        RECT 106.690 189.260 106.950 189.580 ;
        RECT 106.230 187.560 106.490 187.880 ;
        RECT 104.850 187.220 105.110 187.540 ;
        RECT 106.750 186.090 106.890 189.260 ;
        RECT 107.210 186.860 107.350 190.370 ;
        RECT 107.670 189.580 107.810 192.660 ;
        RECT 108.130 190.600 108.270 195.380 ;
        RECT 108.070 190.280 108.330 190.600 ;
        RECT 107.610 189.260 107.870 189.580 ;
        RECT 107.670 187.540 107.810 189.260 ;
        RECT 107.610 187.220 107.870 187.540 ;
        RECT 107.150 186.540 107.410 186.860 ;
        RECT 106.750 185.950 107.350 186.090 ;
        RECT 104.770 185.325 106.650 185.695 ;
        RECT 103.470 183.820 103.730 184.140 ;
        RECT 107.210 183.460 107.350 185.950 ;
        RECT 107.610 185.860 107.870 186.180 ;
        RECT 108.590 186.090 108.730 200.740 ;
        RECT 108.990 200.140 109.250 200.460 ;
        RECT 109.050 194.680 109.190 200.140 ;
        RECT 112.210 199.800 112.470 200.120 ;
        RECT 110.370 199.460 110.630 199.780 ;
        RECT 109.910 195.380 110.170 195.700 ;
        RECT 109.970 194.875 110.110 195.380 ;
        RECT 108.990 194.360 109.250 194.680 ;
        RECT 109.900 194.505 110.180 194.875 ;
        RECT 109.450 192.320 109.710 192.640 ;
        RECT 109.910 192.320 110.170 192.640 ;
        RECT 109.510 189.920 109.650 192.320 ;
        RECT 109.970 191.475 110.110 192.320 ;
        RECT 109.900 191.105 110.180 191.475 ;
        RECT 108.990 189.600 109.250 189.920 ;
        RECT 109.450 189.600 109.710 189.920 ;
        RECT 108.130 185.950 108.730 186.090 ;
        RECT 103.010 183.140 103.270 183.460 ;
        RECT 107.150 183.140 107.410 183.460 ;
        RECT 107.670 183.315 107.810 185.860 ;
        RECT 101.170 178.720 101.430 179.040 ;
        RECT 102.540 178.865 102.820 179.235 ;
        RECT 103.070 178.700 103.210 183.140 ;
        RECT 107.600 182.945 107.880 183.315 ;
        RECT 107.600 182.265 107.880 182.635 ;
        RECT 107.610 182.120 107.870 182.265 ;
        RECT 108.130 181.840 108.270 185.950 ;
        RECT 104.390 181.440 104.650 181.760 ;
        RECT 106.750 181.700 108.270 181.840 ;
        RECT 103.470 180.760 103.730 181.080 ;
        RECT 103.010 178.380 103.270 178.700 ;
        RECT 102.550 176.680 102.810 177.000 ;
        RECT 101.170 176.000 101.430 176.320 ;
        RECT 101.630 176.000 101.890 176.320 ;
        RECT 102.090 176.000 102.350 176.320 ;
        RECT 99.780 173.425 100.060 173.795 ;
        RECT 100.250 173.620 100.510 173.940 ;
        RECT 100.710 173.620 100.970 173.940 ;
        RECT 99.790 173.280 100.050 173.425 ;
        RECT 99.790 172.600 100.050 172.920 ;
        RECT 100.250 172.600 100.510 172.920 ;
        RECT 98.860 172.065 99.140 172.435 ;
        RECT 99.330 172.260 99.590 172.580 ;
        RECT 98.410 170.220 98.670 170.540 ;
        RECT 98.930 167.820 99.070 172.065 ;
        RECT 99.390 170.540 99.530 172.260 ;
        RECT 99.850 171.560 99.990 172.600 ;
        RECT 99.790 171.240 100.050 171.560 ;
        RECT 99.330 170.220 99.590 170.540 ;
        RECT 100.310 170.280 100.450 172.600 ;
        RECT 100.310 170.140 100.910 170.280 ;
        RECT 98.870 167.500 99.130 167.820 ;
        RECT 99.790 167.500 100.050 167.820 ;
        RECT 100.250 167.500 100.510 167.820 ;
        RECT 100.770 167.730 100.910 170.140 ;
        RECT 101.230 168.500 101.370 176.000 ;
        RECT 101.690 175.835 101.830 176.000 ;
        RECT 101.620 175.465 101.900 175.835 ;
        RECT 101.630 175.210 101.890 175.300 ;
        RECT 102.150 175.210 102.290 176.000 ;
        RECT 101.630 175.070 102.290 175.210 ;
        RECT 101.630 174.980 101.890 175.070 ;
        RECT 102.150 173.260 102.290 175.070 ;
        RECT 102.610 174.280 102.750 176.680 ;
        RECT 102.550 173.960 102.810 174.280 ;
        RECT 103.000 174.105 103.280 174.475 ;
        RECT 103.010 173.960 103.270 174.105 ;
        RECT 103.530 173.600 103.670 180.760 ;
        RECT 103.930 180.420 104.190 180.740 ;
        RECT 103.470 173.510 103.730 173.600 ;
        RECT 102.610 173.370 103.730 173.510 ;
        RECT 102.090 172.940 102.350 173.260 ;
        RECT 101.630 172.600 101.890 172.920 ;
        RECT 101.170 168.180 101.430 168.500 ;
        RECT 101.170 167.730 101.430 167.820 ;
        RECT 100.770 167.590 101.430 167.730 ;
        RECT 101.170 167.500 101.430 167.590 ;
        RECT 98.870 166.820 99.130 167.140 ;
        RECT 99.330 166.820 99.590 167.140 ;
        RECT 98.930 166.120 99.070 166.820 ;
        RECT 98.870 165.800 99.130 166.120 ;
        RECT 99.390 164.760 99.530 166.820 ;
        RECT 99.850 165.440 99.990 167.500 ;
        RECT 100.310 166.120 100.450 167.500 ;
        RECT 101.690 167.480 101.830 172.600 ;
        RECT 102.150 170.880 102.290 172.940 ;
        RECT 102.090 170.560 102.350 170.880 ;
        RECT 102.080 170.025 102.360 170.395 ;
        RECT 102.150 168.500 102.290 170.025 ;
        RECT 102.090 168.180 102.350 168.500 ;
        RECT 101.630 167.160 101.890 167.480 ;
        RECT 101.170 167.050 101.430 167.140 ;
        RECT 100.770 166.910 101.430 167.050 ;
        RECT 100.250 165.800 100.510 166.120 ;
        RECT 99.790 165.120 100.050 165.440 ;
        RECT 99.330 164.440 99.590 164.760 ;
        RECT 98.410 164.100 98.670 164.420 ;
        RECT 98.470 163.400 98.610 164.100 ;
        RECT 98.410 163.080 98.670 163.400 ;
        RECT 97.550 157.960 97.690 160.020 ;
        RECT 98.010 159.940 99.070 160.080 ;
        RECT 98.410 159.340 98.670 159.660 ;
        RECT 97.030 157.640 97.290 157.960 ;
        RECT 97.490 157.870 97.750 157.960 ;
        RECT 97.490 157.730 98.150 157.870 ;
        RECT 97.490 157.640 97.750 157.730 ;
        RECT 94.330 147.700 94.930 147.840 ;
        RECT 95.250 155.860 96.310 156.000 ;
        RECT 93.810 146.080 94.070 146.400 ;
        RECT 93.810 140.980 94.070 141.300 ;
        RECT 93.870 135.715 94.010 140.980 ;
        RECT 94.330 138.580 94.470 147.700 ;
        RECT 95.250 145.800 95.390 155.860 ;
        RECT 97.090 152.600 97.230 157.640 ;
        RECT 98.010 157.280 98.150 157.730 ;
        RECT 97.950 156.960 98.210 157.280 ;
        RECT 98.010 155.240 98.150 156.960 ;
        RECT 97.950 154.920 98.210 155.240 ;
        RECT 97.090 152.460 97.690 152.600 ;
        RECT 97.030 151.860 97.290 152.180 ;
        RECT 96.570 150.500 96.830 150.820 ;
        RECT 96.110 149.140 96.370 149.460 ;
        RECT 95.650 148.460 95.910 148.780 ;
        RECT 95.710 146.060 95.850 148.460 ;
        RECT 94.790 145.660 95.390 145.800 ;
        RECT 95.650 145.740 95.910 146.060 ;
        RECT 94.790 140.360 94.930 145.660 ;
        RECT 95.190 143.360 95.450 143.680 ;
        RECT 95.250 141.640 95.390 143.360 ;
        RECT 95.190 141.320 95.450 141.640 ;
        RECT 96.170 140.620 96.310 149.140 ;
        RECT 96.630 146.060 96.770 150.500 ;
        RECT 97.090 146.400 97.230 151.860 ;
        RECT 97.030 146.080 97.290 146.400 ;
        RECT 96.570 145.740 96.830 146.060 ;
        RECT 94.790 140.220 95.390 140.360 ;
        RECT 96.110 140.300 96.370 140.620 ;
        RECT 94.730 139.620 94.990 139.940 ;
        RECT 94.270 138.260 94.530 138.580 ;
        RECT 93.800 135.345 94.080 135.715 ;
        RECT 94.330 135.180 94.470 138.260 ;
        RECT 94.270 134.860 94.530 135.180 ;
        RECT 92.950 133.960 93.550 134.100 ;
        RECT 92.950 129.740 93.090 133.960 ;
        RECT 94.790 130.420 94.930 139.620 ;
        RECT 95.250 138.920 95.390 140.220 ;
        RECT 95.650 139.960 95.910 140.280 ;
        RECT 95.710 139.680 95.850 139.960 ;
        RECT 96.630 139.940 96.770 145.740 ;
        RECT 97.090 144.360 97.230 146.080 ;
        RECT 97.030 144.040 97.290 144.360 ;
        RECT 97.030 143.195 97.290 143.340 ;
        RECT 97.020 142.825 97.300 143.195 ;
        RECT 96.100 139.680 96.380 139.795 ;
        RECT 95.710 139.540 96.380 139.680 ;
        RECT 96.570 139.620 96.830 139.940 ;
        RECT 96.100 139.425 96.380 139.540 ;
        RECT 95.190 138.600 95.450 138.920 ;
        RECT 97.550 138.580 97.690 152.460 ;
        RECT 97.950 146.080 98.210 146.400 ;
        RECT 98.010 145.720 98.150 146.080 ;
        RECT 97.950 145.400 98.210 145.720 ;
        RECT 98.010 143.680 98.150 145.400 ;
        RECT 97.950 143.360 98.210 143.680 ;
        RECT 98.470 143.340 98.610 159.340 ;
        RECT 98.930 150.820 99.070 159.940 ;
        RECT 99.850 156.260 99.990 165.120 ;
        RECT 100.240 164.585 100.520 164.955 ;
        RECT 100.310 164.420 100.450 164.585 ;
        RECT 100.250 164.100 100.510 164.420 ;
        RECT 100.770 162.040 100.910 166.910 ;
        RECT 101.170 166.820 101.430 166.910 ;
        RECT 101.690 166.030 101.830 167.160 ;
        RECT 102.610 167.140 102.750 173.370 ;
        RECT 103.470 173.280 103.730 173.370 ;
        RECT 103.990 173.000 104.130 180.420 ;
        RECT 104.450 179.720 104.590 181.440 ;
        RECT 106.750 180.740 106.890 181.700 ;
        RECT 107.150 181.100 107.410 181.420 ;
        RECT 106.690 180.420 106.950 180.740 ;
        RECT 104.770 179.885 106.650 180.255 ;
        RECT 107.210 179.720 107.350 181.100 ;
        RECT 108.530 180.760 108.790 181.080 ;
        RECT 107.610 180.420 107.870 180.740 ;
        RECT 104.390 179.400 104.650 179.720 ;
        RECT 107.150 179.400 107.410 179.720 ;
        RECT 104.380 178.865 104.660 179.235 ;
        RECT 106.220 178.865 106.500 179.235 ;
        RECT 104.450 173.680 104.590 178.865 ;
        RECT 106.290 178.700 106.430 178.865 ;
        RECT 106.230 178.380 106.490 178.700 ;
        RECT 106.690 178.380 106.950 178.700 ;
        RECT 104.850 177.700 105.110 178.020 ;
        RECT 104.910 176.320 105.050 177.700 ;
        RECT 104.850 176.000 105.110 176.320 ;
        RECT 106.750 176.230 106.890 178.380 ;
        RECT 107.670 177.000 107.810 180.420 ;
        RECT 108.070 178.380 108.330 178.700 ;
        RECT 108.130 177.000 108.270 178.380 ;
        RECT 107.610 176.680 107.870 177.000 ;
        RECT 108.070 176.680 108.330 177.000 ;
        RECT 106.750 176.090 107.810 176.230 ;
        RECT 108.060 176.145 108.340 176.515 ;
        RECT 107.670 175.720 107.810 176.090 ;
        RECT 108.070 176.000 108.330 176.145 ;
        RECT 108.590 175.980 108.730 180.760 ;
        RECT 107.670 175.580 108.270 175.720 ;
        RECT 108.530 175.660 108.790 175.980 ;
        RECT 104.770 174.445 106.650 174.815 ;
        RECT 108.130 174.280 108.270 175.580 ;
        RECT 108.520 174.785 108.800 175.155 ;
        RECT 108.070 173.960 108.330 174.280 ;
        RECT 104.450 173.540 106.890 173.680 ;
        RECT 107.610 173.620 107.870 173.940 ;
        RECT 103.070 172.860 104.130 173.000 ;
        RECT 105.310 172.940 105.570 173.260 ;
        RECT 102.550 166.820 102.810 167.140 ;
        RECT 101.230 165.890 101.830 166.030 ;
        RECT 101.230 165.100 101.370 165.890 ;
        RECT 101.630 165.120 101.890 165.440 ;
        RECT 102.090 165.120 102.350 165.440 ;
        RECT 102.550 165.120 102.810 165.440 ;
        RECT 101.170 164.780 101.430 165.100 ;
        RECT 101.690 162.915 101.830 165.120 ;
        RECT 102.150 163.400 102.290 165.120 ;
        RECT 102.610 163.400 102.750 165.120 ;
        RECT 102.090 163.080 102.350 163.400 ;
        RECT 102.550 163.080 102.810 163.400 ;
        RECT 101.620 162.545 101.900 162.915 ;
        RECT 103.070 162.800 103.210 172.860 ;
        RECT 104.850 172.600 105.110 172.920 ;
        RECT 103.470 172.260 103.730 172.580 ;
        RECT 103.530 169.860 103.670 172.260 ;
        RECT 103.930 170.560 104.190 170.880 ;
        RECT 103.470 169.540 103.730 169.860 ;
        RECT 103.990 168.920 104.130 170.560 ;
        RECT 104.910 169.770 105.050 172.600 ;
        RECT 105.370 171.220 105.510 172.940 ;
        RECT 106.230 172.260 106.490 172.580 ;
        RECT 105.310 170.900 105.570 171.220 ;
        RECT 106.290 170.395 106.430 172.260 ;
        RECT 106.750 170.450 106.890 173.540 ;
        RECT 106.220 170.025 106.500 170.395 ;
        RECT 106.750 170.310 107.350 170.450 ;
        RECT 103.530 168.780 104.130 168.920 ;
        RECT 104.450 169.630 105.050 169.770 ;
        RECT 103.530 164.760 103.670 168.780 ;
        RECT 103.930 168.180 104.190 168.500 ;
        RECT 103.470 164.440 103.730 164.760 ;
        RECT 102.610 162.660 103.210 162.800 ;
        RECT 101.630 162.400 101.890 162.545 ;
        RECT 100.710 161.720 100.970 162.040 ;
        RECT 100.710 158.660 100.970 158.980 ;
        RECT 100.250 157.640 100.510 157.960 ;
        RECT 99.790 155.940 100.050 156.260 ;
        RECT 100.310 152.520 100.450 157.640 ;
        RECT 100.770 157.280 100.910 158.660 ;
        RECT 100.710 156.960 100.970 157.280 ;
        RECT 102.090 156.620 102.350 156.940 ;
        RECT 100.710 153.220 100.970 153.540 ;
        RECT 100.250 152.200 100.510 152.520 ;
        RECT 99.330 151.860 99.590 152.180 ;
        RECT 98.870 150.500 99.130 150.820 ;
        RECT 98.930 148.780 99.070 150.500 ;
        RECT 98.870 148.460 99.130 148.780 ;
        RECT 98.870 147.780 99.130 148.100 ;
        RECT 98.410 143.020 98.670 143.340 ;
        RECT 97.950 140.300 98.210 140.620 ;
        RECT 98.010 138.920 98.150 140.300 ;
        RECT 97.950 138.600 98.210 138.920 ;
        RECT 97.490 138.490 97.750 138.580 ;
        RECT 97.090 138.350 97.750 138.490 ;
        RECT 96.570 135.600 96.830 135.860 ;
        RECT 97.090 135.600 97.230 138.350 ;
        RECT 97.490 138.260 97.750 138.350 ;
        RECT 98.470 137.900 98.610 143.020 ;
        RECT 98.930 138.150 99.070 147.780 ;
        RECT 99.390 146.400 99.530 151.860 ;
        RECT 100.770 149.120 100.910 153.220 ;
        RECT 102.150 151.840 102.290 156.620 ;
        RECT 102.090 151.520 102.350 151.840 ;
        RECT 102.610 151.240 102.750 162.660 ;
        RECT 103.010 162.060 103.270 162.380 ;
        RECT 103.070 160.680 103.210 162.060 ;
        RECT 103.010 160.360 103.270 160.680 ;
        RECT 103.530 159.320 103.670 164.440 ;
        RECT 103.470 159.000 103.730 159.320 ;
        RECT 103.990 156.680 104.130 168.180 ;
        RECT 104.450 167.140 104.590 169.630 ;
        RECT 104.770 169.005 106.650 169.375 ;
        RECT 104.390 166.820 104.650 167.140 ;
        RECT 104.450 165.780 104.590 166.820 ;
        RECT 104.390 165.460 104.650 165.780 ;
        RECT 107.210 165.440 107.350 170.310 ;
        RECT 107.670 169.860 107.810 173.620 ;
        RECT 107.610 169.540 107.870 169.860 ;
        RECT 108.130 168.600 108.270 173.960 ;
        RECT 108.590 173.600 108.730 174.785 ;
        RECT 108.530 173.280 108.790 173.600 ;
        RECT 108.530 170.220 108.790 170.540 ;
        RECT 107.670 168.460 108.270 168.600 ;
        RECT 107.150 165.120 107.410 165.440 ;
        RECT 104.390 164.780 104.650 165.100 ;
        RECT 104.450 161.950 104.590 164.780 ;
        RECT 104.770 163.565 106.650 163.935 ;
        RECT 107.210 163.400 107.350 165.120 ;
        RECT 107.150 163.080 107.410 163.400 ;
        RECT 104.840 162.545 105.120 162.915 ;
        RECT 104.850 162.400 105.110 162.545 ;
        RECT 105.310 162.235 105.570 162.380 ;
        RECT 104.850 161.950 105.110 162.040 ;
        RECT 104.450 161.810 105.110 161.950 ;
        RECT 105.300 161.865 105.580 162.235 ;
        RECT 107.150 162.060 107.410 162.380 ;
        RECT 104.850 161.720 105.110 161.810 ;
        RECT 104.770 158.125 106.650 158.495 ;
        RECT 103.070 156.540 104.130 156.680 ;
        RECT 103.070 154.900 103.210 156.540 ;
        RECT 105.300 156.425 105.580 156.795 ;
        RECT 103.470 155.940 103.730 156.260 ;
        RECT 103.010 154.580 103.270 154.900 ;
        RECT 103.530 154.220 103.670 155.940 ;
        RECT 103.930 154.580 104.190 154.900 ;
        RECT 103.010 153.900 103.270 154.220 ;
        RECT 103.470 153.900 103.730 154.220 ;
        RECT 103.070 152.520 103.210 153.900 ;
        RECT 103.010 152.200 103.270 152.520 ;
        RECT 103.530 151.840 103.670 153.900 ;
        RECT 103.470 151.520 103.730 151.840 ;
        RECT 103.990 151.500 104.130 154.580 ;
        RECT 104.390 154.240 104.650 154.560 ;
        RECT 102.150 151.100 102.750 151.240 ;
        RECT 103.930 151.180 104.190 151.500 ;
        RECT 102.150 149.200 102.290 151.100 ;
        RECT 103.010 150.840 103.270 151.160 ;
        RECT 99.790 148.800 100.050 149.120 ;
        RECT 100.710 148.800 100.970 149.120 ;
        RECT 101.690 149.060 102.290 149.200 ;
        RECT 103.070 149.120 103.210 150.840 ;
        RECT 103.930 150.500 104.190 150.820 ;
        RECT 103.470 149.480 103.730 149.800 ;
        RECT 99.850 146.400 99.990 148.800 ;
        RECT 100.250 147.780 100.510 148.100 ;
        RECT 99.330 146.080 99.590 146.400 ;
        RECT 99.790 146.080 100.050 146.400 ;
        RECT 99.330 142.340 99.590 142.660 ;
        RECT 99.390 140.620 99.530 142.340 ;
        RECT 99.330 140.300 99.590 140.620 ;
        RECT 99.790 139.620 100.050 139.940 ;
        RECT 98.930 138.010 99.530 138.150 ;
        RECT 98.410 137.580 98.670 137.900 ;
        RECT 97.950 136.900 98.210 137.220 ;
        RECT 96.570 135.540 97.690 135.600 ;
        RECT 96.630 135.460 97.690 135.540 ;
        RECT 97.550 135.180 97.690 135.460 ;
        RECT 98.010 135.180 98.150 136.900 ;
        RECT 99.390 135.180 99.530 138.010 ;
        RECT 99.850 135.180 99.990 139.620 ;
        RECT 96.570 134.860 96.830 135.180 ;
        RECT 97.490 134.860 97.750 135.180 ;
        RECT 97.950 134.860 98.210 135.180 ;
        RECT 99.330 134.860 99.590 135.180 ;
        RECT 99.790 134.860 100.050 135.180 ;
        RECT 96.630 132.120 96.770 134.860 ;
        RECT 98.870 134.180 99.130 134.500 ;
        RECT 97.020 133.305 97.300 133.675 ;
        RECT 97.030 133.160 97.290 133.305 ;
        RECT 96.570 131.800 96.830 132.120 ;
        RECT 95.650 131.460 95.910 131.780 ;
        RECT 94.730 130.100 94.990 130.420 ;
        RECT 92.890 129.595 93.150 129.740 ;
        RECT 92.880 129.225 93.160 129.595 ;
        RECT 92.430 128.740 92.690 129.060 ;
        RECT 91.970 127.720 92.230 128.040 ;
        RECT 92.490 127.700 92.630 128.740 ;
        RECT 88.290 127.040 88.550 127.185 ;
        RECT 89.210 127.040 89.470 127.360 ;
        RECT 91.960 127.185 92.240 127.555 ;
        RECT 92.430 127.380 92.690 127.700 ;
        RECT 95.710 127.360 95.850 131.460 ;
        RECT 97.090 128.040 97.230 133.160 ;
        RECT 98.930 132.800 99.070 134.180 ;
        RECT 97.950 132.480 98.210 132.800 ;
        RECT 98.870 132.480 99.130 132.800 ;
        RECT 97.490 129.760 97.750 130.080 ;
        RECT 97.030 127.720 97.290 128.040 ;
        RECT 97.550 127.360 97.690 129.760 ;
        RECT 98.010 129.740 98.150 132.480 ;
        RECT 98.400 131.945 98.680 132.315 ;
        RECT 98.470 130.760 98.610 131.945 ;
        RECT 98.410 130.440 98.670 130.760 ;
        RECT 100.310 130.420 100.450 147.780 ;
        RECT 100.710 146.420 100.970 146.740 ;
        RECT 100.770 143.680 100.910 146.420 ;
        RECT 100.710 143.360 100.970 143.680 ;
        RECT 101.170 142.680 101.430 143.000 ;
        RECT 100.710 141.155 100.970 141.300 ;
        RECT 100.700 140.785 100.980 141.155 ;
        RECT 100.710 137.920 100.970 138.240 ;
        RECT 100.770 135.860 100.910 137.920 ;
        RECT 100.710 135.540 100.970 135.860 ;
        RECT 100.250 130.100 100.510 130.420 ;
        RECT 97.950 129.420 98.210 129.740 ;
        RECT 99.780 127.865 100.060 128.235 ;
        RECT 99.850 127.360 99.990 127.865 ;
        RECT 91.970 127.040 92.230 127.185 ;
        RECT 95.650 127.040 95.910 127.360 ;
        RECT 97.490 127.040 97.750 127.360 ;
        RECT 99.790 127.040 100.050 127.360 ;
        RECT 88.350 126.760 88.490 127.040 ;
        RECT 101.230 127.020 101.370 142.680 ;
        RECT 101.690 139.850 101.830 149.060 ;
        RECT 103.010 148.800 103.270 149.120 ;
        RECT 102.090 148.460 102.350 148.780 ;
        RECT 102.150 147.080 102.290 148.460 ;
        RECT 102.090 146.760 102.350 147.080 ;
        RECT 102.550 145.060 102.810 145.380 ;
        RECT 102.610 143.080 102.750 145.060 ;
        RECT 103.000 143.505 103.280 143.875 ;
        RECT 103.070 143.340 103.210 143.505 ;
        RECT 102.150 142.940 102.750 143.080 ;
        RECT 103.010 143.020 103.270 143.340 ;
        RECT 102.150 140.960 102.290 142.940 ;
        RECT 102.550 142.340 102.810 142.660 ;
        RECT 102.090 140.640 102.350 140.960 ;
        RECT 102.610 140.620 102.750 142.340 ;
        RECT 102.550 140.300 102.810 140.620 ;
        RECT 101.690 139.710 102.750 139.850 ;
        RECT 102.090 136.900 102.350 137.220 ;
        RECT 102.150 136.200 102.290 136.900 ;
        RECT 102.090 136.110 102.350 136.200 ;
        RECT 101.690 135.970 102.350 136.110 ;
        RECT 101.690 130.080 101.830 135.970 ;
        RECT 102.090 135.880 102.350 135.970 ;
        RECT 102.090 132.140 102.350 132.460 ;
        RECT 101.630 129.760 101.890 130.080 ;
        RECT 84.150 126.360 84.410 126.680 ;
        RECT 86.050 126.340 86.190 126.700 ;
        RECT 87.430 126.620 88.490 126.760 ;
        RECT 101.170 126.700 101.430 127.020 ;
        RECT 102.150 126.340 102.290 132.140 ;
        RECT 102.610 128.040 102.750 139.710 ;
        RECT 103.530 138.830 103.670 149.480 ;
        RECT 103.990 143.680 104.130 150.500 ;
        RECT 104.450 149.800 104.590 154.240 ;
        RECT 105.370 154.220 105.510 156.425 ;
        RECT 105.310 153.900 105.570 154.220 ;
        RECT 106.690 154.075 106.950 154.220 ;
        RECT 106.680 153.705 106.960 154.075 ;
        RECT 104.770 152.685 106.650 153.055 ;
        RECT 104.850 151.180 105.110 151.500 ;
        RECT 104.910 149.800 105.050 151.180 ;
        RECT 104.390 149.480 104.650 149.800 ;
        RECT 104.850 149.480 105.110 149.800 ;
        RECT 104.390 148.460 104.650 148.780 ;
        RECT 104.450 145.970 104.590 148.460 ;
        RECT 104.770 147.245 106.650 147.615 ;
        RECT 104.850 145.970 105.110 146.060 ;
        RECT 104.450 145.830 105.110 145.970 ;
        RECT 105.770 145.915 106.030 146.060 ;
        RECT 104.850 145.740 105.110 145.830 ;
        RECT 105.760 145.545 106.040 145.915 ;
        RECT 104.390 145.060 104.650 145.380 ;
        RECT 107.210 145.120 107.350 162.060 ;
        RECT 107.670 157.620 107.810 168.460 ;
        RECT 108.590 168.355 108.730 170.220 ;
        RECT 108.520 167.985 108.800 168.355 ;
        RECT 108.530 162.060 108.790 162.380 ;
        RECT 108.070 161.720 108.330 162.040 ;
        RECT 108.130 160.000 108.270 161.720 ;
        RECT 108.590 160.340 108.730 162.060 ;
        RECT 108.530 160.020 108.790 160.340 ;
        RECT 108.070 159.680 108.330 160.000 ;
        RECT 107.610 157.300 107.870 157.620 ;
        RECT 108.530 156.620 108.790 156.940 ;
        RECT 108.590 154.900 108.730 156.620 ;
        RECT 108.530 154.580 108.790 154.900 ;
        RECT 107.610 153.960 107.870 154.220 ;
        RECT 107.610 153.900 108.270 153.960 ;
        RECT 107.670 153.820 108.270 153.900 ;
        RECT 107.610 153.220 107.870 153.540 ;
        RECT 107.670 145.915 107.810 153.220 ;
        RECT 108.130 150.820 108.270 153.820 ;
        RECT 108.530 151.180 108.790 151.500 ;
        RECT 108.070 150.500 108.330 150.820 ;
        RECT 108.590 147.080 108.730 151.180 ;
        RECT 108.530 146.760 108.790 147.080 ;
        RECT 108.070 146.080 108.330 146.400 ;
        RECT 107.600 145.545 107.880 145.915 ;
        RECT 104.450 144.360 104.590 145.060 ;
        RECT 105.830 144.980 107.350 145.120 ;
        RECT 104.390 144.040 104.650 144.360 ;
        RECT 105.830 143.680 105.970 144.980 ;
        RECT 107.600 144.185 107.880 144.555 ;
        RECT 103.930 143.360 104.190 143.680 ;
        RECT 104.390 143.360 104.650 143.680 ;
        RECT 105.770 143.360 106.030 143.680 ;
        RECT 103.990 141.640 104.130 143.360 ;
        RECT 103.930 141.320 104.190 141.640 ;
        RECT 103.930 139.620 104.190 139.940 ;
        RECT 103.070 138.690 103.670 138.830 ;
        RECT 103.070 136.200 103.210 138.690 ;
        RECT 103.470 137.920 103.730 138.240 ;
        RECT 103.530 137.560 103.670 137.920 ;
        RECT 103.470 137.240 103.730 137.560 ;
        RECT 103.010 135.880 103.270 136.200 ;
        RECT 103.530 135.180 103.670 137.240 ;
        RECT 103.470 134.860 103.730 135.180 ;
        RECT 103.010 134.180 103.270 134.500 ;
        RECT 103.070 132.120 103.210 134.180 ;
        RECT 103.530 133.140 103.670 134.860 ;
        RECT 103.470 132.820 103.730 133.140 ;
        RECT 103.010 131.800 103.270 132.120 ;
        RECT 103.010 129.420 103.270 129.740 ;
        RECT 103.070 128.040 103.210 129.420 ;
        RECT 102.550 127.720 102.810 128.040 ;
        RECT 103.010 127.720 103.270 128.040 ;
        RECT 103.530 127.360 103.670 132.820 ;
        RECT 103.990 129.400 104.130 139.620 ;
        RECT 104.450 136.200 104.590 143.360 ;
        RECT 104.770 141.805 106.650 142.175 ;
        RECT 106.690 140.475 106.950 140.620 ;
        RECT 106.680 140.105 106.960 140.475 ;
        RECT 107.150 136.900 107.410 137.220 ;
        RECT 104.770 136.365 106.650 136.735 ;
        RECT 107.210 136.200 107.350 136.900 ;
        RECT 104.390 135.880 104.650 136.200 ;
        RECT 107.150 135.880 107.410 136.200 ;
        RECT 107.140 135.345 107.420 135.715 ;
        RECT 107.210 135.180 107.350 135.345 ;
        RECT 104.390 134.860 104.650 135.180 ;
        RECT 104.450 132.800 104.590 134.860 ;
        RECT 106.220 134.665 106.500 135.035 ;
        RECT 107.150 134.860 107.410 135.180 ;
        RECT 106.290 133.140 106.430 134.665 ;
        RECT 106.230 132.820 106.490 133.140 ;
        RECT 104.390 132.480 104.650 132.800 ;
        RECT 104.390 131.460 104.650 131.780 ;
        RECT 104.450 130.080 104.590 131.460 ;
        RECT 104.770 130.925 106.650 131.295 ;
        RECT 105.770 130.100 106.030 130.420 ;
        RECT 104.390 129.760 104.650 130.080 ;
        RECT 103.930 129.080 104.190 129.400 ;
        RECT 105.830 127.360 105.970 130.100 ;
        RECT 107.210 129.740 107.350 134.860 ;
        RECT 106.230 129.420 106.490 129.740 ;
        RECT 107.150 129.420 107.410 129.740 ;
        RECT 106.290 128.040 106.430 129.420 ;
        RECT 106.230 127.720 106.490 128.040 ;
        RECT 107.150 127.950 107.410 128.040 ;
        RECT 107.670 127.950 107.810 144.185 ;
        RECT 108.130 143.680 108.270 146.080 ;
        RECT 108.530 145.400 108.790 145.720 ;
        RECT 108.070 143.360 108.330 143.680 ;
        RECT 108.130 141.300 108.270 143.360 ;
        RECT 108.590 143.340 108.730 145.400 ;
        RECT 109.050 145.235 109.190 189.600 ;
        RECT 109.910 188.580 110.170 188.900 ;
        RECT 109.970 187.540 110.110 188.580 ;
        RECT 109.910 187.220 110.170 187.540 ;
        RECT 109.970 185.160 110.110 187.220 ;
        RECT 109.910 184.840 110.170 185.160 ;
        RECT 109.910 183.820 110.170 184.140 ;
        RECT 109.450 183.480 109.710 183.800 ;
        RECT 109.510 182.100 109.650 183.480 ;
        RECT 109.970 182.440 110.110 183.820 ;
        RECT 109.910 182.120 110.170 182.440 ;
        RECT 109.450 181.780 109.710 182.100 ;
        RECT 109.450 181.100 109.710 181.420 ;
        RECT 110.430 181.330 110.570 199.460 ;
        RECT 111.750 197.760 112.010 198.080 ;
        RECT 110.830 196.740 111.090 197.060 ;
        RECT 110.890 196.040 111.030 196.740 ;
        RECT 111.810 196.040 111.950 197.760 ;
        RECT 112.270 197.060 112.410 199.800 ;
        RECT 112.670 199.460 112.930 199.780 ;
        RECT 112.210 196.740 112.470 197.060 ;
        RECT 110.830 195.720 111.090 196.040 ;
        RECT 111.750 195.720 112.010 196.040 ;
        RECT 110.830 194.700 111.090 195.020 ;
        RECT 112.210 194.700 112.470 195.020 ;
        RECT 110.890 193.320 111.030 194.700 ;
        RECT 110.830 193.000 111.090 193.320 ;
        RECT 111.750 193.000 112.010 193.320 ;
        RECT 111.290 192.210 111.550 192.300 ;
        RECT 110.890 192.070 111.550 192.210 ;
        RECT 110.890 187.200 111.030 192.070 ;
        RECT 111.290 191.980 111.550 192.070 ;
        RECT 111.280 191.105 111.560 191.475 ;
        RECT 111.350 187.395 111.490 191.105 ;
        RECT 111.810 190.510 111.950 193.000 ;
        RECT 112.270 192.300 112.410 194.700 ;
        RECT 112.210 191.980 112.470 192.300 ;
        RECT 111.810 190.370 112.410 190.510 ;
        RECT 111.750 189.600 112.010 189.920 ;
        RECT 111.810 188.900 111.950 189.600 ;
        RECT 111.750 188.580 112.010 188.900 ;
        RECT 110.830 186.880 111.090 187.200 ;
        RECT 111.280 187.025 111.560 187.395 ;
        RECT 112.270 187.280 112.410 190.370 ;
        RECT 111.810 187.140 112.410 187.280 ;
        RECT 111.290 186.880 111.550 187.025 ;
        RECT 111.280 185.920 111.560 186.035 ;
        RECT 110.890 185.780 111.560 185.920 ;
        RECT 110.890 181.670 111.030 185.780 ;
        RECT 111.280 185.665 111.560 185.780 ;
        RECT 111.280 183.625 111.560 183.995 ;
        RECT 111.350 183.460 111.490 183.625 ;
        RECT 111.290 183.140 111.550 183.460 ;
        RECT 110.890 181.530 111.490 181.670 ;
        RECT 109.970 181.190 110.570 181.330 ;
        RECT 109.510 180.595 109.650 181.100 ;
        RECT 109.440 180.225 109.720 180.595 ;
        RECT 109.970 177.930 110.110 181.190 ;
        RECT 110.830 180.760 111.090 181.080 ;
        RECT 110.370 180.420 110.630 180.740 ;
        RECT 109.510 177.790 110.110 177.930 ;
        RECT 109.510 160.340 109.650 177.790 ;
        RECT 109.910 176.680 110.170 177.000 ;
        RECT 109.450 160.020 109.710 160.340 ;
        RECT 109.970 154.470 110.110 176.680 ;
        RECT 110.430 172.580 110.570 180.420 ;
        RECT 110.890 177.000 111.030 180.760 ;
        RECT 110.830 176.680 111.090 177.000 ;
        RECT 110.830 175.320 111.090 175.640 ;
        RECT 110.890 173.940 111.030 175.320 ;
        RECT 110.830 173.620 111.090 173.940 ;
        RECT 110.370 172.435 110.630 172.580 ;
        RECT 110.360 172.065 110.640 172.435 ;
        RECT 110.830 172.260 111.090 172.580 ;
        RECT 110.890 170.540 111.030 172.260 ;
        RECT 110.830 170.220 111.090 170.540 ;
        RECT 110.370 164.440 110.630 164.760 ;
        RECT 110.430 162.915 110.570 164.440 ;
        RECT 110.360 162.545 110.640 162.915 ;
        RECT 110.430 159.515 110.570 162.545 ;
        RECT 110.360 159.145 110.640 159.515 ;
        RECT 110.370 158.660 110.630 158.980 ;
        RECT 109.510 154.330 110.110 154.470 ;
        RECT 108.980 144.865 109.260 145.235 ;
        RECT 108.530 143.020 108.790 143.340 ;
        RECT 108.070 140.980 108.330 141.300 ;
        RECT 108.530 140.640 108.790 140.960 ;
        RECT 108.590 138.920 108.730 140.640 ;
        RECT 108.530 138.600 108.790 138.920 ;
        RECT 108.070 134.860 108.330 135.180 ;
        RECT 108.130 134.500 108.270 134.860 ;
        RECT 108.070 134.180 108.330 134.500 ;
        RECT 108.530 134.180 108.790 134.500 ;
        RECT 108.070 131.800 108.330 132.120 ;
        RECT 108.130 129.740 108.270 131.800 ;
        RECT 108.070 129.420 108.330 129.740 ;
        RECT 107.150 127.810 107.810 127.950 ;
        RECT 108.060 127.865 108.340 128.235 ;
        RECT 108.590 128.040 108.730 134.180 ;
        RECT 109.510 133.140 109.650 154.330 ;
        RECT 110.430 153.960 110.570 158.660 ;
        RECT 110.830 155.940 111.090 156.260 ;
        RECT 110.890 154.900 111.030 155.940 ;
        RECT 110.830 154.580 111.090 154.900 ;
        RECT 109.970 153.820 110.570 153.960 ;
        RECT 110.830 153.900 111.090 154.220 ;
        RECT 109.970 151.355 110.110 153.820 ;
        RECT 110.370 153.220 110.630 153.540 ;
        RECT 109.900 150.985 110.180 151.355 ;
        RECT 109.910 149.480 110.170 149.800 ;
        RECT 109.970 147.955 110.110 149.480 ;
        RECT 110.430 148.010 110.570 153.220 ;
        RECT 110.890 152.520 111.030 153.900 ;
        RECT 110.830 152.200 111.090 152.520 ;
        RECT 111.350 151.920 111.490 181.530 ;
        RECT 110.890 151.780 111.490 151.920 ;
        RECT 110.890 148.780 111.030 151.780 ;
        RECT 111.290 151.180 111.550 151.500 ;
        RECT 110.830 148.460 111.090 148.780 ;
        RECT 111.350 148.440 111.490 151.180 ;
        RECT 111.290 148.120 111.550 148.440 ;
        RECT 109.900 147.585 110.180 147.955 ;
        RECT 110.430 147.870 111.030 148.010 ;
        RECT 110.890 147.840 111.030 147.870 ;
        RECT 110.890 147.700 111.490 147.840 ;
        RECT 110.820 146.905 111.100 147.275 ;
        RECT 110.830 146.760 111.090 146.905 ;
        RECT 111.350 146.595 111.490 147.700 ;
        RECT 111.810 146.740 111.950 187.140 ;
        RECT 112.730 181.080 112.870 199.460 ;
        RECT 114.110 198.160 114.250 202.180 ;
        RECT 115.030 200.460 115.170 203.460 ;
        RECT 115.890 203.200 116.150 203.520 ;
        RECT 118.190 203.200 118.450 203.520 ;
        RECT 115.950 201.480 116.090 203.200 ;
        RECT 116.350 202.180 116.610 202.500 ;
        RECT 115.890 201.160 116.150 201.480 ;
        RECT 114.970 200.140 115.230 200.460 ;
        RECT 116.410 200.120 116.550 202.180 ;
        RECT 114.510 199.800 114.770 200.120 ;
        RECT 116.350 199.800 116.610 200.120 ;
        RECT 114.570 198.760 114.710 199.800 ;
        RECT 114.510 198.440 114.770 198.760 ;
        RECT 114.110 198.020 115.630 198.160 ;
        RECT 118.250 198.080 118.390 203.200 ;
        RECT 121.930 201.480 122.070 205.580 ;
        RECT 123.250 204.900 123.510 205.220 ;
        RECT 123.310 203.520 123.450 204.900 ;
        RECT 123.250 203.200 123.510 203.520 ;
        RECT 121.870 201.160 122.130 201.480 ;
        RECT 123.710 200.820 123.970 201.140 ;
        RECT 122.790 200.140 123.050 200.460 ;
        RECT 121.870 199.460 122.130 199.780 ;
        RECT 119.770 198.925 121.650 199.295 ;
        RECT 113.590 197.650 113.850 197.740 ;
        RECT 113.190 197.510 113.850 197.650 ;
        RECT 112.670 180.760 112.930 181.080 ;
        RECT 113.190 180.480 113.330 197.510 ;
        RECT 113.590 197.420 113.850 197.510 ;
        RECT 114.500 195.185 114.780 195.555 ;
        RECT 114.050 193.000 114.310 193.320 ;
        RECT 113.590 192.320 113.850 192.640 ;
        RECT 113.650 189.240 113.790 192.320 ;
        RECT 114.110 190.600 114.250 193.000 ;
        RECT 114.050 190.280 114.310 190.600 ;
        RECT 113.590 188.920 113.850 189.240 ;
        RECT 113.590 187.560 113.850 187.880 ;
        RECT 113.650 186.035 113.790 187.560 ;
        RECT 113.580 185.665 113.860 186.035 ;
        RECT 113.590 183.140 113.850 183.460 ;
        RECT 112.270 180.340 113.330 180.480 ;
        RECT 111.280 146.225 111.560 146.595 ;
        RECT 111.750 146.420 112.010 146.740 ;
        RECT 109.910 145.740 110.170 146.060 ;
        RECT 110.370 145.915 110.630 146.060 ;
        RECT 109.970 138.580 110.110 145.740 ;
        RECT 110.360 145.545 110.640 145.915 ;
        RECT 111.290 145.740 111.550 146.060 ;
        RECT 110.370 145.060 110.630 145.380 ;
        RECT 110.430 144.360 110.570 145.060 ;
        RECT 111.350 144.360 111.490 145.740 ;
        RECT 110.370 144.040 110.630 144.360 ;
        RECT 111.290 144.040 111.550 144.360 ;
        RECT 110.360 143.505 110.640 143.875 ;
        RECT 110.370 143.360 110.630 143.505 ;
        RECT 110.360 142.825 110.640 143.195 ;
        RECT 110.430 141.300 110.570 142.825 ;
        RECT 110.370 140.980 110.630 141.300 ;
        RECT 109.910 138.260 110.170 138.580 ;
        RECT 112.270 134.100 112.410 180.340 ;
        RECT 113.650 179.800 113.790 183.140 ;
        RECT 114.570 181.760 114.710 195.185 ;
        RECT 115.490 192.640 115.630 198.020 ;
        RECT 118.190 197.760 118.450 198.080 ;
        RECT 119.110 197.760 119.370 198.080 ;
        RECT 119.170 197.480 119.310 197.760 ;
        RECT 117.730 197.310 117.990 197.400 ;
        RECT 118.250 197.340 119.310 197.480 ;
        RECT 118.250 197.310 118.390 197.340 ;
        RECT 117.730 197.170 118.390 197.310 ;
        RECT 117.730 197.080 117.990 197.170 ;
        RECT 118.650 196.740 118.910 197.060 ;
        RECT 118.190 195.040 118.450 195.360 ;
        RECT 115.890 194.700 116.150 195.020 ;
        RECT 115.430 192.320 115.690 192.640 ;
        RECT 115.490 189.580 115.630 192.320 ;
        RECT 115.950 189.580 116.090 194.700 ;
        RECT 117.270 194.020 117.530 194.340 ;
        RECT 117.330 191.960 117.470 194.020 ;
        RECT 117.730 192.320 117.990 192.640 ;
        RECT 116.810 191.640 117.070 191.960 ;
        RECT 117.270 191.640 117.530 191.960 ;
        RECT 115.430 189.260 115.690 189.580 ;
        RECT 115.890 189.260 116.150 189.580 ;
        RECT 116.350 188.920 116.610 189.240 ;
        RECT 116.410 188.755 116.550 188.920 ;
        RECT 116.340 188.385 116.620 188.755 ;
        RECT 115.880 187.705 116.160 188.075 ;
        RECT 115.950 187.540 116.090 187.705 ;
        RECT 115.890 187.220 116.150 187.540 ;
        RECT 114.970 186.880 115.230 187.200 ;
        RECT 115.030 183.800 115.170 186.880 ;
        RECT 115.430 184.840 115.690 185.160 ;
        RECT 114.970 183.480 115.230 183.800 ;
        RECT 115.490 183.460 115.630 184.840 ;
        RECT 115.950 184.140 116.090 187.220 ;
        RECT 116.870 186.860 117.010 191.640 ;
        RECT 117.270 188.580 117.530 188.900 ;
        RECT 116.810 186.540 117.070 186.860 ;
        RECT 116.350 186.200 116.610 186.520 ;
        RECT 116.410 185.160 116.550 186.200 ;
        RECT 116.350 184.840 116.610 185.160 ;
        RECT 116.870 184.480 117.010 186.540 ;
        RECT 117.330 186.180 117.470 188.580 ;
        RECT 117.270 185.860 117.530 186.180 ;
        RECT 116.810 184.160 117.070 184.480 ;
        RECT 115.890 183.820 116.150 184.140 ;
        RECT 117.790 183.800 117.930 192.320 ;
        RECT 118.250 189.240 118.390 195.040 ;
        RECT 118.190 188.920 118.450 189.240 ;
        RECT 118.250 187.880 118.390 188.920 ;
        RECT 118.190 187.560 118.450 187.880 ;
        RECT 118.250 187.395 118.390 187.560 ;
        RECT 118.180 187.025 118.460 187.395 ;
        RECT 117.730 183.480 117.990 183.800 ;
        RECT 115.430 183.140 115.690 183.460 ;
        RECT 118.710 182.400 118.850 196.740 ;
        RECT 119.770 193.485 121.650 193.855 ;
        RECT 120.480 192.465 120.760 192.835 ;
        RECT 119.110 188.580 119.370 188.900 ;
        RECT 120.550 188.810 120.690 192.465 ;
        RECT 120.950 192.320 121.210 192.640 ;
        RECT 121.010 192.155 121.150 192.320 ;
        RECT 120.940 191.785 121.220 192.155 ;
        RECT 120.950 191.300 121.210 191.620 ;
        RECT 121.010 190.600 121.150 191.300 ;
        RECT 120.950 190.280 121.210 190.600 ;
        RECT 120.950 188.810 121.210 188.900 ;
        RECT 120.550 188.670 121.210 188.810 ;
        RECT 120.950 188.580 121.210 188.670 ;
        RECT 119.170 187.540 119.310 188.580 ;
        RECT 119.770 188.045 121.650 188.415 ;
        RECT 119.110 187.220 119.370 187.540 ;
        RECT 120.950 186.880 121.210 187.200 ;
        RECT 119.110 186.200 119.370 186.520 ;
        RECT 119.560 186.345 119.840 186.715 ;
        RECT 119.570 186.200 119.830 186.345 ;
        RECT 117.330 182.260 118.850 182.400 ;
        RECT 114.510 181.440 114.770 181.760 ;
        RECT 114.970 180.760 115.230 181.080 ;
        RECT 114.500 180.225 114.780 180.595 ;
        RECT 112.730 179.660 113.790 179.800 ;
        RECT 112.730 166.200 112.870 179.660 ;
        RECT 114.570 179.380 114.710 180.225 ;
        RECT 115.030 179.720 115.170 180.760 ;
        RECT 114.970 179.400 115.230 179.720 ;
        RECT 114.510 179.060 114.770 179.380 ;
        RECT 114.960 179.120 115.240 179.235 ;
        RECT 114.960 178.980 115.630 179.120 ;
        RECT 114.960 178.865 115.240 178.980 ;
        RECT 115.490 178.700 115.630 178.980 ;
        RECT 113.130 178.380 113.390 178.700 ;
        RECT 114.970 178.380 115.230 178.700 ;
        RECT 115.430 178.380 115.690 178.700 ;
        RECT 113.190 177.000 113.330 178.380 ;
        RECT 113.590 178.040 113.850 178.360 ;
        RECT 113.130 176.680 113.390 177.000 ;
        RECT 113.120 174.785 113.400 175.155 ;
        RECT 113.190 173.940 113.330 174.785 ;
        RECT 113.130 173.620 113.390 173.940 ;
        RECT 113.130 172.600 113.390 172.920 ;
        RECT 113.190 167.820 113.330 172.600 ;
        RECT 113.650 171.560 113.790 178.040 ;
        RECT 114.050 176.000 114.310 176.320 ;
        RECT 113.590 171.240 113.850 171.560 ;
        RECT 114.110 170.880 114.250 176.000 ;
        RECT 114.510 175.660 114.770 175.980 ;
        RECT 114.050 170.560 114.310 170.880 ;
        RECT 113.590 170.280 113.850 170.540 ;
        RECT 114.570 170.280 114.710 175.660 ;
        RECT 115.030 174.280 115.170 178.380 ;
        RECT 115.890 178.040 116.150 178.360 ;
        RECT 115.950 177.000 116.090 178.040 ;
        RECT 116.350 177.700 116.610 178.020 ;
        RECT 115.890 176.680 116.150 177.000 ;
        RECT 115.890 174.980 116.150 175.300 ;
        RECT 115.950 174.280 116.090 174.980 ;
        RECT 114.970 173.960 115.230 174.280 ;
        RECT 115.890 173.960 116.150 174.280 ;
        RECT 116.410 172.435 116.550 177.700 ;
        RECT 116.800 176.145 117.080 176.515 ;
        RECT 116.340 172.065 116.620 172.435 ;
        RECT 116.870 171.640 117.010 176.145 ;
        RECT 115.950 171.500 117.010 171.640 ;
        RECT 115.950 170.960 116.090 171.500 ;
        RECT 113.590 170.220 114.710 170.280 ;
        RECT 113.650 170.140 114.710 170.220 ;
        RECT 115.490 170.820 116.090 170.960 ;
        RECT 113.650 168.500 113.790 170.140 ;
        RECT 113.590 168.180 113.850 168.500 ;
        RECT 114.510 167.840 114.770 168.160 ;
        RECT 113.130 167.500 113.390 167.820 ;
        RECT 114.570 167.140 114.710 167.840 ;
        RECT 114.510 166.820 114.770 167.140 ;
        RECT 112.730 166.060 113.330 166.200 ;
        RECT 112.670 165.635 112.930 165.780 ;
        RECT 112.660 165.265 112.940 165.635 ;
        RECT 113.190 160.080 113.330 166.060 ;
        RECT 113.590 165.460 113.850 165.780 ;
        RECT 113.650 162.380 113.790 165.460 ;
        RECT 114.510 165.120 114.770 165.440 ;
        RECT 114.570 163.400 114.710 165.120 ;
        RECT 114.510 163.080 114.770 163.400 ;
        RECT 113.590 162.060 113.850 162.380 ;
        RECT 112.730 159.940 113.330 160.080 ;
        RECT 114.050 160.020 114.310 160.340 ;
        RECT 112.730 152.715 112.870 159.940 ;
        RECT 114.110 156.940 114.250 160.020 ;
        RECT 115.490 157.960 115.630 170.820 ;
        RECT 116.340 170.705 116.620 171.075 ;
        RECT 116.410 170.280 116.550 170.705 ;
        RECT 116.810 170.560 117.070 170.880 ;
        RECT 115.950 170.140 116.550 170.280 ;
        RECT 115.430 157.640 115.690 157.960 ;
        RECT 115.950 157.475 116.090 170.140 ;
        RECT 116.350 169.540 116.610 169.860 ;
        RECT 116.410 164.420 116.550 169.540 ;
        RECT 116.870 168.840 117.010 170.560 ;
        RECT 116.810 168.520 117.070 168.840 ;
        RECT 116.810 167.500 117.070 167.820 ;
        RECT 116.870 165.635 117.010 167.500 ;
        RECT 116.800 165.265 117.080 165.635 ;
        RECT 116.810 164.780 117.070 165.100 ;
        RECT 116.350 164.100 116.610 164.420 ;
        RECT 116.410 162.720 116.550 164.100 ;
        RECT 116.870 163.400 117.010 164.780 ;
        RECT 116.810 163.080 117.070 163.400 ;
        RECT 116.350 162.400 116.610 162.720 ;
        RECT 116.350 157.640 116.610 157.960 ;
        RECT 115.880 157.105 116.160 157.475 ;
        RECT 113.590 156.795 113.850 156.940 ;
        RECT 114.050 156.850 114.310 156.940 ;
        RECT 113.580 156.425 113.860 156.795 ;
        RECT 114.050 156.710 115.170 156.850 ;
        RECT 114.050 156.620 114.310 156.710 ;
        RECT 113.130 155.940 113.390 156.260 ;
        RECT 113.590 155.940 113.850 156.260 ;
        RECT 114.510 155.940 114.770 156.260 ;
        RECT 113.190 155.240 113.330 155.940 ;
        RECT 113.130 154.920 113.390 155.240 ;
        RECT 113.650 154.560 113.790 155.940 ;
        RECT 113.590 154.240 113.850 154.560 ;
        RECT 112.660 152.345 112.940 152.715 ;
        RECT 113.650 152.520 113.790 154.240 ;
        RECT 114.050 153.900 114.310 154.220 ;
        RECT 113.590 152.200 113.850 152.520 ;
        RECT 112.670 151.860 112.930 152.180 ;
        RECT 112.730 148.440 112.870 151.860 ;
        RECT 113.580 151.665 113.860 152.035 ;
        RECT 113.120 150.985 113.400 151.355 ;
        RECT 112.670 148.120 112.930 148.440 ;
        RECT 112.660 147.585 112.940 147.955 ;
        RECT 112.730 137.560 112.870 147.585 ;
        RECT 113.190 146.060 113.330 150.985 ;
        RECT 113.130 145.740 113.390 146.060 ;
        RECT 113.130 143.020 113.390 143.340 ;
        RECT 113.190 141.155 113.330 143.020 ;
        RECT 113.120 140.785 113.400 141.155 ;
        RECT 113.130 140.300 113.390 140.620 ;
        RECT 112.670 137.240 112.930 137.560 ;
        RECT 113.190 136.200 113.330 140.300 ;
        RECT 113.650 139.795 113.790 151.665 ;
        RECT 114.110 148.100 114.250 153.900 ;
        RECT 114.050 147.780 114.310 148.100 ;
        RECT 114.110 140.280 114.250 147.780 ;
        RECT 114.050 139.960 114.310 140.280 ;
        RECT 113.580 139.425 113.860 139.795 ;
        RECT 113.650 138.920 113.790 139.425 ;
        RECT 113.590 138.600 113.850 138.920 ;
        RECT 114.050 138.260 114.310 138.580 ;
        RECT 114.110 136.200 114.250 138.260 ;
        RECT 113.130 135.880 113.390 136.200 ;
        RECT 114.050 135.880 114.310 136.200 ;
        RECT 111.350 133.960 112.870 134.100 ;
        RECT 111.350 133.480 111.490 133.960 ;
        RECT 111.290 133.160 111.550 133.480 ;
        RECT 108.990 132.820 109.250 133.140 ;
        RECT 109.450 132.820 109.710 133.140 ;
        RECT 109.050 130.080 109.190 132.820 ;
        RECT 109.510 130.420 109.650 132.820 ;
        RECT 112.210 131.460 112.470 131.780 ;
        RECT 109.450 130.100 109.710 130.420 ;
        RECT 111.290 130.100 111.550 130.420 ;
        RECT 108.990 129.760 109.250 130.080 ;
        RECT 110.820 129.225 111.100 129.595 ;
        RECT 110.890 129.060 111.030 129.225 ;
        RECT 111.350 129.060 111.490 130.100 ;
        RECT 112.270 129.740 112.410 131.460 ;
        RECT 112.730 130.080 112.870 133.960 ;
        RECT 113.120 132.625 113.400 132.995 ;
        RECT 114.570 132.800 114.710 155.940 ;
        RECT 115.030 152.520 115.170 156.710 ;
        RECT 115.430 156.620 115.690 156.940 ;
        RECT 115.490 154.900 115.630 156.620 ;
        RECT 115.430 154.580 115.690 154.900 ;
        RECT 115.430 153.960 115.690 154.220 ;
        RECT 116.410 153.960 116.550 157.640 ;
        RECT 116.810 157.475 117.070 157.620 ;
        RECT 116.800 157.105 117.080 157.475 ;
        RECT 115.430 153.900 116.550 153.960 ;
        RECT 115.490 153.820 116.550 153.900 ;
        RECT 116.810 153.560 117.070 153.880 ;
        RECT 116.870 152.520 117.010 153.560 ;
        RECT 114.970 152.200 115.230 152.520 ;
        RECT 116.810 152.200 117.070 152.520 ;
        RECT 115.890 148.800 116.150 149.120 ;
        RECT 114.970 148.120 115.230 148.440 ;
        RECT 115.030 146.740 115.170 148.120 ;
        RECT 115.430 147.780 115.690 148.100 ;
        RECT 114.970 146.420 115.230 146.740 ;
        RECT 115.490 144.020 115.630 147.780 ;
        RECT 115.950 146.060 116.090 148.800 ;
        RECT 116.810 146.760 117.070 147.080 ;
        RECT 116.350 146.420 116.610 146.740 ;
        RECT 115.890 145.740 116.150 146.060 ;
        RECT 116.410 145.915 116.550 146.420 ;
        RECT 116.870 146.060 117.010 146.760 ;
        RECT 117.330 146.595 117.470 182.260 ;
        RECT 119.170 179.040 119.310 186.200 ;
        RECT 119.630 183.800 119.770 186.200 ;
        RECT 121.010 186.180 121.150 186.880 ;
        RECT 120.950 185.860 121.210 186.180 ;
        RECT 121.410 185.860 121.670 186.180 ;
        RECT 121.470 184.140 121.610 185.860 ;
        RECT 121.410 183.820 121.670 184.140 ;
        RECT 119.570 183.480 119.830 183.800 ;
        RECT 119.770 182.605 121.650 182.975 ;
        RECT 119.110 178.720 119.370 179.040 ;
        RECT 117.730 178.380 117.990 178.700 ;
        RECT 117.790 175.980 117.930 178.380 ;
        RECT 118.650 177.700 118.910 178.020 ;
        RECT 117.730 175.660 117.990 175.980 ;
        RECT 118.710 175.300 118.850 177.700 ;
        RECT 119.170 177.000 119.310 178.720 ;
        RECT 119.770 177.165 121.650 177.535 ;
        RECT 119.110 176.680 119.370 177.000 ;
        RECT 118.650 174.980 118.910 175.300 ;
        RECT 119.110 172.260 119.370 172.580 ;
        RECT 119.170 171.470 119.310 172.260 ;
        RECT 119.770 171.725 121.650 172.095 ;
        RECT 121.930 171.640 122.070 199.460 ;
        RECT 122.850 198.760 122.990 200.140 ;
        RECT 122.790 198.440 123.050 198.760 ;
        RECT 123.770 197.400 123.910 200.820 ;
        RECT 125.150 200.800 125.290 205.580 ;
        RECT 126.070 202.920 126.210 205.920 ;
        RECT 125.610 202.840 126.210 202.920 ;
        RECT 125.550 202.780 126.210 202.840 ;
        RECT 125.550 202.520 125.810 202.780 ;
        RECT 125.550 201.160 125.810 201.480 ;
        RECT 125.090 200.480 125.350 200.800 ;
        RECT 124.620 197.905 124.900 198.275 ;
        RECT 125.610 198.080 125.750 201.160 ;
        RECT 126.070 200.800 126.210 202.780 ;
        RECT 126.010 200.480 126.270 200.800 ;
        RECT 124.690 197.740 124.830 197.905 ;
        RECT 125.550 197.760 125.810 198.080 ;
        RECT 124.630 197.420 124.890 197.740 ;
        RECT 125.610 197.595 125.750 197.760 ;
        RECT 123.710 197.080 123.970 197.400 ;
        RECT 125.540 197.225 125.820 197.595 ;
        RECT 126.070 197.400 126.210 200.480 ;
        RECT 126.470 199.800 126.730 200.120 ;
        RECT 125.090 194.020 125.350 194.340 ;
        RECT 124.630 192.320 124.890 192.640 ;
        RECT 122.330 191.980 122.590 192.300 ;
        RECT 122.390 187.880 122.530 191.980 ;
        RECT 123.250 191.300 123.510 191.620 ;
        RECT 123.710 191.300 123.970 191.620 ;
        RECT 122.790 189.940 123.050 190.260 ;
        RECT 122.330 187.560 122.590 187.880 ;
        RECT 122.850 183.995 122.990 189.940 ;
        RECT 123.310 189.240 123.450 191.300 ;
        RECT 123.770 190.115 123.910 191.300 ;
        RECT 123.700 189.745 123.980 190.115 ;
        RECT 124.170 189.940 124.430 190.260 ;
        RECT 123.250 188.920 123.510 189.240 ;
        RECT 122.330 183.480 122.590 183.800 ;
        RECT 122.780 183.625 123.060 183.995 ;
        RECT 122.390 173.260 122.530 183.480 ;
        RECT 124.230 182.100 124.370 189.940 ;
        RECT 124.690 189.240 124.830 192.320 ;
        RECT 124.630 188.920 124.890 189.240 ;
        RECT 124.630 186.880 124.890 187.200 ;
        RECT 124.170 181.780 124.430 182.100 ;
        RECT 122.790 181.440 123.050 181.760 ;
        RECT 122.330 172.940 122.590 173.260 ;
        RECT 120.030 171.470 120.290 171.560 ;
        RECT 121.930 171.500 122.530 171.640 ;
        RECT 119.170 171.330 120.290 171.470 ;
        RECT 120.030 171.240 120.290 171.330 ;
        RECT 120.090 170.880 120.230 171.240 ;
        RECT 121.870 170.900 122.130 171.220 ;
        RECT 117.730 170.560 117.990 170.880 ;
        RECT 119.570 170.560 119.830 170.880 ;
        RECT 120.030 170.560 120.290 170.880 ;
        RECT 121.410 170.560 121.670 170.880 ;
        RECT 117.790 169.860 117.930 170.560 ;
        RECT 117.730 169.540 117.990 169.860 ;
        RECT 118.190 169.540 118.450 169.860 ;
        RECT 117.730 167.840 117.990 168.160 ;
        RECT 117.790 166.120 117.930 167.840 ;
        RECT 117.730 165.800 117.990 166.120 ;
        RECT 118.250 165.440 118.390 169.540 ;
        RECT 119.110 168.355 119.370 168.500 ;
        RECT 119.100 167.985 119.380 168.355 ;
        RECT 119.630 167.820 119.770 170.560 ;
        RECT 120.030 169.540 120.290 169.860 ;
        RECT 120.090 168.500 120.230 169.540 ;
        RECT 120.030 168.180 120.290 168.500 ;
        RECT 118.650 167.500 118.910 167.820 ;
        RECT 119.570 167.500 119.830 167.820 ;
        RECT 118.710 166.120 118.850 167.500 ;
        RECT 119.110 166.820 119.370 167.140 ;
        RECT 121.470 167.050 121.610 170.560 ;
        RECT 121.930 169.860 122.070 170.900 ;
        RECT 121.870 169.540 122.130 169.860 ;
        RECT 121.470 166.910 122.070 167.050 ;
        RECT 118.650 165.800 118.910 166.120 ;
        RECT 119.170 166.030 119.310 166.820 ;
        RECT 119.770 166.285 121.650 166.655 ;
        RECT 119.170 165.890 120.690 166.030 ;
        RECT 118.190 165.120 118.450 165.440 ;
        RECT 119.100 165.265 119.380 165.635 ;
        RECT 120.550 165.440 120.690 165.890 ;
        RECT 121.930 165.440 122.070 166.910 ;
        RECT 120.030 165.350 120.290 165.440 ;
        RECT 117.730 162.060 117.990 162.380 ;
        RECT 118.190 162.060 118.450 162.380 ;
        RECT 119.170 162.235 119.310 165.265 ;
        RECT 119.630 165.210 120.290 165.350 ;
        RECT 119.630 162.720 119.770 165.210 ;
        RECT 120.030 165.120 120.290 165.210 ;
        RECT 120.490 165.120 120.750 165.440 ;
        RECT 121.870 165.120 122.130 165.440 ;
        RECT 121.930 164.955 122.070 165.120 ;
        RECT 121.860 164.585 122.140 164.955 ;
        RECT 121.870 162.740 122.130 163.060 ;
        RECT 119.570 162.400 119.830 162.720 ;
        RECT 117.790 153.395 117.930 162.060 ;
        RECT 118.250 158.980 118.390 162.060 ;
        RECT 119.100 161.865 119.380 162.235 ;
        RECT 119.110 161.720 119.370 161.865 ;
        RECT 119.770 160.845 121.650 161.215 ;
        RECT 118.650 160.360 118.910 160.680 ;
        RECT 118.190 158.660 118.450 158.980 ;
        RECT 118.250 154.560 118.390 158.660 ;
        RECT 118.710 157.960 118.850 160.360 ;
        RECT 121.930 159.320 122.070 162.740 ;
        RECT 121.870 159.000 122.130 159.320 ;
        RECT 120.030 158.660 120.290 158.980 ;
        RECT 121.410 158.660 121.670 158.980 ;
        RECT 120.090 157.960 120.230 158.660 ;
        RECT 121.470 157.960 121.610 158.660 ;
        RECT 118.650 157.640 118.910 157.960 ;
        RECT 120.030 157.640 120.290 157.960 ;
        RECT 121.410 157.640 121.670 157.960 ;
        RECT 119.570 157.360 119.830 157.620 ;
        RECT 119.570 157.300 120.690 157.360 ;
        RECT 119.630 157.220 120.690 157.300 ;
        RECT 120.550 156.940 120.690 157.220 ;
        RECT 120.490 156.620 120.750 156.940 ;
        RECT 118.650 155.940 118.910 156.260 ;
        RECT 118.710 154.560 118.850 155.940 ;
        RECT 119.770 155.405 121.650 155.775 ;
        RECT 118.190 154.240 118.450 154.560 ;
        RECT 118.650 154.240 118.910 154.560 ;
        RECT 118.250 153.960 118.390 154.240 ;
        RECT 118.250 153.820 118.850 153.960 ;
        RECT 119.570 153.900 119.830 154.220 ;
        RECT 120.030 154.075 120.290 154.220 ;
        RECT 120.490 154.130 120.750 154.220 ;
        RECT 121.930 154.130 122.070 159.000 ;
        RECT 117.720 153.025 118.000 153.395 ;
        RECT 117.730 151.180 117.990 151.500 ;
        RECT 117.260 146.225 117.540 146.595 ;
        RECT 115.430 143.700 115.690 144.020 ;
        RECT 115.950 143.680 116.090 145.740 ;
        RECT 116.340 145.545 116.620 145.915 ;
        RECT 116.810 145.740 117.070 146.060 ;
        RECT 117.270 145.740 117.530 146.060 ;
        RECT 116.350 145.060 116.610 145.380 ;
        RECT 116.410 143.680 116.550 145.060 ;
        RECT 115.890 143.360 116.150 143.680 ;
        RECT 116.350 143.590 116.610 143.680 ;
        RECT 116.350 143.450 117.010 143.590 ;
        RECT 116.350 143.360 116.610 143.450 ;
        RECT 114.970 143.020 115.230 143.340 ;
        RECT 115.030 138.320 115.170 143.020 ;
        RECT 116.350 142.680 116.610 143.000 ;
        RECT 116.410 140.280 116.550 142.680 ;
        RECT 116.870 140.620 117.010 143.450 ;
        RECT 117.330 143.000 117.470 145.740 ;
        RECT 117.270 142.680 117.530 143.000 ;
        RECT 116.810 140.300 117.070 140.620 ;
        RECT 117.270 140.300 117.530 140.620 ;
        RECT 116.350 139.960 116.610 140.280 ;
        RECT 115.030 138.180 116.090 138.320 ;
        RECT 114.970 134.180 115.230 134.500 ;
        RECT 113.130 132.480 113.390 132.625 ;
        RECT 114.510 132.480 114.770 132.800 ;
        RECT 113.130 131.800 113.390 132.120 ;
        RECT 113.580 131.945 113.860 132.315 ;
        RECT 112.670 129.760 112.930 130.080 ;
        RECT 113.190 129.740 113.330 131.800 ;
        RECT 113.650 130.420 113.790 131.945 ;
        RECT 113.590 130.100 113.850 130.420 ;
        RECT 115.030 130.330 115.170 134.180 ;
        RECT 114.110 130.190 115.170 130.330 ;
        RECT 112.210 129.420 112.470 129.740 ;
        RECT 113.130 129.420 113.390 129.740 ;
        RECT 110.370 128.740 110.630 129.060 ;
        RECT 110.830 128.740 111.090 129.060 ;
        RECT 111.290 128.740 111.550 129.060 ;
        RECT 107.150 127.720 107.410 127.810 ;
        RECT 108.130 127.700 108.270 127.865 ;
        RECT 108.530 127.720 108.790 128.040 ;
        RECT 110.430 127.700 110.570 128.740 ;
        RECT 108.070 127.380 108.330 127.700 ;
        RECT 110.370 127.380 110.630 127.700 ;
        RECT 112.670 127.380 112.930 127.700 ;
        RECT 103.470 127.040 103.730 127.360 ;
        RECT 105.770 127.040 106.030 127.360 ;
        RECT 106.690 126.700 106.950 127.020 ;
        RECT 110.370 126.700 110.630 127.020 ;
        RECT 81.850 126.020 82.110 126.340 ;
        RECT 85.990 126.020 86.250 126.340 ;
        RECT 94.730 126.020 94.990 126.340 ;
        RECT 97.030 126.020 97.290 126.340 ;
        RECT 99.790 126.020 100.050 126.340 ;
        RECT 101.170 126.020 101.430 126.340 ;
        RECT 101.630 126.020 101.890 126.340 ;
        RECT 102.090 126.020 102.350 126.340 ;
        RECT 106.750 126.250 106.890 126.700 ;
        RECT 106.750 126.110 107.350 126.250 ;
        RECT 80.470 125.000 80.730 125.320 ;
        RECT 80.010 124.320 80.270 124.640 ;
        RECT 94.790 124.300 94.930 126.020 ;
        RECT 97.090 125.320 97.230 126.020 ;
        RECT 97.030 125.000 97.290 125.320 ;
        RECT 79.550 123.980 79.810 124.300 ;
        RECT 88.750 123.980 89.010 124.300 ;
        RECT 94.270 123.980 94.530 124.300 ;
        RECT 94.730 123.980 94.990 124.300 ;
        RECT 98.410 123.980 98.670 124.300 ;
        RECT 81.850 123.300 82.110 123.620 ;
        RECT 86.450 123.300 86.710 123.620 ;
        RECT 81.910 122.230 82.050 123.300 ;
        RECT 86.510 122.510 86.650 123.300 ;
        RECT 85.590 122.370 86.650 122.510 ;
        RECT 85.590 122.230 85.730 122.370 ;
        RECT 70.800 120.230 71.080 122.230 ;
        RECT 74.480 120.230 74.760 122.230 ;
        RECT 78.160 120.230 78.440 122.230 ;
        RECT 81.840 120.230 82.120 122.230 ;
        RECT 85.520 120.230 85.800 122.230 ;
        RECT 88.810 121.240 88.950 123.980 ;
        RECT 89.210 123.300 89.470 123.620 ;
        RECT 93.810 123.300 94.070 123.620 ;
        RECT 89.270 122.230 89.410 123.300 ;
        RECT 89.770 122.765 91.650 123.135 ;
        RECT 93.870 122.510 94.010 123.300 ;
        RECT 94.330 122.600 94.470 123.980 ;
        RECT 97.490 123.300 97.750 123.620 ;
        RECT 92.950 122.370 94.010 122.510 ;
        RECT 92.950 122.230 93.090 122.370 ;
        RECT 94.270 122.280 94.530 122.600 ;
        RECT 97.550 122.510 97.690 123.300 ;
        RECT 98.470 122.600 98.610 123.980 ;
        RECT 96.630 122.370 97.690 122.510 ;
        RECT 96.630 122.230 96.770 122.370 ;
        RECT 98.410 122.280 98.670 122.600 ;
        RECT 99.850 122.260 99.990 126.020 ;
        RECT 101.230 124.300 101.370 126.020 ;
        RECT 101.690 124.300 101.830 126.020 ;
        RECT 104.770 125.485 106.650 125.855 ;
        RECT 101.170 123.980 101.430 124.300 ;
        RECT 101.630 123.980 101.890 124.300 ;
        RECT 101.170 123.300 101.430 123.620 ;
        RECT 103.930 123.300 104.190 123.620 ;
        RECT 101.230 122.510 101.370 123.300 ;
        RECT 100.310 122.370 101.370 122.510 ;
        RECT 88.750 120.920 89.010 121.240 ;
        RECT 89.200 120.230 89.480 122.230 ;
        RECT 92.880 120.230 93.160 122.230 ;
        RECT 96.560 120.230 96.840 122.230 ;
        RECT 99.790 121.940 100.050 122.260 ;
        RECT 100.310 122.230 100.450 122.370 ;
        RECT 103.990 122.230 104.130 123.300 ;
        RECT 100.240 120.230 100.520 122.230 ;
        RECT 103.920 120.230 104.200 122.230 ;
        RECT 107.210 121.580 107.350 126.110 ;
        RECT 109.910 126.020 110.170 126.340 ;
        RECT 108.530 124.550 108.790 124.640 ;
        RECT 109.970 124.550 110.110 126.020 ;
        RECT 108.530 124.410 110.110 124.550 ;
        RECT 108.530 124.320 108.790 124.410 ;
        RECT 110.430 124.300 110.570 126.700 ;
        RECT 112.730 126.680 112.870 127.380 ;
        RECT 114.110 127.360 114.250 130.190 ;
        RECT 114.050 127.040 114.310 127.360 ;
        RECT 115.950 127.270 116.090 138.180 ;
        RECT 116.410 138.150 116.550 139.960 ;
        RECT 116.870 138.920 117.010 140.300 ;
        RECT 117.330 138.920 117.470 140.300 ;
        RECT 116.810 138.600 117.070 138.920 ;
        RECT 117.270 138.600 117.530 138.920 ;
        RECT 117.270 138.150 117.530 138.240 ;
        RECT 116.410 138.010 117.530 138.150 ;
        RECT 117.270 137.920 117.530 138.010 ;
        RECT 116.800 136.705 117.080 137.075 ;
        RECT 116.870 135.520 117.010 136.705 ;
        RECT 116.810 135.200 117.070 135.520 ;
        RECT 116.810 131.460 117.070 131.780 ;
        RECT 116.870 129.740 117.010 131.460 ;
        RECT 116.350 129.420 116.610 129.740 ;
        RECT 116.810 129.420 117.070 129.740 ;
        RECT 117.270 129.420 117.530 129.740 ;
        RECT 116.410 128.235 116.550 129.420 ;
        RECT 116.800 128.545 117.080 128.915 ;
        RECT 116.340 127.865 116.620 128.235 ;
        RECT 116.870 128.040 117.010 128.545 ;
        RECT 116.810 127.720 117.070 128.040 ;
        RECT 116.810 127.270 117.070 127.360 ;
        RECT 115.950 127.130 117.070 127.270 ;
        RECT 116.810 127.040 117.070 127.130 ;
        RECT 114.510 126.700 114.770 127.020 ;
        RECT 112.210 126.360 112.470 126.680 ;
        RECT 112.670 126.360 112.930 126.680 ;
        RECT 112.270 125.320 112.410 126.360 ;
        RECT 114.570 125.320 114.710 126.700 ;
        RECT 116.340 125.825 116.620 126.195 ;
        RECT 112.210 125.000 112.470 125.320 ;
        RECT 114.510 125.000 114.770 125.320 ;
        RECT 114.970 124.660 115.230 124.980 ;
        RECT 110.370 123.980 110.630 124.300 ;
        RECT 108.530 123.640 108.790 123.960 ;
        RECT 108.590 122.510 108.730 123.640 ;
        RECT 109.910 123.300 110.170 123.620 ;
        RECT 107.670 122.370 108.730 122.510 ;
        RECT 107.670 122.230 107.810 122.370 ;
        RECT 107.150 121.260 107.410 121.580 ;
        RECT 107.600 120.230 107.880 122.230 ;
        RECT 109.970 122.000 110.110 123.300 ;
        RECT 110.890 122.370 111.490 122.510 ;
        RECT 110.890 122.000 111.030 122.370 ;
        RECT 111.350 122.230 111.490 122.370 ;
        RECT 115.030 122.230 115.170 124.660 ;
        RECT 116.410 122.260 116.550 125.825 ;
        RECT 117.330 124.300 117.470 129.420 ;
        RECT 117.790 125.320 117.930 151.180 ;
        RECT 118.190 147.780 118.450 148.100 ;
        RECT 118.250 146.060 118.390 147.780 ;
        RECT 118.710 146.060 118.850 153.820 ;
        RECT 119.630 151.500 119.770 153.900 ;
        RECT 120.020 153.705 120.300 154.075 ;
        RECT 120.490 153.990 122.070 154.130 ;
        RECT 120.490 153.900 120.750 153.990 ;
        RECT 119.570 151.180 119.830 151.500 ;
        RECT 119.770 149.965 121.650 150.335 ;
        RECT 119.110 148.120 119.370 148.440 ;
        RECT 118.190 145.740 118.450 146.060 ;
        RECT 118.650 145.740 118.910 146.060 ;
        RECT 118.190 145.060 118.450 145.380 ;
        RECT 118.650 145.060 118.910 145.380 ;
        RECT 118.250 140.620 118.390 145.060 ;
        RECT 118.190 140.300 118.450 140.620 ;
        RECT 118.190 139.620 118.450 139.940 ;
        RECT 118.250 138.920 118.390 139.620 ;
        RECT 118.190 138.600 118.450 138.920 ;
        RECT 118.190 137.920 118.450 138.240 ;
        RECT 118.250 136.200 118.390 137.920 ;
        RECT 118.190 135.880 118.450 136.200 ;
        RECT 118.710 129.480 118.850 145.060 ;
        RECT 119.170 138.240 119.310 148.120 ;
        RECT 121.870 147.780 122.130 148.100 ;
        RECT 121.930 146.400 122.070 147.780 ;
        RECT 121.870 146.080 122.130 146.400 ;
        RECT 121.870 145.060 122.130 145.380 ;
        RECT 119.770 144.525 121.650 144.895 ;
        RECT 121.930 143.340 122.070 145.060 ;
        RECT 121.870 143.020 122.130 143.340 ;
        RECT 119.770 139.085 121.650 139.455 ;
        RECT 120.030 138.600 120.290 138.920 ;
        RECT 119.110 137.920 119.370 138.240 ;
        RECT 120.090 137.900 120.230 138.600 ;
        RECT 120.030 137.580 120.290 137.900 ;
        RECT 120.090 137.220 120.230 137.580 ;
        RECT 120.030 136.900 120.290 137.220 ;
        RECT 119.770 133.645 121.650 134.015 ;
        RECT 120.950 132.480 121.210 132.800 ;
        RECT 121.010 132.120 121.150 132.480 ;
        RECT 120.950 131.800 121.210 132.120 ;
        RECT 122.390 130.955 122.530 171.500 ;
        RECT 122.850 170.880 122.990 181.440 ;
        RECT 124.690 180.740 124.830 186.880 ;
        RECT 125.150 186.860 125.290 194.020 ;
        RECT 125.610 193.400 125.750 197.225 ;
        RECT 126.010 197.080 126.270 197.400 ;
        RECT 126.530 194.340 126.670 199.800 ;
        RECT 126.990 195.700 127.130 207.960 ;
        RECT 127.910 205.900 128.050 209.455 ;
        RECT 132.050 208.620 132.190 209.455 ;
        RECT 131.990 208.300 132.250 208.620 ;
        RECT 136.190 207.940 136.330 209.455 ;
        RECT 138.430 208.300 138.690 208.620 ;
        RECT 132.910 207.620 133.170 207.940 ;
        RECT 136.130 207.620 136.390 207.940 ;
        RECT 132.970 206.580 133.110 207.620 ;
        RECT 134.770 207.085 136.650 207.455 ;
        RECT 132.910 206.260 133.170 206.580 ;
        RECT 137.050 206.320 137.310 206.580 ;
        RECT 136.650 206.260 137.310 206.320 ;
        RECT 136.650 206.180 137.250 206.260 ;
        RECT 127.850 205.580 128.110 205.900 ;
        RECT 135.210 205.580 135.470 205.900 ;
        RECT 131.530 205.240 131.790 205.560 ;
        RECT 128.310 204.900 128.570 205.220 ;
        RECT 127.850 198.100 128.110 198.420 ;
        RECT 127.910 197.480 128.050 198.100 ;
        RECT 127.450 197.340 128.050 197.480 ;
        RECT 126.930 195.380 127.190 195.700 ;
        RECT 127.450 195.020 127.590 197.340 ;
        RECT 127.390 194.700 127.650 195.020 ;
        RECT 126.470 194.020 126.730 194.340 ;
        RECT 125.610 193.260 127.130 193.400 ;
        RECT 126.010 191.980 126.270 192.300 ;
        RECT 125.550 191.300 125.810 191.620 ;
        RECT 125.610 187.200 125.750 191.300 ;
        RECT 126.070 189.240 126.210 191.980 ;
        RECT 126.990 191.620 127.130 193.260 ;
        RECT 127.450 192.980 127.590 194.700 ;
        RECT 127.390 192.660 127.650 192.980 ;
        RECT 127.840 192.465 128.120 192.835 ;
        RECT 126.470 191.300 126.730 191.620 ;
        RECT 126.930 191.300 127.190 191.620 ;
        RECT 126.010 188.920 126.270 189.240 ;
        RECT 125.550 186.880 125.810 187.200 ;
        RECT 125.090 186.540 125.350 186.860 ;
        RECT 125.090 184.160 125.350 184.480 ;
        RECT 124.630 180.420 124.890 180.740 ;
        RECT 124.170 178.380 124.430 178.700 ;
        RECT 123.250 177.700 123.510 178.020 ;
        RECT 123.310 175.980 123.450 177.700 ;
        RECT 124.230 177.000 124.370 178.380 ;
        RECT 124.170 176.680 124.430 177.000 ;
        RECT 124.690 176.660 124.830 180.420 ;
        RECT 124.630 176.340 124.890 176.660 ;
        RECT 123.250 175.660 123.510 175.980 ;
        RECT 123.710 174.980 123.970 175.300 ;
        RECT 122.790 170.560 123.050 170.880 ;
        RECT 122.850 167.730 122.990 170.560 ;
        RECT 123.250 167.730 123.510 167.820 ;
        RECT 122.850 167.590 123.510 167.730 ;
        RECT 123.250 167.500 123.510 167.590 ;
        RECT 123.770 167.140 123.910 174.980 ;
        RECT 124.170 173.620 124.430 173.940 ;
        RECT 124.630 173.620 124.890 173.940 ;
        RECT 123.250 166.820 123.510 167.140 ;
        RECT 123.710 166.820 123.970 167.140 ;
        RECT 123.310 166.120 123.450 166.820 ;
        RECT 123.250 165.800 123.510 166.120 ;
        RECT 122.790 161.380 123.050 161.700 ;
        RECT 123.250 161.380 123.510 161.700 ;
        RECT 122.850 155.240 122.990 161.380 ;
        RECT 123.310 157.280 123.450 161.380 ;
        RECT 124.230 160.000 124.370 173.620 ;
        RECT 124.690 171.560 124.830 173.620 ;
        RECT 124.630 171.240 124.890 171.560 ;
        RECT 124.690 165.780 124.830 171.240 ;
        RECT 124.630 165.460 124.890 165.780 ;
        RECT 125.150 163.060 125.290 184.160 ;
        RECT 126.530 182.400 126.670 191.300 ;
        RECT 126.930 190.280 127.190 190.600 ;
        RECT 126.990 184.820 127.130 190.280 ;
        RECT 127.390 189.260 127.650 189.580 ;
        RECT 127.450 187.395 127.590 189.260 ;
        RECT 127.380 187.025 127.660 187.395 ;
        RECT 126.930 184.500 127.190 184.820 ;
        RECT 127.910 184.480 128.050 192.465 ;
        RECT 128.370 190.795 128.510 204.900 ;
        RECT 129.750 202.780 131.270 202.920 ;
        RECT 129.750 201.480 129.890 202.780 ;
        RECT 130.610 202.180 130.870 202.500 ;
        RECT 129.690 201.160 129.950 201.480 ;
        RECT 129.230 200.480 129.490 200.800 ;
        RECT 128.770 199.460 129.030 199.780 ;
        RECT 128.830 198.420 128.970 199.460 ;
        RECT 128.770 198.100 129.030 198.420 ;
        RECT 129.290 196.915 129.430 200.480 ;
        RECT 129.690 197.990 129.950 198.080 ;
        RECT 130.670 197.990 130.810 202.180 ;
        RECT 131.130 201.140 131.270 202.780 ;
        RECT 131.070 200.820 131.330 201.140 ;
        RECT 131.590 200.460 131.730 205.240 ;
        RECT 131.990 203.880 132.250 204.200 ;
        RECT 131.530 200.140 131.790 200.460 ;
        RECT 132.050 200.120 132.190 203.880 ;
        RECT 133.830 203.200 134.090 203.520 ;
        RECT 134.750 203.200 135.010 203.520 ;
        RECT 133.370 202.180 133.630 202.500 ;
        RECT 133.430 201.140 133.570 202.180 ;
        RECT 133.370 200.820 133.630 201.140 ;
        RECT 131.990 199.800 132.250 200.120 ;
        RECT 129.690 197.850 130.810 197.990 ;
        RECT 129.690 197.760 129.950 197.850 ;
        RECT 129.220 196.545 129.500 196.915 ;
        RECT 129.230 194.700 129.490 195.020 ;
        RECT 128.770 193.000 129.030 193.320 ;
        RECT 128.830 192.155 128.970 193.000 ;
        RECT 128.760 191.785 129.040 192.155 ;
        RECT 128.300 190.425 128.580 190.795 ;
        RECT 128.370 189.920 128.510 190.425 ;
        RECT 128.830 190.260 128.970 191.785 ;
        RECT 129.290 190.260 129.430 194.700 ;
        RECT 129.690 194.360 129.950 194.680 ;
        RECT 129.750 193.320 129.890 194.360 ;
        RECT 129.690 193.000 129.950 193.320 ;
        RECT 129.750 192.640 129.890 193.000 ;
        RECT 129.690 192.320 129.950 192.640 ;
        RECT 130.210 191.620 130.350 197.850 ;
        RECT 130.670 196.970 130.810 197.850 ;
        RECT 131.530 197.990 131.790 198.080 ;
        RECT 132.050 197.990 132.190 199.800 ;
        RECT 132.450 199.460 132.710 199.780 ;
        RECT 133.370 199.460 133.630 199.780 ;
        RECT 131.530 197.850 132.190 197.990 ;
        RECT 131.530 197.760 131.790 197.850 ;
        RECT 131.990 197.080 132.250 197.400 ;
        RECT 131.530 196.970 131.790 197.060 ;
        RECT 130.670 196.830 131.790 196.970 ;
        RECT 131.530 196.740 131.790 196.830 ;
        RECT 132.050 195.610 132.190 197.080 ;
        RECT 132.510 196.915 132.650 199.460 ;
        RECT 133.430 198.760 133.570 199.460 ;
        RECT 133.890 198.760 134.030 203.200 ;
        RECT 134.810 202.920 134.950 203.200 ;
        RECT 135.270 203.180 135.410 205.580 ;
        RECT 136.650 204.200 136.790 206.180 ;
        RECT 138.490 205.900 138.630 208.300 ;
        RECT 138.430 205.580 138.690 205.900 ;
        RECT 139.810 205.580 140.070 205.900 ;
        RECT 136.590 203.880 136.850 204.200 ;
        RECT 139.870 203.860 140.010 205.580 ;
        RECT 140.330 204.200 140.470 209.455 ;
        RECT 142.110 207.960 142.370 208.280 ;
        RECT 140.730 207.620 140.990 207.940 ;
        RECT 140.270 203.880 140.530 204.200 ;
        RECT 139.810 203.540 140.070 203.860 ;
        RECT 134.350 202.780 134.950 202.920 ;
        RECT 135.210 202.860 135.470 203.180 ;
        RECT 134.350 201.480 134.490 202.780 ;
        RECT 138.890 202.180 139.150 202.500 ;
        RECT 134.770 201.645 136.650 202.015 ;
        RECT 134.290 201.160 134.550 201.480 ;
        RECT 137.050 200.480 137.310 200.800 ;
        RECT 134.290 200.140 134.550 200.460 ;
        RECT 133.370 198.440 133.630 198.760 ;
        RECT 133.830 198.440 134.090 198.760 ;
        RECT 133.370 197.760 133.630 198.080 ;
        RECT 132.910 197.595 133.170 197.740 ;
        RECT 132.900 197.225 133.180 197.595 ;
        RECT 133.430 197.310 133.570 197.760 ;
        RECT 133.430 197.170 133.600 197.310 ;
        RECT 132.440 196.545 132.720 196.915 ;
        RECT 132.910 196.740 133.170 197.060 ;
        RECT 132.450 195.610 132.710 195.700 ;
        RECT 132.050 195.470 132.710 195.610 ;
        RECT 132.450 195.380 132.710 195.470 ;
        RECT 131.060 194.505 131.340 194.875 ;
        RECT 132.450 194.700 132.710 195.020 ;
        RECT 131.070 194.360 131.330 194.505 ;
        RECT 132.510 192.300 132.650 194.700 ;
        RECT 130.610 191.980 130.870 192.300 ;
        RECT 132.450 192.210 132.710 192.300 ;
        RECT 132.050 192.070 132.710 192.210 ;
        RECT 130.150 191.300 130.410 191.620 ;
        RECT 128.770 189.940 129.030 190.260 ;
        RECT 129.230 189.940 129.490 190.260 ;
        RECT 128.310 189.600 128.570 189.920 ;
        RECT 128.370 187.880 128.510 189.600 ;
        RECT 130.670 189.580 130.810 191.980 ;
        RECT 131.530 191.300 131.790 191.620 ;
        RECT 130.610 189.435 130.870 189.580 ;
        RECT 130.600 189.065 130.880 189.435 ;
        RECT 131.070 189.260 131.330 189.580 ;
        RECT 130.150 188.580 130.410 188.900 ;
        RECT 131.130 188.755 131.270 189.260 ;
        RECT 128.310 187.560 128.570 187.880 ;
        RECT 128.770 186.880 129.030 187.200 ;
        RECT 128.830 184.480 128.970 186.880 ;
        RECT 127.850 184.160 128.110 184.480 ;
        RECT 128.770 184.160 129.030 184.480 ;
        RECT 126.930 183.370 127.190 183.460 ;
        RECT 126.930 183.230 128.510 183.370 ;
        RECT 126.930 183.140 127.190 183.230 ;
        RECT 128.370 182.400 128.510 183.230 ;
        RECT 126.530 182.260 127.130 182.400 ;
        RECT 126.470 181.440 126.730 181.760 ;
        RECT 126.530 179.720 126.670 181.440 ;
        RECT 126.470 179.400 126.730 179.720 ;
        RECT 126.470 178.380 126.730 178.700 ;
        RECT 125.550 177.700 125.810 178.020 ;
        RECT 125.090 162.740 125.350 163.060 ;
        RECT 125.150 162.040 125.290 162.740 ;
        RECT 125.090 161.720 125.350 162.040 ;
        RECT 124.170 159.680 124.430 160.000 ;
        RECT 123.250 156.960 123.510 157.280 ;
        RECT 123.250 155.940 123.510 156.260 ;
        RECT 122.790 154.920 123.050 155.240 ;
        RECT 123.310 154.640 123.450 155.940 ;
        RECT 122.790 154.240 123.050 154.560 ;
        RECT 123.310 154.500 123.910 154.640 ;
        RECT 122.850 151.500 122.990 154.240 ;
        RECT 123.250 153.900 123.510 154.220 ;
        RECT 123.310 152.520 123.450 153.900 ;
        RECT 123.250 152.200 123.510 152.520 ;
        RECT 122.790 151.180 123.050 151.500 ;
        RECT 123.250 144.040 123.510 144.360 ;
        RECT 123.310 141.300 123.450 144.040 ;
        RECT 123.250 140.980 123.510 141.300 ;
        RECT 122.790 140.640 123.050 140.960 ;
        RECT 122.850 138.240 122.990 140.640 ;
        RECT 122.790 137.920 123.050 138.240 ;
        RECT 121.410 130.440 121.670 130.760 ;
        RECT 122.320 130.585 122.600 130.955 ;
        RECT 118.190 129.080 118.450 129.400 ;
        RECT 118.710 129.340 119.310 129.480 ;
        RECT 118.250 128.040 118.390 129.080 ;
        RECT 118.650 128.740 118.910 129.060 ;
        RECT 118.190 127.720 118.450 128.040 ;
        RECT 118.710 127.440 118.850 128.740 ;
        RECT 118.250 127.360 118.850 127.440 ;
        RECT 118.190 127.300 118.850 127.360 ;
        RECT 118.190 127.040 118.450 127.300 ;
        RECT 119.170 126.930 119.310 129.340 ;
        RECT 121.470 129.060 121.610 130.440 ;
        RECT 122.850 130.330 122.990 137.920 ;
        RECT 123.250 136.900 123.510 137.220 ;
        RECT 123.310 135.180 123.450 136.900 ;
        RECT 123.250 134.860 123.510 135.180 ;
        RECT 123.310 132.460 123.450 134.860 ;
        RECT 123.250 132.140 123.510 132.460 ;
        RECT 122.390 130.190 122.990 130.330 ;
        RECT 122.390 129.400 122.530 130.190 ;
        RECT 123.310 130.080 123.450 132.140 ;
        RECT 123.250 129.760 123.510 130.080 ;
        RECT 122.330 129.080 122.590 129.400 ;
        RECT 121.410 128.740 121.670 129.060 ;
        RECT 122.790 128.740 123.050 129.060 ;
        RECT 119.770 128.205 121.650 128.575 ;
        RECT 121.410 127.380 121.670 127.700 ;
        RECT 120.490 126.930 120.750 127.020 ;
        RECT 119.170 126.790 120.750 126.930 ;
        RECT 121.470 126.875 121.610 127.380 ;
        RECT 122.850 127.020 122.990 128.740 ;
        RECT 120.490 126.700 120.750 126.790 ;
        RECT 118.190 126.360 118.450 126.680 ;
        RECT 121.400 126.505 121.680 126.875 ;
        RECT 122.790 126.700 123.050 127.020 ;
        RECT 123.250 126.875 123.510 127.020 ;
        RECT 117.730 125.000 117.990 125.320 ;
        RECT 117.270 123.980 117.530 124.300 ;
        RECT 109.970 121.860 111.030 122.000 ;
        RECT 111.280 120.230 111.560 122.230 ;
        RECT 114.960 120.230 115.240 122.230 ;
        RECT 116.350 121.940 116.610 122.260 ;
        RECT 118.250 121.240 118.390 126.360 ;
        RECT 122.850 124.300 122.990 126.700 ;
        RECT 123.240 126.505 123.520 126.875 ;
        RECT 122.790 123.980 123.050 124.300 ;
        RECT 123.310 123.960 123.450 126.505 ;
        RECT 123.770 125.320 123.910 154.500 ;
        RECT 124.230 152.520 124.370 159.680 ;
        RECT 125.610 159.660 125.750 177.700 ;
        RECT 126.530 177.000 126.670 178.380 ;
        RECT 126.470 176.680 126.730 177.000 ;
        RECT 126.010 176.000 126.270 176.320 ;
        RECT 126.070 171.220 126.210 176.000 ;
        RECT 126.530 173.260 126.670 176.680 ;
        RECT 126.470 172.940 126.730 173.260 ;
        RECT 126.010 170.900 126.270 171.220 ;
        RECT 126.070 168.840 126.210 170.900 ;
        RECT 126.010 168.520 126.270 168.840 ;
        RECT 126.470 167.500 126.730 167.820 ;
        RECT 126.530 165.780 126.670 167.500 ;
        RECT 126.470 165.460 126.730 165.780 ;
        RECT 126.530 162.380 126.670 165.460 ;
        RECT 126.470 162.060 126.730 162.380 ;
        RECT 125.550 159.340 125.810 159.660 ;
        RECT 124.630 154.240 124.890 154.560 ;
        RECT 124.170 152.200 124.430 152.520 ;
        RECT 124.230 148.100 124.370 152.200 ;
        RECT 124.690 152.180 124.830 154.240 ;
        RECT 125.090 154.130 125.350 154.220 ;
        RECT 125.610 154.130 125.750 159.340 ;
        RECT 126.470 159.000 126.730 159.320 ;
        RECT 126.010 158.660 126.270 158.980 ;
        RECT 126.070 157.960 126.210 158.660 ;
        RECT 126.530 157.960 126.670 159.000 ;
        RECT 126.010 157.640 126.270 157.960 ;
        RECT 126.470 157.640 126.730 157.960 ;
        RECT 126.010 156.620 126.270 156.940 ;
        RECT 126.990 156.795 127.130 182.260 ;
        RECT 127.910 182.260 128.510 182.400 ;
        RECT 127.390 161.720 127.650 162.040 ;
        RECT 125.090 153.990 125.750 154.130 ;
        RECT 125.090 153.900 125.350 153.990 ;
        RECT 124.630 151.860 124.890 152.180 ;
        RECT 125.090 151.520 125.350 151.840 ;
        RECT 125.150 150.675 125.290 151.520 ;
        RECT 125.080 150.305 125.360 150.675 ;
        RECT 124.630 148.800 124.890 149.120 ;
        RECT 124.170 147.780 124.430 148.100 ;
        RECT 124.170 145.740 124.430 146.060 ;
        RECT 124.230 141.640 124.370 145.740 ;
        RECT 124.690 144.360 124.830 148.800 ;
        RECT 125.610 146.400 125.750 153.990 ;
        RECT 125.550 146.080 125.810 146.400 ;
        RECT 124.630 144.040 124.890 144.360 ;
        RECT 125.550 143.360 125.810 143.680 ;
        RECT 124.170 141.320 124.430 141.640 ;
        RECT 125.610 140.620 125.750 143.360 ;
        RECT 125.550 140.300 125.810 140.620 ;
        RECT 124.170 138.600 124.430 138.920 ;
        RECT 124.230 133.480 124.370 138.600 ;
        RECT 125.610 137.560 125.750 140.300 ;
        RECT 126.070 138.920 126.210 156.620 ;
        RECT 126.920 156.425 127.200 156.795 ;
        RECT 126.470 153.560 126.730 153.880 ;
        RECT 126.530 150.820 126.670 153.560 ;
        RECT 126.990 151.500 127.130 156.425 ;
        RECT 127.450 154.900 127.590 161.720 ;
        RECT 127.910 157.280 128.050 182.260 ;
        RECT 128.310 178.040 128.570 178.360 ;
        RECT 128.370 175.300 128.510 178.040 ;
        RECT 129.690 177.700 129.950 178.020 ;
        RECT 129.750 177.000 129.890 177.700 ;
        RECT 129.690 176.680 129.950 177.000 ;
        RECT 129.230 175.835 129.490 175.980 ;
        RECT 129.220 175.465 129.500 175.835 ;
        RECT 128.310 174.980 128.570 175.300 ;
        RECT 128.370 165.440 128.510 174.980 ;
        RECT 129.680 172.745 129.960 173.115 ;
        RECT 129.750 171.560 129.890 172.745 ;
        RECT 129.690 171.240 129.950 171.560 ;
        RECT 130.210 170.280 130.350 188.580 ;
        RECT 131.060 188.385 131.340 188.755 ;
        RECT 131.130 187.540 131.270 188.385 ;
        RECT 131.070 187.220 131.330 187.540 ;
        RECT 130.600 184.305 130.880 184.675 ;
        RECT 130.610 184.160 130.870 184.305 ;
        RECT 131.070 183.880 131.330 184.140 ;
        RECT 130.670 183.820 131.330 183.880 ;
        RECT 130.670 183.740 131.270 183.820 ;
        RECT 130.670 182.440 130.810 183.740 ;
        RECT 131.070 183.140 131.330 183.460 ;
        RECT 130.610 182.120 130.870 182.440 ;
        RECT 130.610 180.420 130.870 180.740 ;
        RECT 130.670 171.560 130.810 180.420 ;
        RECT 131.130 179.235 131.270 183.140 ;
        RECT 131.060 178.865 131.340 179.235 ;
        RECT 131.590 178.440 131.730 191.300 ;
        RECT 132.050 187.880 132.190 192.070 ;
        RECT 132.450 191.980 132.710 192.070 ;
        RECT 132.970 188.810 133.110 196.740 ;
        RECT 133.460 196.120 133.600 197.170 ;
        RECT 133.430 195.980 133.600 196.120 ;
        RECT 133.430 194.340 133.570 195.980 ;
        RECT 133.890 195.440 134.030 198.440 ;
        RECT 134.350 198.275 134.490 200.140 ;
        RECT 134.280 198.160 134.560 198.275 ;
        RECT 134.280 198.020 135.410 198.160 ;
        RECT 134.280 197.905 134.560 198.020 ;
        RECT 135.270 197.400 135.410 198.020 ;
        RECT 134.290 197.080 134.550 197.400 ;
        RECT 135.210 197.080 135.470 197.400 ;
        RECT 134.350 195.950 134.490 197.080 ;
        RECT 134.770 196.205 136.650 196.575 ;
        RECT 134.350 195.810 134.950 195.950 ;
        RECT 133.890 195.360 134.490 195.440 ;
        RECT 133.890 195.300 134.550 195.360 ;
        RECT 134.290 195.040 134.550 195.300 ;
        RECT 134.810 194.875 134.950 195.810 ;
        RECT 135.210 195.720 135.470 196.040 ;
        RECT 134.740 194.505 135.020 194.875 ;
        RECT 135.270 194.680 135.410 195.720 ;
        RECT 135.210 194.360 135.470 194.680 ;
        RECT 133.370 194.020 133.630 194.340 ;
        RECT 132.890 188.670 133.110 188.810 ;
        RECT 132.890 187.960 133.030 188.670 ;
        RECT 131.990 187.560 132.250 187.880 ;
        RECT 132.450 187.560 132.710 187.880 ;
        RECT 132.890 187.820 133.110 187.960 ;
        RECT 133.430 187.880 133.570 194.020 ;
        RECT 137.110 193.400 137.250 200.480 ;
        RECT 137.510 199.460 137.770 199.780 ;
        RECT 137.570 198.080 137.710 199.460 ;
        RECT 137.510 197.760 137.770 198.080 ;
        RECT 138.950 197.400 139.090 202.180 ;
        RECT 139.870 201.050 140.010 203.540 ;
        RECT 140.790 203.520 140.930 207.620 ;
        RECT 140.730 203.200 140.990 203.520 ;
        RECT 142.170 203.180 142.310 207.960 ;
        RECT 144.470 206.920 144.610 209.455 ;
        RECT 144.410 206.600 144.670 206.920 ;
        RECT 148.610 206.240 148.750 209.455 ;
        RECT 149.010 206.600 149.270 206.920 ;
        RECT 148.550 205.920 148.810 206.240 ;
        RECT 144.870 205.580 145.130 205.900 ;
        RECT 143.490 205.240 143.750 205.560 ;
        RECT 142.110 202.860 142.370 203.180 ;
        RECT 140.270 201.050 140.530 201.140 ;
        RECT 139.870 200.910 140.530 201.050 ;
        RECT 139.350 199.460 139.610 199.780 ;
        RECT 139.410 198.080 139.550 199.460 ;
        RECT 139.350 197.760 139.610 198.080 ;
        RECT 137.510 197.080 137.770 197.400 ;
        RECT 138.890 197.080 139.150 197.400 ;
        RECT 137.570 196.040 137.710 197.080 ;
        RECT 139.350 196.740 139.610 197.060 ;
        RECT 137.510 195.720 137.770 196.040 ;
        RECT 137.500 195.185 137.780 195.555 ;
        RECT 137.570 194.680 137.710 195.185 ;
        RECT 138.890 195.040 139.150 195.360 ;
        RECT 137.970 194.700 138.230 195.020 ;
        RECT 137.510 194.360 137.770 194.680 ;
        RECT 136.190 193.260 137.250 193.400 ;
        RECT 136.190 192.040 136.330 193.260 ;
        RECT 138.030 192.640 138.170 194.700 ;
        RECT 138.430 194.020 138.690 194.340 ;
        RECT 137.050 192.320 137.310 192.640 ;
        RECT 137.510 192.320 137.770 192.640 ;
        RECT 137.970 192.320 138.230 192.640 ;
        RECT 133.890 191.900 136.330 192.040 ;
        RECT 131.990 184.160 132.250 184.480 ;
        RECT 132.050 183.460 132.190 184.160 ;
        RECT 131.990 183.140 132.250 183.460 ;
        RECT 131.990 180.420 132.250 180.740 ;
        RECT 132.050 179.040 132.190 180.420 ;
        RECT 131.990 178.720 132.250 179.040 ;
        RECT 131.590 178.300 132.190 178.440 ;
        RECT 131.530 177.700 131.790 178.020 ;
        RECT 131.590 176.320 131.730 177.700 ;
        RECT 131.530 176.000 131.790 176.320 ;
        RECT 132.050 175.040 132.190 178.300 ;
        RECT 132.510 177.000 132.650 187.560 ;
        RECT 132.450 176.680 132.710 177.000 ;
        RECT 132.050 174.900 132.650 175.040 ;
        RECT 131.990 173.960 132.250 174.280 ;
        RECT 131.530 173.280 131.790 173.600 ;
        RECT 130.610 171.470 130.870 171.560 ;
        RECT 130.610 171.330 131.270 171.470 ;
        RECT 130.610 171.240 130.870 171.330 ;
        RECT 129.690 169.880 129.950 170.200 ;
        RECT 130.210 170.140 130.810 170.280 ;
        RECT 129.750 168.840 129.890 169.880 ;
        RECT 130.150 169.540 130.410 169.860 ;
        RECT 129.690 168.520 129.950 168.840 ;
        RECT 129.230 167.730 129.490 167.820 ;
        RECT 130.210 167.730 130.350 169.540 ;
        RECT 129.230 167.590 130.350 167.730 ;
        RECT 129.230 167.500 129.490 167.590 ;
        RECT 129.690 166.820 129.950 167.140 ;
        RECT 130.150 166.820 130.410 167.140 ;
        RECT 128.310 165.120 128.570 165.440 ;
        RECT 129.230 164.440 129.490 164.760 ;
        RECT 129.290 162.720 129.430 164.440 ;
        RECT 129.750 163.400 129.890 166.820 ;
        RECT 130.210 165.780 130.350 166.820 ;
        RECT 130.150 165.635 130.410 165.780 ;
        RECT 130.140 165.265 130.420 165.635 ;
        RECT 129.690 163.080 129.950 163.400 ;
        RECT 130.670 162.800 130.810 170.140 ;
        RECT 131.130 167.480 131.270 171.330 ;
        RECT 131.070 167.160 131.330 167.480 ;
        RECT 131.130 164.420 131.270 167.160 ;
        RECT 131.590 165.440 131.730 173.280 ;
        RECT 132.050 171.560 132.190 173.960 ;
        RECT 131.990 171.240 132.250 171.560 ;
        RECT 131.980 167.985 132.260 168.355 ;
        RECT 132.050 167.820 132.190 167.985 ;
        RECT 131.990 167.500 132.250 167.820 ;
        RECT 131.990 166.820 132.250 167.140 ;
        RECT 132.050 165.560 132.190 166.820 ;
        RECT 131.530 165.120 131.790 165.440 ;
        RECT 131.990 165.240 132.250 165.560 ;
        RECT 131.990 164.840 132.250 165.100 ;
        RECT 131.590 164.780 132.250 164.840 ;
        RECT 131.590 164.700 132.190 164.780 ;
        RECT 131.070 164.100 131.330 164.420 ;
        RECT 131.590 163.480 131.730 164.700 ;
        RECT 129.230 162.400 129.490 162.720 ;
        RECT 129.750 162.660 130.810 162.800 ;
        RECT 128.770 161.380 129.030 161.700 ;
        RECT 128.830 160.000 128.970 161.380 ;
        RECT 128.770 159.680 129.030 160.000 ;
        RECT 129.750 159.400 129.890 162.660 ;
        RECT 130.670 160.000 130.810 162.660 ;
        RECT 131.130 163.340 131.730 163.480 ;
        RECT 131.130 162.235 131.270 163.340 ;
        RECT 131.060 161.865 131.340 162.235 ;
        RECT 130.610 159.680 130.870 160.000 ;
        RECT 128.370 159.260 129.890 159.400 ;
        RECT 127.850 156.960 128.110 157.280 ;
        RECT 127.390 154.580 127.650 154.900 ;
        RECT 126.930 151.410 127.190 151.500 ;
        RECT 126.930 151.270 127.590 151.410 ;
        RECT 126.930 151.180 127.190 151.270 ;
        RECT 126.470 150.500 126.730 150.820 ;
        RECT 126.930 148.120 127.190 148.440 ;
        RECT 126.470 147.780 126.730 148.100 ;
        RECT 126.530 144.020 126.670 147.780 ;
        RECT 126.990 144.020 127.130 148.120 ;
        RECT 127.450 146.480 127.590 151.270 ;
        RECT 127.910 148.100 128.050 156.960 ;
        RECT 127.850 147.955 128.110 148.100 ;
        RECT 127.840 147.585 128.120 147.955 ;
        RECT 127.450 146.340 128.050 146.480 ;
        RECT 127.390 145.740 127.650 146.060 ;
        RECT 127.450 144.360 127.590 145.740 ;
        RECT 127.390 144.040 127.650 144.360 ;
        RECT 126.470 143.700 126.730 144.020 ;
        RECT 126.930 143.700 127.190 144.020 ;
        RECT 126.010 138.600 126.270 138.920 ;
        RECT 127.910 138.150 128.050 146.340 ;
        RECT 128.370 144.360 128.510 159.260 ;
        RECT 129.690 158.660 129.950 158.980 ;
        RECT 129.750 157.960 129.890 158.660 ;
        RECT 128.770 157.640 129.030 157.960 ;
        RECT 129.690 157.640 129.950 157.960 ;
        RECT 130.150 157.640 130.410 157.960 ;
        RECT 128.830 157.475 128.970 157.640 ;
        RECT 128.760 157.360 129.040 157.475 ;
        RECT 128.760 157.220 129.890 157.360 ;
        RECT 128.760 157.105 129.040 157.220 ;
        RECT 129.750 156.940 129.890 157.220 ;
        RECT 129.690 156.620 129.950 156.940 ;
        RECT 128.770 153.220 129.030 153.540 ;
        RECT 128.830 151.160 128.970 153.220 ;
        RECT 129.230 152.200 129.490 152.520 ;
        RECT 129.290 151.500 129.430 152.200 ;
        RECT 130.210 151.750 130.350 157.640 ;
        RECT 130.610 153.220 130.870 153.540 ;
        RECT 129.750 151.610 130.350 151.750 ;
        RECT 129.230 151.180 129.490 151.500 ;
        RECT 128.770 150.840 129.030 151.160 ;
        RECT 129.230 150.500 129.490 150.820 ;
        RECT 128.760 148.945 129.040 149.315 ;
        RECT 129.290 149.120 129.430 150.500 ;
        RECT 128.830 146.400 128.970 148.945 ;
        RECT 129.230 148.800 129.490 149.120 ;
        RECT 128.770 146.080 129.030 146.400 ;
        RECT 128.770 145.400 129.030 145.720 ;
        RECT 128.830 144.360 128.970 145.400 ;
        RECT 128.310 144.040 128.570 144.360 ;
        RECT 128.770 144.040 129.030 144.360 ;
        RECT 129.290 143.340 129.430 148.800 ;
        RECT 129.230 143.020 129.490 143.340 ;
        RECT 129.290 140.960 129.430 143.020 ;
        RECT 129.230 140.640 129.490 140.960 ;
        RECT 128.770 138.150 129.030 138.240 ;
        RECT 127.910 138.010 129.030 138.150 ;
        RECT 129.220 138.065 129.500 138.435 ;
        RECT 128.770 137.920 129.030 138.010 ;
        RECT 127.390 137.580 127.650 137.900 ;
        RECT 125.550 137.240 125.810 137.560 ;
        RECT 126.930 137.240 127.190 137.560 ;
        RECT 126.990 136.200 127.130 137.240 ;
        RECT 126.930 135.880 127.190 136.200 ;
        RECT 126.930 134.860 127.190 135.180 ;
        RECT 124.170 133.160 124.430 133.480 ;
        RECT 124.170 132.480 124.430 132.800 ;
        RECT 124.230 125.320 124.370 132.480 ;
        RECT 124.620 130.160 124.900 130.275 ;
        RECT 124.620 130.020 125.290 130.160 ;
        RECT 124.620 129.905 124.900 130.020 ;
        RECT 125.150 127.700 125.290 130.020 ;
        RECT 125.090 127.380 125.350 127.700 ;
        RECT 125.550 126.020 125.810 126.340 ;
        RECT 126.010 126.020 126.270 126.340 ;
        RECT 123.710 125.000 123.970 125.320 ;
        RECT 124.170 125.000 124.430 125.320 ;
        RECT 123.250 123.640 123.510 123.960 ;
        RECT 123.710 123.640 123.970 123.960 ;
        RECT 118.650 123.300 118.910 123.620 ;
        RECT 118.710 122.230 118.850 123.300 ;
        RECT 119.770 122.765 121.650 123.135 ;
        RECT 122.390 122.370 122.990 122.510 ;
        RECT 122.390 122.230 122.530 122.370 ;
        RECT 118.190 120.920 118.450 121.240 ;
        RECT 118.640 120.230 118.920 122.230 ;
        RECT 122.320 120.230 122.600 122.230 ;
        RECT 122.850 122.000 122.990 122.370 ;
        RECT 123.770 122.000 123.910 123.640 ;
        RECT 125.090 123.300 125.350 123.620 ;
        RECT 125.150 122.260 125.290 123.300 ;
        RECT 122.850 121.860 123.910 122.000 ;
        RECT 125.090 121.940 125.350 122.260 ;
        RECT 125.610 121.240 125.750 126.020 ;
        RECT 126.070 122.230 126.210 126.020 ;
        RECT 126.990 124.300 127.130 134.860 ;
        RECT 127.450 126.340 127.590 137.580 ;
        RECT 129.290 137.220 129.430 138.065 ;
        RECT 129.230 136.900 129.490 137.220 ;
        RECT 128.310 134.860 128.570 135.180 ;
        RECT 128.370 132.120 128.510 134.860 ;
        RECT 128.310 131.800 128.570 132.120 ;
        RECT 128.310 130.440 128.570 130.760 ;
        RECT 127.850 129.760 128.110 130.080 ;
        RECT 127.390 126.020 127.650 126.340 ;
        RECT 126.930 123.980 127.190 124.300 ;
        RECT 125.550 120.920 125.810 121.240 ;
        RECT 126.000 120.230 126.280 122.230 ;
        RECT 127.910 121.580 128.050 129.760 ;
        RECT 128.370 127.020 128.510 130.440 ;
        RECT 128.770 129.080 129.030 129.400 ;
        RECT 128.830 127.020 128.970 129.080 ;
        RECT 129.290 128.970 129.430 136.900 ;
        RECT 129.750 135.035 129.890 151.610 ;
        RECT 130.670 148.520 130.810 153.220 ;
        RECT 131.130 149.315 131.270 161.865 ;
        RECT 132.510 157.960 132.650 174.900 ;
        RECT 132.450 157.640 132.710 157.960 ;
        RECT 132.450 156.620 132.710 156.940 ;
        RECT 131.980 151.665 132.260 152.035 ;
        RECT 132.050 151.500 132.190 151.665 ;
        RECT 131.990 151.180 132.250 151.500 ;
        RECT 131.060 149.200 131.340 149.315 ;
        RECT 131.060 149.060 131.730 149.200 ;
        RECT 131.060 148.945 131.340 149.060 ;
        RECT 130.210 148.380 130.810 148.520 ;
        RECT 130.210 138.920 130.350 148.380 ;
        RECT 130.610 147.780 130.870 148.100 ;
        RECT 130.150 138.600 130.410 138.920 ;
        RECT 130.670 135.520 130.810 147.780 ;
        RECT 131.070 145.400 131.330 145.720 ;
        RECT 130.610 135.200 130.870 135.520 ;
        RECT 129.680 134.665 129.960 135.035 ;
        RECT 129.750 133.140 129.890 134.665 ;
        RECT 129.690 132.820 129.950 133.140 ;
        RECT 130.610 132.480 130.870 132.800 ;
        RECT 130.670 132.315 130.810 132.480 ;
        RECT 130.150 131.800 130.410 132.120 ;
        RECT 130.600 131.945 130.880 132.315 ;
        RECT 130.210 130.420 130.350 131.800 ;
        RECT 130.150 130.100 130.410 130.420 ;
        RECT 131.130 130.080 131.270 145.400 ;
        RECT 131.590 144.440 131.730 149.060 ;
        RECT 131.990 148.800 132.250 149.120 ;
        RECT 132.050 148.635 132.190 148.800 ;
        RECT 131.980 148.265 132.260 148.635 ;
        RECT 132.510 148.440 132.650 156.620 ;
        RECT 132.970 151.410 133.110 187.820 ;
        RECT 133.370 187.560 133.630 187.880 ;
        RECT 133.890 186.180 134.030 191.900 ;
        RECT 134.770 190.765 136.650 191.135 ;
        RECT 136.590 190.510 136.850 190.600 ;
        RECT 137.110 190.510 137.250 192.320 ;
        RECT 136.590 190.370 137.250 190.510 ;
        RECT 136.590 190.280 136.850 190.370 ;
        RECT 137.570 189.920 137.710 192.320 ;
        RECT 138.030 191.960 138.170 192.320 ;
        RECT 137.970 191.640 138.230 191.960 ;
        RECT 138.030 190.260 138.170 191.640 ;
        RECT 138.490 190.600 138.630 194.020 ;
        RECT 138.430 190.280 138.690 190.600 ;
        RECT 137.970 189.940 138.230 190.260 ;
        RECT 137.510 189.600 137.770 189.920 ;
        RECT 138.430 188.920 138.690 189.240 ;
        RECT 137.050 188.580 137.310 188.900 ;
        RECT 137.960 188.640 138.240 188.755 ;
        RECT 138.490 188.640 138.630 188.920 ;
        RECT 134.750 187.450 135.010 187.540 ;
        RECT 134.350 187.310 135.010 187.450 ;
        RECT 133.830 185.860 134.090 186.180 ;
        RECT 134.350 185.160 134.490 187.310 ;
        RECT 134.750 187.220 135.010 187.310 ;
        RECT 137.110 187.200 137.250 188.580 ;
        RECT 137.960 188.500 138.630 188.640 ;
        RECT 137.960 188.385 138.240 188.500 ;
        RECT 138.950 187.960 139.090 195.040 ;
        RECT 138.490 187.820 139.090 187.960 ;
        RECT 137.970 187.450 138.230 187.540 ;
        RECT 137.570 187.310 138.230 187.450 ;
        RECT 137.050 186.880 137.310 187.200 ;
        RECT 134.770 185.325 136.650 185.695 ;
        RECT 134.290 184.840 134.550 185.160 ;
        RECT 133.370 183.480 133.630 183.800 ;
        RECT 133.430 179.720 133.570 183.480 ;
        RECT 134.350 182.440 134.490 184.840 ;
        RECT 136.590 184.050 136.850 184.140 ;
        RECT 137.570 184.050 137.710 187.310 ;
        RECT 137.970 187.220 138.230 187.310 ;
        RECT 136.590 183.910 137.710 184.050 ;
        RECT 137.970 184.050 138.230 184.140 ;
        RECT 138.490 184.050 138.630 187.820 ;
        RECT 139.410 184.560 139.550 196.740 ;
        RECT 139.870 195.360 140.010 200.910 ;
        RECT 140.270 200.820 140.530 200.910 ;
        RECT 142.170 200.120 142.310 202.860 ;
        RECT 143.030 202.520 143.290 202.840 ;
        RECT 143.090 200.800 143.230 202.520 ;
        RECT 143.030 200.480 143.290 200.800 ;
        RECT 142.110 199.800 142.370 200.120 ;
        RECT 143.090 198.760 143.230 200.480 ;
        RECT 143.030 198.440 143.290 198.760 ;
        RECT 140.730 197.420 140.990 197.740 ;
        RECT 140.790 195.700 140.930 197.420 ;
        RECT 143.090 196.040 143.230 198.440 ;
        RECT 143.550 197.060 143.690 205.240 ;
        RECT 144.410 202.180 144.670 202.500 ;
        RECT 144.470 200.460 144.610 202.180 ;
        RECT 144.410 200.140 144.670 200.460 ;
        RECT 143.950 199.800 144.210 200.120 ;
        RECT 144.010 198.080 144.150 199.800 ;
        RECT 143.950 197.760 144.210 198.080 ;
        RECT 143.490 196.740 143.750 197.060 ;
        RECT 144.930 196.040 145.070 205.580 ;
        RECT 147.170 204.900 147.430 205.220 ;
        RECT 147.230 203.180 147.370 204.900 ;
        RECT 149.070 204.200 149.210 206.600 ;
        RECT 149.770 204.365 151.650 204.735 ;
        RECT 149.010 203.880 149.270 204.200 ;
        RECT 148.090 203.200 148.350 203.520 ;
        RECT 147.170 202.860 147.430 203.180 ;
        RECT 145.790 202.180 146.050 202.500 ;
        RECT 145.850 200.460 145.990 202.180 ;
        RECT 145.790 200.140 146.050 200.460 ;
        RECT 146.710 199.800 146.970 200.120 ;
        RECT 145.330 199.460 145.590 199.780 ;
        RECT 145.790 199.460 146.050 199.780 ;
        RECT 145.390 197.400 145.530 199.460 ;
        RECT 145.850 198.760 145.990 199.460 ;
        RECT 146.770 198.760 146.910 199.800 ;
        RECT 145.790 198.440 146.050 198.760 ;
        RECT 146.710 198.440 146.970 198.760 ;
        RECT 145.330 197.080 145.590 197.400 ;
        RECT 143.030 195.720 143.290 196.040 ;
        RECT 144.870 195.720 145.130 196.040 ;
        RECT 140.730 195.380 140.990 195.700 ;
        RECT 141.650 195.380 141.910 195.700 ;
        RECT 139.810 195.040 140.070 195.360 ;
        RECT 139.870 192.640 140.010 195.040 ;
        RECT 140.730 194.930 140.990 195.020 ;
        RECT 141.710 194.930 141.850 195.380 ;
        RECT 140.730 194.790 141.850 194.930 ;
        RECT 140.730 194.700 140.990 194.790 ;
        RECT 147.230 194.760 147.370 202.860 ;
        RECT 148.150 197.740 148.290 203.200 ;
        RECT 148.550 202.180 148.810 202.500 ;
        RECT 148.610 198.760 148.750 202.180 ;
        RECT 149.770 198.925 151.650 199.295 ;
        RECT 148.550 198.440 148.810 198.760 ;
        RECT 148.090 197.420 148.350 197.740 ;
        RECT 147.630 196.740 147.890 197.060 ;
        RECT 152.230 196.740 152.490 197.060 ;
        RECT 146.310 194.620 147.370 194.760 ;
        RECT 139.810 192.320 140.070 192.640 ;
        RECT 139.870 189.580 140.010 192.320 ;
        RECT 139.810 189.260 140.070 189.580 ;
        RECT 141.650 188.920 141.910 189.240 ;
        RECT 140.730 186.540 140.990 186.860 ;
        RECT 140.790 185.160 140.930 186.540 ;
        RECT 141.710 186.520 141.850 188.920 ;
        RECT 142.570 186.880 142.830 187.200 ;
        RECT 145.790 186.880 146.050 187.200 ;
        RECT 141.650 186.430 141.910 186.520 ;
        RECT 141.250 186.290 141.910 186.430 ;
        RECT 140.730 184.840 140.990 185.160 ;
        RECT 139.410 184.420 140.470 184.560 ;
        RECT 137.970 183.910 138.630 184.050 ;
        RECT 136.590 183.820 136.850 183.910 ;
        RECT 137.970 183.820 138.230 183.910 ;
        RECT 139.350 183.820 139.610 184.140 ;
        RECT 136.130 183.140 136.390 183.460 ;
        RECT 134.290 182.120 134.550 182.440 ;
        RECT 133.370 179.400 133.630 179.720 ;
        RECT 133.430 178.700 133.570 179.400 ;
        RECT 133.830 179.060 134.090 179.380 ;
        RECT 133.370 178.380 133.630 178.700 ;
        RECT 133.370 176.680 133.630 177.000 ;
        RECT 133.430 153.540 133.570 176.680 ;
        RECT 133.890 174.280 134.030 179.060 ;
        RECT 133.830 173.960 134.090 174.280 ;
        RECT 134.350 168.160 134.490 182.120 ;
        RECT 136.190 182.100 136.330 183.140 ;
        RECT 136.130 181.780 136.390 182.100 ;
        RECT 137.050 181.440 137.310 181.760 ;
        RECT 137.510 181.440 137.770 181.760 ;
        RECT 134.770 179.885 136.650 180.255 ;
        RECT 137.110 179.630 137.250 181.440 ;
        RECT 136.650 179.490 137.250 179.630 ;
        RECT 136.650 178.020 136.790 179.490 ;
        RECT 137.050 178.720 137.310 179.040 ;
        RECT 136.590 177.700 136.850 178.020 ;
        RECT 136.650 175.890 136.790 177.700 ;
        RECT 137.110 176.400 137.250 178.720 ;
        RECT 137.570 177.000 137.710 181.440 ;
        RECT 137.510 176.680 137.770 177.000 ;
        RECT 137.110 176.260 137.710 176.400 ;
        RECT 136.120 175.465 136.400 175.835 ;
        RECT 136.650 175.750 137.250 175.890 ;
        RECT 136.130 175.320 136.390 175.465 ;
        RECT 134.770 174.445 136.650 174.815 ;
        RECT 134.740 173.425 135.020 173.795 ;
        RECT 134.810 173.260 134.950 173.425 ;
        RECT 137.110 173.260 137.250 175.750 ;
        RECT 137.570 174.280 137.710 176.260 ;
        RECT 137.510 173.960 137.770 174.280 ;
        RECT 138.030 173.600 138.170 183.820 ;
        RECT 138.890 183.480 139.150 183.800 ;
        RECT 138.430 176.000 138.690 176.320 ;
        RECT 137.970 173.280 138.230 173.600 ;
        RECT 138.490 173.260 138.630 176.000 ;
        RECT 134.750 173.170 135.010 173.260 ;
        RECT 134.750 173.030 135.870 173.170 ;
        RECT 134.750 172.940 135.010 173.030 ;
        RECT 135.730 172.580 135.870 173.030 ;
        RECT 137.050 172.940 137.310 173.260 ;
        RECT 138.430 172.940 138.690 173.260 ;
        RECT 135.670 172.260 135.930 172.580 ;
        RECT 135.730 170.880 135.870 172.260 ;
        RECT 137.050 171.240 137.310 171.560 ;
        RECT 135.670 170.560 135.930 170.880 ;
        RECT 134.770 169.005 136.650 169.375 ;
        RECT 134.290 167.840 134.550 168.160 ;
        RECT 137.110 166.120 137.250 171.240 ;
        RECT 137.510 170.220 137.770 170.540 ;
        RECT 137.570 168.840 137.710 170.220 ;
        RECT 137.510 168.520 137.770 168.840 ;
        RECT 137.970 166.820 138.230 167.140 ;
        RECT 137.050 165.800 137.310 166.120 ;
        RECT 133.830 165.460 134.090 165.780 ;
        RECT 137.510 165.460 137.770 165.780 ;
        RECT 133.890 164.955 134.030 165.460 ;
        RECT 137.050 165.120 137.310 165.440 ;
        RECT 133.820 164.585 134.100 164.955 ;
        RECT 134.770 163.565 136.650 163.935 ;
        RECT 133.830 163.080 134.090 163.400 ;
        RECT 133.890 160.000 134.030 163.080 ;
        RECT 137.110 162.720 137.250 165.120 ;
        RECT 137.050 162.400 137.310 162.720 ;
        RECT 135.670 161.380 135.930 161.700 ;
        RECT 136.130 161.380 136.390 161.700 ;
        RECT 137.050 161.380 137.310 161.700 ;
        RECT 135.730 160.000 135.870 161.380 ;
        RECT 136.190 160.000 136.330 161.380 ;
        RECT 137.110 160.680 137.250 161.380 ;
        RECT 137.050 160.360 137.310 160.680 ;
        RECT 137.110 160.000 137.250 160.360 ;
        RECT 133.830 159.910 134.090 160.000 ;
        RECT 133.830 159.770 134.490 159.910 ;
        RECT 133.830 159.680 134.090 159.770 ;
        RECT 133.830 155.940 134.090 156.260 ;
        RECT 133.370 153.220 133.630 153.540 ;
        RECT 132.970 151.270 133.570 151.410 ;
        RECT 132.900 149.625 133.180 149.995 ;
        RECT 132.450 148.120 132.710 148.440 ;
        RECT 131.980 147.585 132.260 147.955 ;
        RECT 132.050 147.080 132.190 147.585 ;
        RECT 131.990 146.760 132.250 147.080 ;
        RECT 132.440 146.905 132.720 147.275 ;
        RECT 132.510 146.740 132.650 146.905 ;
        RECT 132.450 146.420 132.710 146.740 ;
        RECT 132.510 146.060 132.650 146.420 ;
        RECT 132.450 145.740 132.710 146.060 ;
        RECT 131.590 144.300 132.190 144.440 ;
        RECT 131.530 143.020 131.790 143.340 ;
        RECT 131.590 133.140 131.730 143.020 ;
        RECT 132.050 140.960 132.190 144.300 ;
        RECT 131.990 140.640 132.250 140.960 ;
        RECT 132.450 137.580 132.710 137.900 ;
        RECT 132.510 135.860 132.650 137.580 ;
        RECT 132.970 136.395 133.110 149.625 ;
        RECT 132.900 136.025 133.180 136.395 ;
        RECT 132.450 135.540 132.710 135.860 ;
        RECT 132.910 135.200 133.170 135.520 ;
        RECT 131.530 132.820 131.790 133.140 ;
        RECT 131.990 132.030 132.250 132.120 ;
        RECT 131.590 131.890 132.250 132.030 ;
        RECT 131.070 129.760 131.330 130.080 ;
        RECT 129.690 129.595 129.950 129.740 ;
        RECT 129.680 129.225 129.960 129.595 ;
        RECT 130.150 129.420 130.410 129.740 ;
        RECT 130.210 128.970 130.350 129.420 ;
        RECT 129.290 128.830 130.350 128.970 ;
        RECT 130.210 128.040 130.350 128.830 ;
        RECT 131.070 128.740 131.330 129.060 ;
        RECT 130.150 127.720 130.410 128.040 ;
        RECT 130.610 127.720 130.870 128.040 ;
        RECT 130.670 127.270 130.810 127.720 ;
        RECT 130.210 127.130 130.810 127.270 ;
        RECT 128.310 126.700 128.570 127.020 ;
        RECT 128.770 126.700 129.030 127.020 ;
        RECT 130.210 124.300 130.350 127.130 ;
        RECT 131.130 126.760 131.270 128.740 ;
        RECT 131.590 127.360 131.730 131.890 ;
        RECT 131.990 131.800 132.250 131.890 ;
        RECT 131.980 129.905 132.260 130.275 ;
        RECT 131.530 127.040 131.790 127.360 ;
        RECT 132.050 127.270 132.190 129.905 ;
        RECT 132.970 127.360 133.110 135.200 ;
        RECT 133.430 130.955 133.570 151.270 ;
        RECT 133.890 143.680 134.030 155.940 ;
        RECT 134.350 154.900 134.490 159.770 ;
        RECT 135.670 159.680 135.930 160.000 ;
        RECT 136.130 159.680 136.390 160.000 ;
        RECT 137.050 159.680 137.310 160.000 ;
        RECT 135.730 159.320 135.870 159.680 ;
        RECT 135.670 159.000 135.930 159.320 ;
        RECT 137.110 158.980 137.250 159.680 ;
        RECT 137.050 158.660 137.310 158.980 ;
        RECT 134.770 158.125 136.650 158.495 ;
        RECT 137.050 157.640 137.310 157.960 ;
        RECT 134.290 154.580 134.550 154.900 ;
        RECT 134.350 149.120 134.490 154.580 ;
        RECT 134.770 152.685 136.650 153.055 ;
        RECT 137.110 151.840 137.250 157.640 ;
        RECT 137.050 151.520 137.310 151.840 ;
        RECT 136.120 150.985 136.400 151.355 ;
        RECT 134.290 148.800 134.550 149.120 ;
        RECT 135.660 148.945 135.940 149.315 ;
        RECT 136.190 149.120 136.330 150.985 ;
        RECT 135.730 148.440 135.870 148.945 ;
        RECT 136.130 148.800 136.390 149.120 ;
        RECT 137.050 148.800 137.310 149.120 ;
        RECT 135.670 148.120 135.930 148.440 ;
        RECT 134.290 147.780 134.550 148.100 ;
        RECT 133.830 143.360 134.090 143.680 ;
        RECT 133.830 140.300 134.090 140.620 ;
        RECT 133.890 134.500 134.030 140.300 ;
        RECT 134.350 138.920 134.490 147.780 ;
        RECT 134.770 147.245 136.650 147.615 ;
        RECT 137.110 146.990 137.250 148.800 ;
        RECT 136.650 146.850 137.250 146.990 ;
        RECT 136.650 146.060 136.790 146.850 ;
        RECT 137.570 146.650 137.710 165.460 ;
        RECT 137.110 146.510 137.710 146.650 ;
        RECT 134.750 145.915 135.010 146.060 ;
        RECT 134.740 145.545 135.020 145.915 ;
        RECT 136.590 145.740 136.850 146.060 ;
        RECT 134.770 141.805 136.650 142.175 ;
        RECT 137.110 140.620 137.250 146.510 ;
        RECT 138.030 143.340 138.170 166.820 ;
        RECT 138.490 155.320 138.630 172.940 ;
        RECT 138.950 162.380 139.090 183.480 ;
        RECT 139.410 181.080 139.550 183.820 ;
        RECT 139.350 180.760 139.610 181.080 ;
        RECT 139.410 176.515 139.550 180.760 ;
        RECT 139.800 178.185 140.080 178.555 ;
        RECT 139.870 178.020 140.010 178.185 ;
        RECT 139.810 177.700 140.070 178.020 ;
        RECT 139.340 176.145 139.620 176.515 ;
        RECT 139.350 175.320 139.610 175.640 ;
        RECT 139.410 168.500 139.550 175.320 ;
        RECT 139.810 172.600 140.070 172.920 ;
        RECT 139.350 168.180 139.610 168.500 ;
        RECT 139.870 167.820 140.010 172.600 ;
        RECT 140.330 170.880 140.470 184.420 ;
        RECT 140.730 181.780 140.990 182.100 ;
        RECT 140.790 175.980 140.930 181.780 ;
        RECT 140.730 175.660 140.990 175.980 ;
        RECT 140.730 174.980 140.990 175.300 ;
        RECT 140.270 170.560 140.530 170.880 ;
        RECT 139.350 167.500 139.610 167.820 ;
        RECT 139.810 167.500 140.070 167.820 ;
        RECT 140.270 167.500 140.530 167.820 ;
        RECT 139.410 166.120 139.550 167.500 ;
        RECT 139.810 166.820 140.070 167.140 ;
        RECT 139.350 165.800 139.610 166.120 ;
        RECT 138.890 162.060 139.150 162.380 ;
        RECT 139.870 161.700 140.010 166.820 ;
        RECT 140.330 164.760 140.470 167.500 ;
        RECT 140.790 167.140 140.930 174.980 ;
        RECT 140.730 166.820 140.990 167.140 ;
        RECT 140.730 165.120 140.990 165.440 ;
        RECT 140.270 164.440 140.530 164.760 ;
        RECT 138.890 161.380 139.150 161.700 ;
        RECT 139.350 161.380 139.610 161.700 ;
        RECT 139.810 161.380 140.070 161.700 ;
        RECT 138.950 160.000 139.090 161.380 ;
        RECT 138.890 159.680 139.150 160.000 ;
        RECT 138.950 156.115 139.090 159.680 ;
        RECT 139.410 156.940 139.550 161.380 ;
        RECT 139.800 157.105 140.080 157.475 ;
        RECT 139.810 156.960 140.070 157.105 ;
        RECT 139.350 156.620 139.610 156.940 ;
        RECT 138.880 155.745 139.160 156.115 ;
        RECT 138.490 155.180 139.550 155.320 ;
        RECT 138.430 154.580 138.690 154.900 ;
        RECT 138.490 148.635 138.630 154.580 ;
        RECT 138.890 151.180 139.150 151.500 ;
        RECT 138.950 150.675 139.090 151.180 ;
        RECT 138.880 150.305 139.160 150.675 ;
        RECT 138.420 148.265 138.700 148.635 ;
        RECT 138.490 148.100 138.630 148.265 ;
        RECT 138.950 148.100 139.090 150.305 ;
        RECT 138.430 147.780 138.690 148.100 ;
        RECT 138.890 147.780 139.150 148.100 ;
        RECT 138.430 146.080 138.690 146.400 ;
        RECT 137.510 143.020 137.770 143.340 ;
        RECT 137.970 143.020 138.230 143.340 ;
        RECT 137.050 140.300 137.310 140.620 ;
        RECT 135.210 139.960 135.470 140.280 ;
        RECT 134.750 139.620 135.010 139.940 ;
        RECT 134.290 138.600 134.550 138.920 ;
        RECT 134.810 137.640 134.950 139.620 ;
        RECT 135.270 138.920 135.410 139.960 ;
        RECT 135.670 139.620 135.930 139.940 ;
        RECT 135.210 138.600 135.470 138.920 ;
        RECT 135.730 137.900 135.870 139.620 ;
        RECT 137.110 138.920 137.250 140.300 ;
        RECT 137.570 138.920 137.710 143.020 ;
        RECT 137.970 141.320 138.230 141.640 ;
        RECT 137.050 138.600 137.310 138.920 ;
        RECT 137.510 138.600 137.770 138.920 ;
        RECT 138.030 138.240 138.170 141.320 ;
        RECT 138.490 140.620 138.630 146.080 ;
        RECT 139.410 146.060 139.550 155.180 ;
        RECT 139.870 154.900 140.010 156.960 ;
        RECT 139.810 154.580 140.070 154.900 ;
        RECT 139.810 153.560 140.070 153.880 ;
        RECT 139.350 145.740 139.610 146.060 ;
        RECT 138.890 142.340 139.150 142.660 ;
        RECT 138.430 140.300 138.690 140.620 ;
        RECT 138.950 140.360 139.090 142.340 ;
        RECT 139.870 141.640 140.010 153.560 ;
        RECT 140.330 144.020 140.470 164.440 ;
        RECT 140.790 160.000 140.930 165.120 ;
        RECT 141.250 160.760 141.390 186.290 ;
        RECT 141.650 186.200 141.910 186.290 ;
        RECT 142.630 184.140 142.770 186.880 ;
        RECT 144.410 186.200 144.670 186.520 ;
        RECT 142.570 183.820 142.830 184.140 ;
        RECT 143.950 183.820 144.210 184.140 ;
        RECT 142.110 183.140 142.370 183.460 ;
        RECT 142.170 179.380 142.310 183.140 ;
        RECT 144.010 181.160 144.150 183.820 ;
        RECT 144.470 183.800 144.610 186.200 ;
        RECT 144.870 185.860 145.130 186.180 ;
        RECT 144.410 183.480 144.670 183.800 ;
        RECT 142.630 181.020 144.150 181.160 ;
        RECT 142.630 180.740 142.770 181.020 ;
        RECT 142.570 180.420 142.830 180.740 ;
        RECT 143.950 180.650 144.210 180.740 ;
        RECT 143.550 180.510 144.210 180.650 ;
        RECT 142.110 179.060 142.370 179.380 ;
        RECT 142.630 178.700 142.770 180.420 ;
        RECT 141.650 178.380 141.910 178.700 ;
        RECT 142.570 178.380 142.830 178.700 ;
        RECT 141.710 176.660 141.850 178.380 ;
        RECT 141.650 176.340 141.910 176.660 ;
        RECT 142.630 176.320 142.770 178.380 ;
        RECT 143.550 178.360 143.690 180.510 ;
        RECT 143.950 180.420 144.210 180.510 ;
        RECT 143.490 178.040 143.750 178.360 ;
        RECT 143.550 176.320 143.690 178.040 ;
        RECT 142.570 176.000 142.830 176.320 ;
        RECT 143.490 176.000 143.750 176.320 ;
        RECT 142.110 173.960 142.370 174.280 ;
        RECT 141.650 170.220 141.910 170.540 ;
        RECT 141.710 161.440 141.850 170.220 ;
        RECT 142.170 162.915 142.310 173.960 ;
        RECT 142.630 167.820 142.770 176.000 ;
        RECT 143.030 175.660 143.290 175.980 ;
        RECT 142.570 167.500 142.830 167.820 ;
        RECT 142.100 162.545 142.380 162.915 ;
        RECT 142.630 162.720 142.770 167.500 ;
        RECT 142.570 162.400 142.830 162.720 ;
        RECT 141.710 161.300 142.770 161.440 ;
        RECT 141.250 160.620 142.310 160.760 ;
        RECT 140.730 159.680 140.990 160.000 ;
        RECT 141.650 159.680 141.910 160.000 ;
        RECT 140.790 151.500 140.930 159.680 ;
        RECT 141.190 159.000 141.450 159.320 ;
        RECT 141.250 154.900 141.390 159.000 ;
        RECT 141.710 157.960 141.850 159.680 ;
        RECT 141.650 157.640 141.910 157.960 ;
        RECT 141.190 154.810 141.450 154.900 ;
        RECT 141.190 154.670 141.850 154.810 ;
        RECT 141.190 154.580 141.450 154.670 ;
        RECT 140.730 151.180 140.990 151.500 ;
        RECT 140.730 148.800 140.990 149.120 ;
        RECT 140.790 146.400 140.930 148.800 ;
        RECT 140.730 146.080 140.990 146.400 ;
        RECT 140.270 143.930 140.530 144.020 ;
        RECT 140.270 143.790 140.930 143.930 ;
        RECT 140.270 143.700 140.530 143.790 ;
        RECT 140.270 142.340 140.530 142.660 ;
        RECT 139.810 141.320 140.070 141.640 ;
        RECT 138.950 140.220 140.010 140.360 ;
        RECT 139.350 139.620 139.610 139.940 ;
        RECT 138.890 138.600 139.150 138.920 ;
        RECT 137.970 137.920 138.230 138.240 ;
        RECT 138.950 137.900 139.090 138.600 ;
        RECT 134.350 137.500 134.950 137.640 ;
        RECT 135.670 137.580 135.930 137.900 ;
        RECT 138.890 137.580 139.150 137.900 ;
        RECT 133.830 134.180 134.090 134.500 ;
        RECT 133.360 130.585 133.640 130.955 ;
        RECT 133.370 130.100 133.630 130.420 ;
        RECT 132.450 127.270 132.710 127.360 ;
        RECT 132.050 127.130 132.710 127.270 ;
        RECT 132.450 127.040 132.710 127.130 ;
        RECT 132.910 127.040 133.170 127.360 ;
        RECT 130.670 126.620 131.270 126.760 ;
        RECT 130.150 123.980 130.410 124.300 ;
        RECT 129.690 123.640 129.950 123.960 ;
        RECT 129.750 122.230 129.890 123.640 ;
        RECT 127.850 121.260 128.110 121.580 ;
        RECT 129.680 120.230 129.960 122.230 ;
        RECT 130.670 121.920 130.810 126.620 ;
        RECT 131.590 124.640 131.730 127.040 ;
        RECT 131.990 125.000 132.250 125.320 ;
        RECT 131.530 124.320 131.790 124.640 ;
        RECT 132.050 122.600 132.190 125.000 ;
        RECT 132.510 123.620 132.650 127.040 ;
        RECT 133.430 124.720 133.570 130.100 ;
        RECT 133.890 129.400 134.030 134.180 ;
        RECT 133.830 129.080 134.090 129.400 ;
        RECT 134.350 127.700 134.490 137.500 ;
        RECT 137.510 136.900 137.770 137.220 ;
        RECT 137.970 136.900 138.230 137.220 ;
        RECT 139.410 136.960 139.550 139.620 ;
        RECT 134.770 136.365 136.650 136.735 ;
        RECT 137.570 135.860 137.710 136.900 ;
        RECT 136.590 135.540 136.850 135.860 ;
        RECT 134.750 134.860 135.010 135.180 ;
        RECT 134.810 134.500 134.950 134.860 ;
        RECT 134.750 134.180 135.010 134.500 ;
        RECT 136.650 132.200 136.790 135.540 ;
        RECT 137.040 135.345 137.320 135.715 ;
        RECT 137.510 135.540 137.770 135.860 ;
        RECT 137.050 135.200 137.310 135.345 ;
        RECT 138.030 133.140 138.170 136.900 ;
        RECT 138.490 136.820 139.550 136.960 ;
        RECT 137.970 132.820 138.230 133.140 ;
        RECT 136.650 132.060 137.250 132.200 ;
        RECT 134.770 130.925 136.650 131.295 ;
        RECT 134.740 129.905 135.020 130.275 ;
        RECT 137.110 130.160 137.250 132.060 ;
        RECT 137.500 131.265 137.780 131.635 ;
        RECT 137.970 131.460 138.230 131.780 ;
        RECT 136.190 130.080 137.250 130.160 ;
        RECT 137.570 130.080 137.710 131.265 ;
        RECT 136.130 130.020 137.250 130.080 ;
        RECT 134.750 129.760 135.010 129.905 ;
        RECT 136.130 129.760 136.390 130.020 ;
        RECT 137.510 129.760 137.770 130.080 ;
        RECT 134.810 129.480 134.950 129.760 ;
        RECT 134.810 129.340 135.410 129.480 ;
        RECT 137.050 129.420 137.310 129.740 ;
        RECT 135.270 128.040 135.410 129.340 ;
        RECT 137.110 128.915 137.250 129.420 ;
        RECT 137.040 128.545 137.320 128.915 ;
        RECT 135.210 127.720 135.470 128.040 ;
        RECT 137.500 127.865 137.780 128.235 ;
        RECT 133.830 127.380 134.090 127.700 ;
        RECT 134.290 127.380 134.550 127.700 ;
        RECT 133.890 125.320 134.030 127.380 ;
        RECT 134.750 127.270 135.010 127.360 ;
        RECT 135.270 127.270 135.410 127.720 ;
        RECT 137.570 127.360 137.710 127.865 ;
        RECT 134.750 127.130 135.410 127.270 ;
        RECT 134.750 127.040 135.010 127.130 ;
        RECT 137.510 127.040 137.770 127.360 ;
        RECT 134.770 125.485 136.650 125.855 ;
        RECT 133.830 125.000 134.090 125.320 ;
        RECT 133.430 124.580 134.490 124.720 ;
        RECT 134.350 124.300 134.490 124.580 ;
        RECT 134.750 124.320 135.010 124.640 ;
        RECT 134.290 123.980 134.550 124.300 ;
        RECT 132.450 123.300 132.710 123.620 ;
        RECT 132.510 122.600 132.650 123.300 ;
        RECT 134.810 122.680 134.950 124.320 ;
        RECT 137.570 124.300 137.710 127.040 ;
        RECT 138.030 126.195 138.170 131.460 ;
        RECT 138.490 127.360 138.630 136.820 ;
        RECT 138.880 135.345 139.160 135.715 ;
        RECT 138.950 134.920 139.090 135.345 ;
        RECT 138.950 134.780 139.550 134.920 ;
        RECT 139.410 134.500 139.550 134.780 ;
        RECT 138.890 134.180 139.150 134.500 ;
        RECT 139.350 134.180 139.610 134.500 ;
        RECT 138.950 133.560 139.090 134.180 ;
        RECT 138.950 133.420 139.550 133.560 ;
        RECT 139.410 132.800 139.550 133.420 ;
        RECT 139.350 132.480 139.610 132.800 ;
        RECT 139.350 131.460 139.610 131.780 ;
        RECT 138.890 130.440 139.150 130.760 ;
        RECT 138.430 127.040 138.690 127.360 ;
        RECT 138.430 126.360 138.690 126.680 ;
        RECT 137.960 125.825 138.240 126.195 ;
        RECT 137.970 124.660 138.230 124.980 ;
        RECT 137.510 123.980 137.770 124.300 ;
        RECT 138.030 122.680 138.170 124.660 ;
        RECT 138.490 124.300 138.630 126.360 ;
        RECT 138.950 125.320 139.090 130.440 ;
        RECT 139.410 125.320 139.550 131.460 ;
        RECT 139.870 127.360 140.010 140.220 ;
        RECT 140.330 138.240 140.470 142.340 ;
        RECT 140.790 141.640 140.930 143.790 ;
        RECT 141.190 142.340 141.450 142.660 ;
        RECT 140.730 141.320 140.990 141.640 ;
        RECT 140.730 139.620 140.990 139.940 ;
        RECT 140.790 138.435 140.930 139.620 ;
        RECT 140.270 137.920 140.530 138.240 ;
        RECT 140.720 138.065 141.000 138.435 ;
        RECT 141.250 137.900 141.390 142.340 ;
        RECT 141.710 138.240 141.850 154.670 ;
        RECT 142.170 153.880 142.310 160.620 ;
        RECT 142.630 160.000 142.770 161.300 ;
        RECT 142.570 159.680 142.830 160.000 ;
        RECT 143.090 159.910 143.230 175.660 ;
        RECT 143.950 173.620 144.210 173.940 ;
        RECT 143.490 172.600 143.750 172.920 ;
        RECT 143.550 170.540 143.690 172.600 ;
        RECT 144.010 171.560 144.150 173.620 ;
        RECT 144.410 173.280 144.670 173.600 ;
        RECT 144.470 171.560 144.610 173.280 ;
        RECT 143.950 171.240 144.210 171.560 ;
        RECT 144.410 171.240 144.670 171.560 ;
        RECT 144.410 170.560 144.670 170.880 ;
        RECT 143.490 170.220 143.750 170.540 ;
        RECT 143.950 164.100 144.210 164.420 ;
        RECT 144.010 160.680 144.150 164.100 ;
        RECT 143.950 160.360 144.210 160.680 ;
        RECT 143.090 159.770 143.690 159.910 ;
        RECT 142.570 158.660 142.830 158.980 ;
        RECT 143.030 158.660 143.290 158.980 ;
        RECT 142.630 157.280 142.770 158.660 ;
        RECT 143.090 157.280 143.230 158.660 ;
        RECT 142.570 156.960 142.830 157.280 ;
        RECT 143.030 156.960 143.290 157.280 ;
        RECT 142.570 155.940 142.830 156.260 ;
        RECT 143.030 155.940 143.290 156.260 ;
        RECT 142.630 155.435 142.770 155.940 ;
        RECT 142.560 155.065 142.840 155.435 ;
        RECT 142.570 153.900 142.830 154.220 ;
        RECT 142.110 153.560 142.370 153.880 ;
        RECT 142.100 151.920 142.380 152.035 ;
        RECT 142.630 151.920 142.770 153.900 ;
        RECT 142.100 151.780 142.770 151.920 ;
        RECT 142.100 151.665 142.380 151.780 ;
        RECT 142.110 151.520 142.370 151.665 ;
        RECT 142.110 150.500 142.370 150.820 ;
        RECT 142.170 140.960 142.310 150.500 ;
        RECT 142.110 140.640 142.370 140.960 ;
        RECT 142.110 139.620 142.370 139.940 ;
        RECT 141.650 137.920 141.910 138.240 ;
        RECT 141.190 137.580 141.450 137.900 ;
        RECT 140.730 137.240 140.990 137.560 ;
        RECT 140.790 136.200 140.930 137.240 ;
        RECT 141.190 136.900 141.450 137.220 ;
        RECT 140.730 135.880 140.990 136.200 ;
        RECT 140.720 133.305 141.000 133.675 ;
        RECT 140.790 132.800 140.930 133.305 ;
        RECT 140.730 132.480 140.990 132.800 ;
        RECT 140.730 131.460 140.990 131.780 ;
        RECT 140.790 129.740 140.930 131.460 ;
        RECT 140.730 129.420 140.990 129.740 ;
        RECT 139.810 127.040 140.070 127.360 ;
        RECT 141.250 125.320 141.390 136.900 ;
        RECT 141.710 135.180 141.850 137.920 ;
        RECT 141.650 134.860 141.910 135.180 ;
        RECT 141.650 133.160 141.910 133.480 ;
        RECT 141.710 131.780 141.850 133.160 ;
        RECT 141.650 131.460 141.910 131.780 ;
        RECT 142.170 130.760 142.310 139.620 ;
        RECT 143.090 138.920 143.230 155.940 ;
        RECT 143.550 143.680 143.690 159.770 ;
        RECT 143.950 159.680 144.210 160.000 ;
        RECT 144.010 155.240 144.150 159.680 ;
        RECT 143.950 154.920 144.210 155.240 ;
        RECT 143.950 150.840 144.210 151.160 ;
        RECT 144.010 149.460 144.150 150.840 ;
        RECT 143.950 149.140 144.210 149.460 ;
        RECT 143.950 147.780 144.210 148.100 ;
        RECT 143.490 143.360 143.750 143.680 ;
        RECT 143.550 141.640 143.690 143.360 ;
        RECT 143.490 141.320 143.750 141.640 ;
        RECT 144.010 140.960 144.150 147.780 ;
        RECT 143.950 140.640 144.210 140.960 ;
        RECT 143.940 140.360 144.220 140.475 ;
        RECT 144.470 140.360 144.610 170.560 ;
        RECT 144.930 156.940 145.070 185.860 ;
        RECT 145.330 183.480 145.590 183.800 ;
        RECT 145.390 182.440 145.530 183.480 ;
        RECT 145.330 182.120 145.590 182.440 ;
        RECT 145.850 181.840 145.990 186.880 ;
        RECT 145.390 181.700 145.990 181.840 ;
        RECT 145.390 173.000 145.530 181.700 ;
        RECT 145.790 179.400 146.050 179.720 ;
        RECT 145.850 173.600 145.990 179.400 ;
        RECT 145.790 173.280 146.050 173.600 ;
        RECT 145.390 172.860 145.990 173.000 ;
        RECT 145.330 169.540 145.590 169.860 ;
        RECT 144.870 156.620 145.130 156.940 ;
        RECT 144.870 154.920 145.130 155.240 ;
        RECT 143.940 140.220 144.610 140.360 ;
        RECT 143.940 140.105 144.220 140.220 ;
        RECT 143.030 138.600 143.290 138.920 ;
        RECT 144.930 137.900 145.070 154.920 ;
        RECT 143.030 137.580 143.290 137.900 ;
        RECT 144.870 137.580 145.130 137.900 ;
        RECT 143.090 135.860 143.230 137.580 ;
        RECT 145.390 137.130 145.530 169.540 ;
        RECT 145.850 157.620 145.990 172.860 ;
        RECT 145.790 157.300 146.050 157.620 ;
        RECT 146.310 156.940 146.450 194.620 ;
        RECT 147.690 194.080 147.830 196.740 ;
        RECT 147.230 193.940 147.830 194.080 ;
        RECT 146.700 191.785 146.980 192.155 ;
        RECT 146.710 191.640 146.970 191.785 ;
        RECT 146.710 189.260 146.970 189.580 ;
        RECT 146.770 187.880 146.910 189.260 ;
        RECT 146.710 187.560 146.970 187.880 ;
        RECT 146.710 185.860 146.970 186.180 ;
        RECT 146.770 170.880 146.910 185.860 ;
        RECT 147.230 175.720 147.370 193.940 ;
        RECT 149.770 193.485 151.650 193.855 ;
        RECT 147.630 192.320 147.890 192.640 ;
        RECT 147.690 190.260 147.830 192.320 ;
        RECT 148.090 191.640 148.350 191.960 ;
        RECT 147.630 189.940 147.890 190.260 ;
        RECT 148.150 187.200 148.290 191.640 ;
        RECT 152.290 190.000 152.430 196.740 ;
        RECT 152.750 192.835 152.890 209.455 ;
        RECT 153.150 199.460 153.410 199.780 ;
        RECT 153.210 198.760 153.350 199.460 ;
        RECT 153.150 198.440 153.410 198.760 ;
        RECT 153.150 194.020 153.410 194.340 ;
        RECT 152.680 192.465 152.960 192.835 ;
        RECT 149.010 189.830 149.270 189.920 ;
        RECT 148.610 189.690 149.270 189.830 ;
        RECT 148.610 188.755 148.750 189.690 ;
        RECT 149.010 189.600 149.270 189.690 ;
        RECT 149.930 189.600 150.190 189.920 ;
        RECT 152.290 189.860 152.890 190.000 ;
        RECT 149.990 189.320 150.130 189.600 ;
        RECT 149.070 189.180 150.130 189.320 ;
        RECT 151.770 189.260 152.030 189.580 ;
        RECT 152.230 189.260 152.490 189.580 ;
        RECT 148.540 188.385 148.820 188.755 ;
        RECT 147.630 186.880 147.890 187.200 ;
        RECT 148.090 186.880 148.350 187.200 ;
        RECT 147.690 183.460 147.830 186.880 ;
        RECT 147.630 183.140 147.890 183.460 ;
        RECT 149.070 182.400 149.210 189.180 ;
        RECT 149.770 188.045 151.650 188.415 ;
        RECT 151.830 187.200 151.970 189.260 ;
        RECT 149.930 186.880 150.190 187.200 ;
        RECT 151.770 186.880 152.030 187.200 ;
        RECT 149.990 183.800 150.130 186.880 ;
        RECT 152.290 185.160 152.430 189.260 ;
        RECT 152.230 184.840 152.490 185.160 ;
        RECT 149.930 183.480 150.190 183.800 ;
        RECT 149.770 182.605 151.650 182.975 ;
        RECT 152.750 182.440 152.890 189.860 ;
        RECT 153.210 189.240 153.350 194.020 ;
        RECT 153.610 189.940 153.870 190.260 ;
        RECT 153.150 188.920 153.410 189.240 ;
        RECT 148.150 182.260 149.210 182.400 ;
        RECT 147.230 175.580 147.830 175.720 ;
        RECT 147.170 174.980 147.430 175.300 ;
        RECT 147.230 173.940 147.370 174.980 ;
        RECT 147.170 173.620 147.430 173.940 ;
        RECT 147.170 172.940 147.430 173.260 ;
        RECT 146.710 170.560 146.970 170.880 ;
        RECT 146.700 165.265 146.980 165.635 ;
        RECT 146.710 165.120 146.970 165.265 ;
        RECT 146.700 162.545 146.980 162.915 ;
        RECT 146.770 160.340 146.910 162.545 ;
        RECT 146.710 160.020 146.970 160.340 ;
        RECT 146.710 157.300 146.970 157.620 ;
        RECT 145.790 156.620 146.050 156.940 ;
        RECT 146.250 156.620 146.510 156.940 ;
        RECT 145.850 152.520 145.990 156.620 ;
        RECT 145.790 152.200 146.050 152.520 ;
        RECT 145.850 151.500 145.990 152.200 ;
        RECT 145.790 151.180 146.050 151.500 ;
        RECT 145.790 150.500 146.050 150.820 ;
        RECT 145.850 149.800 145.990 150.500 ;
        RECT 145.790 149.480 146.050 149.800 ;
        RECT 146.770 149.710 146.910 157.300 ;
        RECT 147.230 152.520 147.370 172.940 ;
        RECT 147.690 154.560 147.830 175.580 ;
        RECT 148.150 170.540 148.290 182.260 ;
        RECT 152.690 182.120 152.950 182.440 ;
        RECT 153.210 181.420 153.350 188.920 ;
        RECT 153.670 187.880 153.810 189.940 ;
        RECT 154.990 188.580 155.250 188.900 ;
        RECT 153.610 187.560 153.870 187.880 ;
        RECT 153.610 185.860 153.870 186.180 ;
        RECT 153.670 184.140 153.810 185.860 ;
        RECT 154.070 184.840 154.330 185.160 ;
        RECT 154.130 184.560 154.270 184.840 ;
        RECT 154.130 184.420 154.730 184.560 ;
        RECT 153.610 183.820 153.870 184.140 ;
        RECT 154.070 182.120 154.330 182.440 ;
        RECT 153.150 181.100 153.410 181.420 ;
        RECT 149.010 180.420 149.270 180.740 ;
        RECT 152.690 180.420 152.950 180.740 ;
        RECT 148.550 178.040 148.810 178.360 ;
        RECT 148.610 177.000 148.750 178.040 ;
        RECT 149.070 177.000 149.210 180.420 ;
        RECT 149.770 177.165 151.650 177.535 ;
        RECT 152.750 177.000 152.890 180.420 ;
        RECT 148.550 176.680 148.810 177.000 ;
        RECT 149.010 176.680 149.270 177.000 ;
        RECT 152.690 176.680 152.950 177.000 ;
        RECT 149.070 173.600 149.210 176.680 ;
        RECT 149.470 176.000 149.730 176.320 ;
        RECT 150.850 176.000 151.110 176.320 ;
        RECT 149.530 174.280 149.670 176.000 ;
        RECT 150.910 175.835 151.050 176.000 ;
        RECT 150.840 175.720 151.120 175.835 ;
        RECT 150.840 175.580 151.970 175.720 ;
        RECT 150.840 175.465 151.120 175.580 ;
        RECT 149.470 173.960 149.730 174.280 ;
        RECT 149.010 173.280 149.270 173.600 ;
        RECT 149.010 172.260 149.270 172.580 ;
        RECT 148.090 170.220 148.350 170.540 ;
        RECT 149.070 168.355 149.210 172.260 ;
        RECT 149.770 171.725 151.650 172.095 ;
        RECT 151.830 170.880 151.970 175.580 ;
        RECT 152.690 172.260 152.950 172.580 ;
        RECT 151.770 170.560 152.030 170.880 ;
        RECT 149.000 167.985 149.280 168.355 ;
        RECT 149.070 167.820 149.210 167.985 ;
        RECT 149.010 167.500 149.270 167.820 ;
        RECT 149.770 166.285 151.650 166.655 ;
        RECT 151.830 166.120 151.970 170.560 ;
        RECT 152.230 166.820 152.490 167.140 ;
        RECT 151.770 165.800 152.030 166.120 ;
        RECT 152.290 165.440 152.430 166.820 ;
        RECT 152.230 165.120 152.490 165.440 ;
        RECT 148.090 164.780 148.350 165.100 ;
        RECT 147.630 154.240 147.890 154.560 ;
        RECT 147.170 152.200 147.430 152.520 ;
        RECT 148.150 149.800 148.290 164.780 ;
        RECT 152.290 163.400 152.430 165.120 ;
        RECT 152.230 163.080 152.490 163.400 ;
        RECT 151.770 161.720 152.030 162.040 ;
        RECT 149.770 160.845 151.650 161.215 ;
        RECT 151.830 160.680 151.970 161.720 ;
        RECT 151.770 160.360 152.030 160.680 ;
        RECT 149.010 156.620 149.270 156.940 ;
        RECT 149.070 154.900 149.210 156.620 ;
        RECT 149.770 155.405 151.650 155.775 ;
        RECT 149.010 154.580 149.270 154.900 ;
        RECT 150.390 154.580 150.650 154.900 ;
        RECT 148.550 154.240 148.810 154.560 ;
        RECT 148.610 151.500 148.750 154.240 ;
        RECT 149.010 152.200 149.270 152.520 ;
        RECT 148.550 151.180 148.810 151.500 ;
        RECT 148.550 150.500 148.810 150.820 ;
        RECT 148.610 149.800 148.750 150.500 ;
        RECT 149.070 149.800 149.210 152.200 ;
        RECT 150.450 151.410 150.590 154.580 ;
        RECT 150.850 151.410 151.110 151.500 ;
        RECT 150.450 151.270 151.110 151.410 ;
        RECT 150.850 151.180 151.110 151.270 ;
        RECT 152.230 150.500 152.490 150.820 ;
        RECT 149.770 149.965 151.650 150.335 ;
        RECT 146.310 149.570 146.910 149.710 ;
        RECT 146.310 144.020 146.450 149.570 ;
        RECT 148.090 149.480 148.350 149.800 ;
        RECT 148.550 149.480 148.810 149.800 ;
        RECT 149.010 149.480 149.270 149.800 ;
        RECT 148.150 149.200 148.290 149.480 ;
        RECT 152.290 149.315 152.430 150.500 ;
        RECT 146.710 148.800 146.970 149.120 ;
        RECT 148.150 149.060 149.210 149.200 ;
        RECT 149.070 149.030 149.210 149.060 ;
        RECT 149.930 149.030 150.190 149.120 ;
        RECT 149.070 148.890 150.190 149.030 ;
        RECT 152.220 148.945 152.500 149.315 ;
        RECT 149.930 148.800 150.190 148.890 ;
        RECT 146.770 146.740 146.910 148.800 ;
        RECT 152.750 148.520 152.890 172.260 ;
        RECT 153.150 170.560 153.410 170.880 ;
        RECT 153.210 168.500 153.350 170.560 ;
        RECT 153.610 169.540 153.870 169.860 ;
        RECT 153.150 168.180 153.410 168.500 ;
        RECT 153.210 166.120 153.350 168.180 ;
        RECT 153.150 165.800 153.410 166.120 ;
        RECT 153.670 165.100 153.810 169.540 ;
        RECT 153.610 164.780 153.870 165.100 ;
        RECT 153.610 164.100 153.870 164.420 ;
        RECT 153.670 149.120 153.810 164.100 ;
        RECT 154.130 156.940 154.270 182.120 ;
        RECT 154.070 156.620 154.330 156.940 ;
        RECT 154.130 151.500 154.270 156.620 ;
        RECT 154.070 151.180 154.330 151.500 ;
        RECT 153.610 148.800 153.870 149.120 ;
        RECT 151.770 148.120 152.030 148.440 ;
        RECT 152.290 148.380 152.890 148.520 ;
        RECT 146.710 146.420 146.970 146.740 ;
        RECT 149.770 144.525 151.650 144.895 ;
        RECT 146.250 143.700 146.510 144.020 ;
        RECT 146.310 141.640 146.450 143.700 ;
        RECT 151.830 143.680 151.970 148.120 ;
        RECT 151.770 143.360 152.030 143.680 ;
        RECT 149.010 142.340 149.270 142.660 ;
        RECT 146.250 141.320 146.510 141.640 ;
        RECT 148.550 140.300 148.810 140.620 ;
        RECT 145.780 139.425 146.060 139.795 ;
        RECT 144.930 136.990 145.530 137.130 ;
        RECT 143.030 135.540 143.290 135.860 ;
        RECT 142.570 134.180 142.830 134.500 ;
        RECT 142.630 132.800 142.770 134.180 ;
        RECT 143.090 133.140 143.230 135.540 ;
        RECT 144.410 135.035 144.670 135.180 ;
        RECT 144.400 134.665 144.680 135.035 ;
        RECT 143.490 134.180 143.750 134.500 ;
        RECT 143.030 132.820 143.290 133.140 ;
        RECT 142.570 132.480 142.830 132.800 ;
        RECT 142.110 130.440 142.370 130.760 ;
        RECT 143.550 130.080 143.690 134.180 ;
        RECT 143.950 132.820 144.210 133.140 ;
        RECT 143.490 129.760 143.750 130.080 ;
        RECT 142.570 129.595 142.830 129.740 ;
        RECT 142.560 129.225 142.840 129.595 ;
        RECT 143.030 129.420 143.290 129.740 ;
        RECT 141.650 127.040 141.910 127.360 ;
        RECT 138.890 125.000 139.150 125.320 ;
        RECT 139.350 125.000 139.610 125.320 ;
        RECT 141.190 125.000 141.450 125.320 ;
        RECT 138.430 123.980 138.690 124.300 ;
        RECT 139.810 123.980 140.070 124.300 ;
        RECT 131.990 122.280 132.250 122.600 ;
        RECT 132.450 122.280 132.710 122.600 ;
        RECT 133.430 122.540 134.950 122.680 ;
        RECT 137.110 122.540 138.170 122.680 ;
        RECT 133.430 122.230 133.570 122.540 ;
        RECT 137.110 122.230 137.250 122.540 ;
        RECT 130.610 121.600 130.870 121.920 ;
        RECT 133.360 120.230 133.640 122.230 ;
        RECT 137.040 120.230 137.320 122.230 ;
        RECT 138.490 121.580 138.630 123.980 ;
        RECT 139.870 122.600 140.010 123.980 ;
        RECT 139.810 122.280 140.070 122.600 ;
        RECT 140.790 122.540 141.390 122.680 ;
        RECT 141.710 122.600 141.850 127.040 ;
        RECT 142.570 126.020 142.830 126.340 ;
        RECT 142.630 125.400 142.770 126.020 ;
        RECT 142.170 125.260 142.770 125.400 ;
        RECT 143.090 125.320 143.230 129.420 ;
        RECT 143.550 127.360 143.690 129.760 ;
        RECT 143.490 127.040 143.750 127.360 ;
        RECT 143.480 126.505 143.760 126.875 ;
        RECT 144.010 126.680 144.150 132.820 ;
        RECT 144.930 132.800 145.070 136.990 ;
        RECT 145.850 134.500 145.990 139.425 ;
        RECT 148.610 136.200 148.750 140.300 ;
        RECT 149.070 137.900 149.210 142.340 ;
        RECT 151.830 141.300 151.970 143.360 ;
        RECT 152.290 143.340 152.430 148.380 ;
        RECT 152.690 147.780 152.950 148.100 ;
        RECT 152.230 143.020 152.490 143.340 ;
        RECT 151.770 140.980 152.030 141.300 ;
        RECT 151.830 140.620 151.970 140.980 ;
        RECT 152.750 140.620 152.890 147.780 ;
        RECT 153.150 143.020 153.410 143.340 ;
        RECT 151.770 140.300 152.030 140.620 ;
        RECT 152.690 140.300 152.950 140.620 ;
        RECT 149.770 139.085 151.650 139.455 ;
        RECT 149.010 137.580 149.270 137.900 ;
        RECT 149.070 136.200 149.210 137.580 ;
        RECT 151.830 137.220 151.970 140.300 ;
        RECT 152.230 139.960 152.490 140.280 ;
        RECT 152.290 138.240 152.430 139.960 ;
        RECT 152.230 137.920 152.490 138.240 ;
        RECT 151.770 136.900 152.030 137.220 ;
        RECT 148.550 135.880 148.810 136.200 ;
        RECT 149.010 135.880 149.270 136.200 ;
        RECT 152.290 135.520 152.430 137.920 ;
        RECT 153.210 137.900 153.350 143.020 ;
        RECT 154.590 140.620 154.730 184.420 ;
        RECT 155.050 181.420 155.190 188.580 ;
        RECT 154.990 181.100 155.250 181.420 ;
        RECT 155.450 175.320 155.710 175.640 ;
        RECT 154.990 167.840 155.250 168.160 ;
        RECT 155.050 164.420 155.190 167.840 ;
        RECT 154.990 164.100 155.250 164.420 ;
        RECT 154.530 140.300 154.790 140.620 ;
        RECT 153.150 137.580 153.410 137.900 ;
        RECT 152.230 135.200 152.490 135.520 ;
        RECT 153.670 135.460 155.190 135.600 ;
        RECT 153.670 135.180 153.810 135.460 ;
        RECT 148.550 134.860 148.810 135.180 ;
        RECT 153.610 134.860 153.870 135.180 ;
        RECT 145.790 134.180 146.050 134.500 ;
        RECT 145.850 132.800 145.990 134.180 ;
        RECT 144.870 132.480 145.130 132.800 ;
        RECT 145.790 132.480 146.050 132.800 ;
        RECT 144.410 131.460 144.670 131.780 ;
        RECT 144.470 130.955 144.610 131.460 ;
        RECT 144.400 130.585 144.680 130.955 ;
        RECT 144.930 129.740 145.070 132.480 ;
        RECT 145.790 131.800 146.050 132.120 ;
        RECT 145.330 131.460 145.590 131.780 ;
        RECT 145.390 130.760 145.530 131.460 ;
        RECT 145.330 130.440 145.590 130.760 ;
        RECT 144.870 129.420 145.130 129.740 ;
        RECT 144.410 127.720 144.670 128.040 ;
        RECT 140.790 122.230 140.930 122.540 ;
        RECT 138.430 121.260 138.690 121.580 ;
        RECT 140.720 120.230 141.000 122.230 ;
        RECT 141.250 122.000 141.390 122.540 ;
        RECT 141.650 122.280 141.910 122.600 ;
        RECT 142.170 122.000 142.310 125.260 ;
        RECT 143.030 125.000 143.290 125.320 ;
        RECT 143.550 124.300 143.690 126.505 ;
        RECT 143.950 126.360 144.210 126.680 ;
        RECT 143.940 125.825 144.220 126.195 ;
        RECT 144.010 124.300 144.150 125.825 ;
        RECT 143.490 123.980 143.750 124.300 ;
        RECT 143.950 123.980 144.210 124.300 ;
        RECT 144.470 122.230 144.610 127.720 ;
        RECT 144.930 126.680 145.070 129.420 ;
        RECT 145.320 129.225 145.600 129.595 ;
        RECT 145.390 128.040 145.530 129.225 ;
        RECT 145.850 129.060 145.990 131.800 ;
        RECT 147.170 131.460 147.430 131.780 ;
        RECT 148.090 131.635 148.350 131.780 ;
        RECT 146.240 130.585 146.520 130.955 ;
        RECT 146.310 130.080 146.450 130.585 ;
        RECT 146.250 129.760 146.510 130.080 ;
        RECT 145.790 128.740 146.050 129.060 ;
        RECT 146.250 128.740 146.510 129.060 ;
        RECT 145.330 127.720 145.590 128.040 ;
        RECT 146.310 127.555 146.450 128.740 ;
        RECT 146.700 128.545 146.980 128.915 ;
        RECT 146.240 127.185 146.520 127.555 ;
        RECT 146.770 127.360 146.910 128.545 ;
        RECT 146.710 127.040 146.970 127.360 ;
        RECT 144.870 126.360 145.130 126.680 ;
        RECT 147.230 126.080 147.370 131.460 ;
        RECT 148.080 131.265 148.360 131.635 ;
        RECT 147.630 129.080 147.890 129.400 ;
        RECT 148.090 129.080 148.350 129.400 ;
        RECT 147.690 127.360 147.830 129.080 ;
        RECT 148.150 128.040 148.290 129.080 ;
        RECT 148.090 127.720 148.350 128.040 ;
        RECT 147.630 127.040 147.890 127.360 ;
        RECT 147.230 125.940 148.290 126.080 ;
        RECT 148.150 122.230 148.290 125.940 ;
        RECT 148.610 123.620 148.750 134.860 ;
        RECT 152.690 134.750 152.950 134.840 ;
        RECT 152.690 134.610 153.350 134.750 ;
        RECT 152.690 134.520 152.950 134.610 ;
        RECT 151.770 134.180 152.030 134.500 ;
        RECT 149.770 133.645 151.650 134.015 ;
        RECT 149.010 133.160 149.270 133.480 ;
        RECT 149.070 129.595 149.210 133.160 ;
        RECT 149.930 131.460 150.190 131.780 ;
        RECT 150.390 131.460 150.650 131.780 ;
        RECT 149.990 130.160 150.130 131.460 ;
        RECT 150.450 130.760 150.590 131.460 ;
        RECT 150.390 130.440 150.650 130.760 ;
        RECT 150.850 130.160 151.110 130.420 ;
        RECT 149.990 130.100 151.110 130.160 ;
        RECT 149.990 130.020 151.050 130.100 ;
        RECT 149.000 129.480 149.280 129.595 ;
        RECT 149.000 129.340 150.590 129.480 ;
        RECT 149.000 129.225 149.280 129.340 ;
        RECT 150.450 129.060 150.590 129.340 ;
        RECT 150.390 128.740 150.650 129.060 ;
        RECT 149.770 128.205 151.650 128.575 ;
        RECT 149.010 123.640 149.270 123.960 ;
        RECT 148.550 123.300 148.810 123.620 ;
        RECT 149.070 122.600 149.210 123.640 ;
        RECT 149.770 122.765 151.650 123.135 ;
        RECT 149.010 122.280 149.270 122.600 ;
        RECT 151.830 122.230 151.970 134.180 ;
        RECT 152.230 131.460 152.490 131.780 ;
        RECT 152.290 124.300 152.430 131.460 ;
        RECT 153.210 129.740 153.350 134.610 ;
        RECT 154.070 134.520 154.330 134.840 ;
        RECT 153.610 133.160 153.870 133.480 ;
        RECT 153.150 129.420 153.410 129.740 ;
        RECT 153.150 127.040 153.410 127.360 ;
        RECT 153.210 125.320 153.350 127.040 ;
        RECT 153.150 125.000 153.410 125.320 ;
        RECT 153.670 124.640 153.810 133.160 ;
        RECT 154.130 127.700 154.270 134.520 ;
        RECT 154.530 134.180 154.790 134.500 ;
        RECT 154.590 129.740 154.730 134.180 ;
        RECT 154.530 129.420 154.790 129.740 ;
        RECT 155.050 127.700 155.190 135.460 ;
        RECT 155.510 133.140 155.650 175.320 ;
        RECT 155.910 171.240 156.170 171.560 ;
        RECT 155.970 133.140 156.110 171.240 ;
        RECT 155.450 132.820 155.710 133.140 ;
        RECT 155.910 132.820 156.170 133.140 ;
        RECT 155.450 131.800 155.710 132.120 ;
        RECT 154.070 127.380 154.330 127.700 ;
        RECT 154.990 127.380 155.250 127.700 ;
        RECT 153.610 124.320 153.870 124.640 ;
        RECT 152.230 123.980 152.490 124.300 ;
        RECT 155.510 122.230 155.650 131.800 ;
        RECT 141.250 121.860 142.310 122.000 ;
        RECT 144.400 120.230 144.680 122.230 ;
        RECT 148.080 120.230 148.360 122.230 ;
        RECT 151.760 120.230 152.040 122.230 ;
        RECT 155.440 120.230 155.720 122.230 ;
        RECT 77.570 79.080 78.630 80.080 ;
        RECT 114.570 79.080 115.630 80.080 ;
        RECT 151.570 79.080 152.630 80.080 ;
        RECT 77.600 30.000 78.600 79.080 ;
        RECT 114.600 30.000 115.600 79.080 ;
        RECT 151.600 30.000 152.600 79.080 ;
        RECT 35.990 24.045 36.350 24.345 ;
        RECT 36.020 21.995 36.320 24.045 ;
        RECT 35.990 21.695 36.350 21.995 ;
        RECT 36.020 19.745 36.320 21.695 ;
        RECT 35.990 19.445 36.350 19.745 ;
        RECT 35.370 18.345 35.670 18.375 ;
        RECT 34.290 18.045 35.670 18.345 ;
        RECT 35.370 18.015 35.670 18.045 ;
      LAYER via2 ;
        RECT 122.015 216.515 122.385 216.885 ;
        RECT 113.825 214.925 114.175 215.275 ;
        RECT 118.315 215.015 118.690 215.390 ;
        RECT 110.265 214.165 110.735 214.635 ;
        RECT 126.520 214.220 126.880 214.580 ;
        RECT 127.830 214.230 128.175 214.575 ;
        RECT 131.935 214.235 132.270 214.570 ;
        RECT 135.990 214.190 136.415 214.615 ;
        RECT 140.230 214.230 140.575 214.575 ;
        RECT 144.295 214.195 144.705 214.605 ;
        RECT 148.510 214.210 148.890 214.590 ;
        RECT 152.595 214.195 153.005 214.605 ;
        RECT 74.770 207.130 75.050 207.410 ;
        RECT 75.170 207.130 75.450 207.410 ;
        RECT 75.570 207.130 75.850 207.410 ;
        RECT 75.970 207.130 76.250 207.410 ;
        RECT 76.370 207.130 76.650 207.410 ;
        RECT 89.770 204.410 90.050 204.690 ;
        RECT 90.170 204.410 90.450 204.690 ;
        RECT 90.570 204.410 90.850 204.690 ;
        RECT 90.970 204.410 91.250 204.690 ;
        RECT 91.370 204.410 91.650 204.690 ;
        RECT 92.420 203.390 92.700 203.670 ;
        RECT 74.770 201.690 75.050 201.970 ;
        RECT 75.170 201.690 75.450 201.970 ;
        RECT 75.570 201.690 75.850 201.970 ;
        RECT 75.970 201.690 76.250 201.970 ;
        RECT 76.370 201.690 76.650 201.970 ;
        RECT 78.160 198.630 78.440 198.910 ;
        RECT 74.770 196.250 75.050 196.530 ;
        RECT 75.170 196.250 75.450 196.530 ;
        RECT 75.570 196.250 75.850 196.530 ;
        RECT 75.970 196.250 76.250 196.530 ;
        RECT 76.370 196.250 76.650 196.530 ;
        RECT 81.380 194.550 81.660 194.830 ;
        RECT 74.770 190.810 75.050 191.090 ;
        RECT 75.170 190.810 75.450 191.090 ;
        RECT 75.570 190.810 75.850 191.090 ;
        RECT 75.970 190.810 76.250 191.090 ;
        RECT 76.370 190.810 76.650 191.090 ;
        RECT 74.770 185.370 75.050 185.650 ;
        RECT 75.170 185.370 75.450 185.650 ;
        RECT 75.570 185.370 75.850 185.650 ;
        RECT 75.970 185.370 76.250 185.650 ;
        RECT 76.370 185.370 76.650 185.650 ;
        RECT 74.770 179.930 75.050 180.210 ;
        RECT 75.170 179.930 75.450 180.210 ;
        RECT 75.570 179.930 75.850 180.210 ;
        RECT 75.970 179.930 76.250 180.210 ;
        RECT 76.370 179.930 76.650 180.210 ;
        RECT 81.380 191.830 81.660 192.110 ;
        RECT 74.770 174.490 75.050 174.770 ;
        RECT 75.170 174.490 75.450 174.770 ;
        RECT 75.570 174.490 75.850 174.770 ;
        RECT 75.970 174.490 76.250 174.770 ;
        RECT 76.370 174.490 76.650 174.770 ;
        RECT 74.770 169.050 75.050 169.330 ;
        RECT 75.170 169.050 75.450 169.330 ;
        RECT 75.570 169.050 75.850 169.330 ;
        RECT 75.970 169.050 76.250 169.330 ;
        RECT 76.370 169.050 76.650 169.330 ;
        RECT 77.240 164.630 77.520 164.910 ;
        RECT 74.770 163.610 75.050 163.890 ;
        RECT 75.170 163.610 75.450 163.890 ;
        RECT 75.570 163.610 75.850 163.890 ;
        RECT 75.970 163.610 76.250 163.890 ;
        RECT 76.370 163.610 76.650 163.890 ;
        RECT 74.770 158.170 75.050 158.450 ;
        RECT 75.170 158.170 75.450 158.450 ;
        RECT 75.570 158.170 75.850 158.450 ;
        RECT 75.970 158.170 76.250 158.450 ;
        RECT 76.370 158.170 76.650 158.450 ;
        RECT 74.770 152.730 75.050 153.010 ;
        RECT 75.170 152.730 75.450 153.010 ;
        RECT 75.570 152.730 75.850 153.010 ;
        RECT 75.970 152.730 76.250 153.010 ;
        RECT 76.370 152.730 76.650 153.010 ;
        RECT 74.770 147.290 75.050 147.570 ;
        RECT 75.170 147.290 75.450 147.570 ;
        RECT 75.570 147.290 75.850 147.570 ;
        RECT 75.970 147.290 76.250 147.570 ;
        RECT 76.370 147.290 76.650 147.570 ;
        RECT 74.770 141.850 75.050 142.130 ;
        RECT 75.170 141.850 75.450 142.130 ;
        RECT 75.570 141.850 75.850 142.130 ;
        RECT 75.970 141.850 76.250 142.130 ;
        RECT 76.370 141.850 76.650 142.130 ;
        RECT 74.770 136.410 75.050 136.690 ;
        RECT 75.170 136.410 75.450 136.690 ;
        RECT 75.570 136.410 75.850 136.690 ;
        RECT 75.970 136.410 76.250 136.690 ;
        RECT 76.370 136.410 76.650 136.690 ;
        RECT 74.480 132.670 74.760 132.950 ;
        RECT 74.770 130.970 75.050 131.250 ;
        RECT 75.170 130.970 75.450 131.250 ;
        RECT 75.570 130.970 75.850 131.250 ;
        RECT 75.970 130.970 76.250 131.250 ;
        RECT 76.370 130.970 76.650 131.250 ;
        RECT 81.380 183.670 81.660 183.950 ;
        RECT 84.140 198.630 84.420 198.910 ;
        RECT 82.300 184.350 82.580 184.630 ;
        RECT 78.620 159.190 78.900 159.470 ;
        RECT 80.920 165.310 81.200 165.590 ;
        RECT 85.520 189.790 85.800 190.070 ;
        RECT 89.770 198.970 90.050 199.250 ;
        RECT 90.170 198.970 90.450 199.250 ;
        RECT 90.570 198.970 90.850 199.250 ;
        RECT 90.970 198.970 91.250 199.250 ;
        RECT 91.370 198.970 91.650 199.250 ;
        RECT 88.280 192.510 88.560 192.790 ;
        RECT 89.770 193.530 90.050 193.810 ;
        RECT 90.170 193.530 90.450 193.810 ;
        RECT 90.570 193.530 90.850 193.810 ;
        RECT 90.970 193.530 91.250 193.810 ;
        RECT 91.370 193.530 91.650 193.810 ;
        RECT 90.580 192.510 90.860 192.790 ;
        RECT 91.040 190.470 91.320 190.750 ;
        RECT 89.660 189.790 89.940 190.070 ;
        RECT 92.420 194.550 92.700 194.830 ;
        RECT 93.340 195.230 93.620 195.510 ;
        RECT 88.280 187.070 88.560 187.350 ;
        RECT 89.770 188.090 90.050 188.370 ;
        RECT 90.170 188.090 90.450 188.370 ;
        RECT 90.570 188.090 90.850 188.370 ;
        RECT 90.970 188.090 91.250 188.370 ;
        RECT 91.370 188.090 91.650 188.370 ;
        RECT 82.300 156.470 82.580 156.750 ;
        RECT 80.920 144.910 81.200 145.190 ;
        RECT 94.260 189.110 94.540 189.390 ;
        RECT 89.770 182.650 90.050 182.930 ;
        RECT 90.170 182.650 90.450 182.930 ;
        RECT 90.570 182.650 90.850 182.930 ;
        RECT 90.970 182.650 91.250 182.930 ;
        RECT 91.370 182.650 91.650 182.930 ;
        RECT 87.360 174.830 87.640 175.110 ;
        RECT 88.280 174.150 88.560 174.430 ;
        RECT 89.770 177.210 90.050 177.490 ;
        RECT 90.170 177.210 90.450 177.490 ;
        RECT 90.570 177.210 90.850 177.490 ;
        RECT 90.970 177.210 91.250 177.490 ;
        RECT 91.370 177.210 91.650 177.490 ;
        RECT 91.040 172.790 91.320 173.070 ;
        RECT 86.900 170.070 87.180 170.350 ;
        RECT 89.770 171.770 90.050 172.050 ;
        RECT 90.170 171.770 90.450 172.050 ;
        RECT 90.570 171.770 90.850 172.050 ;
        RECT 90.970 171.770 91.250 172.050 ;
        RECT 91.370 171.770 91.650 172.050 ;
        RECT 89.660 170.750 89.940 171.030 ;
        RECT 86.440 169.390 86.720 169.670 ;
        RECT 85.520 168.030 85.800 168.310 ;
        RECT 91.040 170.070 91.320 170.350 ;
        RECT 93.340 175.510 93.620 175.790 ;
        RECT 100.240 202.710 100.520 202.990 ;
        RECT 99.320 195.230 99.600 195.510 ;
        RECT 99.780 194.550 100.060 194.830 ;
        RECT 98.860 189.790 99.140 190.070 ;
        RECT 97.940 188.430 98.220 188.710 ;
        RECT 100.700 197.270 100.980 197.550 ;
        RECT 99.780 187.750 100.060 188.030 ;
        RECT 98.400 187.070 98.680 187.350 ;
        RECT 99.780 183.670 100.060 183.950 ;
        RECT 99.320 182.310 99.600 182.590 ;
        RECT 102.540 186.390 102.820 186.670 ;
        RECT 104.770 207.130 105.050 207.410 ;
        RECT 105.170 207.130 105.450 207.410 ;
        RECT 105.570 207.130 105.850 207.410 ;
        RECT 105.970 207.130 106.250 207.410 ;
        RECT 106.370 207.130 106.650 207.410 ;
        RECT 104.840 202.710 105.120 202.990 ;
        RECT 104.770 201.690 105.050 201.970 ;
        RECT 105.170 201.690 105.450 201.970 ;
        RECT 105.570 201.690 105.850 201.970 ;
        RECT 105.970 201.690 106.250 201.970 ;
        RECT 106.370 201.690 106.650 201.970 ;
        RECT 113.120 203.390 113.400 203.670 ;
        RECT 119.770 204.410 120.050 204.690 ;
        RECT 120.170 204.410 120.450 204.690 ;
        RECT 120.570 204.410 120.850 204.690 ;
        RECT 120.970 204.410 121.250 204.690 ;
        RECT 121.370 204.410 121.650 204.690 ;
        RECT 103.460 196.590 103.740 196.870 ;
        RECT 103.460 195.230 103.740 195.510 ;
        RECT 97.020 176.190 97.300 176.470 ;
        RECT 90.580 169.390 90.860 169.670 ;
        RECT 89.770 166.330 90.050 166.610 ;
        RECT 90.170 166.330 90.450 166.610 ;
        RECT 90.570 166.330 90.850 166.610 ;
        RECT 90.970 166.330 91.250 166.610 ;
        RECT 91.370 166.330 91.650 166.610 ;
        RECT 94.260 173.470 94.540 173.750 ;
        RECT 95.640 174.830 95.920 175.110 ;
        RECT 89.770 160.890 90.050 161.170 ;
        RECT 90.170 160.890 90.450 161.170 ;
        RECT 90.570 160.890 90.850 161.170 ;
        RECT 90.970 160.890 91.250 161.170 ;
        RECT 91.370 160.890 91.650 161.170 ;
        RECT 76.780 129.270 77.060 129.550 ;
        RECT 74.770 125.530 75.050 125.810 ;
        RECT 75.170 125.530 75.450 125.810 ;
        RECT 75.570 125.530 75.850 125.810 ;
        RECT 75.970 125.530 76.250 125.810 ;
        RECT 76.370 125.530 76.650 125.810 ;
        RECT 89.770 155.450 90.050 155.730 ;
        RECT 90.170 155.450 90.450 155.730 ;
        RECT 90.570 155.450 90.850 155.730 ;
        RECT 90.970 155.450 91.250 155.730 ;
        RECT 91.370 155.450 91.650 155.730 ;
        RECT 88.740 144.910 89.020 145.190 ;
        RECT 89.770 150.010 90.050 150.290 ;
        RECT 90.170 150.010 90.450 150.290 ;
        RECT 90.570 150.010 90.850 150.290 ;
        RECT 90.970 150.010 91.250 150.290 ;
        RECT 91.370 150.010 91.650 150.290 ;
        RECT 89.770 144.570 90.050 144.850 ;
        RECT 90.170 144.570 90.450 144.850 ;
        RECT 90.570 144.570 90.850 144.850 ;
        RECT 90.970 144.570 91.250 144.850 ;
        RECT 91.370 144.570 91.650 144.850 ;
        RECT 89.770 139.130 90.050 139.410 ;
        RECT 90.170 139.130 90.450 139.410 ;
        RECT 90.570 139.130 90.850 139.410 ;
        RECT 90.970 139.130 91.250 139.410 ;
        RECT 91.370 139.130 91.650 139.410 ;
        RECT 90.120 136.750 90.400 137.030 ;
        RECT 92.880 145.590 93.160 145.870 ;
        RECT 92.420 142.870 92.700 143.150 ;
        RECT 92.420 140.150 92.700 140.430 ;
        RECT 85.520 132.670 85.800 132.950 ;
        RECT 89.770 133.690 90.050 133.970 ;
        RECT 90.170 133.690 90.450 133.970 ;
        RECT 90.570 133.690 90.850 133.970 ;
        RECT 90.970 133.690 91.250 133.970 ;
        RECT 91.370 133.690 91.650 133.970 ;
        RECT 88.280 127.230 88.560 127.510 ;
        RECT 89.770 128.250 90.050 128.530 ;
        RECT 90.170 128.250 90.450 128.530 ;
        RECT 90.570 128.250 90.850 128.530 ;
        RECT 90.970 128.250 91.250 128.530 ;
        RECT 91.370 128.250 91.650 128.530 ;
        RECT 97.480 161.910 97.760 162.190 ;
        RECT 98.400 177.550 98.680 177.830 ;
        RECT 104.770 196.250 105.050 196.530 ;
        RECT 105.170 196.250 105.450 196.530 ;
        RECT 105.570 196.250 105.850 196.530 ;
        RECT 105.970 196.250 106.250 196.530 ;
        RECT 106.370 196.250 106.650 196.530 ;
        RECT 106.680 194.550 106.960 194.830 ;
        RECT 104.380 191.830 104.660 192.110 ;
        RECT 104.770 190.810 105.050 191.090 ;
        RECT 105.170 190.810 105.450 191.090 ;
        RECT 105.570 190.810 105.850 191.090 ;
        RECT 105.970 190.810 106.250 191.090 ;
        RECT 106.370 190.810 106.650 191.090 ;
        RECT 107.140 190.470 107.420 190.750 ;
        RECT 105.300 189.790 105.580 190.070 ;
        RECT 106.220 189.790 106.500 190.070 ;
        RECT 104.770 185.370 105.050 185.650 ;
        RECT 105.170 185.370 105.450 185.650 ;
        RECT 105.570 185.370 105.850 185.650 ;
        RECT 105.970 185.370 106.250 185.650 ;
        RECT 106.370 185.370 106.650 185.650 ;
        RECT 109.900 194.550 110.180 194.830 ;
        RECT 109.900 191.150 110.180 191.430 ;
        RECT 102.540 178.910 102.820 179.190 ;
        RECT 107.600 182.990 107.880 183.270 ;
        RECT 107.600 182.310 107.880 182.590 ;
        RECT 99.780 173.470 100.060 173.750 ;
        RECT 98.860 172.110 99.140 172.390 ;
        RECT 101.620 175.510 101.900 175.790 ;
        RECT 103.000 174.150 103.280 174.430 ;
        RECT 102.080 170.070 102.360 170.350 ;
        RECT 93.800 135.390 94.080 135.670 ;
        RECT 97.020 142.870 97.300 143.150 ;
        RECT 96.100 139.470 96.380 139.750 ;
        RECT 100.240 164.630 100.520 164.910 ;
        RECT 104.770 179.930 105.050 180.210 ;
        RECT 105.170 179.930 105.450 180.210 ;
        RECT 105.570 179.930 105.850 180.210 ;
        RECT 105.970 179.930 106.250 180.210 ;
        RECT 106.370 179.930 106.650 180.210 ;
        RECT 104.380 178.910 104.660 179.190 ;
        RECT 106.220 178.910 106.500 179.190 ;
        RECT 108.060 176.190 108.340 176.470 ;
        RECT 104.770 174.490 105.050 174.770 ;
        RECT 105.170 174.490 105.450 174.770 ;
        RECT 105.570 174.490 105.850 174.770 ;
        RECT 105.970 174.490 106.250 174.770 ;
        RECT 106.370 174.490 106.650 174.770 ;
        RECT 108.520 174.830 108.800 175.110 ;
        RECT 101.620 162.590 101.900 162.870 ;
        RECT 106.220 170.070 106.500 170.350 ;
        RECT 104.770 169.050 105.050 169.330 ;
        RECT 105.170 169.050 105.450 169.330 ;
        RECT 105.570 169.050 105.850 169.330 ;
        RECT 105.970 169.050 106.250 169.330 ;
        RECT 106.370 169.050 106.650 169.330 ;
        RECT 104.770 163.610 105.050 163.890 ;
        RECT 105.170 163.610 105.450 163.890 ;
        RECT 105.570 163.610 105.850 163.890 ;
        RECT 105.970 163.610 106.250 163.890 ;
        RECT 106.370 163.610 106.650 163.890 ;
        RECT 104.840 162.590 105.120 162.870 ;
        RECT 105.300 161.910 105.580 162.190 ;
        RECT 104.770 158.170 105.050 158.450 ;
        RECT 105.170 158.170 105.450 158.450 ;
        RECT 105.570 158.170 105.850 158.450 ;
        RECT 105.970 158.170 106.250 158.450 ;
        RECT 106.370 158.170 106.650 158.450 ;
        RECT 105.300 156.470 105.580 156.750 ;
        RECT 97.020 133.350 97.300 133.630 ;
        RECT 92.880 129.270 93.160 129.550 ;
        RECT 91.960 127.230 92.240 127.510 ;
        RECT 98.400 131.990 98.680 132.270 ;
        RECT 100.700 140.830 100.980 141.110 ;
        RECT 99.780 127.910 100.060 128.190 ;
        RECT 103.000 143.550 103.280 143.830 ;
        RECT 106.680 153.750 106.960 154.030 ;
        RECT 104.770 152.730 105.050 153.010 ;
        RECT 105.170 152.730 105.450 153.010 ;
        RECT 105.570 152.730 105.850 153.010 ;
        RECT 105.970 152.730 106.250 153.010 ;
        RECT 106.370 152.730 106.650 153.010 ;
        RECT 104.770 147.290 105.050 147.570 ;
        RECT 105.170 147.290 105.450 147.570 ;
        RECT 105.570 147.290 105.850 147.570 ;
        RECT 105.970 147.290 106.250 147.570 ;
        RECT 106.370 147.290 106.650 147.570 ;
        RECT 105.760 145.590 106.040 145.870 ;
        RECT 108.520 168.030 108.800 168.310 ;
        RECT 107.600 145.590 107.880 145.870 ;
        RECT 107.600 144.230 107.880 144.510 ;
        RECT 104.770 141.850 105.050 142.130 ;
        RECT 105.170 141.850 105.450 142.130 ;
        RECT 105.570 141.850 105.850 142.130 ;
        RECT 105.970 141.850 106.250 142.130 ;
        RECT 106.370 141.850 106.650 142.130 ;
        RECT 106.680 140.150 106.960 140.430 ;
        RECT 104.770 136.410 105.050 136.690 ;
        RECT 105.170 136.410 105.450 136.690 ;
        RECT 105.570 136.410 105.850 136.690 ;
        RECT 105.970 136.410 106.250 136.690 ;
        RECT 106.370 136.410 106.650 136.690 ;
        RECT 107.140 135.390 107.420 135.670 ;
        RECT 106.220 134.710 106.500 134.990 ;
        RECT 104.770 130.970 105.050 131.250 ;
        RECT 105.170 130.970 105.450 131.250 ;
        RECT 105.570 130.970 105.850 131.250 ;
        RECT 105.970 130.970 106.250 131.250 ;
        RECT 106.370 130.970 106.650 131.250 ;
        RECT 111.280 191.150 111.560 191.430 ;
        RECT 111.280 187.070 111.560 187.350 ;
        RECT 111.280 185.710 111.560 185.990 ;
        RECT 111.280 183.670 111.560 183.950 ;
        RECT 109.440 180.270 109.720 180.550 ;
        RECT 110.360 172.110 110.640 172.390 ;
        RECT 110.360 162.590 110.640 162.870 ;
        RECT 110.360 159.190 110.640 159.470 ;
        RECT 108.980 144.910 109.260 145.190 ;
        RECT 108.060 127.910 108.340 128.190 ;
        RECT 109.900 151.030 110.180 151.310 ;
        RECT 109.900 147.630 110.180 147.910 ;
        RECT 110.820 146.950 111.100 147.230 ;
        RECT 119.770 198.970 120.050 199.250 ;
        RECT 120.170 198.970 120.450 199.250 ;
        RECT 120.570 198.970 120.850 199.250 ;
        RECT 120.970 198.970 121.250 199.250 ;
        RECT 121.370 198.970 121.650 199.250 ;
        RECT 114.500 195.230 114.780 195.510 ;
        RECT 113.580 185.710 113.860 185.990 ;
        RECT 111.280 146.270 111.560 146.550 ;
        RECT 110.360 145.590 110.640 145.870 ;
        RECT 110.360 143.550 110.640 143.830 ;
        RECT 110.360 142.870 110.640 143.150 ;
        RECT 116.340 188.430 116.620 188.710 ;
        RECT 115.880 187.750 116.160 188.030 ;
        RECT 118.180 187.070 118.460 187.350 ;
        RECT 119.770 193.530 120.050 193.810 ;
        RECT 120.170 193.530 120.450 193.810 ;
        RECT 120.570 193.530 120.850 193.810 ;
        RECT 120.970 193.530 121.250 193.810 ;
        RECT 121.370 193.530 121.650 193.810 ;
        RECT 120.480 192.510 120.760 192.790 ;
        RECT 120.940 191.830 121.220 192.110 ;
        RECT 119.770 188.090 120.050 188.370 ;
        RECT 120.170 188.090 120.450 188.370 ;
        RECT 120.570 188.090 120.850 188.370 ;
        RECT 120.970 188.090 121.250 188.370 ;
        RECT 121.370 188.090 121.650 188.370 ;
        RECT 119.560 186.390 119.840 186.670 ;
        RECT 114.500 180.270 114.780 180.550 ;
        RECT 114.960 178.910 115.240 179.190 ;
        RECT 113.120 174.830 113.400 175.110 ;
        RECT 116.800 176.190 117.080 176.470 ;
        RECT 116.340 172.110 116.620 172.390 ;
        RECT 112.660 165.310 112.940 165.590 ;
        RECT 116.340 170.750 116.620 171.030 ;
        RECT 116.800 165.310 117.080 165.590 ;
        RECT 115.880 157.150 116.160 157.430 ;
        RECT 113.580 156.470 113.860 156.750 ;
        RECT 112.660 152.390 112.940 152.670 ;
        RECT 113.580 151.710 113.860 151.990 ;
        RECT 113.120 151.030 113.400 151.310 ;
        RECT 112.660 147.630 112.940 147.910 ;
        RECT 113.120 140.830 113.400 141.110 ;
        RECT 113.580 139.470 113.860 139.750 ;
        RECT 110.820 129.270 111.100 129.550 ;
        RECT 113.120 132.670 113.400 132.950 ;
        RECT 116.800 157.150 117.080 157.430 ;
        RECT 119.770 182.650 120.050 182.930 ;
        RECT 120.170 182.650 120.450 182.930 ;
        RECT 120.570 182.650 120.850 182.930 ;
        RECT 120.970 182.650 121.250 182.930 ;
        RECT 121.370 182.650 121.650 182.930 ;
        RECT 119.770 177.210 120.050 177.490 ;
        RECT 120.170 177.210 120.450 177.490 ;
        RECT 120.570 177.210 120.850 177.490 ;
        RECT 120.970 177.210 121.250 177.490 ;
        RECT 121.370 177.210 121.650 177.490 ;
        RECT 119.770 171.770 120.050 172.050 ;
        RECT 120.170 171.770 120.450 172.050 ;
        RECT 120.570 171.770 120.850 172.050 ;
        RECT 120.970 171.770 121.250 172.050 ;
        RECT 121.370 171.770 121.650 172.050 ;
        RECT 124.620 197.950 124.900 198.230 ;
        RECT 125.540 197.270 125.820 197.550 ;
        RECT 123.700 189.790 123.980 190.070 ;
        RECT 122.780 183.670 123.060 183.950 ;
        RECT 119.100 168.030 119.380 168.310 ;
        RECT 119.770 166.330 120.050 166.610 ;
        RECT 120.170 166.330 120.450 166.610 ;
        RECT 120.570 166.330 120.850 166.610 ;
        RECT 120.970 166.330 121.250 166.610 ;
        RECT 121.370 166.330 121.650 166.610 ;
        RECT 119.100 165.310 119.380 165.590 ;
        RECT 121.860 164.630 122.140 164.910 ;
        RECT 119.100 161.910 119.380 162.190 ;
        RECT 119.770 160.890 120.050 161.170 ;
        RECT 120.170 160.890 120.450 161.170 ;
        RECT 120.570 160.890 120.850 161.170 ;
        RECT 120.970 160.890 121.250 161.170 ;
        RECT 121.370 160.890 121.650 161.170 ;
        RECT 119.770 155.450 120.050 155.730 ;
        RECT 120.170 155.450 120.450 155.730 ;
        RECT 120.570 155.450 120.850 155.730 ;
        RECT 120.970 155.450 121.250 155.730 ;
        RECT 121.370 155.450 121.650 155.730 ;
        RECT 117.720 153.070 118.000 153.350 ;
        RECT 117.260 146.270 117.540 146.550 ;
        RECT 116.340 145.590 116.620 145.870 ;
        RECT 113.580 131.990 113.860 132.270 ;
        RECT 89.770 122.810 90.050 123.090 ;
        RECT 90.170 122.810 90.450 123.090 ;
        RECT 90.570 122.810 90.850 123.090 ;
        RECT 90.970 122.810 91.250 123.090 ;
        RECT 91.370 122.810 91.650 123.090 ;
        RECT 104.770 125.530 105.050 125.810 ;
        RECT 105.170 125.530 105.450 125.810 ;
        RECT 105.570 125.530 105.850 125.810 ;
        RECT 105.970 125.530 106.250 125.810 ;
        RECT 106.370 125.530 106.650 125.810 ;
        RECT 116.800 136.750 117.080 137.030 ;
        RECT 116.800 128.590 117.080 128.870 ;
        RECT 116.340 127.910 116.620 128.190 ;
        RECT 116.340 125.870 116.620 126.150 ;
        RECT 120.020 153.750 120.300 154.030 ;
        RECT 119.770 150.010 120.050 150.290 ;
        RECT 120.170 150.010 120.450 150.290 ;
        RECT 120.570 150.010 120.850 150.290 ;
        RECT 120.970 150.010 121.250 150.290 ;
        RECT 121.370 150.010 121.650 150.290 ;
        RECT 119.770 144.570 120.050 144.850 ;
        RECT 120.170 144.570 120.450 144.850 ;
        RECT 120.570 144.570 120.850 144.850 ;
        RECT 120.970 144.570 121.250 144.850 ;
        RECT 121.370 144.570 121.650 144.850 ;
        RECT 119.770 139.130 120.050 139.410 ;
        RECT 120.170 139.130 120.450 139.410 ;
        RECT 120.570 139.130 120.850 139.410 ;
        RECT 120.970 139.130 121.250 139.410 ;
        RECT 121.370 139.130 121.650 139.410 ;
        RECT 119.770 133.690 120.050 133.970 ;
        RECT 120.170 133.690 120.450 133.970 ;
        RECT 120.570 133.690 120.850 133.970 ;
        RECT 120.970 133.690 121.250 133.970 ;
        RECT 121.370 133.690 121.650 133.970 ;
        RECT 134.770 207.130 135.050 207.410 ;
        RECT 135.170 207.130 135.450 207.410 ;
        RECT 135.570 207.130 135.850 207.410 ;
        RECT 135.970 207.130 136.250 207.410 ;
        RECT 136.370 207.130 136.650 207.410 ;
        RECT 127.840 192.510 128.120 192.790 ;
        RECT 127.380 187.070 127.660 187.350 ;
        RECT 129.220 196.590 129.500 196.870 ;
        RECT 128.760 191.830 129.040 192.110 ;
        RECT 128.300 190.470 128.580 190.750 ;
        RECT 134.770 201.690 135.050 201.970 ;
        RECT 135.170 201.690 135.450 201.970 ;
        RECT 135.570 201.690 135.850 201.970 ;
        RECT 135.970 201.690 136.250 201.970 ;
        RECT 136.370 201.690 136.650 201.970 ;
        RECT 132.900 197.270 133.180 197.550 ;
        RECT 132.440 196.590 132.720 196.870 ;
        RECT 131.060 194.550 131.340 194.830 ;
        RECT 130.600 189.110 130.880 189.390 ;
        RECT 122.320 130.630 122.600 130.910 ;
        RECT 119.770 128.250 120.050 128.530 ;
        RECT 120.170 128.250 120.450 128.530 ;
        RECT 120.570 128.250 120.850 128.530 ;
        RECT 120.970 128.250 121.250 128.530 ;
        RECT 121.370 128.250 121.650 128.530 ;
        RECT 121.400 126.550 121.680 126.830 ;
        RECT 123.240 126.550 123.520 126.830 ;
        RECT 125.080 150.350 125.360 150.630 ;
        RECT 126.920 156.470 127.200 156.750 ;
        RECT 129.220 175.510 129.500 175.790 ;
        RECT 129.680 172.790 129.960 173.070 ;
        RECT 131.060 188.430 131.340 188.710 ;
        RECT 130.600 184.350 130.880 184.630 ;
        RECT 131.060 178.910 131.340 179.190 ;
        RECT 134.280 197.950 134.560 198.230 ;
        RECT 134.770 196.250 135.050 196.530 ;
        RECT 135.170 196.250 135.450 196.530 ;
        RECT 135.570 196.250 135.850 196.530 ;
        RECT 135.970 196.250 136.250 196.530 ;
        RECT 136.370 196.250 136.650 196.530 ;
        RECT 134.740 194.550 135.020 194.830 ;
        RECT 137.500 195.230 137.780 195.510 ;
        RECT 130.140 165.310 130.420 165.590 ;
        RECT 131.980 168.030 132.260 168.310 ;
        RECT 131.060 161.910 131.340 162.190 ;
        RECT 127.840 147.630 128.120 147.910 ;
        RECT 128.760 157.150 129.040 157.430 ;
        RECT 128.760 148.990 129.040 149.270 ;
        RECT 129.220 138.110 129.500 138.390 ;
        RECT 124.620 129.950 124.900 130.230 ;
        RECT 119.770 122.810 120.050 123.090 ;
        RECT 120.170 122.810 120.450 123.090 ;
        RECT 120.570 122.810 120.850 123.090 ;
        RECT 120.970 122.810 121.250 123.090 ;
        RECT 121.370 122.810 121.650 123.090 ;
        RECT 131.980 151.710 132.260 151.990 ;
        RECT 131.060 148.990 131.340 149.270 ;
        RECT 129.680 134.710 129.960 134.990 ;
        RECT 130.600 131.990 130.880 132.270 ;
        RECT 131.980 148.310 132.260 148.590 ;
        RECT 134.770 190.810 135.050 191.090 ;
        RECT 135.170 190.810 135.450 191.090 ;
        RECT 135.570 190.810 135.850 191.090 ;
        RECT 135.970 190.810 136.250 191.090 ;
        RECT 136.370 190.810 136.650 191.090 ;
        RECT 137.960 188.430 138.240 188.710 ;
        RECT 134.770 185.370 135.050 185.650 ;
        RECT 135.170 185.370 135.450 185.650 ;
        RECT 135.570 185.370 135.850 185.650 ;
        RECT 135.970 185.370 136.250 185.650 ;
        RECT 136.370 185.370 136.650 185.650 ;
        RECT 149.770 204.410 150.050 204.690 ;
        RECT 150.170 204.410 150.450 204.690 ;
        RECT 150.570 204.410 150.850 204.690 ;
        RECT 150.970 204.410 151.250 204.690 ;
        RECT 151.370 204.410 151.650 204.690 ;
        RECT 149.770 198.970 150.050 199.250 ;
        RECT 150.170 198.970 150.450 199.250 ;
        RECT 150.570 198.970 150.850 199.250 ;
        RECT 150.970 198.970 151.250 199.250 ;
        RECT 151.370 198.970 151.650 199.250 ;
        RECT 134.770 179.930 135.050 180.210 ;
        RECT 135.170 179.930 135.450 180.210 ;
        RECT 135.570 179.930 135.850 180.210 ;
        RECT 135.970 179.930 136.250 180.210 ;
        RECT 136.370 179.930 136.650 180.210 ;
        RECT 136.120 175.510 136.400 175.790 ;
        RECT 134.770 174.490 135.050 174.770 ;
        RECT 135.170 174.490 135.450 174.770 ;
        RECT 135.570 174.490 135.850 174.770 ;
        RECT 135.970 174.490 136.250 174.770 ;
        RECT 136.370 174.490 136.650 174.770 ;
        RECT 134.740 173.470 135.020 173.750 ;
        RECT 134.770 169.050 135.050 169.330 ;
        RECT 135.170 169.050 135.450 169.330 ;
        RECT 135.570 169.050 135.850 169.330 ;
        RECT 135.970 169.050 136.250 169.330 ;
        RECT 136.370 169.050 136.650 169.330 ;
        RECT 133.820 164.630 134.100 164.910 ;
        RECT 134.770 163.610 135.050 163.890 ;
        RECT 135.170 163.610 135.450 163.890 ;
        RECT 135.570 163.610 135.850 163.890 ;
        RECT 135.970 163.610 136.250 163.890 ;
        RECT 136.370 163.610 136.650 163.890 ;
        RECT 132.900 149.670 133.180 149.950 ;
        RECT 131.980 147.630 132.260 147.910 ;
        RECT 132.440 146.950 132.720 147.230 ;
        RECT 132.900 136.070 133.180 136.350 ;
        RECT 129.680 129.270 129.960 129.550 ;
        RECT 131.980 129.950 132.260 130.230 ;
        RECT 134.770 158.170 135.050 158.450 ;
        RECT 135.170 158.170 135.450 158.450 ;
        RECT 135.570 158.170 135.850 158.450 ;
        RECT 135.970 158.170 136.250 158.450 ;
        RECT 136.370 158.170 136.650 158.450 ;
        RECT 134.770 152.730 135.050 153.010 ;
        RECT 135.170 152.730 135.450 153.010 ;
        RECT 135.570 152.730 135.850 153.010 ;
        RECT 135.970 152.730 136.250 153.010 ;
        RECT 136.370 152.730 136.650 153.010 ;
        RECT 136.120 151.030 136.400 151.310 ;
        RECT 135.660 148.990 135.940 149.270 ;
        RECT 134.770 147.290 135.050 147.570 ;
        RECT 135.170 147.290 135.450 147.570 ;
        RECT 135.570 147.290 135.850 147.570 ;
        RECT 135.970 147.290 136.250 147.570 ;
        RECT 136.370 147.290 136.650 147.570 ;
        RECT 134.740 145.590 135.020 145.870 ;
        RECT 134.770 141.850 135.050 142.130 ;
        RECT 135.170 141.850 135.450 142.130 ;
        RECT 135.570 141.850 135.850 142.130 ;
        RECT 135.970 141.850 136.250 142.130 ;
        RECT 136.370 141.850 136.650 142.130 ;
        RECT 139.800 178.230 140.080 178.510 ;
        RECT 139.340 176.190 139.620 176.470 ;
        RECT 139.800 157.150 140.080 157.430 ;
        RECT 138.880 155.790 139.160 156.070 ;
        RECT 138.880 150.350 139.160 150.630 ;
        RECT 138.420 148.310 138.700 148.590 ;
        RECT 142.100 162.590 142.380 162.870 ;
        RECT 133.360 130.630 133.640 130.910 ;
        RECT 134.770 136.410 135.050 136.690 ;
        RECT 135.170 136.410 135.450 136.690 ;
        RECT 135.570 136.410 135.850 136.690 ;
        RECT 135.970 136.410 136.250 136.690 ;
        RECT 136.370 136.410 136.650 136.690 ;
        RECT 137.040 135.390 137.320 135.670 ;
        RECT 134.770 130.970 135.050 131.250 ;
        RECT 135.170 130.970 135.450 131.250 ;
        RECT 135.570 130.970 135.850 131.250 ;
        RECT 135.970 130.970 136.250 131.250 ;
        RECT 136.370 130.970 136.650 131.250 ;
        RECT 134.740 129.950 135.020 130.230 ;
        RECT 137.500 131.310 137.780 131.590 ;
        RECT 137.040 128.590 137.320 128.870 ;
        RECT 137.500 127.910 137.780 128.190 ;
        RECT 134.770 125.530 135.050 125.810 ;
        RECT 135.170 125.530 135.450 125.810 ;
        RECT 135.570 125.530 135.850 125.810 ;
        RECT 135.970 125.530 136.250 125.810 ;
        RECT 136.370 125.530 136.650 125.810 ;
        RECT 138.880 135.390 139.160 135.670 ;
        RECT 137.960 125.870 138.240 126.150 ;
        RECT 140.720 138.110 141.000 138.390 ;
        RECT 142.560 155.110 142.840 155.390 ;
        RECT 142.100 151.710 142.380 151.990 ;
        RECT 140.720 133.350 141.000 133.630 ;
        RECT 143.940 140.150 144.220 140.430 ;
        RECT 146.700 191.830 146.980 192.110 ;
        RECT 149.770 193.530 150.050 193.810 ;
        RECT 150.170 193.530 150.450 193.810 ;
        RECT 150.570 193.530 150.850 193.810 ;
        RECT 150.970 193.530 151.250 193.810 ;
        RECT 151.370 193.530 151.650 193.810 ;
        RECT 152.680 192.510 152.960 192.790 ;
        RECT 148.540 188.430 148.820 188.710 ;
        RECT 149.770 188.090 150.050 188.370 ;
        RECT 150.170 188.090 150.450 188.370 ;
        RECT 150.570 188.090 150.850 188.370 ;
        RECT 150.970 188.090 151.250 188.370 ;
        RECT 151.370 188.090 151.650 188.370 ;
        RECT 149.770 182.650 150.050 182.930 ;
        RECT 150.170 182.650 150.450 182.930 ;
        RECT 150.570 182.650 150.850 182.930 ;
        RECT 150.970 182.650 151.250 182.930 ;
        RECT 151.370 182.650 151.650 182.930 ;
        RECT 146.700 165.310 146.980 165.590 ;
        RECT 146.700 162.590 146.980 162.870 ;
        RECT 149.770 177.210 150.050 177.490 ;
        RECT 150.170 177.210 150.450 177.490 ;
        RECT 150.570 177.210 150.850 177.490 ;
        RECT 150.970 177.210 151.250 177.490 ;
        RECT 151.370 177.210 151.650 177.490 ;
        RECT 150.840 175.510 151.120 175.790 ;
        RECT 149.770 171.770 150.050 172.050 ;
        RECT 150.170 171.770 150.450 172.050 ;
        RECT 150.570 171.770 150.850 172.050 ;
        RECT 150.970 171.770 151.250 172.050 ;
        RECT 151.370 171.770 151.650 172.050 ;
        RECT 149.000 168.030 149.280 168.310 ;
        RECT 149.770 166.330 150.050 166.610 ;
        RECT 150.170 166.330 150.450 166.610 ;
        RECT 150.570 166.330 150.850 166.610 ;
        RECT 150.970 166.330 151.250 166.610 ;
        RECT 151.370 166.330 151.650 166.610 ;
        RECT 149.770 160.890 150.050 161.170 ;
        RECT 150.170 160.890 150.450 161.170 ;
        RECT 150.570 160.890 150.850 161.170 ;
        RECT 150.970 160.890 151.250 161.170 ;
        RECT 151.370 160.890 151.650 161.170 ;
        RECT 149.770 155.450 150.050 155.730 ;
        RECT 150.170 155.450 150.450 155.730 ;
        RECT 150.570 155.450 150.850 155.730 ;
        RECT 150.970 155.450 151.250 155.730 ;
        RECT 151.370 155.450 151.650 155.730 ;
        RECT 149.770 150.010 150.050 150.290 ;
        RECT 150.170 150.010 150.450 150.290 ;
        RECT 150.570 150.010 150.850 150.290 ;
        RECT 150.970 150.010 151.250 150.290 ;
        RECT 151.370 150.010 151.650 150.290 ;
        RECT 152.220 148.990 152.500 149.270 ;
        RECT 149.770 144.570 150.050 144.850 ;
        RECT 150.170 144.570 150.450 144.850 ;
        RECT 150.570 144.570 150.850 144.850 ;
        RECT 150.970 144.570 151.250 144.850 ;
        RECT 151.370 144.570 151.650 144.850 ;
        RECT 145.780 139.470 146.060 139.750 ;
        RECT 144.400 134.710 144.680 134.990 ;
        RECT 142.560 129.270 142.840 129.550 ;
        RECT 143.480 126.550 143.760 126.830 ;
        RECT 149.770 139.130 150.050 139.410 ;
        RECT 150.170 139.130 150.450 139.410 ;
        RECT 150.570 139.130 150.850 139.410 ;
        RECT 150.970 139.130 151.250 139.410 ;
        RECT 151.370 139.130 151.650 139.410 ;
        RECT 144.400 130.630 144.680 130.910 ;
        RECT 143.940 125.870 144.220 126.150 ;
        RECT 145.320 129.270 145.600 129.550 ;
        RECT 146.240 130.630 146.520 130.910 ;
        RECT 146.700 128.590 146.980 128.870 ;
        RECT 146.240 127.230 146.520 127.510 ;
        RECT 148.080 131.310 148.360 131.590 ;
        RECT 149.770 133.690 150.050 133.970 ;
        RECT 150.170 133.690 150.450 133.970 ;
        RECT 150.570 133.690 150.850 133.970 ;
        RECT 150.970 133.690 151.250 133.970 ;
        RECT 151.370 133.690 151.650 133.970 ;
        RECT 149.000 129.270 149.280 129.550 ;
        RECT 149.770 128.250 150.050 128.530 ;
        RECT 150.170 128.250 150.450 128.530 ;
        RECT 150.570 128.250 150.850 128.530 ;
        RECT 150.970 128.250 151.250 128.530 ;
        RECT 151.370 128.250 151.650 128.530 ;
        RECT 149.770 122.810 150.050 123.090 ;
        RECT 150.170 122.810 150.450 123.090 ;
        RECT 150.570 122.810 150.850 123.090 ;
        RECT 150.970 122.810 151.250 123.090 ;
        RECT 151.370 122.810 151.650 123.090 ;
      LAYER met3 ;
        RECT 127.805 221.495 128.200 221.500 ;
        RECT 127.780 221.110 128.225 221.495 ;
        RECT 125.375 216.910 125.785 216.935 ;
        RECT 121.990 216.490 125.790 216.910 ;
        RECT 126.495 216.900 126.905 216.905 ;
        RECT 126.470 216.500 126.930 216.900 ;
        RECT 125.375 216.465 125.785 216.490 ;
        RECT 120.495 215.415 120.910 215.440 ;
        RECT 110.245 215.360 110.755 215.385 ;
        RECT 110.240 214.140 110.760 215.360 ;
        RECT 116.605 215.300 116.995 215.325 ;
        RECT 113.800 214.900 117.000 215.300 ;
        RECT 118.290 214.990 120.915 215.415 ;
        RECT 120.495 214.965 120.910 214.990 ;
        RECT 116.605 214.875 116.995 214.900 ;
        RECT 126.495 214.195 126.905 216.500 ;
        RECT 127.805 214.205 128.200 221.110 ;
        RECT 131.910 220.490 132.295 220.495 ;
        RECT 131.885 220.115 132.320 220.490 ;
        RECT 131.910 214.210 132.295 220.115 ;
        RECT 135.965 214.165 136.440 219.340 ;
        RECT 140.205 217.995 140.600 218.000 ;
        RECT 140.180 217.610 140.625 217.995 ;
        RECT 140.205 214.205 140.600 217.610 ;
        RECT 144.270 216.825 144.730 216.830 ;
        RECT 144.245 216.375 144.755 216.825 ;
        RECT 144.270 214.170 144.730 216.375 ;
        RECT 152.570 215.625 153.030 215.630 ;
        RECT 148.485 215.610 148.915 215.615 ;
        RECT 148.460 215.190 148.940 215.610 ;
        RECT 148.485 214.185 148.915 215.190 ;
        RECT 152.545 215.175 153.055 215.625 ;
        RECT 152.570 214.170 153.030 215.175 ;
        RECT 74.720 207.105 76.700 207.435 ;
        RECT 104.720 207.105 106.700 207.435 ;
        RECT 134.720 207.105 136.700 207.435 ;
        RECT 89.720 204.385 91.700 204.715 ;
        RECT 119.720 204.385 121.700 204.715 ;
        RECT 149.720 204.385 151.700 204.715 ;
        RECT 92.395 203.680 92.725 203.695 ;
        RECT 100.420 203.680 100.800 203.690 ;
        RECT 92.395 203.380 100.800 203.680 ;
        RECT 92.395 203.365 92.725 203.380 ;
        RECT 100.420 203.370 100.800 203.380 ;
        RECT 111.460 203.680 111.840 203.690 ;
        RECT 113.095 203.680 113.425 203.695 ;
        RECT 111.460 203.380 113.425 203.680 ;
        RECT 111.460 203.370 111.840 203.380 ;
        RECT 113.095 203.365 113.425 203.380 ;
        RECT 100.215 203.000 100.545 203.015 ;
        RECT 104.815 203.000 105.145 203.015 ;
        RECT 100.215 202.700 105.145 203.000 ;
        RECT 100.215 202.685 100.545 202.700 ;
        RECT 104.815 202.685 105.145 202.700 ;
        RECT 74.720 201.665 76.700 201.995 ;
        RECT 104.720 201.665 106.700 201.995 ;
        RECT 134.720 201.665 136.700 201.995 ;
        RECT 89.720 198.945 91.700 199.275 ;
        RECT 119.720 198.945 121.700 199.275 ;
        RECT 149.720 198.945 151.700 199.275 ;
        RECT 78.135 198.920 78.465 198.935 ;
        RECT 84.115 198.920 84.445 198.935 ;
        RECT 78.135 198.620 84.445 198.920 ;
        RECT 78.135 198.605 78.465 198.620 ;
        RECT 84.115 198.605 84.445 198.620 ;
        RECT 124.595 198.240 124.925 198.255 ;
        RECT 134.255 198.240 134.585 198.255 ;
        RECT 124.595 197.940 134.585 198.240 ;
        RECT 124.595 197.925 124.925 197.940 ;
        RECT 134.255 197.925 134.585 197.940 ;
        RECT 100.675 197.560 101.005 197.575 ;
        RECT 114.220 197.560 114.600 197.570 ;
        RECT 100.675 197.260 114.600 197.560 ;
        RECT 100.675 197.245 101.005 197.260 ;
        RECT 114.220 197.250 114.600 197.260 ;
        RECT 125.515 197.560 125.845 197.575 ;
        RECT 132.875 197.560 133.205 197.575 ;
        RECT 125.515 197.260 133.205 197.560 ;
        RECT 125.515 197.245 125.845 197.260 ;
        RECT 132.875 197.245 133.205 197.260 ;
        RECT 98.580 196.880 98.960 196.890 ;
        RECT 103.435 196.880 103.765 196.895 ;
        RECT 98.580 196.580 103.765 196.880 ;
        RECT 98.580 196.570 98.960 196.580 ;
        RECT 103.435 196.565 103.765 196.580 ;
        RECT 124.340 196.880 124.720 196.890 ;
        RECT 129.195 196.880 129.525 196.895 ;
        RECT 124.340 196.580 129.525 196.880 ;
        RECT 124.340 196.570 124.720 196.580 ;
        RECT 129.195 196.565 129.525 196.580 ;
        RECT 132.415 196.880 132.745 196.895 ;
        RECT 133.540 196.880 133.920 196.890 ;
        RECT 132.415 196.580 133.920 196.880 ;
        RECT 132.415 196.565 132.745 196.580 ;
        RECT 133.540 196.570 133.920 196.580 ;
        RECT 74.720 196.225 76.700 196.555 ;
        RECT 104.720 196.225 106.700 196.555 ;
        RECT 134.720 196.225 136.700 196.555 ;
        RECT 93.315 195.520 93.645 195.535 ;
        RECT 99.295 195.520 99.625 195.535 ;
        RECT 93.315 195.220 99.625 195.520 ;
        RECT 93.315 195.205 93.645 195.220 ;
        RECT 99.295 195.205 99.625 195.220 ;
        RECT 103.435 195.520 103.765 195.535 ;
        RECT 114.475 195.520 114.805 195.535 ;
        RECT 137.475 195.520 137.805 195.535 ;
        RECT 103.435 195.220 137.805 195.520 ;
        RECT 103.435 195.205 103.765 195.220 ;
        RECT 114.475 195.205 114.805 195.220 ;
        RECT 137.475 195.205 137.805 195.220 ;
        RECT 81.355 194.840 81.685 194.855 ;
        RECT 92.395 194.840 92.725 194.855 ;
        RECT 81.355 194.540 92.725 194.840 ;
        RECT 81.355 194.525 81.685 194.540 ;
        RECT 92.395 194.525 92.725 194.540 ;
        RECT 99.755 194.840 100.085 194.855 ;
        RECT 106.655 194.840 106.985 194.855 ;
        RECT 109.875 194.840 110.205 194.855 ;
        RECT 99.755 194.540 110.205 194.840 ;
        RECT 99.755 194.525 100.085 194.540 ;
        RECT 106.655 194.525 106.985 194.540 ;
        RECT 109.875 194.525 110.205 194.540 ;
        RECT 131.035 194.840 131.365 194.855 ;
        RECT 134.715 194.840 135.045 194.855 ;
        RECT 131.035 194.540 135.045 194.840 ;
        RECT 131.035 194.525 131.365 194.540 ;
        RECT 134.715 194.525 135.045 194.540 ;
        RECT 89.720 193.505 91.700 193.835 ;
        RECT 119.720 193.505 121.700 193.835 ;
        RECT 149.720 193.505 151.700 193.835 ;
        RECT 88.255 192.800 88.585 192.815 ;
        RECT 90.555 192.800 90.885 192.815 ;
        RECT 120.455 192.800 120.785 192.815 ;
        RECT 88.255 192.500 90.885 192.800 ;
        RECT 88.255 192.485 88.585 192.500 ;
        RECT 90.555 192.485 90.885 192.500 ;
        RECT 103.220 192.500 120.785 192.800 ;
        RECT 81.355 192.120 81.685 192.135 ;
        RECT 103.220 192.120 103.520 192.500 ;
        RECT 120.455 192.485 120.785 192.500 ;
        RECT 127.815 192.800 128.145 192.815 ;
        RECT 152.655 192.800 152.985 192.815 ;
        RECT 127.815 192.500 152.985 192.800 ;
        RECT 127.815 192.485 128.145 192.500 ;
        RECT 152.655 192.485 152.985 192.500 ;
        RECT 81.355 191.820 103.520 192.120 ;
        RECT 104.355 192.120 104.685 192.135 ;
        RECT 120.915 192.120 121.245 192.135 ;
        RECT 104.355 191.820 121.245 192.120 ;
        RECT 81.355 191.805 81.685 191.820 ;
        RECT 104.355 191.805 104.685 191.820 ;
        RECT 120.915 191.805 121.245 191.820 ;
        RECT 128.735 192.120 129.065 192.135 ;
        RECT 146.675 192.120 147.005 192.135 ;
        RECT 128.735 191.820 147.005 192.120 ;
        RECT 128.735 191.805 129.065 191.820 ;
        RECT 146.675 191.805 147.005 191.820 ;
        RECT 109.875 191.440 110.205 191.455 ;
        RECT 111.255 191.440 111.585 191.455 ;
        RECT 109.875 191.140 111.585 191.440 ;
        RECT 109.875 191.125 110.205 191.140 ;
        RECT 111.255 191.125 111.585 191.140 ;
        RECT 74.720 190.785 76.700 191.115 ;
        RECT 104.720 190.785 106.700 191.115 ;
        RECT 134.720 190.785 136.700 191.115 ;
        RECT 91.015 190.760 91.345 190.775 ;
        RECT 107.115 190.760 107.445 190.775 ;
        RECT 128.275 190.760 128.605 190.775 ;
        RECT 91.015 190.460 99.840 190.760 ;
        RECT 91.015 190.445 91.345 190.460 ;
        RECT 85.495 190.080 85.825 190.095 ;
        RECT 89.635 190.080 89.965 190.095 ;
        RECT 98.835 190.080 99.165 190.095 ;
        RECT 85.495 189.780 99.165 190.080 ;
        RECT 99.540 190.080 99.840 190.460 ;
        RECT 107.115 190.460 128.605 190.760 ;
        RECT 107.115 190.445 107.445 190.460 ;
        RECT 128.275 190.445 128.605 190.460 ;
        RECT 105.275 190.080 105.605 190.095 ;
        RECT 99.540 189.780 105.605 190.080 ;
        RECT 85.495 189.765 85.825 189.780 ;
        RECT 89.635 189.765 89.965 189.780 ;
        RECT 98.835 189.765 99.165 189.780 ;
        RECT 105.275 189.765 105.605 189.780 ;
        RECT 106.195 190.080 106.525 190.095 ;
        RECT 123.675 190.080 124.005 190.095 ;
        RECT 106.195 189.780 124.005 190.080 ;
        RECT 106.195 189.765 106.525 189.780 ;
        RECT 123.675 189.765 124.005 189.780 ;
        RECT 94.235 189.400 94.565 189.415 ;
        RECT 130.575 189.400 130.905 189.415 ;
        RECT 94.235 189.100 130.905 189.400 ;
        RECT 94.235 189.085 94.565 189.100 ;
        RECT 130.575 189.085 130.905 189.100 ;
        RECT 97.915 188.720 98.245 188.735 ;
        RECT 116.315 188.720 116.645 188.735 ;
        RECT 97.915 188.420 116.645 188.720 ;
        RECT 97.915 188.405 98.245 188.420 ;
        RECT 116.315 188.405 116.645 188.420 ;
        RECT 131.035 188.720 131.365 188.735 ;
        RECT 137.935 188.720 138.265 188.735 ;
        RECT 148.515 188.720 148.845 188.735 ;
        RECT 131.035 188.420 148.845 188.720 ;
        RECT 131.035 188.405 131.365 188.420 ;
        RECT 137.935 188.405 138.265 188.420 ;
        RECT 148.515 188.405 148.845 188.420 ;
        RECT 89.720 188.065 91.700 188.395 ;
        RECT 119.720 188.065 121.700 188.395 ;
        RECT 149.720 188.065 151.700 188.395 ;
        RECT 99.755 188.040 100.085 188.055 ;
        RECT 115.855 188.040 116.185 188.055 ;
        RECT 99.755 187.740 116.185 188.040 ;
        RECT 99.755 187.725 100.085 187.740 ;
        RECT 115.855 187.725 116.185 187.740 ;
        RECT 88.255 187.360 88.585 187.375 ;
        RECT 98.375 187.360 98.705 187.375 ;
        RECT 111.255 187.360 111.585 187.375 ;
        RECT 88.255 187.060 111.585 187.360 ;
        RECT 88.255 187.045 88.585 187.060 ;
        RECT 98.375 187.045 98.705 187.060 ;
        RECT 111.255 187.045 111.585 187.060 ;
        RECT 118.155 187.360 118.485 187.375 ;
        RECT 127.355 187.360 127.685 187.375 ;
        RECT 118.155 187.060 127.685 187.360 ;
        RECT 118.155 187.045 118.485 187.060 ;
        RECT 127.355 187.045 127.685 187.060 ;
        RECT 102.515 186.680 102.845 186.695 ;
        RECT 119.535 186.680 119.865 186.695 ;
        RECT 102.515 186.380 119.865 186.680 ;
        RECT 102.515 186.365 102.845 186.380 ;
        RECT 119.535 186.365 119.865 186.380 ;
        RECT 111.255 186.000 111.585 186.015 ;
        RECT 113.555 186.000 113.885 186.015 ;
        RECT 111.255 185.700 113.885 186.000 ;
        RECT 111.255 185.685 111.585 185.700 ;
        RECT 113.555 185.685 113.885 185.700 ;
        RECT 74.720 185.345 76.700 185.675 ;
        RECT 104.720 185.345 106.700 185.675 ;
        RECT 134.720 185.345 136.700 185.675 ;
        RECT 82.275 184.640 82.605 184.655 ;
        RECT 130.575 184.640 130.905 184.655 ;
        RECT 82.275 184.340 130.905 184.640 ;
        RECT 82.275 184.325 82.605 184.340 ;
        RECT 130.575 184.325 130.905 184.340 ;
        RECT 81.355 183.960 81.685 183.975 ;
        RECT 99.755 183.960 100.085 183.975 ;
        RECT 111.255 183.960 111.585 183.975 ;
        RECT 81.355 183.660 111.585 183.960 ;
        RECT 81.355 183.645 81.685 183.660 ;
        RECT 99.755 183.645 100.085 183.660 ;
        RECT 111.255 183.645 111.585 183.660 ;
        RECT 122.755 183.960 123.085 183.975 ;
        RECT 138.140 183.960 138.520 183.970 ;
        RECT 122.755 183.660 138.520 183.960 ;
        RECT 122.755 183.645 123.085 183.660 ;
        RECT 138.140 183.650 138.520 183.660 ;
        RECT 107.575 183.280 107.905 183.295 ;
        RECT 112.380 183.280 112.760 183.290 ;
        RECT 107.575 182.980 112.760 183.280 ;
        RECT 107.575 182.965 107.905 182.980 ;
        RECT 112.380 182.970 112.760 182.980 ;
        RECT 89.720 182.625 91.700 182.955 ;
        RECT 119.720 182.625 121.700 182.955 ;
        RECT 149.720 182.625 151.700 182.955 ;
        RECT 99.295 182.600 99.625 182.615 ;
        RECT 107.575 182.600 107.905 182.615 ;
        RECT 99.295 182.300 107.905 182.600 ;
        RECT 99.295 182.285 99.625 182.300 ;
        RECT 107.575 182.285 107.905 182.300 ;
        RECT 109.415 180.560 109.745 180.575 ;
        RECT 114.475 180.560 114.805 180.575 ;
        RECT 109.415 180.260 114.805 180.560 ;
        RECT 109.415 180.245 109.745 180.260 ;
        RECT 114.475 180.245 114.805 180.260 ;
        RECT 74.720 179.905 76.700 180.235 ;
        RECT 104.720 179.905 106.700 180.235 ;
        RECT 134.720 179.905 136.700 180.235 ;
        RECT 102.515 179.200 102.845 179.215 ;
        RECT 104.355 179.200 104.685 179.215 ;
        RECT 102.515 178.900 104.685 179.200 ;
        RECT 102.515 178.885 102.845 178.900 ;
        RECT 104.355 178.885 104.685 178.900 ;
        RECT 106.195 179.200 106.525 179.215 ;
        RECT 114.935 179.200 115.265 179.215 ;
        RECT 106.195 178.900 115.265 179.200 ;
        RECT 106.195 178.885 106.525 178.900 ;
        RECT 114.935 178.885 115.265 178.900 ;
        RECT 131.035 179.200 131.365 179.215 ;
        RECT 131.700 179.200 132.080 179.210 ;
        RECT 131.035 178.900 132.080 179.200 ;
        RECT 131.035 178.885 131.365 178.900 ;
        RECT 131.700 178.890 132.080 178.900 ;
        RECT 139.775 178.520 140.105 178.535 ;
        RECT 110.580 178.220 140.105 178.520 ;
        RECT 98.375 177.840 98.705 177.855 ;
        RECT 110.580 177.840 110.880 178.220 ;
        RECT 139.775 178.205 140.105 178.220 ;
        RECT 98.375 177.540 110.880 177.840 ;
        RECT 98.375 177.525 98.705 177.540 ;
        RECT 89.720 177.185 91.700 177.515 ;
        RECT 119.720 177.185 121.700 177.515 ;
        RECT 149.720 177.185 151.700 177.515 ;
        RECT 96.995 176.480 97.325 176.495 ;
        RECT 108.035 176.480 108.365 176.495 ;
        RECT 96.995 176.180 108.365 176.480 ;
        RECT 96.995 176.165 97.325 176.180 ;
        RECT 108.035 176.165 108.365 176.180 ;
        RECT 116.775 176.480 117.105 176.495 ;
        RECT 139.315 176.480 139.645 176.495 ;
        RECT 116.775 176.180 139.645 176.480 ;
        RECT 116.775 176.165 117.105 176.180 ;
        RECT 139.315 176.165 139.645 176.180 ;
        RECT 93.315 175.800 93.645 175.815 ;
        RECT 101.595 175.800 101.925 175.815 ;
        RECT 129.195 175.810 129.525 175.815 ;
        RECT 128.940 175.800 129.525 175.810 ;
        RECT 93.315 175.500 108.810 175.800 ;
        RECT 128.740 175.500 129.525 175.800 ;
        RECT 93.315 175.485 93.645 175.500 ;
        RECT 101.595 175.485 101.925 175.500 ;
        RECT 108.510 175.135 108.810 175.500 ;
        RECT 128.940 175.490 129.525 175.500 ;
        RECT 129.195 175.485 129.525 175.490 ;
        RECT 136.095 175.800 136.425 175.815 ;
        RECT 150.815 175.800 151.145 175.815 ;
        RECT 136.095 175.500 151.145 175.800 ;
        RECT 136.095 175.485 136.425 175.500 ;
        RECT 150.815 175.485 151.145 175.500 ;
        RECT 87.335 175.120 87.665 175.135 ;
        RECT 95.615 175.120 95.945 175.135 ;
        RECT 87.335 174.820 95.945 175.120 ;
        RECT 87.335 174.805 87.665 174.820 ;
        RECT 95.615 174.805 95.945 174.820 ;
        RECT 108.495 174.805 108.825 175.135 ;
        RECT 112.380 175.120 112.760 175.130 ;
        RECT 113.095 175.120 113.425 175.135 ;
        RECT 112.380 174.820 113.425 175.120 ;
        RECT 112.380 174.810 112.760 174.820 ;
        RECT 113.095 174.805 113.425 174.820 ;
        RECT 74.720 174.465 76.700 174.795 ;
        RECT 104.720 174.465 106.700 174.795 ;
        RECT 134.720 174.465 136.700 174.795 ;
        RECT 88.255 174.440 88.585 174.455 ;
        RECT 102.975 174.440 103.305 174.455 ;
        RECT 88.255 174.140 103.305 174.440 ;
        RECT 88.255 174.125 88.585 174.140 ;
        RECT 102.975 174.125 103.305 174.140 ;
        RECT 94.235 173.760 94.565 173.775 ;
        RECT 99.755 173.760 100.085 173.775 ;
        RECT 134.715 173.760 135.045 173.775 ;
        RECT 94.235 173.460 97.310 173.760 ;
        RECT 94.235 173.445 94.565 173.460 ;
        RECT 91.015 173.080 91.345 173.095 ;
        RECT 97.010 173.080 97.310 173.460 ;
        RECT 99.755 173.460 135.045 173.760 ;
        RECT 99.755 173.445 100.085 173.460 ;
        RECT 134.715 173.445 135.045 173.460 ;
        RECT 129.655 173.080 129.985 173.095 ;
        RECT 91.015 172.780 92.480 173.080 ;
        RECT 97.010 172.780 129.985 173.080 ;
        RECT 91.015 172.765 91.345 172.780 ;
        RECT 89.720 171.745 91.700 172.075 ;
        RECT 89.635 171.040 89.965 171.055 ;
        RECT 92.180 171.040 92.480 172.780 ;
        RECT 129.655 172.765 129.985 172.780 ;
        RECT 98.835 172.400 99.165 172.415 ;
        RECT 110.335 172.400 110.665 172.415 ;
        RECT 98.835 172.100 110.665 172.400 ;
        RECT 98.835 172.085 99.165 172.100 ;
        RECT 110.335 172.085 110.665 172.100 ;
        RECT 116.315 172.085 116.645 172.415 ;
        RECT 116.330 171.055 116.630 172.085 ;
        RECT 119.720 171.745 121.700 172.075 ;
        RECT 149.720 171.745 151.700 172.075 ;
        RECT 89.635 170.740 92.480 171.040 ;
        RECT 89.635 170.725 89.965 170.740 ;
        RECT 116.315 170.725 116.645 171.055 ;
        RECT 86.875 170.360 87.205 170.375 ;
        RECT 91.015 170.360 91.345 170.375 ;
        RECT 86.875 170.060 91.345 170.360 ;
        RECT 86.875 170.045 87.205 170.060 ;
        RECT 91.015 170.045 91.345 170.060 ;
        RECT 102.055 170.360 102.385 170.375 ;
        RECT 106.195 170.360 106.525 170.375 ;
        RECT 102.055 170.060 106.525 170.360 ;
        RECT 102.055 170.045 102.385 170.060 ;
        RECT 106.195 170.045 106.525 170.060 ;
        RECT 86.415 169.680 86.745 169.695 ;
        RECT 90.555 169.680 90.885 169.695 ;
        RECT 86.415 169.380 90.885 169.680 ;
        RECT 86.415 169.365 86.745 169.380 ;
        RECT 90.555 169.365 90.885 169.380 ;
        RECT 74.720 169.025 76.700 169.355 ;
        RECT 104.720 169.025 106.700 169.355 ;
        RECT 134.720 169.025 136.700 169.355 ;
        RECT 85.495 168.320 85.825 168.335 ;
        RECT 108.495 168.320 108.825 168.335 ;
        RECT 85.495 168.020 108.825 168.320 ;
        RECT 85.495 168.005 85.825 168.020 ;
        RECT 108.495 168.005 108.825 168.020 ;
        RECT 119.075 168.320 119.405 168.335 ;
        RECT 131.955 168.320 132.285 168.335 ;
        RECT 148.975 168.320 149.305 168.335 ;
        RECT 119.075 168.020 149.305 168.320 ;
        RECT 119.075 168.005 119.405 168.020 ;
        RECT 131.955 168.005 132.285 168.020 ;
        RECT 148.975 168.005 149.305 168.020 ;
        RECT 89.720 166.305 91.700 166.635 ;
        RECT 119.720 166.305 121.700 166.635 ;
        RECT 149.720 166.305 151.700 166.635 ;
        RECT 80.895 165.600 81.225 165.615 ;
        RECT 112.635 165.600 112.965 165.615 ;
        RECT 80.895 165.300 112.965 165.600 ;
        RECT 80.895 165.285 81.225 165.300 ;
        RECT 112.635 165.285 112.965 165.300 ;
        RECT 116.775 165.600 117.105 165.615 ;
        RECT 119.075 165.600 119.405 165.615 ;
        RECT 116.775 165.300 119.405 165.600 ;
        RECT 116.775 165.285 117.105 165.300 ;
        RECT 119.075 165.285 119.405 165.300 ;
        RECT 130.115 165.600 130.445 165.615 ;
        RECT 146.675 165.600 147.005 165.615 ;
        RECT 130.115 165.300 147.005 165.600 ;
        RECT 130.115 165.285 130.445 165.300 ;
        RECT 146.675 165.285 147.005 165.300 ;
        RECT 77.215 164.920 77.545 164.935 ;
        RECT 100.215 164.920 100.545 164.935 ;
        RECT 77.215 164.620 100.545 164.920 ;
        RECT 77.215 164.605 77.545 164.620 ;
        RECT 100.215 164.605 100.545 164.620 ;
        RECT 121.835 164.920 122.165 164.935 ;
        RECT 133.795 164.920 134.125 164.935 ;
        RECT 121.835 164.620 134.125 164.920 ;
        RECT 121.835 164.605 122.165 164.620 ;
        RECT 133.795 164.605 134.125 164.620 ;
        RECT 74.720 163.585 76.700 163.915 ;
        RECT 104.720 163.585 106.700 163.915 ;
        RECT 134.720 163.585 136.700 163.915 ;
        RECT 101.595 162.880 101.925 162.895 ;
        RECT 104.815 162.880 105.145 162.895 ;
        RECT 101.595 162.580 105.145 162.880 ;
        RECT 101.595 162.565 101.925 162.580 ;
        RECT 104.815 162.565 105.145 162.580 ;
        RECT 110.335 162.880 110.665 162.895 ;
        RECT 142.075 162.880 142.405 162.895 ;
        RECT 146.675 162.880 147.005 162.895 ;
        RECT 110.335 162.580 147.005 162.880 ;
        RECT 110.335 162.565 110.665 162.580 ;
        RECT 142.075 162.565 142.405 162.580 ;
        RECT 146.675 162.565 147.005 162.580 ;
        RECT 97.455 162.200 97.785 162.215 ;
        RECT 105.275 162.200 105.605 162.215 ;
        RECT 97.455 161.900 105.605 162.200 ;
        RECT 97.455 161.885 97.785 161.900 ;
        RECT 105.275 161.885 105.605 161.900 ;
        RECT 119.075 162.200 119.405 162.215 ;
        RECT 131.035 162.200 131.365 162.215 ;
        RECT 119.075 161.900 131.365 162.200 ;
        RECT 119.075 161.885 119.405 161.900 ;
        RECT 131.035 161.885 131.365 161.900 ;
        RECT 89.720 160.865 91.700 161.195 ;
        RECT 119.720 160.865 121.700 161.195 ;
        RECT 149.720 160.865 151.700 161.195 ;
        RECT 78.595 159.480 78.925 159.495 ;
        RECT 110.335 159.480 110.665 159.495 ;
        RECT 78.595 159.180 110.665 159.480 ;
        RECT 78.595 159.165 78.925 159.180 ;
        RECT 110.335 159.165 110.665 159.180 ;
        RECT 74.720 158.145 76.700 158.475 ;
        RECT 104.720 158.145 106.700 158.475 ;
        RECT 134.720 158.145 136.700 158.475 ;
        RECT 97.660 157.440 98.040 157.450 ;
        RECT 115.855 157.440 116.185 157.455 ;
        RECT 97.660 157.140 116.185 157.440 ;
        RECT 97.660 157.130 98.040 157.140 ;
        RECT 115.855 157.125 116.185 157.140 ;
        RECT 116.775 157.440 117.105 157.455 ;
        RECT 128.735 157.440 129.065 157.455 ;
        RECT 116.775 157.140 129.065 157.440 ;
        RECT 116.775 157.125 117.105 157.140 ;
        RECT 128.735 157.125 129.065 157.140 ;
        RECT 138.140 157.440 138.520 157.450 ;
        RECT 139.775 157.440 140.105 157.455 ;
        RECT 138.140 157.140 140.105 157.440 ;
        RECT 138.140 157.130 138.520 157.140 ;
        RECT 139.775 157.125 140.105 157.140 ;
        RECT 82.275 156.760 82.605 156.775 ;
        RECT 105.275 156.760 105.605 156.775 ;
        RECT 82.275 156.460 105.605 156.760 ;
        RECT 82.275 156.445 82.605 156.460 ;
        RECT 105.275 156.445 105.605 156.460 ;
        RECT 113.555 156.760 113.885 156.775 ;
        RECT 126.895 156.760 127.225 156.775 ;
        RECT 113.555 156.460 127.225 156.760 ;
        RECT 113.555 156.445 113.885 156.460 ;
        RECT 126.895 156.445 127.225 156.460 ;
        RECT 137.220 156.080 137.600 156.090 ;
        RECT 138.855 156.080 139.185 156.095 ;
        RECT 137.220 155.780 139.185 156.080 ;
        RECT 137.220 155.770 137.600 155.780 ;
        RECT 138.855 155.765 139.185 155.780 ;
        RECT 89.720 155.425 91.700 155.755 ;
        RECT 119.720 155.425 121.700 155.755 ;
        RECT 149.720 155.425 151.700 155.755 ;
        RECT 141.820 155.400 142.200 155.410 ;
        RECT 142.535 155.400 142.865 155.415 ;
        RECT 141.820 155.100 142.865 155.400 ;
        RECT 141.820 155.090 142.200 155.100 ;
        RECT 142.535 155.085 142.865 155.100 ;
        RECT 106.655 154.040 106.985 154.055 ;
        RECT 119.995 154.040 120.325 154.055 ;
        RECT 106.655 153.740 120.325 154.040 ;
        RECT 106.655 153.725 106.985 153.740 ;
        RECT 119.995 153.725 120.325 153.740 ;
        RECT 116.980 153.360 117.360 153.370 ;
        RECT 117.695 153.360 118.025 153.375 ;
        RECT 116.980 153.060 118.025 153.360 ;
        RECT 116.980 153.050 117.360 153.060 ;
        RECT 117.695 153.045 118.025 153.060 ;
        RECT 74.720 152.705 76.700 153.035 ;
        RECT 104.720 152.705 106.700 153.035 ;
        RECT 134.720 152.705 136.700 153.035 ;
        RECT 112.635 152.365 112.965 152.695 ;
        RECT 112.650 152.000 112.950 152.365 ;
        RECT 113.555 152.000 113.885 152.015 ;
        RECT 112.650 151.700 113.885 152.000 ;
        RECT 113.555 151.685 113.885 151.700 ;
        RECT 131.955 152.000 132.285 152.015 ;
        RECT 142.075 152.000 142.405 152.015 ;
        RECT 131.955 151.700 142.405 152.000 ;
        RECT 131.955 151.685 132.285 151.700 ;
        RECT 142.075 151.685 142.405 151.700 ;
        RECT 109.875 151.320 110.205 151.335 ;
        RECT 113.095 151.320 113.425 151.335 ;
        RECT 109.875 151.020 113.425 151.320 ;
        RECT 109.875 151.005 110.205 151.020 ;
        RECT 113.095 151.005 113.425 151.020 ;
        RECT 136.095 151.320 136.425 151.335 ;
        RECT 137.220 151.320 137.600 151.330 ;
        RECT 136.095 151.020 137.600 151.320 ;
        RECT 136.095 151.005 136.425 151.020 ;
        RECT 137.220 151.010 137.600 151.020 ;
        RECT 125.055 150.640 125.385 150.655 ;
        RECT 138.855 150.640 139.185 150.655 ;
        RECT 125.055 150.340 139.185 150.640 ;
        RECT 125.055 150.325 125.385 150.340 ;
        RECT 138.855 150.325 139.185 150.340 ;
        RECT 89.720 149.985 91.700 150.315 ;
        RECT 119.720 149.985 121.700 150.315 ;
        RECT 149.720 149.985 151.700 150.315 ;
        RECT 131.700 149.960 132.080 149.970 ;
        RECT 132.875 149.960 133.205 149.975 ;
        RECT 131.700 149.660 133.205 149.960 ;
        RECT 131.700 149.650 132.080 149.660 ;
        RECT 132.875 149.645 133.205 149.660 ;
        RECT 128.735 149.280 129.065 149.295 ;
        RECT 131.035 149.280 131.365 149.295 ;
        RECT 128.735 148.980 131.365 149.280 ;
        RECT 128.735 148.965 129.065 148.980 ;
        RECT 131.035 148.965 131.365 148.980 ;
        RECT 135.635 149.280 135.965 149.295 ;
        RECT 152.195 149.280 152.525 149.295 ;
        RECT 135.635 148.980 152.525 149.280 ;
        RECT 135.635 148.965 135.965 148.980 ;
        RECT 152.195 148.965 152.525 148.980 ;
        RECT 131.955 148.600 132.285 148.615 ;
        RECT 138.395 148.600 138.725 148.615 ;
        RECT 131.955 148.300 138.725 148.600 ;
        RECT 131.955 148.285 132.285 148.300 ;
        RECT 138.395 148.285 138.725 148.300 ;
        RECT 109.875 147.920 110.205 147.935 ;
        RECT 112.635 147.920 112.965 147.935 ;
        RECT 109.875 147.620 112.965 147.920 ;
        RECT 109.875 147.605 110.205 147.620 ;
        RECT 112.635 147.605 112.965 147.620 ;
        RECT 127.815 147.920 128.145 147.935 ;
        RECT 131.955 147.920 132.285 147.935 ;
        RECT 127.815 147.620 132.285 147.920 ;
        RECT 127.815 147.605 128.145 147.620 ;
        RECT 131.955 147.605 132.285 147.620 ;
        RECT 74.720 147.265 76.700 147.595 ;
        RECT 104.720 147.265 106.700 147.595 ;
        RECT 134.720 147.265 136.700 147.595 ;
        RECT 110.795 147.240 111.125 147.255 ;
        RECT 132.415 147.240 132.745 147.255 ;
        RECT 110.795 146.940 132.745 147.240 ;
        RECT 110.795 146.925 111.125 146.940 ;
        RECT 132.415 146.925 132.745 146.940 ;
        RECT 111.255 146.560 111.585 146.575 ;
        RECT 110.580 146.260 111.585 146.560 ;
        RECT 110.580 145.895 110.880 146.260 ;
        RECT 111.255 146.245 111.585 146.260 ;
        RECT 117.235 146.560 117.565 146.575 ;
        RECT 117.900 146.560 118.280 146.570 ;
        RECT 117.235 146.260 118.280 146.560 ;
        RECT 117.235 146.245 117.565 146.260 ;
        RECT 117.900 146.250 118.280 146.260 ;
        RECT 92.855 145.880 93.185 145.895 ;
        RECT 105.735 145.880 106.065 145.895 ;
        RECT 107.575 145.880 107.905 145.895 ;
        RECT 92.855 145.580 106.065 145.880 ;
        RECT 92.855 145.565 93.185 145.580 ;
        RECT 105.735 145.565 106.065 145.580 ;
        RECT 106.900 145.580 107.905 145.880 ;
        RECT 80.895 145.200 81.225 145.215 ;
        RECT 88.715 145.200 89.045 145.215 ;
        RECT 80.895 144.900 89.045 145.200 ;
        RECT 80.895 144.885 81.225 144.900 ;
        RECT 88.715 144.885 89.045 144.900 ;
        RECT 89.720 144.545 91.700 144.875 ;
        RECT 106.900 144.520 107.200 145.580 ;
        RECT 107.575 145.565 107.905 145.580 ;
        RECT 110.335 145.580 110.880 145.895 ;
        RECT 116.315 145.880 116.645 145.895 ;
        RECT 134.715 145.880 135.045 145.895 ;
        RECT 116.315 145.580 135.045 145.880 ;
        RECT 110.335 145.565 110.665 145.580 ;
        RECT 116.315 145.565 116.645 145.580 ;
        RECT 134.715 145.565 135.045 145.580 ;
        RECT 107.780 145.200 108.160 145.210 ;
        RECT 108.955 145.200 109.285 145.215 ;
        RECT 107.780 144.900 109.285 145.200 ;
        RECT 107.780 144.890 108.160 144.900 ;
        RECT 108.955 144.885 109.285 144.900 ;
        RECT 119.720 144.545 121.700 144.875 ;
        RECT 149.720 144.545 151.700 144.875 ;
        RECT 107.575 144.520 107.905 144.535 ;
        RECT 106.900 144.220 107.905 144.520 ;
        RECT 107.575 144.205 107.905 144.220 ;
        RECT 102.975 143.840 103.305 143.855 ;
        RECT 110.335 143.840 110.665 143.855 ;
        RECT 102.975 143.540 110.665 143.840 ;
        RECT 102.975 143.525 103.305 143.540 ;
        RECT 110.335 143.525 110.665 143.540 ;
        RECT 92.395 143.160 92.725 143.175 ;
        RECT 96.995 143.160 97.325 143.175 ;
        RECT 110.335 143.160 110.665 143.175 ;
        RECT 92.395 142.860 110.665 143.160 ;
        RECT 92.395 142.845 92.725 142.860 ;
        RECT 96.995 142.845 97.325 142.860 ;
        RECT 110.335 142.845 110.665 142.860 ;
        RECT 74.720 141.825 76.700 142.155 ;
        RECT 104.720 141.825 106.700 142.155 ;
        RECT 134.720 141.825 136.700 142.155 ;
        RECT 100.675 141.120 101.005 141.135 ;
        RECT 113.095 141.120 113.425 141.135 ;
        RECT 100.675 140.820 113.425 141.120 ;
        RECT 100.675 140.805 101.005 140.820 ;
        RECT 113.095 140.805 113.425 140.820 ;
        RECT 92.395 140.440 92.725 140.455 ;
        RECT 106.655 140.440 106.985 140.455 ;
        RECT 143.915 140.450 144.245 140.455 ;
        RECT 92.395 140.140 106.985 140.440 ;
        RECT 92.395 140.125 92.725 140.140 ;
        RECT 106.655 140.125 106.985 140.140 ;
        RECT 143.660 140.440 144.245 140.450 ;
        RECT 143.660 140.140 144.470 140.440 ;
        RECT 143.660 140.130 144.245 140.140 ;
        RECT 143.915 140.125 144.245 140.130 ;
        RECT 96.075 139.760 96.405 139.775 ;
        RECT 113.555 139.760 113.885 139.775 ;
        RECT 96.075 139.460 113.885 139.760 ;
        RECT 96.075 139.445 96.405 139.460 ;
        RECT 113.555 139.445 113.885 139.460 ;
        RECT 128.940 139.760 129.320 139.770 ;
        RECT 145.755 139.760 146.085 139.775 ;
        RECT 128.940 139.460 146.085 139.760 ;
        RECT 128.940 139.450 129.320 139.460 ;
        RECT 145.755 139.445 146.085 139.460 ;
        RECT 89.720 139.105 91.700 139.435 ;
        RECT 119.720 139.105 121.700 139.435 ;
        RECT 149.720 139.105 151.700 139.435 ;
        RECT 129.195 138.400 129.525 138.415 ;
        RECT 140.695 138.400 141.025 138.415 ;
        RECT 129.195 138.100 141.025 138.400 ;
        RECT 129.195 138.085 129.525 138.100 ;
        RECT 140.695 138.085 141.025 138.100 ;
        RECT 90.095 137.040 90.425 137.055 ;
        RECT 116.775 137.050 117.105 137.055 ;
        RECT 97.660 137.040 98.040 137.050 ;
        RECT 90.095 136.740 98.040 137.040 ;
        RECT 90.095 136.725 90.425 136.740 ;
        RECT 97.660 136.730 98.040 136.740 ;
        RECT 116.775 137.040 117.360 137.050 ;
        RECT 116.775 136.740 117.560 137.040 ;
        RECT 116.775 136.730 117.360 136.740 ;
        RECT 116.775 136.725 117.105 136.730 ;
        RECT 74.720 136.385 76.700 136.715 ;
        RECT 104.720 136.385 106.700 136.715 ;
        RECT 134.720 136.385 136.700 136.715 ;
        RECT 132.875 136.360 133.205 136.375 ;
        RECT 132.875 136.060 133.880 136.360 ;
        RECT 132.875 136.045 133.205 136.060 ;
        RECT 93.775 135.680 94.105 135.695 ;
        RECT 107.115 135.680 107.445 135.695 ;
        RECT 93.775 135.380 107.445 135.680 ;
        RECT 133.580 135.680 133.880 136.060 ;
        RECT 137.015 135.680 137.345 135.695 ;
        RECT 138.855 135.680 139.185 135.695 ;
        RECT 133.580 135.380 139.185 135.680 ;
        RECT 93.775 135.365 94.105 135.380 ;
        RECT 107.115 135.365 107.445 135.380 ;
        RECT 137.015 135.365 137.345 135.380 ;
        RECT 138.855 135.365 139.185 135.380 ;
        RECT 106.195 135.000 106.525 135.015 ;
        RECT 107.780 135.000 108.160 135.010 ;
        RECT 106.195 134.700 108.160 135.000 ;
        RECT 106.195 134.685 106.525 134.700 ;
        RECT 107.780 134.690 108.160 134.700 ;
        RECT 129.655 135.000 129.985 135.015 ;
        RECT 144.375 135.000 144.705 135.015 ;
        RECT 129.655 134.700 144.705 135.000 ;
        RECT 129.655 134.685 129.985 134.700 ;
        RECT 144.375 134.685 144.705 134.700 ;
        RECT 89.720 133.665 91.700 133.995 ;
        RECT 119.720 133.665 121.700 133.995 ;
        RECT 149.720 133.665 151.700 133.995 ;
        RECT 96.995 133.640 97.325 133.655 ;
        RECT 100.420 133.640 100.800 133.650 ;
        RECT 96.995 133.340 100.800 133.640 ;
        RECT 96.995 133.325 97.325 133.340 ;
        RECT 100.420 133.330 100.800 133.340 ;
        RECT 140.695 133.640 141.025 133.655 ;
        RECT 141.820 133.640 142.200 133.650 ;
        RECT 140.695 133.340 142.200 133.640 ;
        RECT 140.695 133.325 141.025 133.340 ;
        RECT 141.820 133.330 142.200 133.340 ;
        RECT 74.455 132.960 74.785 132.975 ;
        RECT 85.495 132.960 85.825 132.975 ;
        RECT 113.095 132.960 113.425 132.975 ;
        RECT 74.455 132.660 81.900 132.960 ;
        RECT 74.455 132.645 74.785 132.660 ;
        RECT 81.600 132.280 81.900 132.660 ;
        RECT 85.495 132.660 113.425 132.960 ;
        RECT 85.495 132.645 85.825 132.660 ;
        RECT 113.095 132.645 113.425 132.660 ;
        RECT 98.375 132.290 98.705 132.295 ;
        RECT 98.375 132.280 98.960 132.290 ;
        RECT 113.555 132.280 113.885 132.295 ;
        RECT 114.220 132.280 114.600 132.290 ;
        RECT 130.575 132.280 130.905 132.295 ;
        RECT 81.600 131.980 99.160 132.280 ;
        RECT 113.555 131.980 130.905 132.280 ;
        RECT 98.375 131.970 98.960 131.980 ;
        RECT 98.375 131.965 98.705 131.970 ;
        RECT 113.555 131.965 113.885 131.980 ;
        RECT 114.220 131.970 114.600 131.980 ;
        RECT 130.575 131.965 130.905 131.980 ;
        RECT 137.475 131.600 137.805 131.615 ;
        RECT 148.055 131.600 148.385 131.615 ;
        RECT 137.475 131.300 148.385 131.600 ;
        RECT 137.475 131.285 137.805 131.300 ;
        RECT 148.055 131.285 148.385 131.300 ;
        RECT 74.720 130.945 76.700 131.275 ;
        RECT 104.720 130.945 106.700 131.275 ;
        RECT 134.720 130.945 136.700 131.275 ;
        RECT 122.295 130.920 122.625 130.935 ;
        RECT 133.335 130.920 133.665 130.935 ;
        RECT 122.295 130.605 122.840 130.920 ;
        RECT 122.540 130.240 122.840 130.605 ;
        RECT 132.660 130.620 133.665 130.920 ;
        RECT 124.595 130.240 124.925 130.255 ;
        RECT 109.660 129.940 124.925 130.240 ;
        RECT 76.755 129.560 77.085 129.575 ;
        RECT 92.855 129.560 93.185 129.575 ;
        RECT 76.755 129.260 93.185 129.560 ;
        RECT 76.755 129.245 77.085 129.260 ;
        RECT 92.855 129.245 93.185 129.260 ;
        RECT 89.720 128.225 91.700 128.555 ;
        RECT 99.755 128.200 100.085 128.215 ;
        RECT 108.035 128.200 108.365 128.215 ;
        RECT 109.660 128.200 109.960 129.940 ;
        RECT 124.595 129.925 124.925 129.940 ;
        RECT 131.955 130.240 132.285 130.255 ;
        RECT 132.660 130.240 132.960 130.620 ;
        RECT 133.335 130.605 133.665 130.620 ;
        RECT 144.375 130.920 144.705 130.935 ;
        RECT 146.215 130.920 146.545 130.935 ;
        RECT 144.375 130.620 146.545 130.920 ;
        RECT 144.375 130.605 144.705 130.620 ;
        RECT 146.215 130.605 146.545 130.620 ;
        RECT 131.955 129.940 132.960 130.240 ;
        RECT 133.540 130.240 133.920 130.250 ;
        RECT 134.715 130.240 135.045 130.255 ;
        RECT 133.540 129.940 135.045 130.240 ;
        RECT 131.955 129.925 132.285 129.940 ;
        RECT 133.540 129.930 133.920 129.940 ;
        RECT 134.715 129.925 135.045 129.940 ;
        RECT 110.795 129.560 111.125 129.575 ;
        RECT 111.460 129.560 111.840 129.570 ;
        RECT 129.655 129.560 129.985 129.575 ;
        RECT 110.795 129.260 129.985 129.560 ;
        RECT 110.795 129.245 111.125 129.260 ;
        RECT 111.460 129.250 111.840 129.260 ;
        RECT 129.655 129.245 129.985 129.260 ;
        RECT 142.535 129.560 142.865 129.575 ;
        RECT 145.295 129.560 145.625 129.575 ;
        RECT 148.975 129.560 149.305 129.575 ;
        RECT 142.535 129.260 149.305 129.560 ;
        RECT 142.535 129.245 142.865 129.260 ;
        RECT 145.295 129.245 145.625 129.260 ;
        RECT 148.975 129.245 149.305 129.260 ;
        RECT 116.775 128.880 117.105 128.895 ;
        RECT 117.900 128.880 118.280 128.890 ;
        RECT 116.775 128.580 118.280 128.880 ;
        RECT 116.775 128.565 117.105 128.580 ;
        RECT 117.900 128.570 118.280 128.580 ;
        RECT 137.015 128.880 137.345 128.895 ;
        RECT 146.675 128.880 147.005 128.895 ;
        RECT 137.015 128.580 147.005 128.880 ;
        RECT 137.015 128.565 137.345 128.580 ;
        RECT 146.675 128.565 147.005 128.580 ;
        RECT 119.720 128.225 121.700 128.555 ;
        RECT 149.720 128.225 151.700 128.555 ;
        RECT 99.755 127.900 109.960 128.200 ;
        RECT 116.315 128.200 116.645 128.215 ;
        RECT 116.980 128.200 117.360 128.210 ;
        RECT 116.315 127.900 117.360 128.200 ;
        RECT 99.755 127.885 100.085 127.900 ;
        RECT 108.035 127.885 108.365 127.900 ;
        RECT 116.315 127.885 116.645 127.900 ;
        RECT 116.980 127.890 117.360 127.900 ;
        RECT 137.475 128.200 137.805 128.215 ;
        RECT 143.660 128.200 144.040 128.210 ;
        RECT 137.475 127.900 144.040 128.200 ;
        RECT 137.475 127.885 137.805 127.900 ;
        RECT 143.660 127.890 144.040 127.900 ;
        RECT 88.255 127.520 88.585 127.535 ;
        RECT 91.935 127.520 92.265 127.535 ;
        RECT 146.215 127.520 146.545 127.535 ;
        RECT 88.255 127.220 146.545 127.520 ;
        RECT 88.255 127.205 88.585 127.220 ;
        RECT 91.935 127.205 92.265 127.220 ;
        RECT 146.215 127.205 146.545 127.220 ;
        RECT 117.900 126.840 118.280 126.850 ;
        RECT 121.375 126.840 121.705 126.855 ;
        RECT 117.900 126.540 121.705 126.840 ;
        RECT 117.900 126.530 118.280 126.540 ;
        RECT 121.375 126.525 121.705 126.540 ;
        RECT 123.215 126.840 123.545 126.855 ;
        RECT 143.455 126.850 143.785 126.855 ;
        RECT 124.340 126.840 124.720 126.850 ;
        RECT 143.455 126.840 144.040 126.850 ;
        RECT 123.215 126.540 124.720 126.840 ;
        RECT 143.230 126.540 144.040 126.840 ;
        RECT 123.215 126.525 123.545 126.540 ;
        RECT 124.340 126.530 124.720 126.540 ;
        RECT 143.455 126.530 144.040 126.540 ;
        RECT 143.455 126.525 143.785 126.530 ;
        RECT 116.315 126.160 116.645 126.175 ;
        RECT 116.980 126.160 117.360 126.170 ;
        RECT 116.315 125.860 117.360 126.160 ;
        RECT 116.315 125.845 116.645 125.860 ;
        RECT 116.980 125.850 117.360 125.860 ;
        RECT 137.935 126.160 138.265 126.175 ;
        RECT 143.915 126.160 144.245 126.175 ;
        RECT 137.935 125.860 144.245 126.160 ;
        RECT 137.935 125.845 138.265 125.860 ;
        RECT 143.915 125.845 144.245 125.860 ;
        RECT 74.720 125.505 76.700 125.835 ;
        RECT 104.720 125.505 106.700 125.835 ;
        RECT 134.720 125.505 136.700 125.835 ;
        RECT 89.720 122.785 91.700 123.115 ;
        RECT 119.720 122.785 121.700 123.115 ;
        RECT 149.720 122.785 151.700 123.115 ;
      LAYER via3 ;
        RECT 127.810 221.110 128.195 221.495 ;
        RECT 125.375 216.495 125.785 216.905 ;
        RECT 126.500 216.500 126.900 216.900 ;
        RECT 110.245 214.845 110.755 215.355 ;
        RECT 116.605 214.905 116.995 215.295 ;
        RECT 120.495 214.995 120.910 215.410 ;
        RECT 131.915 220.115 132.290 220.490 ;
        RECT 136.040 218.940 136.360 219.260 ;
        RECT 140.210 217.610 140.595 217.995 ;
        RECT 144.275 216.375 144.725 216.825 ;
        RECT 148.490 215.190 148.910 215.610 ;
        RECT 152.575 215.175 153.025 215.625 ;
        RECT 74.750 207.110 75.070 207.430 ;
        RECT 75.150 207.110 75.470 207.430 ;
        RECT 75.550 207.110 75.870 207.430 ;
        RECT 75.950 207.110 76.270 207.430 ;
        RECT 76.350 207.110 76.670 207.430 ;
        RECT 104.750 207.110 105.070 207.430 ;
        RECT 105.150 207.110 105.470 207.430 ;
        RECT 105.550 207.110 105.870 207.430 ;
        RECT 105.950 207.110 106.270 207.430 ;
        RECT 106.350 207.110 106.670 207.430 ;
        RECT 134.750 207.110 135.070 207.430 ;
        RECT 135.150 207.110 135.470 207.430 ;
        RECT 135.550 207.110 135.870 207.430 ;
        RECT 135.950 207.110 136.270 207.430 ;
        RECT 136.350 207.110 136.670 207.430 ;
        RECT 89.750 204.390 90.070 204.710 ;
        RECT 90.150 204.390 90.470 204.710 ;
        RECT 90.550 204.390 90.870 204.710 ;
        RECT 90.950 204.390 91.270 204.710 ;
        RECT 91.350 204.390 91.670 204.710 ;
        RECT 119.750 204.390 120.070 204.710 ;
        RECT 120.150 204.390 120.470 204.710 ;
        RECT 120.550 204.390 120.870 204.710 ;
        RECT 120.950 204.390 121.270 204.710 ;
        RECT 121.350 204.390 121.670 204.710 ;
        RECT 149.750 204.390 150.070 204.710 ;
        RECT 150.150 204.390 150.470 204.710 ;
        RECT 150.550 204.390 150.870 204.710 ;
        RECT 150.950 204.390 151.270 204.710 ;
        RECT 151.350 204.390 151.670 204.710 ;
        RECT 100.450 203.370 100.770 203.690 ;
        RECT 111.490 203.370 111.810 203.690 ;
        RECT 74.750 201.670 75.070 201.990 ;
        RECT 75.150 201.670 75.470 201.990 ;
        RECT 75.550 201.670 75.870 201.990 ;
        RECT 75.950 201.670 76.270 201.990 ;
        RECT 76.350 201.670 76.670 201.990 ;
        RECT 104.750 201.670 105.070 201.990 ;
        RECT 105.150 201.670 105.470 201.990 ;
        RECT 105.550 201.670 105.870 201.990 ;
        RECT 105.950 201.670 106.270 201.990 ;
        RECT 106.350 201.670 106.670 201.990 ;
        RECT 134.750 201.670 135.070 201.990 ;
        RECT 135.150 201.670 135.470 201.990 ;
        RECT 135.550 201.670 135.870 201.990 ;
        RECT 135.950 201.670 136.270 201.990 ;
        RECT 136.350 201.670 136.670 201.990 ;
        RECT 89.750 198.950 90.070 199.270 ;
        RECT 90.150 198.950 90.470 199.270 ;
        RECT 90.550 198.950 90.870 199.270 ;
        RECT 90.950 198.950 91.270 199.270 ;
        RECT 91.350 198.950 91.670 199.270 ;
        RECT 119.750 198.950 120.070 199.270 ;
        RECT 120.150 198.950 120.470 199.270 ;
        RECT 120.550 198.950 120.870 199.270 ;
        RECT 120.950 198.950 121.270 199.270 ;
        RECT 121.350 198.950 121.670 199.270 ;
        RECT 149.750 198.950 150.070 199.270 ;
        RECT 150.150 198.950 150.470 199.270 ;
        RECT 150.550 198.950 150.870 199.270 ;
        RECT 150.950 198.950 151.270 199.270 ;
        RECT 151.350 198.950 151.670 199.270 ;
        RECT 114.250 197.250 114.570 197.570 ;
        RECT 98.610 196.570 98.930 196.890 ;
        RECT 124.370 196.570 124.690 196.890 ;
        RECT 133.570 196.570 133.890 196.890 ;
        RECT 74.750 196.230 75.070 196.550 ;
        RECT 75.150 196.230 75.470 196.550 ;
        RECT 75.550 196.230 75.870 196.550 ;
        RECT 75.950 196.230 76.270 196.550 ;
        RECT 76.350 196.230 76.670 196.550 ;
        RECT 104.750 196.230 105.070 196.550 ;
        RECT 105.150 196.230 105.470 196.550 ;
        RECT 105.550 196.230 105.870 196.550 ;
        RECT 105.950 196.230 106.270 196.550 ;
        RECT 106.350 196.230 106.670 196.550 ;
        RECT 134.750 196.230 135.070 196.550 ;
        RECT 135.150 196.230 135.470 196.550 ;
        RECT 135.550 196.230 135.870 196.550 ;
        RECT 135.950 196.230 136.270 196.550 ;
        RECT 136.350 196.230 136.670 196.550 ;
        RECT 89.750 193.510 90.070 193.830 ;
        RECT 90.150 193.510 90.470 193.830 ;
        RECT 90.550 193.510 90.870 193.830 ;
        RECT 90.950 193.510 91.270 193.830 ;
        RECT 91.350 193.510 91.670 193.830 ;
        RECT 119.750 193.510 120.070 193.830 ;
        RECT 120.150 193.510 120.470 193.830 ;
        RECT 120.550 193.510 120.870 193.830 ;
        RECT 120.950 193.510 121.270 193.830 ;
        RECT 121.350 193.510 121.670 193.830 ;
        RECT 149.750 193.510 150.070 193.830 ;
        RECT 150.150 193.510 150.470 193.830 ;
        RECT 150.550 193.510 150.870 193.830 ;
        RECT 150.950 193.510 151.270 193.830 ;
        RECT 151.350 193.510 151.670 193.830 ;
        RECT 74.750 190.790 75.070 191.110 ;
        RECT 75.150 190.790 75.470 191.110 ;
        RECT 75.550 190.790 75.870 191.110 ;
        RECT 75.950 190.790 76.270 191.110 ;
        RECT 76.350 190.790 76.670 191.110 ;
        RECT 104.750 190.790 105.070 191.110 ;
        RECT 105.150 190.790 105.470 191.110 ;
        RECT 105.550 190.790 105.870 191.110 ;
        RECT 105.950 190.790 106.270 191.110 ;
        RECT 106.350 190.790 106.670 191.110 ;
        RECT 134.750 190.790 135.070 191.110 ;
        RECT 135.150 190.790 135.470 191.110 ;
        RECT 135.550 190.790 135.870 191.110 ;
        RECT 135.950 190.790 136.270 191.110 ;
        RECT 136.350 190.790 136.670 191.110 ;
        RECT 89.750 188.070 90.070 188.390 ;
        RECT 90.150 188.070 90.470 188.390 ;
        RECT 90.550 188.070 90.870 188.390 ;
        RECT 90.950 188.070 91.270 188.390 ;
        RECT 91.350 188.070 91.670 188.390 ;
        RECT 119.750 188.070 120.070 188.390 ;
        RECT 120.150 188.070 120.470 188.390 ;
        RECT 120.550 188.070 120.870 188.390 ;
        RECT 120.950 188.070 121.270 188.390 ;
        RECT 121.350 188.070 121.670 188.390 ;
        RECT 149.750 188.070 150.070 188.390 ;
        RECT 150.150 188.070 150.470 188.390 ;
        RECT 150.550 188.070 150.870 188.390 ;
        RECT 150.950 188.070 151.270 188.390 ;
        RECT 151.350 188.070 151.670 188.390 ;
        RECT 74.750 185.350 75.070 185.670 ;
        RECT 75.150 185.350 75.470 185.670 ;
        RECT 75.550 185.350 75.870 185.670 ;
        RECT 75.950 185.350 76.270 185.670 ;
        RECT 76.350 185.350 76.670 185.670 ;
        RECT 104.750 185.350 105.070 185.670 ;
        RECT 105.150 185.350 105.470 185.670 ;
        RECT 105.550 185.350 105.870 185.670 ;
        RECT 105.950 185.350 106.270 185.670 ;
        RECT 106.350 185.350 106.670 185.670 ;
        RECT 134.750 185.350 135.070 185.670 ;
        RECT 135.150 185.350 135.470 185.670 ;
        RECT 135.550 185.350 135.870 185.670 ;
        RECT 135.950 185.350 136.270 185.670 ;
        RECT 136.350 185.350 136.670 185.670 ;
        RECT 138.170 183.650 138.490 183.970 ;
        RECT 112.410 182.970 112.730 183.290 ;
        RECT 89.750 182.630 90.070 182.950 ;
        RECT 90.150 182.630 90.470 182.950 ;
        RECT 90.550 182.630 90.870 182.950 ;
        RECT 90.950 182.630 91.270 182.950 ;
        RECT 91.350 182.630 91.670 182.950 ;
        RECT 119.750 182.630 120.070 182.950 ;
        RECT 120.150 182.630 120.470 182.950 ;
        RECT 120.550 182.630 120.870 182.950 ;
        RECT 120.950 182.630 121.270 182.950 ;
        RECT 121.350 182.630 121.670 182.950 ;
        RECT 149.750 182.630 150.070 182.950 ;
        RECT 150.150 182.630 150.470 182.950 ;
        RECT 150.550 182.630 150.870 182.950 ;
        RECT 150.950 182.630 151.270 182.950 ;
        RECT 151.350 182.630 151.670 182.950 ;
        RECT 74.750 179.910 75.070 180.230 ;
        RECT 75.150 179.910 75.470 180.230 ;
        RECT 75.550 179.910 75.870 180.230 ;
        RECT 75.950 179.910 76.270 180.230 ;
        RECT 76.350 179.910 76.670 180.230 ;
        RECT 104.750 179.910 105.070 180.230 ;
        RECT 105.150 179.910 105.470 180.230 ;
        RECT 105.550 179.910 105.870 180.230 ;
        RECT 105.950 179.910 106.270 180.230 ;
        RECT 106.350 179.910 106.670 180.230 ;
        RECT 134.750 179.910 135.070 180.230 ;
        RECT 135.150 179.910 135.470 180.230 ;
        RECT 135.550 179.910 135.870 180.230 ;
        RECT 135.950 179.910 136.270 180.230 ;
        RECT 136.350 179.910 136.670 180.230 ;
        RECT 131.730 178.890 132.050 179.210 ;
        RECT 89.750 177.190 90.070 177.510 ;
        RECT 90.150 177.190 90.470 177.510 ;
        RECT 90.550 177.190 90.870 177.510 ;
        RECT 90.950 177.190 91.270 177.510 ;
        RECT 91.350 177.190 91.670 177.510 ;
        RECT 119.750 177.190 120.070 177.510 ;
        RECT 120.150 177.190 120.470 177.510 ;
        RECT 120.550 177.190 120.870 177.510 ;
        RECT 120.950 177.190 121.270 177.510 ;
        RECT 121.350 177.190 121.670 177.510 ;
        RECT 149.750 177.190 150.070 177.510 ;
        RECT 150.150 177.190 150.470 177.510 ;
        RECT 150.550 177.190 150.870 177.510 ;
        RECT 150.950 177.190 151.270 177.510 ;
        RECT 151.350 177.190 151.670 177.510 ;
        RECT 128.970 175.490 129.290 175.810 ;
        RECT 112.410 174.810 112.730 175.130 ;
        RECT 74.750 174.470 75.070 174.790 ;
        RECT 75.150 174.470 75.470 174.790 ;
        RECT 75.550 174.470 75.870 174.790 ;
        RECT 75.950 174.470 76.270 174.790 ;
        RECT 76.350 174.470 76.670 174.790 ;
        RECT 104.750 174.470 105.070 174.790 ;
        RECT 105.150 174.470 105.470 174.790 ;
        RECT 105.550 174.470 105.870 174.790 ;
        RECT 105.950 174.470 106.270 174.790 ;
        RECT 106.350 174.470 106.670 174.790 ;
        RECT 134.750 174.470 135.070 174.790 ;
        RECT 135.150 174.470 135.470 174.790 ;
        RECT 135.550 174.470 135.870 174.790 ;
        RECT 135.950 174.470 136.270 174.790 ;
        RECT 136.350 174.470 136.670 174.790 ;
        RECT 89.750 171.750 90.070 172.070 ;
        RECT 90.150 171.750 90.470 172.070 ;
        RECT 90.550 171.750 90.870 172.070 ;
        RECT 90.950 171.750 91.270 172.070 ;
        RECT 91.350 171.750 91.670 172.070 ;
        RECT 119.750 171.750 120.070 172.070 ;
        RECT 120.150 171.750 120.470 172.070 ;
        RECT 120.550 171.750 120.870 172.070 ;
        RECT 120.950 171.750 121.270 172.070 ;
        RECT 121.350 171.750 121.670 172.070 ;
        RECT 149.750 171.750 150.070 172.070 ;
        RECT 150.150 171.750 150.470 172.070 ;
        RECT 150.550 171.750 150.870 172.070 ;
        RECT 150.950 171.750 151.270 172.070 ;
        RECT 151.350 171.750 151.670 172.070 ;
        RECT 74.750 169.030 75.070 169.350 ;
        RECT 75.150 169.030 75.470 169.350 ;
        RECT 75.550 169.030 75.870 169.350 ;
        RECT 75.950 169.030 76.270 169.350 ;
        RECT 76.350 169.030 76.670 169.350 ;
        RECT 104.750 169.030 105.070 169.350 ;
        RECT 105.150 169.030 105.470 169.350 ;
        RECT 105.550 169.030 105.870 169.350 ;
        RECT 105.950 169.030 106.270 169.350 ;
        RECT 106.350 169.030 106.670 169.350 ;
        RECT 134.750 169.030 135.070 169.350 ;
        RECT 135.150 169.030 135.470 169.350 ;
        RECT 135.550 169.030 135.870 169.350 ;
        RECT 135.950 169.030 136.270 169.350 ;
        RECT 136.350 169.030 136.670 169.350 ;
        RECT 89.750 166.310 90.070 166.630 ;
        RECT 90.150 166.310 90.470 166.630 ;
        RECT 90.550 166.310 90.870 166.630 ;
        RECT 90.950 166.310 91.270 166.630 ;
        RECT 91.350 166.310 91.670 166.630 ;
        RECT 119.750 166.310 120.070 166.630 ;
        RECT 120.150 166.310 120.470 166.630 ;
        RECT 120.550 166.310 120.870 166.630 ;
        RECT 120.950 166.310 121.270 166.630 ;
        RECT 121.350 166.310 121.670 166.630 ;
        RECT 149.750 166.310 150.070 166.630 ;
        RECT 150.150 166.310 150.470 166.630 ;
        RECT 150.550 166.310 150.870 166.630 ;
        RECT 150.950 166.310 151.270 166.630 ;
        RECT 151.350 166.310 151.670 166.630 ;
        RECT 74.750 163.590 75.070 163.910 ;
        RECT 75.150 163.590 75.470 163.910 ;
        RECT 75.550 163.590 75.870 163.910 ;
        RECT 75.950 163.590 76.270 163.910 ;
        RECT 76.350 163.590 76.670 163.910 ;
        RECT 104.750 163.590 105.070 163.910 ;
        RECT 105.150 163.590 105.470 163.910 ;
        RECT 105.550 163.590 105.870 163.910 ;
        RECT 105.950 163.590 106.270 163.910 ;
        RECT 106.350 163.590 106.670 163.910 ;
        RECT 134.750 163.590 135.070 163.910 ;
        RECT 135.150 163.590 135.470 163.910 ;
        RECT 135.550 163.590 135.870 163.910 ;
        RECT 135.950 163.590 136.270 163.910 ;
        RECT 136.350 163.590 136.670 163.910 ;
        RECT 89.750 160.870 90.070 161.190 ;
        RECT 90.150 160.870 90.470 161.190 ;
        RECT 90.550 160.870 90.870 161.190 ;
        RECT 90.950 160.870 91.270 161.190 ;
        RECT 91.350 160.870 91.670 161.190 ;
        RECT 119.750 160.870 120.070 161.190 ;
        RECT 120.150 160.870 120.470 161.190 ;
        RECT 120.550 160.870 120.870 161.190 ;
        RECT 120.950 160.870 121.270 161.190 ;
        RECT 121.350 160.870 121.670 161.190 ;
        RECT 149.750 160.870 150.070 161.190 ;
        RECT 150.150 160.870 150.470 161.190 ;
        RECT 150.550 160.870 150.870 161.190 ;
        RECT 150.950 160.870 151.270 161.190 ;
        RECT 151.350 160.870 151.670 161.190 ;
        RECT 74.750 158.150 75.070 158.470 ;
        RECT 75.150 158.150 75.470 158.470 ;
        RECT 75.550 158.150 75.870 158.470 ;
        RECT 75.950 158.150 76.270 158.470 ;
        RECT 76.350 158.150 76.670 158.470 ;
        RECT 104.750 158.150 105.070 158.470 ;
        RECT 105.150 158.150 105.470 158.470 ;
        RECT 105.550 158.150 105.870 158.470 ;
        RECT 105.950 158.150 106.270 158.470 ;
        RECT 106.350 158.150 106.670 158.470 ;
        RECT 134.750 158.150 135.070 158.470 ;
        RECT 135.150 158.150 135.470 158.470 ;
        RECT 135.550 158.150 135.870 158.470 ;
        RECT 135.950 158.150 136.270 158.470 ;
        RECT 136.350 158.150 136.670 158.470 ;
        RECT 97.690 157.130 98.010 157.450 ;
        RECT 138.170 157.130 138.490 157.450 ;
        RECT 137.250 155.770 137.570 156.090 ;
        RECT 89.750 155.430 90.070 155.750 ;
        RECT 90.150 155.430 90.470 155.750 ;
        RECT 90.550 155.430 90.870 155.750 ;
        RECT 90.950 155.430 91.270 155.750 ;
        RECT 91.350 155.430 91.670 155.750 ;
        RECT 119.750 155.430 120.070 155.750 ;
        RECT 120.150 155.430 120.470 155.750 ;
        RECT 120.550 155.430 120.870 155.750 ;
        RECT 120.950 155.430 121.270 155.750 ;
        RECT 121.350 155.430 121.670 155.750 ;
        RECT 149.750 155.430 150.070 155.750 ;
        RECT 150.150 155.430 150.470 155.750 ;
        RECT 150.550 155.430 150.870 155.750 ;
        RECT 150.950 155.430 151.270 155.750 ;
        RECT 151.350 155.430 151.670 155.750 ;
        RECT 141.850 155.090 142.170 155.410 ;
        RECT 117.010 153.050 117.330 153.370 ;
        RECT 74.750 152.710 75.070 153.030 ;
        RECT 75.150 152.710 75.470 153.030 ;
        RECT 75.550 152.710 75.870 153.030 ;
        RECT 75.950 152.710 76.270 153.030 ;
        RECT 76.350 152.710 76.670 153.030 ;
        RECT 104.750 152.710 105.070 153.030 ;
        RECT 105.150 152.710 105.470 153.030 ;
        RECT 105.550 152.710 105.870 153.030 ;
        RECT 105.950 152.710 106.270 153.030 ;
        RECT 106.350 152.710 106.670 153.030 ;
        RECT 134.750 152.710 135.070 153.030 ;
        RECT 135.150 152.710 135.470 153.030 ;
        RECT 135.550 152.710 135.870 153.030 ;
        RECT 135.950 152.710 136.270 153.030 ;
        RECT 136.350 152.710 136.670 153.030 ;
        RECT 137.250 151.010 137.570 151.330 ;
        RECT 89.750 149.990 90.070 150.310 ;
        RECT 90.150 149.990 90.470 150.310 ;
        RECT 90.550 149.990 90.870 150.310 ;
        RECT 90.950 149.990 91.270 150.310 ;
        RECT 91.350 149.990 91.670 150.310 ;
        RECT 119.750 149.990 120.070 150.310 ;
        RECT 120.150 149.990 120.470 150.310 ;
        RECT 120.550 149.990 120.870 150.310 ;
        RECT 120.950 149.990 121.270 150.310 ;
        RECT 121.350 149.990 121.670 150.310 ;
        RECT 149.750 149.990 150.070 150.310 ;
        RECT 150.150 149.990 150.470 150.310 ;
        RECT 150.550 149.990 150.870 150.310 ;
        RECT 150.950 149.990 151.270 150.310 ;
        RECT 151.350 149.990 151.670 150.310 ;
        RECT 131.730 149.650 132.050 149.970 ;
        RECT 74.750 147.270 75.070 147.590 ;
        RECT 75.150 147.270 75.470 147.590 ;
        RECT 75.550 147.270 75.870 147.590 ;
        RECT 75.950 147.270 76.270 147.590 ;
        RECT 76.350 147.270 76.670 147.590 ;
        RECT 104.750 147.270 105.070 147.590 ;
        RECT 105.150 147.270 105.470 147.590 ;
        RECT 105.550 147.270 105.870 147.590 ;
        RECT 105.950 147.270 106.270 147.590 ;
        RECT 106.350 147.270 106.670 147.590 ;
        RECT 134.750 147.270 135.070 147.590 ;
        RECT 135.150 147.270 135.470 147.590 ;
        RECT 135.550 147.270 135.870 147.590 ;
        RECT 135.950 147.270 136.270 147.590 ;
        RECT 136.350 147.270 136.670 147.590 ;
        RECT 117.930 146.250 118.250 146.570 ;
        RECT 89.750 144.550 90.070 144.870 ;
        RECT 90.150 144.550 90.470 144.870 ;
        RECT 90.550 144.550 90.870 144.870 ;
        RECT 90.950 144.550 91.270 144.870 ;
        RECT 91.350 144.550 91.670 144.870 ;
        RECT 107.810 144.890 108.130 145.210 ;
        RECT 119.750 144.550 120.070 144.870 ;
        RECT 120.150 144.550 120.470 144.870 ;
        RECT 120.550 144.550 120.870 144.870 ;
        RECT 120.950 144.550 121.270 144.870 ;
        RECT 121.350 144.550 121.670 144.870 ;
        RECT 149.750 144.550 150.070 144.870 ;
        RECT 150.150 144.550 150.470 144.870 ;
        RECT 150.550 144.550 150.870 144.870 ;
        RECT 150.950 144.550 151.270 144.870 ;
        RECT 151.350 144.550 151.670 144.870 ;
        RECT 74.750 141.830 75.070 142.150 ;
        RECT 75.150 141.830 75.470 142.150 ;
        RECT 75.550 141.830 75.870 142.150 ;
        RECT 75.950 141.830 76.270 142.150 ;
        RECT 76.350 141.830 76.670 142.150 ;
        RECT 104.750 141.830 105.070 142.150 ;
        RECT 105.150 141.830 105.470 142.150 ;
        RECT 105.550 141.830 105.870 142.150 ;
        RECT 105.950 141.830 106.270 142.150 ;
        RECT 106.350 141.830 106.670 142.150 ;
        RECT 134.750 141.830 135.070 142.150 ;
        RECT 135.150 141.830 135.470 142.150 ;
        RECT 135.550 141.830 135.870 142.150 ;
        RECT 135.950 141.830 136.270 142.150 ;
        RECT 136.350 141.830 136.670 142.150 ;
        RECT 143.690 140.130 144.010 140.450 ;
        RECT 128.970 139.450 129.290 139.770 ;
        RECT 89.750 139.110 90.070 139.430 ;
        RECT 90.150 139.110 90.470 139.430 ;
        RECT 90.550 139.110 90.870 139.430 ;
        RECT 90.950 139.110 91.270 139.430 ;
        RECT 91.350 139.110 91.670 139.430 ;
        RECT 119.750 139.110 120.070 139.430 ;
        RECT 120.150 139.110 120.470 139.430 ;
        RECT 120.550 139.110 120.870 139.430 ;
        RECT 120.950 139.110 121.270 139.430 ;
        RECT 121.350 139.110 121.670 139.430 ;
        RECT 149.750 139.110 150.070 139.430 ;
        RECT 150.150 139.110 150.470 139.430 ;
        RECT 150.550 139.110 150.870 139.430 ;
        RECT 150.950 139.110 151.270 139.430 ;
        RECT 151.350 139.110 151.670 139.430 ;
        RECT 97.690 136.730 98.010 137.050 ;
        RECT 117.010 136.730 117.330 137.050 ;
        RECT 74.750 136.390 75.070 136.710 ;
        RECT 75.150 136.390 75.470 136.710 ;
        RECT 75.550 136.390 75.870 136.710 ;
        RECT 75.950 136.390 76.270 136.710 ;
        RECT 76.350 136.390 76.670 136.710 ;
        RECT 104.750 136.390 105.070 136.710 ;
        RECT 105.150 136.390 105.470 136.710 ;
        RECT 105.550 136.390 105.870 136.710 ;
        RECT 105.950 136.390 106.270 136.710 ;
        RECT 106.350 136.390 106.670 136.710 ;
        RECT 134.750 136.390 135.070 136.710 ;
        RECT 135.150 136.390 135.470 136.710 ;
        RECT 135.550 136.390 135.870 136.710 ;
        RECT 135.950 136.390 136.270 136.710 ;
        RECT 136.350 136.390 136.670 136.710 ;
        RECT 107.810 134.690 108.130 135.010 ;
        RECT 89.750 133.670 90.070 133.990 ;
        RECT 90.150 133.670 90.470 133.990 ;
        RECT 90.550 133.670 90.870 133.990 ;
        RECT 90.950 133.670 91.270 133.990 ;
        RECT 91.350 133.670 91.670 133.990 ;
        RECT 119.750 133.670 120.070 133.990 ;
        RECT 120.150 133.670 120.470 133.990 ;
        RECT 120.550 133.670 120.870 133.990 ;
        RECT 120.950 133.670 121.270 133.990 ;
        RECT 121.350 133.670 121.670 133.990 ;
        RECT 149.750 133.670 150.070 133.990 ;
        RECT 150.150 133.670 150.470 133.990 ;
        RECT 150.550 133.670 150.870 133.990 ;
        RECT 150.950 133.670 151.270 133.990 ;
        RECT 151.350 133.670 151.670 133.990 ;
        RECT 100.450 133.330 100.770 133.650 ;
        RECT 141.850 133.330 142.170 133.650 ;
        RECT 98.610 131.970 98.930 132.290 ;
        RECT 114.250 131.970 114.570 132.290 ;
        RECT 74.750 130.950 75.070 131.270 ;
        RECT 75.150 130.950 75.470 131.270 ;
        RECT 75.550 130.950 75.870 131.270 ;
        RECT 75.950 130.950 76.270 131.270 ;
        RECT 76.350 130.950 76.670 131.270 ;
        RECT 104.750 130.950 105.070 131.270 ;
        RECT 105.150 130.950 105.470 131.270 ;
        RECT 105.550 130.950 105.870 131.270 ;
        RECT 105.950 130.950 106.270 131.270 ;
        RECT 106.350 130.950 106.670 131.270 ;
        RECT 134.750 130.950 135.070 131.270 ;
        RECT 135.150 130.950 135.470 131.270 ;
        RECT 135.550 130.950 135.870 131.270 ;
        RECT 135.950 130.950 136.270 131.270 ;
        RECT 136.350 130.950 136.670 131.270 ;
        RECT 89.750 128.230 90.070 128.550 ;
        RECT 90.150 128.230 90.470 128.550 ;
        RECT 90.550 128.230 90.870 128.550 ;
        RECT 90.950 128.230 91.270 128.550 ;
        RECT 91.350 128.230 91.670 128.550 ;
        RECT 133.570 129.930 133.890 130.250 ;
        RECT 111.490 129.250 111.810 129.570 ;
        RECT 117.930 128.570 118.250 128.890 ;
        RECT 119.750 128.230 120.070 128.550 ;
        RECT 120.150 128.230 120.470 128.550 ;
        RECT 120.550 128.230 120.870 128.550 ;
        RECT 120.950 128.230 121.270 128.550 ;
        RECT 121.350 128.230 121.670 128.550 ;
        RECT 149.750 128.230 150.070 128.550 ;
        RECT 150.150 128.230 150.470 128.550 ;
        RECT 150.550 128.230 150.870 128.550 ;
        RECT 150.950 128.230 151.270 128.550 ;
        RECT 151.350 128.230 151.670 128.550 ;
        RECT 117.010 127.890 117.330 128.210 ;
        RECT 143.690 127.890 144.010 128.210 ;
        RECT 117.930 126.530 118.250 126.850 ;
        RECT 124.370 126.530 124.690 126.850 ;
        RECT 143.690 126.530 144.010 126.850 ;
        RECT 117.010 125.850 117.330 126.170 ;
        RECT 74.750 125.510 75.070 125.830 ;
        RECT 75.150 125.510 75.470 125.830 ;
        RECT 75.550 125.510 75.870 125.830 ;
        RECT 75.950 125.510 76.270 125.830 ;
        RECT 76.350 125.510 76.670 125.830 ;
        RECT 104.750 125.510 105.070 125.830 ;
        RECT 105.150 125.510 105.470 125.830 ;
        RECT 105.550 125.510 105.870 125.830 ;
        RECT 105.950 125.510 106.270 125.830 ;
        RECT 106.350 125.510 106.670 125.830 ;
        RECT 134.750 125.510 135.070 125.830 ;
        RECT 135.150 125.510 135.470 125.830 ;
        RECT 135.550 125.510 135.870 125.830 ;
        RECT 135.950 125.510 136.270 125.830 ;
        RECT 136.350 125.510 136.670 125.830 ;
        RECT 89.750 122.790 90.070 123.110 ;
        RECT 90.150 122.790 90.470 123.110 ;
        RECT 90.550 122.790 90.870 123.110 ;
        RECT 90.950 122.790 91.270 123.110 ;
        RECT 91.350 122.790 91.670 123.110 ;
        RECT 119.750 122.790 120.070 123.110 ;
        RECT 120.150 122.790 120.470 123.110 ;
        RECT 120.550 122.790 120.870 123.110 ;
        RECT 120.950 122.790 121.270 123.110 ;
        RECT 121.350 122.790 121.670 123.110 ;
        RECT 149.750 122.790 150.070 123.110 ;
        RECT 150.150 122.790 150.470 123.110 ;
        RECT 150.550 122.790 150.870 123.110 ;
        RECT 150.950 122.790 151.270 123.110 ;
        RECT 151.350 122.790 151.670 123.110 ;
      LAYER met4 ;
        RECT 3.990 222.190 4.290 224.760 ;
        RECT 7.670 222.190 7.970 224.760 ;
        RECT 11.350 222.190 11.650 224.760 ;
        RECT 15.030 222.190 15.330 224.760 ;
        RECT 18.710 222.190 19.010 224.760 ;
        RECT 22.390 222.190 22.690 224.760 ;
        RECT 26.070 222.190 26.370 224.760 ;
        RECT 29.750 222.190 30.050 224.760 ;
        RECT 33.430 222.190 33.730 224.760 ;
        RECT 37.110 222.190 37.410 224.760 ;
        RECT 40.790 222.190 41.090 224.760 ;
        RECT 44.470 222.190 44.770 224.760 ;
        RECT 48.150 222.190 48.450 224.760 ;
        RECT 51.830 222.190 52.130 224.760 ;
        RECT 55.510 222.190 55.810 224.760 ;
        RECT 59.190 222.190 59.490 224.760 ;
        RECT 62.870 222.190 63.170 224.760 ;
        RECT 66.550 222.190 66.850 224.760 ;
        RECT 70.230 222.190 70.530 224.760 ;
        RECT 73.910 222.190 74.210 224.760 ;
        RECT 77.590 222.190 77.890 224.760 ;
        RECT 81.270 222.190 81.570 224.760 ;
        RECT 84.950 222.190 85.250 224.760 ;
        RECT 88.630 223.440 88.930 224.760 ;
        RECT 92.310 223.440 92.610 224.760 ;
        RECT 95.990 223.440 96.290 224.760 ;
        RECT 99.670 223.440 99.970 224.760 ;
        RECT 103.350 223.440 103.650 224.760 ;
        RECT 107.030 223.440 107.330 224.760 ;
        RECT 110.710 223.440 111.010 224.760 ;
        RECT 10.500 220.760 29.000 222.190 ;
        RECT 10.500 219.630 19.000 220.760 ;
        RECT 20.500 219.630 29.000 220.760 ;
        RECT 114.390 216.550 114.690 224.760 ;
        RECT 118.070 216.550 118.370 224.760 ;
        RECT 121.750 218.150 122.050 224.760 ;
        RECT 112.650 216.250 114.690 216.550 ;
        RECT 116.650 216.250 118.370 216.550 ;
        RECT 120.550 217.850 122.050 218.150 ;
        RECT 110.240 215.250 110.760 215.360 ;
        RECT 112.650 215.250 112.950 216.250 ;
        RECT 116.650 215.300 116.950 216.250 ;
        RECT 120.550 215.415 120.850 217.850 ;
        RECT 125.430 216.910 125.730 224.760 ;
        RECT 129.110 222.450 129.410 224.760 ;
        RECT 126.550 222.150 129.410 222.450 ;
        RECT 125.370 216.490 125.790 216.910 ;
        RECT 126.550 216.905 126.850 222.150 ;
        RECT 127.805 221.450 128.200 221.500 ;
        RECT 132.790 221.450 133.090 224.760 ;
        RECT 127.805 221.150 133.090 221.450 ;
        RECT 127.805 221.105 128.200 221.150 ;
        RECT 131.910 220.450 132.295 220.495 ;
        RECT 136.470 220.450 136.770 224.760 ;
        RECT 131.910 220.150 136.770 220.450 ;
        RECT 131.910 220.110 132.295 220.150 ;
        RECT 136.035 219.250 136.365 219.265 ;
        RECT 140.150 219.250 140.450 224.760 ;
        RECT 136.035 218.950 140.450 219.250 ;
        RECT 136.035 218.935 136.365 218.950 ;
        RECT 140.205 217.950 140.600 218.000 ;
        RECT 143.830 217.950 144.130 224.760 ;
        RECT 147.510 224.085 147.810 224.760 ;
        RECT 140.205 217.650 144.130 217.950 ;
        RECT 140.205 217.605 140.600 217.650 ;
        RECT 126.495 216.495 126.905 216.905 ;
        RECT 144.270 216.765 144.730 216.830 ;
        RECT 147.495 216.765 147.825 224.085 ;
        RECT 144.270 216.435 147.825 216.765 ;
        RECT 144.270 216.370 144.730 216.435 ;
        RECT 148.485 215.550 148.915 215.615 ;
        RECT 151.190 215.550 151.490 224.760 ;
        RECT 110.240 214.950 112.950 215.250 ;
        RECT 110.240 214.840 110.760 214.950 ;
        RECT 116.600 214.900 117.000 215.300 ;
        RECT 120.490 214.990 120.915 215.415 ;
        RECT 148.485 215.250 151.490 215.550 ;
        RECT 152.570 215.550 153.030 215.630 ;
        RECT 154.870 215.550 155.170 224.760 ;
        RECT 152.570 215.250 155.170 215.550 ;
        RECT 148.485 215.185 148.915 215.250 ;
        RECT 152.570 215.170 153.030 215.250 ;
        RECT 74.710 122.710 76.710 207.510 ;
        RECT 89.710 122.710 91.710 207.510 ;
        RECT 100.445 203.365 100.775 203.695 ;
        RECT 98.605 196.565 98.935 196.895 ;
        RECT 97.685 157.125 98.015 157.455 ;
        RECT 97.700 137.055 98.000 157.125 ;
        RECT 97.685 136.725 98.015 137.055 ;
        RECT 98.620 132.295 98.920 196.565 ;
        RECT 100.460 133.655 100.760 203.365 ;
        RECT 100.445 133.325 100.775 133.655 ;
        RECT 98.605 131.965 98.935 132.295 ;
        RECT 104.710 122.710 106.710 207.510 ;
        RECT 111.485 203.365 111.815 203.695 ;
        RECT 107.805 144.885 108.135 145.215 ;
        RECT 107.820 135.015 108.120 144.885 ;
        RECT 107.805 134.685 108.135 135.015 ;
        RECT 111.500 129.575 111.800 203.365 ;
        RECT 114.245 197.245 114.575 197.575 ;
        RECT 112.405 182.965 112.735 183.295 ;
        RECT 112.420 175.135 112.720 182.965 ;
        RECT 112.405 174.805 112.735 175.135 ;
        RECT 114.260 132.295 114.560 197.245 ;
        RECT 117.005 153.045 117.335 153.375 ;
        RECT 117.020 137.055 117.320 153.045 ;
        RECT 117.925 146.245 118.255 146.575 ;
        RECT 117.005 136.725 117.335 137.055 ;
        RECT 114.245 131.965 114.575 132.295 ;
        RECT 111.485 129.245 111.815 129.575 ;
        RECT 117.940 128.895 118.240 146.245 ;
        RECT 117.925 128.565 118.255 128.895 ;
        RECT 117.005 127.885 117.335 128.215 ;
        RECT 117.020 126.175 117.320 127.885 ;
        RECT 117.940 126.855 118.240 128.565 ;
        RECT 117.925 126.525 118.255 126.855 ;
        RECT 117.005 125.845 117.335 126.175 ;
        RECT 119.710 122.710 121.710 207.510 ;
        RECT 124.365 196.565 124.695 196.895 ;
        RECT 133.565 196.565 133.895 196.895 ;
        RECT 124.380 126.855 124.680 196.565 ;
        RECT 131.725 178.885 132.055 179.215 ;
        RECT 128.965 175.485 129.295 175.815 ;
        RECT 128.980 139.775 129.280 175.485 ;
        RECT 131.740 149.975 132.040 178.885 ;
        RECT 131.725 149.645 132.055 149.975 ;
        RECT 128.965 139.445 129.295 139.775 ;
        RECT 133.580 130.255 133.880 196.565 ;
        RECT 133.565 129.925 133.895 130.255 ;
        RECT 124.365 126.525 124.695 126.855 ;
        RECT 134.710 122.710 136.710 207.510 ;
        RECT 138.165 183.645 138.495 183.975 ;
        RECT 138.180 157.455 138.480 183.645 ;
        RECT 138.165 157.125 138.495 157.455 ;
        RECT 137.245 155.765 137.575 156.095 ;
        RECT 137.260 151.335 137.560 155.765 ;
        RECT 141.845 155.085 142.175 155.415 ;
        RECT 137.245 151.005 137.575 151.335 ;
        RECT 141.860 133.655 142.160 155.085 ;
        RECT 143.685 140.125 144.015 140.455 ;
        RECT 141.845 133.325 142.175 133.655 ;
        RECT 143.700 128.215 144.000 140.125 ;
        RECT 143.685 127.885 144.015 128.215 ;
        RECT 143.700 126.855 144.000 127.885 ;
        RECT 143.685 126.525 144.015 126.855 ;
        RECT 149.710 122.710 151.710 207.510 ;
        RECT 5.415 30.685 6.425 30.690 ;
        RECT 2.500 29.685 6.425 30.685 ;
        RECT 5.415 29.680 6.425 29.685 ;
        RECT 134.480 1.000 135.080 2.440 ;
        RECT 156.560 1.000 157.160 2.440 ;
  END
END tt_um_algofoogle_tt06_grab_bag
END LIBRARY

