Cosimulation of Anton's VGA digital test block with 3 R2R DACs, using Verilator and d_cosim in ngspice-42

*.lib /home/matt/work/asic-workshop/shuttle-2404/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.lib /home/anton/.volare/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* https://sourceforge.net/p/ngspice/ngspice/ci/master/tree/examples/xspice/verilator/

* The digital portion of the circuit is specified in compiled Verilog.
* list the inputs and outputs.
* NOTE: We name bus signals individually, in the order they're defined in the Verilog:
adut 
+ [ clk rst_n in7 in6 in5 in4 in3 in2 in1 in0 ] 
+ [ 
+ hsync vsync hblank vblank 
+ r7 r6 r5 r4 r3 r2 r1 r0 
+ g7 g6 g5 g4 g3 g2 g1 g0
+ b7 b6 b5 b4 b3 b2 b1 b0 
+ dr7 dg7 db7 
+ dr6 dg6 db6 
+ m7 m6 m5 m4 m3 m2 m1 m0 
+ o_reset o_visible
+ c7 c6 c5 c4 c3 c2 c1 c0 
+ o_clk
+ x7 x6 x5 x4 x3 x2 x1 x0 
+ o_clk2 o_zero o_one
+] null dut
.model dut d_cosim simulation="./spicewrap.so"

* connect the driver to the R2R dac
* had to edit spice exported by xschem to add the subckt and ends

.include "../xschem/simulation/r2r.spice" 
*.include "../mag/r2r.spice" 

xr2r_R red      r7 r6 r5 r4 r3 r2 r1 r0 GND GND r2r
xr2r_G green    g7 g6 g5 g4 g3 g2 g1 g0 GND GND r2r
xr2r_B blue     b7 b6 b5 b4 b3 b2 b1 b0 GND GND r2r

* simulate tt output path
Cr1 red             GND 2.5p
Rr1 red             red_pin_out 500
Cr2 red_pin_out     GND 2.5p

Cg1 green           GND 2.5p
Rg1 green           green_pin_out 500
Cg2 green_pin_out   GND 2.5p

Cb1 blue            GND 2.5p
Rb1 blue            blue_pin_out 500
Cb2 blue_pin_out    GND 2.5p

**** End of the ADC and its subcircuits.  Begin test circuit ****

.param vcc=1.8
vcc vcc 0 {vcc}

* Digital clock signal

aclock 0 clk clock
.model clock d_osc cntl_array=[-1 1] freq_array=[25Meg 25Meg]

* reset signal

Vreset rst_n GND PULSE 1.8 0 1n 20p 20p 1u 500u

* DAC input value
Vin0 in0 GND PULSE 0 1.8 2u 0p 0p 20n 40n
Vin1 in1 GND PULSE 0 1.8 2u 0p 0p 40n 80n
Vin2 in2 GND PULSE 0 1.8 2u 0p 0p 80n 160n
Vin3 in3 GND PULSE 0 1.8 2u 0p 0p 160n 320n
Vin4 in4 GND PULSE 0 1.8 2u 0p 0p 320n 640n
Vin5 in5 GND PULSE 0 1.8 2u 0p 0p 640n 1280n
Vin6 in6 GND PULSE 0 1.8 2u 0p 0p 1280n 2560n
Vin7 in7 GND PULSE 0 1.8 2u 0p 0p 2560n 5120n

.control
tran 2n 30u
* plot in0
* plot in1
* plot in2
* plot rst_n
* plot clk
* plot red_pin_out
* plot hsync
* plot vsync
* plot hblank
* plot vblank
* plot dr7
* plot dg7
* plot db7
* plot dr6
* plot dg6
* plot db6
.endc
.end
