VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_algofoogle_tt06_grab_bag
  CLASS BLOCK ;
  FOREIGN tt_um_algofoogle_tt06_grab_bag ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.480000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 423.736481 ;
    ANTENNADIFFAREA 564.607666 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 423.736481 ;
    ANTENNADIFFAREA 564.607666 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 423.736481 ;
    ANTENNADIFFAREA 564.607666 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.480000 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 670.274109 ;
    ANTENNADIFFAREA 954.641174 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 10.500 5.000 12.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 35.910 213.435 150.370 215.040 ;
      LAYER pwell ;
        RECT 36.105 212.235 37.475 213.045 ;
        RECT 37.485 212.235 42.995 213.045 ;
        RECT 43.005 212.235 44.835 213.045 ;
        RECT 47.500 212.915 48.420 213.145 ;
        RECT 44.955 212.235 48.420 212.915 ;
        RECT 48.995 212.320 49.425 213.105 ;
        RECT 49.445 212.235 54.955 213.045 ;
        RECT 55.885 212.915 57.230 213.145 ;
        RECT 55.885 212.235 57.715 212.915 ;
        RECT 58.655 212.235 61.395 212.915 ;
        RECT 61.875 212.320 62.305 213.105 ;
        RECT 63.730 212.915 65.075 213.145 ;
        RECT 63.245 212.235 65.075 212.915 ;
        RECT 66.015 212.235 68.755 212.915 ;
        RECT 68.765 212.235 70.595 213.045 ;
        RECT 70.605 212.915 71.950 213.145 ;
        RECT 70.605 212.235 72.435 212.915 ;
        RECT 72.445 212.235 73.795 213.145 ;
        RECT 74.755 212.320 75.185 213.105 ;
        RECT 78.450 212.915 79.795 213.145 ;
        RECT 75.215 212.235 77.955 212.915 ;
        RECT 77.965 212.235 79.795 212.915 ;
        RECT 80.735 212.235 83.475 212.915 ;
        RECT 83.485 212.235 85.315 213.045 ;
        RECT 85.325 212.915 86.670 213.145 ;
        RECT 85.325 212.235 87.155 212.915 ;
        RECT 87.635 212.320 88.065 213.105 ;
        RECT 88.095 212.235 90.835 212.915 ;
        RECT 90.845 212.235 96.355 213.045 ;
        RECT 96.365 212.235 98.195 213.045 ;
        RECT 98.215 212.235 99.565 213.145 ;
        RECT 100.515 212.320 100.945 213.105 ;
        RECT 101.625 212.915 105.555 213.145 ;
        RECT 101.140 212.235 105.555 212.915 ;
        RECT 105.565 212.235 111.075 213.045 ;
        RECT 111.085 212.235 112.915 213.045 ;
        RECT 113.395 212.320 113.825 213.105 ;
        RECT 113.845 212.915 114.775 213.145 ;
        RECT 113.845 212.235 117.745 212.915 ;
        RECT 117.985 212.235 121.655 213.045 ;
        RECT 122.125 212.235 123.495 213.015 ;
        RECT 123.505 212.235 126.255 213.045 ;
        RECT 126.275 212.320 126.705 213.105 ;
        RECT 126.725 212.235 128.095 213.015 ;
        RECT 128.105 212.235 129.475 213.045 ;
        RECT 129.485 212.235 130.855 213.015 ;
        RECT 130.865 212.235 132.695 213.045 ;
        RECT 132.705 212.235 134.075 213.015 ;
        RECT 134.085 212.235 135.455 213.015 ;
        RECT 135.465 212.235 136.835 213.045 ;
        RECT 136.845 212.235 138.215 213.015 ;
        RECT 139.155 212.320 139.585 213.105 ;
        RECT 139.605 212.945 140.550 213.145 ;
        RECT 139.605 212.265 142.355 212.945 ;
        RECT 139.605 212.235 140.550 212.265 ;
        RECT 36.245 212.025 36.415 212.235 ;
        RECT 37.625 212.025 37.795 212.235 ;
        RECT 43.145 212.045 43.315 212.235 ;
        RECT 44.985 212.045 45.155 212.235 ;
        RECT 45.905 212.025 46.075 212.215 ;
        RECT 46.365 212.025 46.535 212.215 ;
        RECT 48.660 212.075 48.780 212.185 ;
        RECT 49.585 212.045 49.755 212.235 ;
        RECT 53.735 212.070 53.895 212.180 ;
        RECT 54.645 212.025 54.815 212.215 ;
        RECT 55.115 212.080 55.275 212.190 ;
        RECT 57.405 212.045 57.575 212.235 ;
        RECT 57.875 212.080 58.035 212.190 ;
        RECT 61.085 212.045 61.255 212.235 ;
        RECT 61.540 212.075 61.660 212.185 ;
        RECT 62.475 212.070 62.635 212.190 ;
        RECT 63.385 212.025 63.555 212.235 ;
        RECT 65.235 212.080 65.395 212.190 ;
        RECT 66.145 212.025 66.315 212.215 ;
        RECT 66.610 212.025 66.780 212.215 ;
        RECT 68.445 212.045 68.615 212.235 ;
        RECT 68.905 212.025 69.075 212.235 ;
        RECT 69.375 212.070 69.535 212.180 ;
        RECT 70.285 212.025 70.455 212.215 ;
        RECT 72.125 212.045 72.295 212.235 ;
        RECT 72.590 212.045 72.760 212.235 ;
        RECT 73.505 212.025 73.675 212.215 ;
        RECT 73.975 212.080 74.135 212.190 ;
        RECT 76.725 212.025 76.895 212.215 ;
        RECT 77.645 212.045 77.815 212.235 ;
        RECT 78.105 212.045 78.275 212.235 ;
        RECT 79.480 212.075 79.600 212.185 ;
        RECT 79.945 212.045 80.115 212.215 ;
        RECT 79.965 212.025 80.115 212.045 ;
        RECT 82.245 212.025 82.415 212.215 ;
        RECT 83.165 212.045 83.335 212.235 ;
        RECT 83.625 212.045 83.795 212.235 ;
        RECT 86.845 212.045 87.015 212.235 ;
        RECT 87.305 212.185 87.475 212.215 ;
        RECT 87.300 212.075 87.475 212.185 ;
        RECT 87.305 212.025 87.475 212.075 ;
        RECT 88.225 212.025 88.395 212.215 ;
        RECT 90.525 212.045 90.695 212.235 ;
        RECT 90.985 212.025 91.155 212.235 ;
        RECT 93.745 212.025 93.915 212.215 ;
        RECT 95.125 212.025 95.295 212.215 ;
        RECT 96.505 212.045 96.675 212.235 ;
        RECT 99.265 212.045 99.435 212.235 ;
        RECT 101.140 212.215 101.250 212.235 ;
        RECT 99.735 212.080 99.895 212.190 ;
        RECT 101.080 212.045 101.250 212.215 ;
        RECT 102.485 212.025 102.655 212.215 ;
        RECT 105.705 212.045 105.875 212.235 ;
        RECT 109.855 212.070 110.015 212.180 ;
        RECT 110.765 212.025 110.935 212.215 ;
        RECT 111.225 212.045 111.395 212.235 ;
        RECT 113.060 212.075 113.180 212.185 ;
        RECT 114.260 212.025 114.430 212.235 ;
        RECT 118.125 212.025 118.295 212.235 ;
        RECT 120.885 212.025 121.055 212.215 ;
        RECT 121.800 212.075 121.920 212.185 ;
        RECT 122.265 212.045 122.435 212.235 ;
        RECT 123.645 212.045 123.815 212.235 ;
        RECT 123.920 212.025 124.090 212.215 ;
        RECT 126.865 212.045 127.035 212.235 ;
        RECT 128.245 212.045 128.415 212.235 ;
        RECT 130.545 212.045 130.715 212.235 ;
        RECT 131.005 212.045 131.175 212.235 ;
        RECT 131.190 212.025 131.360 212.215 ;
        RECT 131.925 212.025 132.095 212.215 ;
        RECT 133.765 212.045 133.935 212.235 ;
        RECT 135.145 212.045 135.315 212.235 ;
        RECT 135.605 212.045 135.775 212.235 ;
        RECT 137.895 212.045 138.065 212.235 ;
        RECT 138.375 212.080 138.535 212.190 ;
        RECT 139.740 212.075 139.860 212.185 ;
        RECT 140.205 212.025 140.375 212.215 ;
        RECT 141.585 212.025 141.755 212.215 ;
        RECT 142.040 212.045 142.210 212.265 ;
        RECT 142.365 212.235 143.735 213.015 ;
        RECT 144.205 212.235 145.575 213.015 ;
        RECT 145.585 212.235 147.415 213.045 ;
        RECT 147.425 212.235 148.795 213.015 ;
        RECT 148.805 212.235 150.175 213.045 ;
        RECT 143.415 212.045 143.585 212.235 ;
        RECT 143.880 212.075 144.000 212.185 ;
        RECT 145.255 212.045 145.425 212.235 ;
        RECT 145.725 212.045 145.895 212.235 ;
        RECT 148.475 212.045 148.645 212.235 ;
        RECT 149.865 212.025 150.035 212.235 ;
        RECT 36.105 211.215 37.475 212.025 ;
        RECT 37.485 211.345 44.795 212.025 ;
        RECT 41.000 211.125 41.910 211.345 ;
        RECT 43.445 211.115 44.795 211.345 ;
        RECT 44.855 211.115 46.205 212.025 ;
        RECT 46.225 211.345 53.535 212.025 ;
        RECT 54.505 211.345 61.815 212.025 ;
        RECT 49.740 211.125 50.650 211.345 ;
        RECT 52.185 211.115 53.535 211.345 ;
        RECT 58.020 211.125 58.930 211.345 ;
        RECT 60.465 211.115 61.815 211.345 ;
        RECT 61.875 211.155 62.305 211.940 ;
        RECT 63.245 211.345 65.075 212.025 ;
        RECT 65.085 211.245 66.455 212.025 ;
        RECT 66.465 211.115 67.815 212.025 ;
        RECT 67.845 211.245 69.215 212.025 ;
        RECT 70.245 211.115 73.355 212.025 ;
        RECT 73.465 211.115 76.575 212.025 ;
        RECT 76.585 211.215 79.335 212.025 ;
        RECT 79.965 211.205 81.895 212.025 ;
        RECT 82.105 211.345 84.855 212.025 ;
        RECT 80.945 211.115 81.895 211.205 ;
        RECT 83.925 211.115 84.855 211.345 ;
        RECT 84.875 211.115 87.605 212.025 ;
        RECT 87.635 211.155 88.065 211.940 ;
        RECT 88.085 211.115 90.490 212.025 ;
        RECT 90.845 211.215 93.595 212.025 ;
        RECT 93.605 211.245 94.975 212.025 ;
        RECT 94.985 211.345 102.295 212.025 ;
        RECT 102.345 211.345 109.655 212.025 ;
        RECT 98.500 211.125 99.410 211.345 ;
        RECT 100.945 211.115 102.295 211.345 ;
        RECT 105.860 211.125 106.770 211.345 ;
        RECT 108.305 211.115 109.655 211.345 ;
        RECT 110.625 211.115 113.375 212.025 ;
        RECT 113.395 211.155 113.825 211.940 ;
        RECT 113.845 211.345 117.745 212.025 ;
        RECT 113.845 211.115 114.775 211.345 ;
        RECT 117.985 211.115 120.735 212.025 ;
        RECT 120.745 211.115 123.495 212.025 ;
        RECT 123.505 211.345 127.405 212.025 ;
        RECT 127.875 211.345 131.775 212.025 ;
        RECT 131.785 211.345 139.095 212.025 ;
        RECT 123.505 211.115 124.435 211.345 ;
        RECT 130.845 211.115 131.775 211.345 ;
        RECT 135.300 211.125 136.210 211.345 ;
        RECT 137.745 211.115 139.095 211.345 ;
        RECT 139.155 211.155 139.585 211.940 ;
        RECT 140.065 211.245 141.435 212.025 ;
        RECT 141.445 211.345 148.755 212.025 ;
        RECT 144.960 211.125 145.870 211.345 ;
        RECT 147.405 211.115 148.755 211.345 ;
        RECT 148.805 211.215 150.175 212.025 ;
      LAYER nwell ;
        RECT 35.910 207.995 150.370 210.825 ;
      LAYER pwell ;
        RECT 36.105 206.795 37.475 207.605 ;
        RECT 37.485 206.795 41.155 207.605 ;
        RECT 41.165 206.795 42.535 207.605 ;
        RECT 42.560 206.795 44.375 207.705 ;
        RECT 44.845 206.795 46.215 207.575 ;
        RECT 46.685 206.795 48.055 207.575 ;
        RECT 48.995 206.880 49.425 207.665 ;
        RECT 49.445 206.795 54.955 207.605 ;
        RECT 54.965 206.795 57.715 207.605 ;
        RECT 57.765 207.475 59.115 207.705 ;
        RECT 60.650 207.475 61.560 207.695 ;
        RECT 57.765 206.795 65.075 207.475 ;
        RECT 65.085 206.795 66.915 207.475 ;
        RECT 66.925 206.795 72.435 207.605 ;
        RECT 72.445 206.795 73.795 207.705 ;
        RECT 74.755 206.880 75.185 207.665 ;
        RECT 75.205 206.795 77.955 207.705 ;
        RECT 77.975 206.795 79.325 207.705 ;
        RECT 81.315 207.475 82.245 207.705 ;
        RECT 80.410 206.795 82.245 207.475 ;
        RECT 83.585 206.795 86.695 207.705 ;
        RECT 86.715 206.795 90.835 207.705 ;
        RECT 90.845 206.795 92.195 207.705 ;
        RECT 92.225 206.795 97.735 207.605 ;
        RECT 98.665 206.795 100.015 207.705 ;
        RECT 100.515 206.880 100.945 207.665 ;
        RECT 101.505 206.795 103.715 207.705 ;
        RECT 103.725 206.795 105.555 207.605 ;
        RECT 106.025 206.795 107.395 207.575 ;
        RECT 107.405 206.795 110.155 207.605 ;
        RECT 110.825 207.475 114.755 207.705 ;
        RECT 110.340 206.795 114.755 207.475 ;
        RECT 114.765 207.475 115.695 207.705 ;
        RECT 114.765 206.795 118.665 207.475 ;
        RECT 118.905 206.795 120.275 207.575 ;
        RECT 120.285 206.795 121.655 207.575 ;
        RECT 122.585 206.795 125.335 207.705 ;
        RECT 126.275 206.880 126.705 207.665 ;
        RECT 126.725 207.505 127.680 207.705 ;
        RECT 126.725 206.825 129.005 207.505 ;
        RECT 133.145 207.475 134.075 207.705 ;
        RECT 126.725 206.795 127.680 206.825 ;
        RECT 36.245 206.585 36.415 206.795 ;
        RECT 37.625 206.585 37.795 206.795 ;
        RECT 41.305 206.585 41.475 206.795 ;
        RECT 42.685 206.585 42.855 206.795 ;
        RECT 44.520 206.635 44.640 206.745 ;
        RECT 44.985 206.585 45.155 206.795 ;
        RECT 46.360 206.635 46.480 206.745 ;
        RECT 46.825 206.605 46.995 206.795 ;
        RECT 48.215 206.640 48.375 206.750 ;
        RECT 49.585 206.605 49.755 206.795 ;
        RECT 52.345 206.585 52.515 206.775 ;
        RECT 55.105 206.605 55.275 206.795 ;
        RECT 57.865 206.585 58.035 206.775 ;
        RECT 61.540 206.635 61.660 206.745 ;
        RECT 62.475 206.630 62.635 206.740 ;
        RECT 64.765 206.585 64.935 206.795 ;
        RECT 65.225 206.585 65.395 206.775 ;
        RECT 66.605 206.585 66.775 206.795 ;
        RECT 67.065 206.605 67.235 206.795 ;
        RECT 70.285 206.585 70.455 206.775 ;
        RECT 71.660 206.585 71.830 206.775 ;
        RECT 72.590 206.605 72.760 206.795 ;
        RECT 73.045 206.585 73.215 206.775 ;
        RECT 73.975 206.640 74.135 206.750 ;
        RECT 76.720 206.635 76.840 206.745 ;
        RECT 77.195 206.585 77.365 206.775 ;
        RECT 77.645 206.605 77.815 206.795 ;
        RECT 78.105 206.605 78.275 206.795 ;
        RECT 80.410 206.775 80.575 206.795 ;
        RECT 78.565 206.585 78.735 206.775 ;
        RECT 79.495 206.640 79.655 206.750 ;
        RECT 80.405 206.605 80.575 206.775 ;
        RECT 82.715 206.640 82.875 206.750 ;
        RECT 83.625 206.605 83.795 206.795 ;
        RECT 85.010 206.585 85.180 206.775 ;
        RECT 85.465 206.605 85.635 206.775 ;
        RECT 88.685 206.605 88.855 206.795 ;
        RECT 90.525 206.605 90.695 206.795 ;
        RECT 90.990 206.605 91.160 206.795 ;
        RECT 91.900 206.605 92.070 206.775 ;
        RECT 85.470 206.585 85.635 206.605 ;
        RECT 91.900 206.585 92.045 206.605 ;
        RECT 92.365 206.585 92.535 206.795 ;
        RECT 97.885 206.585 98.055 206.775 ;
        RECT 98.810 206.605 98.980 206.795 ;
        RECT 103.400 206.775 103.570 206.795 ;
        RECT 100.180 206.635 100.300 206.745 ;
        RECT 101.100 206.635 101.220 206.745 ;
        RECT 103.400 206.605 103.575 206.775 ;
        RECT 103.865 206.605 104.035 206.795 ;
        RECT 105.700 206.635 105.820 206.745 ;
        RECT 107.085 206.605 107.255 206.795 ;
        RECT 107.545 206.605 107.715 206.795 ;
        RECT 110.340 206.775 110.450 206.795 ;
        RECT 103.405 206.585 103.575 206.605 ;
        RECT 108.925 206.585 109.095 206.775 ;
        RECT 110.280 206.605 110.450 206.775 ;
        RECT 112.615 206.630 112.775 206.740 ;
        RECT 113.985 206.585 114.155 206.775 ;
        RECT 115.180 206.605 115.350 206.795 ;
        RECT 116.745 206.585 116.915 206.775 ;
        RECT 119.505 206.585 119.675 206.775 ;
        RECT 119.955 206.605 120.125 206.795 ;
        RECT 120.435 206.605 120.605 206.795 ;
        RECT 121.815 206.640 121.975 206.750 ;
        RECT 122.255 206.585 122.425 206.775 ;
        RECT 122.725 206.605 122.895 206.795 ;
        RECT 123.635 206.585 123.805 206.775 ;
        RECT 125.495 206.640 125.655 206.750 ;
        RECT 127.510 206.585 127.680 206.775 ;
        RECT 128.240 206.635 128.360 206.745 ;
        RECT 128.710 206.605 128.880 206.825 ;
        RECT 130.175 206.795 134.075 207.475 ;
        RECT 134.085 206.795 135.915 207.605 ;
        RECT 136.385 206.795 138.215 207.475 ;
        RECT 138.225 206.795 143.735 207.605 ;
        RECT 143.745 206.795 147.415 207.605 ;
        RECT 147.425 206.795 148.795 207.605 ;
        RECT 148.805 206.795 150.175 207.605 ;
        RECT 129.175 206.640 129.335 206.750 ;
        RECT 130.085 206.585 130.255 206.775 ;
        RECT 130.545 206.585 130.715 206.775 ;
        RECT 133.305 206.585 133.475 206.775 ;
        RECT 133.490 206.605 133.660 206.795 ;
        RECT 134.225 206.605 134.395 206.795 ;
        RECT 134.685 206.585 134.855 206.775 ;
        RECT 136.060 206.635 136.180 206.745 ;
        RECT 137.905 206.605 138.075 206.795 ;
        RECT 138.365 206.605 138.535 206.795 ;
        RECT 139.740 206.635 139.860 206.745 ;
        RECT 140.205 206.585 140.375 206.775 ;
        RECT 141.585 206.585 141.755 206.775 ;
        RECT 143.885 206.605 144.055 206.795 ;
        RECT 147.565 206.605 147.735 206.795 ;
        RECT 149.865 206.585 150.035 206.795 ;
        RECT 36.105 205.775 37.475 206.585 ;
        RECT 37.485 205.775 41.155 206.585 ;
        RECT 41.165 205.775 42.535 206.585 ;
        RECT 42.545 205.905 44.835 206.585 ;
        RECT 44.845 205.905 52.155 206.585 ;
        RECT 43.915 205.675 44.835 205.905 ;
        RECT 48.360 205.685 49.270 205.905 ;
        RECT 50.805 205.675 52.155 205.905 ;
        RECT 52.205 205.775 57.715 206.585 ;
        RECT 57.725 205.775 61.395 206.585 ;
        RECT 61.875 205.715 62.305 206.500 ;
        RECT 63.245 205.905 65.075 206.585 ;
        RECT 63.245 205.675 64.590 205.905 ;
        RECT 65.095 205.675 66.445 206.585 ;
        RECT 66.465 205.775 70.135 206.585 ;
        RECT 70.145 205.775 71.515 206.585 ;
        RECT 71.545 205.675 72.895 206.585 ;
        RECT 72.905 205.775 76.575 206.585 ;
        RECT 77.045 205.805 78.415 206.585 ;
        RECT 78.425 205.775 83.935 206.585 ;
        RECT 83.945 205.675 85.295 206.585 ;
        RECT 85.470 205.905 87.305 206.585 ;
        RECT 86.375 205.675 87.305 205.905 ;
        RECT 87.635 205.715 88.065 206.500 ;
        RECT 88.190 205.905 92.045 206.585 ;
        RECT 88.190 205.675 91.520 205.905 ;
        RECT 92.225 205.775 97.735 206.585 ;
        RECT 97.745 205.775 103.255 206.585 ;
        RECT 103.265 205.775 108.775 206.585 ;
        RECT 108.785 205.775 112.455 206.585 ;
        RECT 113.395 205.715 113.825 206.500 ;
        RECT 113.845 205.675 116.595 206.585 ;
        RECT 116.605 205.675 119.355 206.585 ;
        RECT 119.365 205.775 121.195 206.585 ;
        RECT 121.205 205.805 122.575 206.585 ;
        RECT 122.585 205.805 123.955 206.585 ;
        RECT 124.195 205.905 128.095 206.585 ;
        RECT 128.565 205.905 130.395 206.585 ;
        RECT 127.165 205.675 128.095 205.905 ;
        RECT 130.405 205.775 133.155 206.585 ;
        RECT 133.165 205.805 134.535 206.585 ;
        RECT 134.545 205.775 138.215 206.585 ;
        RECT 139.155 205.715 139.585 206.500 ;
        RECT 140.065 205.805 141.435 206.585 ;
        RECT 141.445 205.905 148.755 206.585 ;
        RECT 144.960 205.685 145.870 205.905 ;
        RECT 147.405 205.675 148.755 205.905 ;
        RECT 148.805 205.775 150.175 206.585 ;
      LAYER nwell ;
        RECT 35.910 202.555 150.370 205.385 ;
      LAYER pwell ;
        RECT 36.105 201.355 37.475 202.165 ;
        RECT 37.485 201.355 39.315 202.165 ;
        RECT 39.345 201.355 40.695 202.265 ;
        RECT 42.075 202.035 42.995 202.265 ;
        RECT 44.055 202.035 44.985 202.265 ;
        RECT 40.705 201.355 42.995 202.035 ;
        RECT 43.150 201.355 44.985 202.035 ;
        RECT 45.500 201.355 48.975 202.265 ;
        RECT 48.995 201.440 49.425 202.225 ;
        RECT 49.465 201.355 50.815 202.265 ;
        RECT 54.340 202.035 55.250 202.255 ;
        RECT 56.785 202.035 58.135 202.265 ;
        RECT 61.845 202.035 62.775 202.265 ;
        RECT 50.825 201.355 58.135 202.035 ;
        RECT 58.875 201.355 62.775 202.035 ;
        RECT 62.865 201.355 65.865 202.265 ;
        RECT 66.005 201.355 67.355 202.265 ;
        RECT 70.900 202.035 71.810 202.255 ;
        RECT 73.345 202.035 74.695 202.265 ;
        RECT 67.385 201.355 74.695 202.035 ;
        RECT 74.755 201.440 75.185 202.225 ;
        RECT 75.205 201.355 78.875 202.165 ;
        RECT 79.345 201.355 82.095 202.265 ;
        RECT 82.105 201.355 85.775 202.165 ;
        RECT 86.245 201.355 89.165 202.265 ;
        RECT 89.465 201.355 92.215 202.265 ;
        RECT 92.225 201.355 97.735 202.165 ;
        RECT 97.745 201.355 100.495 202.265 ;
        RECT 100.515 201.440 100.945 202.225 ;
        RECT 100.965 201.355 104.075 202.265 ;
        RECT 104.185 201.355 106.935 202.265 ;
        RECT 106.945 201.355 112.455 202.165 ;
        RECT 112.465 201.355 114.295 202.165 ;
        RECT 114.305 201.355 117.055 202.265 ;
        RECT 117.065 201.355 122.575 202.165 ;
        RECT 123.505 201.355 126.255 202.265 ;
        RECT 126.275 201.440 126.705 202.225 ;
        RECT 126.725 202.035 130.655 202.265 ;
        RECT 126.725 201.355 131.140 202.035 ;
        RECT 131.325 201.355 132.695 202.135 ;
        RECT 132.705 201.355 134.075 202.165 ;
        RECT 137.600 202.035 138.510 202.255 ;
        RECT 140.045 202.035 141.395 202.265 ;
        RECT 134.085 201.355 141.395 202.035 ;
        RECT 141.445 202.035 142.375 202.265 ;
        RECT 141.445 201.355 145.345 202.035 ;
        RECT 145.585 201.355 147.415 202.165 ;
        RECT 147.425 201.355 148.795 202.135 ;
        RECT 148.805 201.355 150.175 202.165 ;
        RECT 36.245 201.145 36.415 201.355 ;
        RECT 37.625 201.145 37.795 201.355 ;
        RECT 39.460 201.165 39.630 201.355 ;
        RECT 40.845 201.165 41.015 201.355 ;
        RECT 43.150 201.335 43.315 201.355 ;
        RECT 48.660 201.335 48.830 201.355 ;
        RECT 41.300 201.195 41.420 201.305 ;
        RECT 41.770 201.145 41.940 201.335 ;
        RECT 43.145 201.165 43.315 201.335 ;
        RECT 43.610 201.145 43.780 201.335 ;
        RECT 46.825 201.145 46.995 201.335 ;
        RECT 48.640 201.165 48.830 201.335 ;
        RECT 49.580 201.165 49.750 201.355 ;
        RECT 50.965 201.165 51.135 201.355 ;
        RECT 48.700 201.145 48.810 201.165 ;
        RECT 53.265 201.145 53.435 201.335 ;
        RECT 55.100 201.195 55.220 201.305 ;
        RECT 55.575 201.145 55.745 201.335 ;
        RECT 56.940 201.195 57.060 201.305 ;
        RECT 57.415 201.145 57.585 201.335 ;
        RECT 58.320 201.195 58.440 201.305 ;
        RECT 61.545 201.145 61.715 201.335 ;
        RECT 62.190 201.165 62.360 201.355 ;
        RECT 62.440 201.165 62.610 201.335 ;
        RECT 62.925 201.165 63.095 201.355 ;
        RECT 67.070 201.335 67.240 201.355 ;
        RECT 67.065 201.165 67.240 201.335 ;
        RECT 67.525 201.165 67.695 201.355 ;
        RECT 62.500 201.145 62.610 201.165 ;
        RECT 67.065 201.145 67.235 201.165 ;
        RECT 71.665 201.145 71.835 201.335 ;
        RECT 72.125 201.145 72.295 201.335 ;
        RECT 75.345 201.165 75.515 201.355 ;
        RECT 79.020 201.195 79.140 201.305 ;
        RECT 79.485 201.145 79.655 201.355 ;
        RECT 80.865 201.145 81.035 201.335 ;
        RECT 82.245 201.165 82.415 201.355 ;
        RECT 86.390 201.335 86.560 201.355 ;
        RECT 83.625 201.145 83.795 201.335 ;
        RECT 85.920 201.195 86.040 201.305 ;
        RECT 86.380 201.165 86.560 201.335 ;
        RECT 86.380 201.145 86.550 201.165 ;
        RECT 88.235 201.145 88.405 201.335 ;
        RECT 89.605 201.165 89.775 201.355 ;
        RECT 90.985 201.145 91.155 201.335 ;
        RECT 91.445 201.145 91.615 201.335 ;
        RECT 92.365 201.165 92.535 201.355 ;
        RECT 94.210 201.145 94.380 201.335 ;
        RECT 97.425 201.145 97.595 201.335 ;
        RECT 97.885 201.165 98.055 201.355 ;
        RECT 100.645 201.145 100.815 201.335 ;
        RECT 103.865 201.145 104.035 201.355 ;
        RECT 106.625 201.165 106.795 201.355 ;
        RECT 107.085 201.165 107.255 201.355 ;
        RECT 109.385 201.145 109.555 201.335 ;
        RECT 112.145 201.145 112.315 201.335 ;
        RECT 112.605 201.165 112.775 201.355 ;
        RECT 114.445 201.165 114.615 201.355 ;
        RECT 117.205 201.165 117.375 201.355 ;
        RECT 120.885 201.145 121.055 201.335 ;
        RECT 121.345 201.145 121.515 201.335 ;
        RECT 122.735 201.200 122.895 201.310 ;
        RECT 123.645 201.165 123.815 201.355 ;
        RECT 131.030 201.335 131.140 201.355 ;
        RECT 125.020 201.195 125.140 201.305 ;
        RECT 125.480 201.145 125.650 201.335 ;
        RECT 131.030 201.165 131.200 201.335 ;
        RECT 132.375 201.165 132.545 201.355 ;
        RECT 132.845 201.165 133.015 201.355 ;
        RECT 133.765 201.145 133.935 201.335 ;
        RECT 134.225 201.145 134.395 201.355 ;
        RECT 137.905 201.145 138.075 201.335 ;
        RECT 139.745 201.145 139.915 201.335 ;
        RECT 141.860 201.165 142.030 201.355 ;
        RECT 145.265 201.145 145.435 201.335 ;
        RECT 145.725 201.165 145.895 201.355 ;
        RECT 148.475 201.165 148.645 201.355 ;
        RECT 149.865 201.145 150.035 201.355 ;
        RECT 36.105 200.335 37.475 201.145 ;
        RECT 37.485 200.335 41.155 201.145 ;
        RECT 41.625 200.235 43.455 201.145 ;
        RECT 43.465 200.235 46.385 201.145 ;
        RECT 46.685 200.465 48.515 201.145 ;
        RECT 48.700 200.465 53.115 201.145 ;
        RECT 49.185 200.235 53.115 200.465 ;
        RECT 53.125 200.335 54.955 201.145 ;
        RECT 55.425 200.365 56.795 201.145 ;
        RECT 57.265 200.365 58.635 201.145 ;
        RECT 58.775 200.235 61.775 201.145 ;
        RECT 61.875 200.275 62.305 201.060 ;
        RECT 62.500 200.465 66.915 201.145 ;
        RECT 62.985 200.235 66.915 200.465 ;
        RECT 66.925 200.335 70.595 201.145 ;
        RECT 70.605 200.365 71.975 201.145 ;
        RECT 71.985 200.465 79.295 201.145 ;
        RECT 75.500 200.245 76.410 200.465 ;
        RECT 77.945 200.235 79.295 200.465 ;
        RECT 79.345 200.335 80.715 201.145 ;
        RECT 80.725 200.235 83.475 201.145 ;
        RECT 83.485 200.335 86.235 201.145 ;
        RECT 86.265 200.235 87.615 201.145 ;
        RECT 87.635 200.275 88.065 201.060 ;
        RECT 88.085 200.365 89.455 201.145 ;
        RECT 89.465 200.465 91.295 201.145 ;
        RECT 91.305 200.335 94.055 201.145 ;
        RECT 94.065 200.235 96.985 201.145 ;
        RECT 97.325 200.235 100.495 201.145 ;
        RECT 100.505 200.235 103.715 201.145 ;
        RECT 103.725 200.335 109.235 201.145 ;
        RECT 109.245 200.335 111.995 201.145 ;
        RECT 112.005 200.365 113.375 201.145 ;
        RECT 113.395 200.275 113.825 201.060 ;
        RECT 113.885 200.465 121.195 201.145 ;
        RECT 113.885 200.235 115.235 200.465 ;
        RECT 116.770 200.245 117.680 200.465 ;
        RECT 121.205 200.335 124.875 201.145 ;
        RECT 125.365 200.235 126.715 201.145 ;
        RECT 126.765 200.465 134.075 201.145 ;
        RECT 126.765 200.235 128.115 200.465 ;
        RECT 129.650 200.245 130.560 200.465 ;
        RECT 134.085 200.335 137.755 201.145 ;
        RECT 137.765 200.335 139.135 201.145 ;
        RECT 139.155 200.275 139.585 201.060 ;
        RECT 139.605 200.335 145.115 201.145 ;
        RECT 145.125 200.335 148.795 201.145 ;
        RECT 148.805 200.335 150.175 201.145 ;
      LAYER nwell ;
        RECT 35.910 197.115 150.370 199.945 ;
      LAYER pwell ;
        RECT 36.105 195.915 37.475 196.725 ;
        RECT 37.485 195.915 41.155 196.725 ;
        RECT 41.185 195.915 42.535 196.825 ;
        RECT 44.125 196.735 45.075 196.825 ;
        RECT 42.545 195.915 43.915 196.725 ;
        RECT 44.125 195.915 46.055 196.735 ;
        RECT 46.225 195.915 48.975 196.725 ;
        RECT 48.995 196.000 49.425 196.785 ;
        RECT 50.105 196.595 54.035 196.825 ;
        RECT 49.620 195.915 54.035 196.595 ;
        RECT 54.965 195.915 56.335 196.695 ;
        RECT 56.345 195.915 57.715 196.695 ;
        RECT 57.725 195.915 59.095 196.695 ;
        RECT 59.565 195.915 62.485 196.825 ;
        RECT 63.245 195.915 65.075 196.595 ;
        RECT 66.005 195.915 67.835 196.595 ;
        RECT 67.845 195.915 73.355 196.725 ;
        RECT 73.365 195.915 74.735 196.725 ;
        RECT 74.755 196.000 75.185 196.785 ;
        RECT 75.205 195.915 80.715 196.725 ;
        RECT 80.725 195.915 83.475 196.725 ;
        RECT 84.995 196.595 85.925 196.825 ;
        RECT 84.090 195.915 85.925 196.595 ;
        RECT 86.245 195.915 89.165 196.825 ;
        RECT 89.465 195.915 92.385 196.825 ;
        RECT 92.685 195.915 98.195 196.725 ;
        RECT 98.205 195.915 100.035 196.725 ;
        RECT 100.515 196.000 100.945 196.785 ;
        RECT 100.965 195.915 104.635 196.825 ;
        RECT 104.645 196.595 105.565 196.825 ;
        RECT 104.645 195.915 106.935 196.595 ;
        RECT 107.865 195.915 109.215 196.825 ;
        RECT 109.255 195.915 110.605 196.825 ;
        RECT 110.625 195.915 112.455 196.725 ;
        RECT 112.925 195.915 114.295 196.695 ;
        RECT 114.305 196.595 115.235 196.825 ;
        RECT 114.305 195.915 118.205 196.595 ;
        RECT 119.365 195.915 121.195 196.595 ;
        RECT 121.205 195.915 123.955 196.725 ;
        RECT 123.965 195.915 125.335 196.695 ;
        RECT 126.275 196.000 126.705 196.785 ;
        RECT 126.725 195.915 130.200 196.825 ;
        RECT 130.405 195.915 135.915 196.725 ;
        RECT 135.925 195.915 137.295 196.725 ;
        RECT 137.305 195.915 138.675 196.695 ;
        RECT 142.660 196.595 143.570 196.815 ;
        RECT 145.105 196.595 146.455 196.825 ;
        RECT 139.145 195.915 146.455 196.595 ;
        RECT 146.505 195.915 148.335 196.725 ;
        RECT 148.805 195.915 150.175 196.725 ;
        RECT 36.245 195.705 36.415 195.915 ;
        RECT 37.625 195.705 37.795 195.915 ;
        RECT 39.465 195.705 39.635 195.895 ;
        RECT 42.220 195.725 42.390 195.915 ;
        RECT 42.685 195.725 42.855 195.915 ;
        RECT 45.905 195.895 46.055 195.915 ;
        RECT 45.905 195.725 46.075 195.895 ;
        RECT 46.365 195.725 46.535 195.915 ;
        RECT 49.620 195.895 49.730 195.915 ;
        RECT 46.825 195.705 46.995 195.895 ;
        RECT 49.560 195.725 49.730 195.895 ;
        RECT 50.495 195.705 50.665 195.895 ;
        RECT 50.965 195.705 51.135 195.895 ;
        RECT 53.265 195.705 53.435 195.895 ;
        RECT 53.725 195.705 53.895 195.895 ;
        RECT 54.195 195.760 54.355 195.870 ;
        RECT 55.115 195.725 55.285 195.915 ;
        RECT 57.395 195.725 57.565 195.915 ;
        RECT 57.875 195.750 58.035 195.860 ;
        RECT 58.775 195.725 58.945 195.915 ;
        RECT 59.710 195.895 59.880 195.915 ;
        RECT 59.240 195.755 59.360 195.865 ;
        RECT 59.705 195.725 59.880 195.895 ;
        RECT 59.705 195.705 59.875 195.725 ;
        RECT 60.175 195.705 60.345 195.895 ;
        RECT 61.540 195.755 61.660 195.865 ;
        RECT 62.465 195.705 62.635 195.895 ;
        RECT 62.920 195.755 63.040 195.865 ;
        RECT 64.765 195.725 64.935 195.915 ;
        RECT 65.235 195.760 65.395 195.870 ;
        RECT 66.145 195.725 66.315 195.915 ;
        RECT 67.985 195.725 68.155 195.915 ;
        RECT 70.745 195.705 70.915 195.895 ;
        RECT 72.580 195.755 72.700 195.865 ;
        RECT 73.505 195.725 73.675 195.915 ;
        RECT 75.345 195.725 75.515 195.915 ;
        RECT 80.865 195.895 81.035 195.915 ;
        RECT 84.090 195.895 84.255 195.915 ;
        RECT 36.105 194.895 37.475 195.705 ;
        RECT 37.485 194.895 39.315 195.705 ;
        RECT 39.325 195.025 46.635 195.705 ;
        RECT 42.840 194.805 43.750 195.025 ;
        RECT 45.285 194.795 46.635 195.025 ;
        RECT 46.685 194.895 49.435 195.705 ;
        RECT 49.445 194.925 50.815 195.705 ;
        RECT 50.825 194.895 52.195 195.705 ;
        RECT 52.215 194.795 53.565 195.705 ;
        RECT 53.585 194.795 57.645 195.705 ;
        RECT 58.655 194.795 60.005 195.705 ;
        RECT 60.025 194.925 61.395 195.705 ;
        RECT 61.875 194.835 62.305 195.620 ;
        RECT 62.325 195.025 70.595 195.705 ;
        RECT 69.145 194.795 70.595 195.025 ;
        RECT 70.605 194.895 72.435 195.705 ;
        RECT 72.905 195.675 73.840 195.705 ;
        RECT 75.800 195.675 75.970 195.895 ;
        RECT 77.645 195.705 77.815 195.895 ;
        RECT 78.105 195.705 78.275 195.895 ;
        RECT 80.855 195.725 81.035 195.895 ;
        RECT 80.855 195.705 81.025 195.725 ;
        RECT 81.325 195.705 81.495 195.895 ;
        RECT 83.620 195.755 83.740 195.865 ;
        RECT 84.085 195.725 84.255 195.895 ;
        RECT 85.000 195.755 85.120 195.865 ;
        RECT 85.475 195.705 85.645 195.895 ;
        RECT 86.390 195.725 86.560 195.915 ;
        RECT 86.855 195.750 87.015 195.860 ;
        RECT 88.220 195.755 88.340 195.865 ;
        RECT 88.685 195.705 88.855 195.895 ;
        RECT 89.610 195.725 89.780 195.915 ;
        RECT 91.420 195.725 91.590 195.895 ;
        RECT 92.825 195.725 92.995 195.915 ;
        RECT 91.480 195.705 91.590 195.725 ;
        RECT 96.045 195.705 96.215 195.895 ;
        RECT 98.345 195.725 98.515 195.915 ;
        RECT 98.780 195.725 98.950 195.895 ;
        RECT 100.180 195.755 100.300 195.865 ;
        RECT 101.105 195.725 101.275 195.915 ;
        RECT 98.840 195.705 98.950 195.725 ;
        RECT 103.410 195.705 103.580 195.895 ;
        RECT 105.695 195.705 105.865 195.895 ;
        RECT 106.625 195.725 106.795 195.915 ;
        RECT 107.095 195.760 107.255 195.870 ;
        RECT 108.930 195.725 109.100 195.915 ;
        RECT 110.305 195.895 110.475 195.915 ;
        RECT 110.305 195.725 110.500 195.895 ;
        RECT 110.765 195.725 110.935 195.915 ;
        RECT 112.605 195.865 112.775 195.895 ;
        RECT 113.075 195.865 113.245 195.915 ;
        RECT 112.600 195.755 112.775 195.865 ;
        RECT 113.060 195.755 113.245 195.865 ;
        RECT 112.605 195.725 112.775 195.755 ;
        RECT 113.075 195.725 113.245 195.755 ;
        RECT 110.330 195.705 110.440 195.725 ;
        RECT 112.605 195.705 112.770 195.725 ;
        RECT 113.985 195.705 114.155 195.895 ;
        RECT 114.720 195.725 114.890 195.915 ;
        RECT 115.365 195.705 115.535 195.895 ;
        RECT 118.595 195.760 118.755 195.870 ;
        RECT 119.505 195.725 119.675 195.915 ;
        RECT 121.345 195.895 121.515 195.915 ;
        RECT 121.345 195.725 121.540 195.895 ;
        RECT 121.800 195.755 121.920 195.865 ;
        RECT 124.115 195.725 124.285 195.915 ;
        RECT 121.370 195.705 121.480 195.725 ;
        RECT 125.020 195.705 125.190 195.895 ;
        RECT 125.495 195.760 125.655 195.870 ;
        RECT 126.870 195.725 127.040 195.915 ;
        RECT 127.785 195.705 127.955 195.895 ;
        RECT 128.245 195.705 128.415 195.895 ;
        RECT 130.545 195.725 130.715 195.915 ;
        RECT 131.935 195.750 132.095 195.860 ;
        RECT 136.065 195.725 136.235 195.915 ;
        RECT 136.250 195.705 136.420 195.895 ;
        RECT 136.985 195.725 137.155 195.895 ;
        RECT 137.445 195.725 137.615 195.915 ;
        RECT 138.820 195.755 138.940 195.865 ;
        RECT 139.285 195.725 139.455 195.915 ;
        RECT 137.005 195.705 137.155 195.725 ;
        RECT 139.745 195.705 139.915 195.895 ;
        RECT 146.645 195.725 146.815 195.915 ;
        RECT 147.105 195.705 147.275 195.895 ;
        RECT 148.480 195.755 148.600 195.865 ;
        RECT 149.865 195.705 150.035 195.915 ;
        RECT 72.905 195.475 75.970 195.675 ;
        RECT 72.905 194.995 76.115 195.475 ;
        RECT 72.905 194.795 73.855 194.995 ;
        RECT 75.185 194.795 76.115 194.995 ;
        RECT 76.125 194.795 77.940 195.705 ;
        RECT 77.965 194.895 79.795 195.705 ;
        RECT 79.805 194.925 81.175 195.705 ;
        RECT 81.185 194.895 84.855 195.705 ;
        RECT 85.325 194.925 86.695 195.705 ;
        RECT 87.635 194.835 88.065 195.620 ;
        RECT 88.545 194.795 91.295 195.705 ;
        RECT 91.480 195.025 95.895 195.705 ;
        RECT 91.965 194.795 95.895 195.025 ;
        RECT 95.905 194.895 98.655 195.705 ;
        RECT 98.840 195.025 103.255 195.705 ;
        RECT 99.325 194.795 103.255 195.025 ;
        RECT 103.265 194.795 104.615 195.705 ;
        RECT 104.645 194.925 106.015 195.705 ;
        RECT 106.025 195.025 110.440 195.705 ;
        RECT 110.935 195.025 112.770 195.705 ;
        RECT 106.025 194.795 109.955 195.025 ;
        RECT 110.935 194.795 111.865 195.025 ;
        RECT 113.395 194.835 113.825 195.620 ;
        RECT 113.855 194.795 115.205 195.705 ;
        RECT 115.225 194.895 117.055 195.705 ;
        RECT 117.065 195.025 121.480 195.705 ;
        RECT 117.065 194.795 120.995 195.025 ;
        RECT 122.415 194.795 125.335 195.705 ;
        RECT 125.355 194.795 128.085 195.705 ;
        RECT 128.105 194.895 131.775 195.705 ;
        RECT 132.935 195.025 136.835 195.705 ;
        RECT 135.905 194.795 136.835 195.025 ;
        RECT 137.005 194.885 138.935 195.705 ;
        RECT 137.985 194.795 138.935 194.885 ;
        RECT 139.155 194.835 139.585 195.620 ;
        RECT 139.605 195.025 146.915 195.705 ;
        RECT 143.120 194.805 144.030 195.025 ;
        RECT 145.565 194.795 146.915 195.025 ;
        RECT 146.965 194.895 148.795 195.705 ;
        RECT 148.805 194.895 150.175 195.705 ;
      LAYER nwell ;
        RECT 35.910 191.675 150.370 194.505 ;
      LAYER pwell ;
        RECT 36.105 190.475 37.475 191.285 ;
        RECT 37.485 190.475 41.155 191.285 ;
        RECT 42.085 190.475 43.915 191.385 ;
        RECT 43.925 190.475 47.595 191.285 ;
        RECT 47.605 190.475 48.975 191.285 ;
        RECT 48.995 190.560 49.425 191.345 ;
        RECT 49.445 190.475 51.275 191.285 ;
        RECT 51.750 191.155 53.130 191.385 ;
        RECT 54.920 191.155 56.295 191.385 ;
        RECT 51.750 190.705 56.295 191.155 ;
        RECT 51.750 190.475 54.910 190.705 ;
        RECT 36.245 190.265 36.415 190.475 ;
        RECT 37.625 190.265 37.795 190.475 ;
        RECT 41.295 190.430 41.465 190.455 ;
        RECT 41.295 190.320 41.475 190.430 ;
        RECT 41.295 190.265 41.465 190.320 ;
        RECT 41.775 190.265 41.945 190.455 ;
        RECT 43.145 190.265 43.315 190.455 ;
        RECT 43.600 190.285 43.770 190.475 ;
        RECT 44.065 190.285 44.235 190.475 ;
        RECT 44.990 190.265 45.160 190.455 ;
        RECT 47.745 190.285 47.915 190.475 ;
        RECT 49.585 190.285 49.755 190.475 ;
        RECT 50.505 190.265 50.675 190.455 ;
        RECT 50.965 190.265 51.135 190.455 ;
        RECT 51.420 190.315 51.540 190.425 ;
        RECT 56.020 190.285 56.190 190.705 ;
        RECT 56.345 190.475 60.015 191.385 ;
        RECT 60.485 190.475 61.855 191.255 ;
        RECT 61.865 191.155 65.795 191.385 ;
        RECT 61.865 190.475 66.280 191.155 ;
        RECT 66.465 190.475 68.295 191.155 ;
        RECT 68.305 190.475 73.815 191.285 ;
        RECT 74.755 190.560 75.185 191.345 ;
        RECT 75.215 190.475 77.945 191.385 ;
        RECT 77.965 190.475 79.795 191.385 ;
        RECT 79.805 190.475 81.175 191.255 ;
        RECT 81.185 190.475 86.695 191.285 ;
        RECT 87.950 190.475 91.605 191.385 ;
        RECT 91.765 190.475 94.515 191.385 ;
        RECT 95.445 190.475 96.815 191.255 ;
        RECT 96.825 190.475 100.300 191.385 ;
        RECT 100.515 190.560 100.945 191.345 ;
        RECT 101.290 190.475 104.945 191.385 ;
        RECT 105.105 191.155 106.030 191.385 ;
        RECT 105.105 190.475 108.775 191.155 ;
        RECT 108.805 190.475 110.155 191.385 ;
        RECT 110.825 191.155 114.755 191.385 ;
        RECT 110.340 190.475 114.755 191.155 ;
        RECT 114.845 190.475 117.845 191.385 ;
        RECT 118.905 190.475 120.275 191.255 ;
        RECT 120.285 190.475 121.655 191.255 ;
        RECT 121.665 190.475 125.335 191.285 ;
        RECT 126.275 190.560 126.705 191.345 ;
        RECT 127.645 190.475 129.015 191.255 ;
        RECT 129.035 190.475 131.765 191.385 ;
        RECT 131.785 191.155 132.705 191.385 ;
        RECT 131.785 190.475 134.075 191.155 ;
        RECT 134.095 190.475 135.445 191.385 ;
        RECT 135.465 190.475 136.835 191.285 ;
        RECT 136.845 190.475 138.215 191.255 ;
        RECT 138.225 191.155 142.155 191.385 ;
        RECT 138.225 190.475 142.640 191.155 ;
        RECT 142.825 190.475 144.655 191.385 ;
        RECT 144.665 190.475 148.335 191.285 ;
        RECT 148.805 190.475 150.175 191.285 ;
        RECT 56.490 190.455 56.660 190.475 ;
        RECT 56.480 190.285 56.660 190.455 ;
        RECT 56.480 190.265 56.650 190.285 ;
        RECT 57.865 190.265 58.035 190.455 ;
        RECT 60.175 190.425 60.345 190.455 ;
        RECT 59.700 190.315 59.820 190.425 ;
        RECT 60.160 190.315 60.345 190.425 ;
        RECT 60.175 190.265 60.345 190.315 ;
        RECT 61.535 190.285 61.705 190.475 ;
        RECT 66.170 190.455 66.280 190.475 ;
        RECT 62.465 190.265 62.635 190.455 ;
        RECT 66.170 190.285 66.340 190.455 ;
        RECT 67.985 190.285 68.155 190.475 ;
        RECT 68.445 190.285 68.615 190.475 ;
        RECT 72.585 190.265 72.755 190.455 ;
        RECT 73.045 190.265 73.215 190.455 ;
        RECT 73.975 190.320 74.135 190.430 ;
        RECT 75.345 190.285 75.515 190.475 ;
        RECT 79.480 190.455 79.650 190.475 ;
        RECT 76.265 190.265 76.435 190.455 ;
        RECT 76.730 190.265 76.900 190.455 ;
        RECT 79.475 190.285 79.650 190.455 ;
        RECT 79.475 190.265 79.645 190.285 ;
        RECT 79.945 190.265 80.115 190.455 ;
        RECT 80.855 190.285 81.025 190.475 ;
        RECT 81.325 190.285 81.495 190.475 ;
        RECT 91.445 190.455 91.605 190.475 ;
        RECT 83.635 190.310 83.795 190.420 ;
        RECT 86.855 190.320 87.015 190.430 ;
        RECT 87.305 190.265 87.475 190.455 ;
        RECT 91.440 190.285 91.615 190.455 ;
        RECT 91.440 190.265 91.610 190.285 ;
        RECT 91.905 190.265 92.075 190.475 ;
        RECT 94.675 190.320 94.835 190.430 ;
        RECT 96.495 190.285 96.665 190.475 ;
        RECT 96.970 190.285 97.140 190.475 ;
        RECT 104.785 190.455 104.945 190.475 ;
        RECT 97.425 190.265 97.595 190.455 ;
        RECT 98.805 190.265 98.975 190.455 ;
        RECT 100.640 190.265 100.810 190.455 ;
        RECT 102.025 190.265 102.195 190.455 ;
        RECT 104.785 190.285 104.955 190.455 ;
        RECT 105.250 190.285 105.420 190.475 ;
        RECT 105.715 190.310 105.875 190.420 ;
        RECT 107.535 190.265 107.705 190.455 ;
        RECT 108.005 190.265 108.175 190.455 ;
        RECT 108.920 190.285 109.090 190.475 ;
        RECT 110.340 190.455 110.450 190.475 ;
        RECT 110.280 190.285 110.450 190.455 ;
        RECT 113.985 190.265 114.155 190.455 ;
        RECT 114.905 190.285 115.075 190.475 ;
        RECT 116.750 190.265 116.920 190.455 ;
        RECT 118.135 190.320 118.295 190.430 ;
        RECT 119.055 190.285 119.225 190.475 ;
        RECT 120.435 190.425 120.605 190.475 ;
        RECT 120.420 190.315 120.605 190.425 ;
        RECT 120.435 190.285 120.605 190.315 ;
        RECT 120.885 190.265 121.055 190.455 ;
        RECT 121.805 190.285 121.975 190.475 ;
        RECT 125.495 190.320 125.655 190.430 ;
        RECT 126.875 190.320 127.035 190.430 ;
        RECT 128.695 190.285 128.865 190.475 ;
        RECT 131.465 190.265 131.635 190.475 ;
        RECT 131.925 190.265 132.095 190.455 ;
        RECT 133.765 190.285 133.935 190.475 ;
        RECT 134.225 190.285 134.395 190.475 ;
        RECT 134.685 190.285 134.855 190.455 ;
        RECT 135.605 190.285 135.775 190.475 ;
        RECT 134.705 190.265 134.855 190.285 ;
        RECT 136.985 190.265 137.155 190.475 ;
        RECT 142.530 190.455 142.640 190.475 ;
        RECT 138.820 190.315 138.940 190.425 ;
        RECT 139.745 190.265 139.915 190.455 ;
        RECT 141.130 190.265 141.300 190.455 ;
        RECT 142.530 190.285 142.700 190.455 ;
        RECT 142.970 190.285 143.140 190.475 ;
        RECT 144.805 190.285 144.975 190.475 ;
        RECT 146.185 190.285 146.355 190.455 ;
        RECT 146.185 190.265 146.335 190.285 ;
        RECT 146.645 190.265 146.815 190.455 ;
        RECT 148.480 190.315 148.600 190.425 ;
        RECT 149.865 190.265 150.035 190.475 ;
        RECT 36.105 189.455 37.475 190.265 ;
        RECT 37.485 189.455 40.235 190.265 ;
        RECT 40.245 189.485 41.615 190.265 ;
        RECT 41.625 189.485 42.995 190.265 ;
        RECT 43.020 189.355 44.835 190.265 ;
        RECT 44.845 189.355 48.515 190.265 ;
        RECT 48.525 189.585 50.815 190.265 ;
        RECT 48.525 189.355 49.445 189.585 ;
        RECT 50.825 189.455 56.335 190.265 ;
        RECT 56.365 189.355 57.715 190.265 ;
        RECT 57.725 189.455 59.555 190.265 ;
        RECT 60.025 189.485 61.395 190.265 ;
        RECT 61.875 189.395 62.305 190.180 ;
        RECT 62.325 189.455 63.695 190.265 ;
        RECT 63.790 189.585 72.895 190.265 ;
        RECT 72.905 189.455 74.275 190.265 ;
        RECT 74.285 189.585 76.575 190.265 ;
        RECT 74.285 189.355 75.205 189.585 ;
        RECT 76.585 189.355 78.415 190.265 ;
        RECT 78.425 189.485 79.795 190.265 ;
        RECT 79.805 189.455 83.475 190.265 ;
        RECT 84.405 189.355 87.615 190.265 ;
        RECT 87.635 189.395 88.065 190.180 ;
        RECT 88.280 189.355 91.755 190.265 ;
        RECT 91.765 189.455 97.275 190.265 ;
        RECT 97.285 189.455 98.655 190.265 ;
        RECT 98.680 189.355 100.495 190.265 ;
        RECT 100.525 189.355 101.875 190.265 ;
        RECT 101.885 189.455 105.555 190.265 ;
        RECT 106.485 189.485 107.855 190.265 ;
        RECT 107.865 189.455 113.375 190.265 ;
        RECT 113.395 189.395 113.825 190.180 ;
        RECT 113.845 189.455 116.595 190.265 ;
        RECT 116.605 189.355 120.275 190.265 ;
        RECT 120.745 189.585 129.850 190.265 ;
        RECT 129.945 189.585 131.775 190.265 ;
        RECT 131.785 189.455 134.535 190.265 ;
        RECT 134.705 189.445 136.635 190.265 ;
        RECT 136.845 189.455 138.675 190.265 ;
        RECT 135.685 189.355 136.635 189.445 ;
        RECT 139.155 189.395 139.585 190.180 ;
        RECT 139.615 189.355 140.965 190.265 ;
        RECT 140.985 189.355 143.905 190.265 ;
        RECT 144.405 189.445 146.335 190.265 ;
        RECT 146.505 189.455 148.335 190.265 ;
        RECT 148.805 189.455 150.175 190.265 ;
        RECT 144.405 189.355 145.355 189.445 ;
      LAYER nwell ;
        RECT 35.910 186.235 150.370 189.065 ;
      LAYER pwell ;
        RECT 36.105 185.035 37.475 185.845 ;
        RECT 37.485 185.035 42.995 185.845 ;
        RECT 43.005 185.035 45.755 185.845 ;
        RECT 45.845 185.035 48.845 185.945 ;
        RECT 48.995 185.120 49.425 185.905 ;
        RECT 49.445 185.745 50.390 185.945 ;
        RECT 49.445 185.065 52.195 185.745 ;
        RECT 49.445 185.035 50.390 185.065 ;
        RECT 36.245 184.825 36.415 185.035 ;
        RECT 37.625 184.825 37.795 185.035 ;
        RECT 43.145 185.015 43.315 185.035 ;
        RECT 43.145 184.845 43.320 185.015 ;
        RECT 44.985 184.845 45.155 185.015 ;
        RECT 45.905 184.845 46.075 185.035 ;
        RECT 43.150 184.825 43.320 184.845 ;
        RECT 44.990 184.825 45.155 184.845 ;
        RECT 36.105 184.015 37.475 184.825 ;
        RECT 37.485 184.015 42.995 184.825 ;
        RECT 43.005 183.915 44.835 184.825 ;
        RECT 44.990 184.145 46.825 184.825 ;
        RECT 45.895 183.915 46.825 184.145 ;
        RECT 47.145 184.795 48.090 184.825 ;
        RECT 49.580 184.795 49.750 185.015 ;
        RECT 50.055 184.870 50.215 184.980 ;
        RECT 50.960 184.795 51.130 185.015 ;
        RECT 51.880 184.845 52.050 185.065 ;
        RECT 52.205 185.035 57.715 185.845 ;
        RECT 58.015 185.035 60.935 185.945 ;
        RECT 67.765 185.715 69.215 185.945 ;
        RECT 60.945 185.035 69.215 185.715 ;
        RECT 69.225 185.035 72.895 185.845 ;
        RECT 72.905 185.035 74.720 185.945 ;
        RECT 74.755 185.120 75.185 185.905 ;
        RECT 78.720 185.715 79.630 185.935 ;
        RECT 81.165 185.715 82.515 185.945 ;
        RECT 75.205 185.035 82.515 185.715 ;
        RECT 82.565 185.035 86.235 185.845 ;
        RECT 86.245 185.035 87.615 185.845 ;
        RECT 87.625 185.035 88.995 185.815 ;
        RECT 89.005 185.035 94.515 185.845 ;
        RECT 95.185 185.715 99.115 185.945 ;
        RECT 94.700 185.035 99.115 185.715 ;
        RECT 99.125 185.035 100.495 185.845 ;
        RECT 100.515 185.120 100.945 185.905 ;
        RECT 101.625 185.715 105.555 185.945 ;
        RECT 101.140 185.035 105.555 185.715 ;
        RECT 105.565 185.715 109.495 185.945 ;
        RECT 110.825 185.715 114.755 185.945 ;
        RECT 105.565 185.035 109.980 185.715 ;
        RECT 52.345 184.845 52.515 185.035 ;
        RECT 60.620 185.015 60.790 185.035 ;
        RECT 52.160 184.795 53.115 184.825 ;
        RECT 53.260 184.795 53.430 185.015 ;
        RECT 55.565 184.825 55.735 185.015 ;
        RECT 58.325 184.845 58.495 185.015 ;
        RECT 60.620 184.845 60.795 185.015 ;
        RECT 61.085 184.845 61.255 185.035 ;
        RECT 62.475 184.870 62.635 184.980 ;
        RECT 58.330 184.825 58.495 184.845 ;
        RECT 60.625 184.825 60.795 184.845 ;
        RECT 64.295 184.825 64.465 185.015 ;
        RECT 64.765 184.825 64.935 185.015 ;
        RECT 69.365 184.845 69.535 185.035 ;
        RECT 70.285 184.825 70.455 185.015 ;
        RECT 74.425 184.845 74.595 185.035 ;
        RECT 75.345 184.845 75.515 185.035 ;
        RECT 75.805 184.825 75.975 185.015 ;
        RECT 77.655 184.825 77.825 185.015 ;
        RECT 79.025 184.825 79.195 185.015 ;
        RECT 82.705 184.845 82.875 185.035 ;
        RECT 83.625 184.845 83.795 185.015 ;
        RECT 83.625 184.825 83.775 184.845 ;
        RECT 85.005 184.825 85.175 185.015 ;
        RECT 85.465 184.825 85.635 185.015 ;
        RECT 86.385 184.845 86.555 185.035 ;
        RECT 87.300 184.875 87.420 184.985 ;
        RECT 88.675 184.845 88.845 185.035 ;
        RECT 89.145 184.845 89.315 185.035 ;
        RECT 94.700 185.015 94.810 185.035 ;
        RECT 91.440 184.825 91.610 185.015 ;
        RECT 91.905 184.825 92.075 185.015 ;
        RECT 94.640 184.845 94.810 185.015 ;
        RECT 96.035 184.825 96.205 185.015 ;
        RECT 96.505 184.845 96.675 185.015 ;
        RECT 99.265 184.845 99.435 185.035 ;
        RECT 101.140 185.015 101.250 185.035 ;
        RECT 109.870 185.015 109.980 185.035 ;
        RECT 110.340 185.035 114.755 185.715 ;
        RECT 114.765 185.035 119.295 185.945 ;
        RECT 120.285 185.715 121.420 185.945 ;
        RECT 124.555 185.715 125.485 185.945 ;
        RECT 120.285 185.035 123.495 185.715 ;
        RECT 123.650 185.035 125.485 185.715 ;
        RECT 126.275 185.120 126.705 185.905 ;
        RECT 128.095 185.715 129.015 185.945 ;
        RECT 126.725 185.035 129.015 185.715 ;
        RECT 129.225 185.855 130.175 185.945 ;
        RECT 129.225 185.035 131.155 185.855 ;
        RECT 132.695 185.715 133.615 185.945 ;
        RECT 131.325 185.035 133.615 185.715 ;
        RECT 133.625 185.035 134.995 185.815 ;
        RECT 135.005 185.035 136.835 185.845 ;
        RECT 136.845 185.035 140.905 185.945 ;
        RECT 141.055 185.035 145.115 185.945 ;
        RECT 145.125 185.715 146.045 185.945 ;
        RECT 145.125 185.035 147.415 185.715 ;
        RECT 147.425 185.035 148.795 185.845 ;
        RECT 148.805 185.035 150.175 185.845 ;
        RECT 110.340 185.015 110.450 185.035 ;
        RECT 101.080 184.845 101.250 185.015 ;
        RECT 104.325 184.845 104.495 185.015 ;
        RECT 96.515 184.825 96.675 184.845 ;
        RECT 104.325 184.825 104.485 184.845 ;
        RECT 105.695 184.825 105.865 185.015 ;
        RECT 106.175 184.870 106.335 184.980 ;
        RECT 107.080 184.825 107.250 185.015 ;
        RECT 108.440 184.845 108.610 185.015 ;
        RECT 109.870 184.845 110.040 185.015 ;
        RECT 110.280 184.845 110.450 185.015 ;
        RECT 113.060 184.875 113.180 184.985 ;
        RECT 108.500 184.825 108.610 184.845 ;
        RECT 113.985 184.825 114.155 185.015 ;
        RECT 114.910 184.845 115.080 185.035 ;
        RECT 115.825 184.825 115.995 185.015 ;
        RECT 117.215 184.825 117.385 185.015 ;
        RECT 54.460 184.795 55.415 184.825 ;
        RECT 47.145 184.115 49.895 184.795 ;
        RECT 50.835 184.115 53.115 184.795 ;
        RECT 53.135 184.115 55.415 184.795 ;
        RECT 47.145 183.915 48.090 184.115 ;
        RECT 52.160 183.915 53.115 184.115 ;
        RECT 54.460 183.915 55.415 184.115 ;
        RECT 55.425 184.015 58.175 184.825 ;
        RECT 58.330 184.145 60.165 184.825 ;
        RECT 59.235 183.915 60.165 184.145 ;
        RECT 60.485 184.015 61.855 184.825 ;
        RECT 61.875 183.955 62.305 184.740 ;
        RECT 63.245 184.045 64.615 184.825 ;
        RECT 64.625 184.015 70.135 184.825 ;
        RECT 70.145 184.015 75.655 184.825 ;
        RECT 75.665 184.015 77.495 184.825 ;
        RECT 77.505 184.045 78.875 184.825 ;
        RECT 78.895 183.915 81.625 184.825 ;
        RECT 81.845 184.005 83.775 184.825 ;
        RECT 81.845 183.915 82.795 184.005 ;
        RECT 83.955 183.915 85.305 184.825 ;
        RECT 85.325 184.015 87.155 184.825 ;
        RECT 87.635 183.955 88.065 184.740 ;
        RECT 88.280 183.915 91.755 184.825 ;
        RECT 91.765 183.915 94.975 184.825 ;
        RECT 94.985 184.045 96.355 184.825 ;
        RECT 96.515 183.915 100.170 184.825 ;
        RECT 100.830 183.915 104.485 184.825 ;
        RECT 104.645 184.045 106.015 184.825 ;
        RECT 106.965 183.915 108.315 184.825 ;
        RECT 108.500 184.145 112.915 184.825 ;
        RECT 108.985 183.915 112.915 184.145 ;
        RECT 113.395 183.955 113.825 184.740 ;
        RECT 113.845 184.145 115.675 184.825 ;
        RECT 115.685 184.015 117.055 184.825 ;
        RECT 117.065 184.045 118.435 184.825 ;
        RECT 118.585 184.795 118.755 185.015 ;
        RECT 119.515 184.880 119.675 184.990 ;
        RECT 121.805 184.825 121.975 185.015 ;
        RECT 123.185 184.845 123.355 185.035 ;
        RECT 123.650 185.015 123.815 185.035 ;
        RECT 123.645 184.845 123.815 185.015 ;
        RECT 124.115 184.870 124.275 184.980 ;
        RECT 125.035 184.825 125.205 185.015 ;
        RECT 125.940 184.875 126.060 184.985 ;
        RECT 126.400 184.875 126.520 184.985 ;
        RECT 126.865 184.825 127.035 185.035 ;
        RECT 131.005 185.015 131.155 185.035 ;
        RECT 129.615 184.825 129.785 185.015 ;
        RECT 130.085 184.825 130.255 185.015 ;
        RECT 131.005 184.845 131.175 185.015 ;
        RECT 131.465 184.845 131.635 185.035 ;
        RECT 132.380 184.825 132.550 185.015 ;
        RECT 132.845 184.825 133.015 185.015 ;
        RECT 133.775 184.845 133.945 185.035 ;
        RECT 135.145 185.015 135.315 185.035 ;
        RECT 135.135 184.845 135.315 185.015 ;
        RECT 135.135 184.825 135.305 184.845 ;
        RECT 135.605 184.825 135.775 185.015 ;
        RECT 136.985 184.845 137.155 185.035 ;
        RECT 142.505 184.825 142.675 185.015 ;
        RECT 143.875 184.825 144.045 185.015 ;
        RECT 144.345 184.825 144.515 185.015 ;
        RECT 144.805 184.845 144.975 185.035 ;
        RECT 147.105 184.845 147.275 185.035 ;
        RECT 147.565 184.845 147.735 185.035 ;
        RECT 148.035 184.870 148.195 184.980 ;
        RECT 149.865 184.825 150.035 185.035 ;
        RECT 120.710 184.795 121.655 184.825 ;
        RECT 118.585 184.595 121.655 184.795 ;
        RECT 118.445 184.115 121.655 184.595 ;
        RECT 121.665 184.145 123.955 184.825 ;
        RECT 118.445 183.915 119.375 184.115 ;
        RECT 120.710 183.915 121.655 184.115 ;
        RECT 123.035 183.915 123.955 184.145 ;
        RECT 124.885 184.045 126.255 184.825 ;
        RECT 126.725 184.145 128.555 184.825 ;
        RECT 128.565 184.045 129.935 184.825 ;
        RECT 129.945 184.015 131.315 184.825 ;
        RECT 131.345 183.915 132.695 184.825 ;
        RECT 132.715 183.915 134.065 184.825 ;
        RECT 134.085 184.045 135.455 184.825 ;
        RECT 135.465 184.015 139.135 184.825 ;
        RECT 139.155 183.955 139.585 184.740 ;
        RECT 139.735 183.915 142.735 184.825 ;
        RECT 142.825 184.045 144.195 184.825 ;
        RECT 144.205 184.015 147.875 184.825 ;
        RECT 148.805 184.015 150.175 184.825 ;
      LAYER nwell ;
        RECT 35.910 180.795 150.370 183.625 ;
      LAYER pwell ;
        RECT 36.105 179.595 37.475 180.405 ;
        RECT 37.485 179.595 42.995 180.405 ;
        RECT 43.005 179.595 44.375 180.405 ;
        RECT 44.385 179.595 45.755 180.375 ;
        RECT 45.765 179.595 47.135 180.375 ;
        RECT 47.145 179.595 48.975 180.505 ;
        RECT 48.995 179.680 49.425 180.465 ;
        RECT 51.250 180.305 52.195 180.505 ;
        RECT 49.445 179.625 52.195 180.305 ;
        RECT 36.245 179.385 36.415 179.595 ;
        RECT 37.625 179.385 37.795 179.595 ;
        RECT 43.145 179.405 43.315 179.595 ;
        RECT 44.535 179.405 44.705 179.595 ;
        RECT 44.985 179.385 45.155 179.575 ;
        RECT 45.915 179.405 46.085 179.595 ;
        RECT 46.820 179.435 46.940 179.545 ;
        RECT 36.105 178.575 37.475 179.385 ;
        RECT 37.485 178.705 44.795 179.385 ;
        RECT 41.000 178.485 41.910 178.705 ;
        RECT 43.445 178.475 44.795 178.705 ;
        RECT 44.845 178.575 46.675 179.385 ;
        RECT 47.290 179.355 47.460 179.595 ;
        RECT 49.590 179.405 49.760 179.625 ;
        RECT 51.250 179.595 52.195 179.625 ;
        RECT 52.205 179.595 55.875 180.405 ;
        RECT 56.805 179.595 58.175 180.375 ;
        RECT 58.185 179.595 61.855 180.405 ;
        RECT 68.685 180.275 70.135 180.505 ;
        RECT 61.865 179.595 70.135 180.275 ;
        RECT 70.145 179.595 73.815 180.405 ;
        RECT 74.755 179.680 75.185 180.465 ;
        RECT 75.205 179.595 81.025 180.505 ;
        RECT 81.185 179.595 86.695 180.405 ;
        RECT 86.705 179.595 88.075 180.405 ;
        RECT 88.085 179.595 91.295 180.505 ;
        RECT 91.305 179.595 94.055 180.505 ;
        RECT 94.065 179.595 95.435 180.375 ;
        RECT 95.445 179.595 97.275 180.405 ;
        RECT 97.745 179.595 100.495 180.505 ;
        RECT 100.515 179.680 100.945 180.465 ;
        RECT 100.965 179.595 104.635 180.405 ;
        RECT 104.645 180.275 108.575 180.505 ;
        RECT 104.645 179.595 109.060 180.275 ;
        RECT 109.245 179.595 111.995 180.505 ;
        RECT 112.005 179.595 113.375 180.375 ;
        RECT 113.385 179.595 114.755 180.375 ;
        RECT 114.765 179.595 116.135 180.375 ;
        RECT 116.145 179.595 117.515 180.375 ;
        RECT 119.330 180.305 120.275 180.505 ;
        RECT 117.525 179.625 120.275 180.305 ;
        RECT 51.885 179.385 52.055 179.575 ;
        RECT 52.345 179.545 52.515 179.595 ;
        RECT 52.340 179.435 52.515 179.545 ;
        RECT 52.345 179.405 52.515 179.435 ;
        RECT 53.715 179.385 53.885 179.575 ;
        RECT 54.185 179.385 54.355 179.575 ;
        RECT 56.035 179.440 56.195 179.550 ;
        RECT 56.955 179.405 57.125 179.595 ;
        RECT 58.325 179.575 58.495 179.595 ;
        RECT 57.860 179.435 57.980 179.545 ;
        RECT 58.325 179.405 58.505 179.575 ;
        RECT 58.335 179.385 58.505 179.405 ;
        RECT 59.715 179.385 59.885 179.575 ;
        RECT 61.095 179.430 61.255 179.540 ;
        RECT 62.005 179.405 62.175 179.595 ;
        RECT 62.465 179.385 62.635 179.575 ;
        RECT 70.285 179.405 70.455 179.595 ;
        RECT 70.745 179.385 70.915 179.575 ;
        RECT 73.975 179.440 74.135 179.550 ;
        RECT 75.345 179.405 75.515 179.595 ;
        RECT 76.275 179.430 76.435 179.540 ;
        RECT 81.325 179.405 81.495 179.595 ;
        RECT 82.705 179.385 82.875 179.575 ;
        RECT 83.165 179.385 83.335 179.575 ;
        RECT 86.845 179.405 87.015 179.595 ;
        RECT 88.225 179.405 88.395 179.595 ;
        RECT 92.825 179.405 92.995 179.575 ;
        RECT 93.745 179.405 93.915 179.595 ;
        RECT 95.115 179.405 95.285 179.595 ;
        RECT 95.585 179.405 95.755 179.595 ;
        RECT 97.420 179.435 97.540 179.545 ;
        RECT 97.885 179.405 98.055 179.595 ;
        RECT 101.105 179.405 101.275 179.595 ;
        RECT 108.950 179.575 109.060 179.595 ;
        RECT 92.825 179.385 92.985 179.405 ;
        RECT 102.025 179.385 102.195 179.575 ;
        RECT 102.485 179.405 102.655 179.575 ;
        RECT 106.625 179.405 106.795 179.575 ;
        RECT 108.950 179.405 109.120 179.575 ;
        RECT 102.495 179.385 102.655 179.405 ;
        RECT 106.630 179.385 106.795 179.405 ;
        RECT 109.835 179.385 110.005 179.575 ;
        RECT 110.315 179.385 110.485 179.575 ;
        RECT 111.685 179.385 111.855 179.595 ;
        RECT 112.155 179.405 112.325 179.595 ;
        RECT 113.985 179.385 114.155 179.575 ;
        RECT 114.435 179.405 114.605 179.595 ;
        RECT 115.815 179.405 115.985 179.595 ;
        RECT 116.295 179.405 116.465 179.595 ;
        RECT 117.670 179.405 117.840 179.625 ;
        RECT 119.330 179.595 120.275 179.625 ;
        RECT 120.285 179.595 121.655 180.375 ;
        RECT 121.665 179.595 125.335 180.405 ;
        RECT 126.275 179.680 126.705 180.465 ;
        RECT 126.925 180.415 127.875 180.505 ;
        RECT 126.925 179.595 128.855 180.415 ;
        RECT 129.025 179.595 130.395 180.405 ;
        RECT 130.425 179.595 131.775 180.505 ;
        RECT 132.705 180.305 133.650 180.505 ;
        RECT 135.465 180.305 136.410 180.505 ;
        RECT 140.950 180.305 141.895 180.505 ;
        RECT 132.705 179.625 135.455 180.305 ;
        RECT 135.465 179.625 138.215 180.305 ;
        RECT 139.145 179.625 141.895 180.305 ;
        RECT 142.565 180.275 146.495 180.505 ;
        RECT 132.705 179.595 133.650 179.625 ;
        RECT 119.500 179.385 119.670 179.575 ;
        RECT 119.965 179.385 120.135 179.575 ;
        RECT 120.435 179.405 120.605 179.595 ;
        RECT 121.805 179.405 121.975 179.595 ;
        RECT 128.705 179.575 128.855 179.595 ;
        RECT 125.495 179.440 125.655 179.550 ;
        RECT 128.705 179.405 128.875 179.575 ;
        RECT 129.165 179.405 129.335 179.595 ;
        RECT 130.545 179.425 130.715 179.575 ;
        RECT 131.015 179.430 131.175 179.540 ;
        RECT 49.865 179.355 50.815 179.385 ;
        RECT 47.145 178.675 50.815 179.355 ;
        RECT 49.865 178.475 50.815 178.675 ;
        RECT 50.835 178.475 52.185 179.385 ;
        RECT 52.665 178.605 54.035 179.385 ;
        RECT 54.045 178.575 57.715 179.385 ;
        RECT 58.185 178.605 59.555 179.385 ;
        RECT 59.565 178.605 60.935 179.385 ;
        RECT 61.875 178.515 62.305 179.300 ;
        RECT 62.325 178.705 70.595 179.385 ;
        RECT 69.145 178.475 70.595 178.705 ;
        RECT 70.605 178.575 76.115 179.385 ;
        RECT 77.175 178.475 83.015 179.385 ;
        RECT 83.025 178.575 86.695 179.385 ;
        RECT 87.635 178.515 88.065 179.300 ;
        RECT 89.330 178.475 92.985 179.385 ;
        RECT 93.230 178.705 102.335 179.385 ;
        RECT 102.495 178.475 106.150 179.385 ;
        RECT 106.630 178.705 108.465 179.385 ;
        RECT 107.535 178.475 108.465 178.705 ;
        RECT 108.785 178.605 110.155 179.385 ;
        RECT 110.165 178.605 111.535 179.385 ;
        RECT 111.545 178.575 113.375 179.385 ;
        RECT 113.395 178.515 113.825 179.300 ;
        RECT 113.845 178.575 116.595 179.385 ;
        RECT 116.895 178.475 119.815 179.385 ;
        RECT 119.825 178.705 128.930 179.385 ;
        RECT 129.945 178.475 130.835 179.425 ;
        RECT 131.460 179.405 131.630 179.595 ;
        RECT 131.930 179.355 132.100 179.575 ;
        RECT 135.140 179.405 135.310 179.625 ;
        RECT 135.465 179.595 136.410 179.625 ;
        RECT 135.605 179.385 135.775 179.575 ;
        RECT 137.900 179.405 138.070 179.625 ;
        RECT 138.375 179.440 138.535 179.550 ;
        RECT 139.290 179.405 139.460 179.625 ;
        RECT 140.950 179.595 141.895 179.625 ;
        RECT 142.080 179.595 146.495 180.275 ;
        RECT 146.525 179.595 147.875 180.505 ;
        RECT 148.805 179.595 150.175 180.405 ;
        RECT 142.080 179.575 142.190 179.595 ;
        RECT 139.740 179.435 139.860 179.545 ;
        RECT 140.205 179.385 140.375 179.575 ;
        RECT 142.020 179.405 142.190 179.575 ;
        RECT 146.640 179.405 146.810 179.595 ;
        RECT 147.565 179.385 147.735 179.575 ;
        RECT 148.035 179.440 148.195 179.550 ;
        RECT 149.865 179.385 150.035 179.595 ;
        RECT 134.505 179.355 135.455 179.385 ;
        RECT 131.785 178.675 135.455 179.355 ;
        RECT 135.465 178.705 139.135 179.385 ;
        RECT 134.505 178.475 135.455 178.675 ;
        RECT 138.205 178.475 139.135 178.705 ;
        RECT 139.155 178.515 139.585 179.300 ;
        RECT 140.065 178.705 147.375 179.385 ;
        RECT 143.580 178.485 144.490 178.705 ;
        RECT 146.025 178.475 147.375 178.705 ;
        RECT 147.425 178.575 148.795 179.385 ;
        RECT 148.805 178.575 150.175 179.385 ;
      LAYER nwell ;
        RECT 35.910 175.355 150.370 178.185 ;
      LAYER pwell ;
        RECT 36.105 174.155 37.475 174.965 ;
        RECT 37.485 174.155 40.235 174.965 ;
        RECT 40.245 174.155 41.595 175.065 ;
        RECT 41.625 174.155 44.375 174.965 ;
        RECT 44.385 174.835 48.315 175.065 ;
        RECT 44.385 174.155 48.800 174.835 ;
        RECT 48.995 174.240 49.425 175.025 ;
        RECT 49.445 174.865 50.390 175.065 ;
        RECT 49.445 174.185 52.195 174.865 ;
        RECT 49.445 174.155 50.390 174.185 ;
        RECT 36.245 173.945 36.415 174.155 ;
        RECT 37.625 173.945 37.795 174.155 ;
        RECT 40.390 173.965 40.560 174.155 ;
        RECT 41.315 173.990 41.475 174.100 ;
        RECT 41.765 173.965 41.935 174.155 ;
        RECT 48.690 174.135 48.800 174.155 ;
        RECT 43.600 173.945 43.770 174.135 ;
        RECT 44.065 173.945 44.235 174.135 ;
        RECT 47.285 173.945 47.455 174.135 ;
        RECT 47.755 173.945 47.925 174.135 ;
        RECT 48.690 173.965 48.860 174.135 ;
        RECT 49.120 173.945 49.290 174.135 ;
        RECT 50.515 173.945 50.685 174.135 ;
        RECT 51.880 173.965 52.050 174.185 ;
        RECT 52.205 174.155 53.575 174.935 ;
        RECT 53.585 174.835 55.035 175.065 ;
        RECT 53.585 174.155 61.855 174.835 ;
        RECT 61.950 174.155 71.055 174.835 ;
        RECT 71.065 174.155 74.735 174.965 ;
        RECT 74.755 174.240 75.185 175.025 ;
        RECT 75.205 174.155 80.715 174.965 ;
        RECT 80.725 174.155 82.555 174.965 ;
        RECT 84.075 174.835 85.005 175.065 ;
        RECT 86.375 174.835 87.305 175.065 ;
        RECT 83.170 174.155 85.005 174.835 ;
        RECT 85.470 174.155 87.305 174.835 ;
        RECT 87.820 174.155 91.295 175.065 ;
        RECT 91.595 174.155 94.515 175.065 ;
        RECT 94.525 174.155 95.895 174.965 ;
        RECT 95.905 174.835 99.835 175.065 ;
        RECT 95.905 174.155 100.320 174.835 ;
        RECT 100.515 174.240 100.945 175.025 ;
        RECT 52.355 173.965 52.525 174.155 ;
        RECT 53.255 173.945 53.425 174.135 ;
        RECT 53.720 173.995 53.840 174.105 ;
        RECT 54.195 173.945 54.365 174.135 ;
        RECT 56.475 173.945 56.645 174.135 ;
        RECT 56.945 173.945 57.115 174.135 ;
        RECT 60.625 173.945 60.795 174.135 ;
        RECT 61.545 173.965 61.715 174.155 ;
        RECT 62.465 173.945 62.635 174.135 ;
        RECT 63.845 173.945 64.015 174.135 ;
        RECT 70.745 173.965 70.915 174.155 ;
        RECT 71.205 173.965 71.375 174.155 ;
        RECT 72.120 173.995 72.240 174.105 ;
        RECT 72.595 173.945 72.765 174.135 ;
        RECT 73.965 173.945 74.135 174.135 ;
        RECT 75.345 173.965 75.515 174.155 ;
        RECT 80.865 173.965 81.035 174.155 ;
        RECT 83.170 174.135 83.335 174.155 ;
        RECT 85.470 174.135 85.635 174.155 ;
        RECT 81.325 173.945 81.495 174.135 ;
        RECT 82.700 173.995 82.820 174.105 ;
        RECT 83.165 173.965 83.335 174.135 ;
        RECT 85.005 173.945 85.175 174.135 ;
        RECT 85.465 173.965 85.635 174.135 ;
        RECT 86.380 173.945 86.550 174.135 ;
        RECT 88.225 173.965 88.395 174.135 ;
        RECT 90.980 173.965 91.150 174.155 ;
        RECT 88.235 173.945 88.395 173.965 ;
        RECT 92.370 173.945 92.540 174.135 ;
        RECT 94.200 173.965 94.370 174.155 ;
        RECT 94.665 173.965 94.835 174.155 ;
        RECT 100.210 174.135 100.320 174.155 ;
        RECT 101.115 174.155 104.770 175.065 ;
        RECT 105.395 174.155 108.315 175.065 ;
        RECT 108.325 174.155 111.535 175.065 ;
        RECT 111.545 174.155 114.295 174.965 ;
        RECT 114.965 174.835 118.895 175.065 ;
        RECT 114.480 174.155 118.895 174.835 ;
        RECT 118.905 174.155 120.720 175.065 ;
        RECT 120.745 174.155 122.575 175.065 ;
        RECT 123.045 174.155 126.255 175.065 ;
        RECT 126.275 174.240 126.705 175.025 ;
        RECT 126.745 174.155 128.095 175.065 ;
        RECT 131.620 174.835 132.530 175.055 ;
        RECT 134.065 174.835 135.835 175.065 ;
        RECT 128.105 174.155 135.835 174.835 ;
        RECT 136.385 174.155 137.755 174.935 ;
        RECT 137.775 174.155 139.125 175.065 ;
        RECT 139.145 174.155 144.655 174.965 ;
        RECT 144.665 174.155 148.335 174.965 ;
        RECT 148.805 174.155 150.175 174.965 ;
        RECT 101.115 174.135 101.275 174.155 ;
        RECT 95.585 173.945 95.755 174.135 ;
        RECT 99.260 173.995 99.380 174.105 ;
        RECT 99.725 173.965 99.895 174.135 ;
        RECT 100.210 173.965 100.380 174.135 ;
        RECT 101.105 173.965 101.275 174.135 ;
        RECT 99.735 173.945 99.895 173.965 ;
        RECT 103.860 173.945 104.030 174.135 ;
        RECT 105.255 173.990 105.415 174.100 ;
        RECT 108.000 173.965 108.170 174.155 ;
        RECT 108.465 173.945 108.635 174.155 ;
        RECT 108.925 173.945 109.095 174.135 ;
        RECT 111.685 173.965 111.855 174.155 ;
        RECT 114.480 174.135 114.590 174.155 ;
        RECT 112.615 173.990 112.775 174.100 ;
        RECT 113.985 173.945 114.155 174.135 ;
        RECT 114.420 173.965 114.590 174.135 ;
        RECT 115.820 173.995 115.940 174.105 ;
        RECT 116.295 173.945 116.465 174.135 ;
        RECT 117.665 173.945 117.835 174.135 ;
        RECT 119.500 173.995 119.620 174.105 ;
        RECT 119.965 173.945 120.135 174.135 ;
        RECT 120.425 173.965 120.595 174.155 ;
        RECT 120.890 173.965 121.060 174.155 ;
        RECT 121.805 173.945 121.975 174.135 ;
        RECT 122.720 173.995 122.840 174.105 ;
        RECT 123.185 173.965 123.355 174.155 ;
        RECT 127.325 173.945 127.495 174.135 ;
        RECT 127.780 173.965 127.950 174.155 ;
        RECT 128.245 173.965 128.415 174.155 ;
        RECT 132.845 173.945 133.015 174.135 ;
        RECT 136.060 173.995 136.180 174.105 ;
        RECT 136.525 173.945 136.695 174.155 ;
        RECT 138.825 174.135 138.995 174.155 ;
        RECT 138.815 173.965 138.995 174.135 ;
        RECT 139.285 173.965 139.455 174.155 ;
        RECT 138.815 173.945 138.985 173.965 ;
        RECT 139.745 173.945 139.915 174.135 ;
        RECT 143.885 173.945 144.055 174.135 ;
        RECT 144.805 173.965 144.975 174.155 ;
        RECT 147.565 173.945 147.735 174.135 ;
        RECT 148.480 173.995 148.600 174.105 ;
        RECT 149.865 173.945 150.035 174.155 ;
        RECT 36.105 173.135 37.475 173.945 ;
        RECT 37.485 173.135 41.155 173.945 ;
        RECT 42.085 173.035 43.915 173.945 ;
        RECT 43.925 173.135 45.295 173.945 ;
        RECT 45.305 173.265 47.595 173.945 ;
        RECT 45.305 173.035 46.225 173.265 ;
        RECT 47.605 173.165 48.975 173.945 ;
        RECT 49.005 173.035 50.355 173.945 ;
        RECT 50.365 173.165 51.735 173.945 ;
        RECT 52.205 173.165 53.575 173.945 ;
        RECT 54.045 173.165 55.415 173.945 ;
        RECT 55.425 173.165 56.795 173.945 ;
        RECT 56.805 173.135 60.475 173.945 ;
        RECT 60.485 173.135 61.855 173.945 ;
        RECT 61.875 173.075 62.305 173.860 ;
        RECT 62.325 173.135 63.695 173.945 ;
        RECT 63.705 173.265 71.975 173.945 ;
        RECT 70.525 173.035 71.975 173.265 ;
        RECT 72.445 173.165 73.815 173.945 ;
        RECT 73.825 173.265 81.135 173.945 ;
        RECT 77.340 173.045 78.250 173.265 ;
        RECT 79.785 173.035 81.135 173.265 ;
        RECT 81.185 173.135 84.855 173.945 ;
        RECT 84.865 173.135 86.235 173.945 ;
        RECT 86.265 173.035 87.615 173.945 ;
        RECT 87.635 173.075 88.065 173.860 ;
        RECT 88.235 173.035 91.890 173.945 ;
        RECT 92.225 173.035 95.145 173.945 ;
        RECT 95.445 173.135 99.115 173.945 ;
        RECT 99.735 173.035 103.390 173.945 ;
        RECT 103.745 173.035 105.095 173.945 ;
        RECT 106.025 173.035 108.775 173.945 ;
        RECT 108.785 173.135 112.455 173.945 ;
        RECT 113.395 173.075 113.825 173.860 ;
        RECT 113.845 173.135 115.675 173.945 ;
        RECT 116.145 173.165 117.515 173.945 ;
        RECT 117.525 173.135 119.355 173.945 ;
        RECT 119.840 173.035 121.655 173.945 ;
        RECT 121.665 173.135 127.175 173.945 ;
        RECT 127.185 173.135 132.695 173.945 ;
        RECT 132.705 173.135 136.375 173.945 ;
        RECT 136.385 173.135 137.755 173.945 ;
        RECT 137.765 173.165 139.135 173.945 ;
        RECT 139.155 173.075 139.585 173.860 ;
        RECT 139.605 173.035 143.665 173.945 ;
        RECT 143.745 173.135 147.415 173.945 ;
        RECT 147.425 173.135 148.795 173.945 ;
        RECT 148.805 173.135 150.175 173.945 ;
      LAYER nwell ;
        RECT 35.910 169.915 150.370 172.745 ;
      LAYER pwell ;
        RECT 36.105 168.715 37.475 169.525 ;
        RECT 37.485 168.715 40.235 169.525 ;
        RECT 40.705 168.715 42.535 169.625 ;
        RECT 43.685 169.535 44.635 169.625 ;
        RECT 42.705 168.715 44.635 169.535 ;
        RECT 44.865 168.715 46.215 169.625 ;
        RECT 46.225 169.395 47.145 169.625 ;
        RECT 46.225 168.715 48.515 169.395 ;
        RECT 48.995 168.800 49.425 169.585 ;
        RECT 49.445 168.715 54.955 169.525 ;
        RECT 54.965 168.715 60.475 169.525 ;
        RECT 60.945 168.715 62.315 169.495 ;
        RECT 69.145 169.395 70.595 169.625 ;
        RECT 62.325 168.715 70.595 169.395 ;
        RECT 70.605 168.715 74.275 169.525 ;
        RECT 74.755 168.800 75.185 169.585 ;
        RECT 75.205 169.425 76.155 169.625 ;
        RECT 77.485 169.425 78.415 169.625 ;
        RECT 75.205 168.945 78.415 169.425 ;
        RECT 75.205 168.745 78.270 168.945 ;
        RECT 75.205 168.715 76.140 168.745 ;
        RECT 36.245 168.505 36.415 168.715 ;
        RECT 37.625 168.505 37.795 168.715 ;
        RECT 40.380 168.555 40.500 168.665 ;
        RECT 40.850 168.525 41.020 168.715 ;
        RECT 42.705 168.695 42.855 168.715 ;
        RECT 41.300 168.555 41.420 168.665 ;
        RECT 36.105 167.695 37.475 168.505 ;
        RECT 37.485 167.695 41.155 168.505 ;
        RECT 41.770 168.475 41.940 168.695 ;
        RECT 42.685 168.525 42.855 168.695 ;
        RECT 44.985 168.505 45.155 168.695 ;
        RECT 45.900 168.525 46.070 168.715 ;
        RECT 48.205 168.525 48.375 168.715 ;
        RECT 48.660 168.555 48.780 168.665 ;
        RECT 49.585 168.525 49.755 168.715 ;
        RECT 52.345 168.505 52.515 168.695 ;
        RECT 55.105 168.525 55.275 168.715 ;
        RECT 57.870 168.505 58.040 168.695 ;
        RECT 60.620 168.555 60.740 168.665 ;
        RECT 61.095 168.525 61.265 168.715 ;
        RECT 62.465 168.505 62.635 168.715 ;
        RECT 69.825 168.505 69.995 168.695 ;
        RECT 70.745 168.525 70.915 168.715 ;
        RECT 71.215 168.505 71.385 168.695 ;
        RECT 72.585 168.505 72.755 168.695 ;
        RECT 74.420 168.555 74.540 168.665 ;
        RECT 75.810 168.505 75.980 168.695 ;
        RECT 78.100 168.525 78.270 168.745 ;
        RECT 78.425 168.715 83.935 169.525 ;
        RECT 83.945 168.715 87.615 169.525 ;
        RECT 87.625 168.715 90.545 169.625 ;
        RECT 91.135 168.715 94.055 169.625 ;
        RECT 95.115 169.395 96.045 169.625 ;
        RECT 94.210 168.715 96.045 169.395 ;
        RECT 96.365 168.715 100.035 169.525 ;
        RECT 100.515 168.800 100.945 169.585 ;
        RECT 100.965 168.715 103.715 169.625 ;
        RECT 103.725 168.715 107.395 169.525 ;
        RECT 107.425 168.715 108.775 169.625 ;
        RECT 109.075 168.715 111.995 169.625 ;
        RECT 113.055 169.395 113.985 169.625 ;
        RECT 112.150 168.715 113.985 169.395 ;
        RECT 114.305 168.715 115.675 169.495 ;
        RECT 115.685 168.715 121.195 169.525 ;
        RECT 121.205 168.715 123.035 169.525 ;
        RECT 123.065 168.715 124.415 169.625 ;
        RECT 124.425 168.715 126.255 169.525 ;
        RECT 126.275 168.800 126.705 169.585 ;
        RECT 126.725 168.715 129.935 169.625 ;
        RECT 129.945 168.715 135.455 169.525 ;
        RECT 135.465 168.715 137.295 169.525 ;
        RECT 139.570 169.425 140.515 169.625 ;
        RECT 137.765 168.745 140.515 169.425 ;
        RECT 144.040 169.395 144.950 169.615 ;
        RECT 146.485 169.395 147.835 169.625 ;
        RECT 78.565 168.525 78.735 168.715 ;
        RECT 79.025 168.505 79.195 168.695 ;
        RECT 80.405 168.505 80.575 168.695 ;
        RECT 84.085 168.525 84.255 168.715 ;
        RECT 85.920 168.555 86.040 168.665 ;
        RECT 87.295 168.505 87.465 168.695 ;
        RECT 87.770 168.525 87.940 168.715 ;
        RECT 91.440 168.505 91.610 168.695 ;
        RECT 91.905 168.505 92.075 168.695 ;
        RECT 93.740 168.525 93.910 168.715 ;
        RECT 94.210 168.695 94.375 168.715 ;
        RECT 96.505 168.695 96.675 168.715 ;
        RECT 94.205 168.525 94.375 168.695 ;
        RECT 96.500 168.525 96.675 168.695 ;
        RECT 96.965 168.525 97.135 168.695 ;
        RECT 100.180 168.555 100.300 168.665 ;
        RECT 96.500 168.505 96.670 168.525 ;
        RECT 96.975 168.505 97.135 168.525 ;
        RECT 101.105 168.505 101.275 168.715 ;
        RECT 103.865 168.505 104.035 168.715 ;
        RECT 107.540 168.525 107.710 168.715 ;
        RECT 111.680 168.695 111.850 168.715 ;
        RECT 112.150 168.695 112.315 168.715 ;
        RECT 110.295 168.505 110.465 168.695 ;
        RECT 111.675 168.525 111.850 168.695 ;
        RECT 111.675 168.505 111.845 168.525 ;
        RECT 112.145 168.505 112.315 168.695 ;
        RECT 113.985 168.505 114.155 168.695 ;
        RECT 115.355 168.525 115.525 168.715 ;
        RECT 115.825 168.525 115.995 168.715 ;
        RECT 118.575 168.505 118.745 168.695 ;
        RECT 119.055 168.505 119.225 168.695 ;
        RECT 120.435 168.550 120.595 168.660 ;
        RECT 121.345 168.525 121.515 168.715 ;
        RECT 122.260 168.505 122.430 168.695 ;
        RECT 124.100 168.525 124.270 168.715 ;
        RECT 124.565 168.525 124.735 168.715 ;
        RECT 124.565 168.505 124.715 168.525 ;
        RECT 125.025 168.505 125.195 168.695 ;
        RECT 126.865 168.525 127.035 168.715 ;
        RECT 128.250 168.505 128.420 168.695 ;
        RECT 129.625 168.505 129.795 168.695 ;
        RECT 130.085 168.525 130.255 168.715 ;
        RECT 131.460 168.555 131.580 168.665 ;
        RECT 131.925 168.505 132.095 168.695 ;
        RECT 135.605 168.525 135.775 168.715 ;
        RECT 137.440 168.555 137.560 168.665 ;
        RECT 137.910 168.525 138.080 168.745 ;
        RECT 139.570 168.715 140.515 168.745 ;
        RECT 140.525 168.715 147.835 169.395 ;
        RECT 148.805 168.715 150.175 169.525 ;
        RECT 139.740 168.555 139.860 168.665 ;
        RECT 43.900 168.475 44.835 168.505 ;
        RECT 41.770 168.275 44.835 168.475 ;
        RECT 41.625 167.795 44.835 168.275 ;
        RECT 44.845 167.825 52.155 168.505 ;
        RECT 41.625 167.595 42.555 167.795 ;
        RECT 43.885 167.595 44.835 167.795 ;
        RECT 48.360 167.605 49.270 167.825 ;
        RECT 50.805 167.595 52.155 167.825 ;
        RECT 52.205 167.695 57.715 168.505 ;
        RECT 57.725 167.595 60.645 168.505 ;
        RECT 61.875 167.635 62.305 168.420 ;
        RECT 62.325 167.825 69.635 168.505 ;
        RECT 65.840 167.605 66.750 167.825 ;
        RECT 68.285 167.595 69.635 167.825 ;
        RECT 69.685 167.695 71.055 168.505 ;
        RECT 71.065 167.725 72.435 168.505 ;
        RECT 72.445 167.825 75.655 168.505 ;
        RECT 74.520 167.595 75.655 167.825 ;
        RECT 75.665 167.595 78.585 168.505 ;
        RECT 78.895 167.595 80.245 168.505 ;
        RECT 80.265 167.695 85.775 168.505 ;
        RECT 86.245 167.725 87.615 168.505 ;
        RECT 87.635 167.635 88.065 168.420 ;
        RECT 88.280 167.595 91.755 168.505 ;
        RECT 91.765 167.695 93.595 168.505 ;
        RECT 93.895 167.595 96.815 168.505 ;
        RECT 96.975 167.595 100.630 168.505 ;
        RECT 100.965 167.595 103.715 168.505 ;
        RECT 103.725 167.695 109.235 168.505 ;
        RECT 109.245 167.725 110.615 168.505 ;
        RECT 110.625 167.725 111.995 168.505 ;
        RECT 112.005 167.695 113.375 168.505 ;
        RECT 113.395 167.635 113.825 168.420 ;
        RECT 113.845 167.695 117.515 168.505 ;
        RECT 117.525 167.725 118.895 168.505 ;
        RECT 118.905 167.725 120.275 168.505 ;
        RECT 121.225 167.595 122.575 168.505 ;
        RECT 122.785 167.685 124.715 168.505 ;
        RECT 122.785 167.595 123.735 167.685 ;
        RECT 124.885 167.595 128.095 168.505 ;
        RECT 128.105 167.595 129.455 168.505 ;
        RECT 129.485 167.695 131.315 168.505 ;
        RECT 131.785 167.825 139.095 168.505 ;
        RECT 135.300 167.605 136.210 167.825 ;
        RECT 137.745 167.595 139.095 167.825 ;
        RECT 139.155 167.635 139.585 168.420 ;
        RECT 140.205 168.275 140.375 168.695 ;
        RECT 140.665 168.525 140.835 168.715 ;
        RECT 144.345 168.505 144.515 168.695 ;
        RECT 146.185 168.505 146.355 168.695 ;
        RECT 148.035 168.560 148.195 168.670 ;
        RECT 149.865 168.505 150.035 168.715 ;
        RECT 141.485 168.275 144.195 168.505 ;
        RECT 140.100 167.825 144.195 168.275 ;
        RECT 144.205 167.825 146.035 168.505 ;
        RECT 140.100 167.595 141.475 167.825 ;
        RECT 143.245 167.595 144.195 167.825 ;
        RECT 144.690 167.595 146.035 167.825 ;
        RECT 146.045 167.695 148.795 168.505 ;
        RECT 148.805 167.695 150.175 168.505 ;
      LAYER nwell ;
        RECT 35.910 164.475 150.370 167.305 ;
      LAYER pwell ;
        RECT 36.105 163.275 37.475 164.085 ;
        RECT 37.485 163.275 42.995 164.085 ;
        RECT 43.005 163.275 44.835 164.185 ;
        RECT 44.845 163.275 46.215 164.055 ;
        RECT 46.225 163.275 48.975 164.085 ;
        RECT 48.995 163.360 49.425 164.145 ;
        RECT 49.445 163.275 53.115 164.085 ;
        RECT 53.125 163.955 57.055 164.185 ;
        RECT 53.125 163.275 57.540 163.955 ;
        RECT 57.725 163.275 59.095 164.085 ;
        RECT 59.105 163.275 60.475 164.055 ;
        RECT 61.145 163.955 65.075 164.185 ;
        RECT 65.745 163.955 69.675 164.185 ;
        RECT 60.660 163.275 65.075 163.955 ;
        RECT 65.260 163.275 69.675 163.955 ;
        RECT 70.245 163.275 73.355 164.185 ;
        RECT 73.365 163.275 74.735 164.085 ;
        RECT 74.755 163.360 75.185 164.145 ;
        RECT 75.215 163.275 77.945 164.185 ;
        RECT 77.965 163.275 83.475 164.085 ;
        RECT 83.485 163.275 84.855 164.085 ;
        RECT 85.915 163.955 86.845 164.185 ;
        RECT 85.010 163.275 86.845 163.955 ;
        RECT 87.315 163.275 90.970 164.185 ;
        RECT 91.595 163.275 94.515 164.185 ;
        RECT 94.985 163.275 98.460 164.185 ;
        RECT 98.665 163.275 100.495 164.085 ;
        RECT 100.515 163.360 100.945 164.145 ;
        RECT 101.625 163.955 105.555 164.185 ;
        RECT 101.140 163.275 105.555 163.955 ;
        RECT 105.565 163.275 106.935 164.085 ;
        RECT 106.945 163.275 108.315 164.055 ;
        RECT 108.325 163.275 111.535 164.185 ;
        RECT 111.545 163.955 114.370 164.185 ;
        RECT 125.105 164.095 126.055 164.185 ;
        RECT 111.545 163.275 115.075 163.955 ;
        RECT 115.225 163.275 120.735 164.085 ;
        RECT 121.665 163.275 123.035 164.055 ;
        RECT 124.125 163.275 126.055 164.095 ;
        RECT 126.275 163.360 126.705 164.145 ;
        RECT 126.745 163.275 128.095 164.185 ;
        RECT 128.105 163.275 133.615 164.085 ;
        RECT 133.625 163.275 137.295 164.085 ;
        RECT 137.305 163.275 138.675 164.085 ;
        RECT 138.685 163.985 139.640 164.185 ;
        RECT 138.685 163.305 140.965 163.985 ;
        RECT 138.685 163.275 139.640 163.305 ;
        RECT 36.245 163.065 36.415 163.275 ;
        RECT 37.625 163.065 37.795 163.275 ;
        RECT 39.460 163.115 39.580 163.225 ;
        RECT 39.925 163.065 40.095 163.255 ;
        RECT 44.520 163.085 44.690 163.275 ;
        RECT 45.905 163.085 46.075 163.275 ;
        RECT 46.365 163.085 46.535 163.275 ;
        RECT 47.285 163.065 47.455 163.255 ;
        RECT 49.585 163.085 49.755 163.275 ;
        RECT 57.430 163.255 57.540 163.275 ;
        RECT 50.040 163.115 50.160 163.225 ;
        RECT 51.415 163.065 51.585 163.255 ;
        RECT 51.860 163.085 52.030 163.255 ;
        RECT 56.485 163.085 56.655 163.255 ;
        RECT 57.430 163.085 57.600 163.255 ;
        RECT 57.865 163.085 58.035 163.275 ;
        RECT 51.920 163.065 52.030 163.085 ;
        RECT 56.505 163.065 56.655 163.085 ;
        RECT 58.785 163.065 58.955 163.255 ;
        RECT 59.245 163.085 59.415 163.275 ;
        RECT 60.660 163.255 60.770 163.275 ;
        RECT 65.260 163.255 65.370 163.275 ;
        RECT 60.175 163.065 60.345 163.255 ;
        RECT 60.600 163.085 60.770 163.255 ;
        RECT 61.540 163.115 61.660 163.225 ;
        RECT 62.465 163.065 62.635 163.255 ;
        RECT 63.845 163.065 64.015 163.255 ;
        RECT 65.200 163.085 65.370 163.255 ;
        RECT 66.600 163.115 66.720 163.225 ;
        RECT 67.065 163.065 67.235 163.255 ;
        RECT 69.820 163.115 69.940 163.225 ;
        RECT 70.285 163.085 70.455 163.275 ;
        RECT 70.305 163.065 70.455 163.085 ;
        RECT 72.585 163.065 72.755 163.255 ;
        RECT 73.505 163.085 73.675 163.275 ;
        RECT 77.645 163.085 77.815 163.275 ;
        RECT 78.105 163.065 78.275 163.275 ;
        RECT 83.625 163.065 83.795 163.275 ;
        RECT 85.010 163.255 85.175 163.275 ;
        RECT 87.315 163.255 87.475 163.275 ;
        RECT 85.005 163.085 85.175 163.255 ;
        RECT 86.395 163.065 86.565 163.255 ;
        RECT 87.305 163.085 87.475 163.255 ;
        RECT 88.225 163.065 88.395 163.255 ;
        RECT 91.900 163.065 92.070 163.255 ;
        RECT 93.285 163.065 93.455 163.255 ;
        RECT 94.200 163.085 94.370 163.275 ;
        RECT 94.660 163.115 94.780 163.225 ;
        RECT 95.130 163.085 95.300 163.275 ;
        RECT 96.960 163.115 97.080 163.225 ;
        RECT 98.805 163.085 98.975 163.275 ;
        RECT 101.140 163.255 101.250 163.275 ;
        RECT 99.725 163.065 99.895 163.255 ;
        RECT 100.195 163.110 100.355 163.220 ;
        RECT 101.080 163.085 101.275 163.255 ;
        RECT 101.105 163.065 101.275 163.085 ;
        RECT 105.235 163.065 105.405 163.255 ;
        RECT 105.705 163.065 105.875 163.275 ;
        RECT 107.995 163.085 108.165 163.275 ;
        RECT 108.465 163.085 108.635 163.275 ;
        RECT 114.875 163.255 115.075 163.275 ;
        RECT 109.385 163.085 109.555 163.255 ;
        RECT 113.985 163.085 114.155 163.255 ;
        RECT 114.905 163.085 115.075 163.255 ;
        RECT 115.365 163.085 115.535 163.275 ;
        RECT 109.395 163.065 109.555 163.085 ;
        RECT 113.995 163.065 114.155 163.085 ;
        RECT 118.125 163.065 118.295 163.255 ;
        RECT 120.895 163.120 121.055 163.230 ;
        RECT 121.815 163.085 121.985 163.275 ;
        RECT 124.125 163.255 124.275 163.275 ;
        RECT 123.195 163.120 123.355 163.230 ;
        RECT 36.105 162.255 37.475 163.065 ;
        RECT 37.485 162.255 39.315 163.065 ;
        RECT 39.785 162.385 47.095 163.065 ;
        RECT 43.300 162.165 44.210 162.385 ;
        RECT 45.745 162.155 47.095 162.385 ;
        RECT 47.145 162.255 49.895 163.065 ;
        RECT 50.365 162.285 51.735 163.065 ;
        RECT 51.920 162.385 56.335 163.065 ;
        RECT 52.405 162.155 56.335 162.385 ;
        RECT 56.505 162.245 58.435 163.065 ;
        RECT 58.645 162.255 60.015 163.065 ;
        RECT 60.025 162.285 61.395 163.065 ;
        RECT 57.485 162.155 58.435 162.245 ;
        RECT 61.875 162.195 62.305 162.980 ;
        RECT 62.335 162.155 63.685 163.065 ;
        RECT 63.705 162.255 66.455 163.065 ;
        RECT 66.965 162.155 70.135 163.065 ;
        RECT 70.305 162.245 72.235 163.065 ;
        RECT 72.445 162.255 77.955 163.065 ;
        RECT 77.965 162.255 83.475 163.065 ;
        RECT 83.485 162.255 86.235 163.065 ;
        RECT 86.245 162.285 87.615 163.065 ;
        RECT 71.285 162.155 72.235 162.245 ;
        RECT 87.635 162.195 88.065 162.980 ;
        RECT 88.085 162.255 91.755 163.065 ;
        RECT 91.785 162.155 93.135 163.065 ;
        RECT 93.145 162.255 96.815 163.065 ;
        RECT 97.285 162.155 100.035 163.065 ;
        RECT 100.965 162.155 104.175 163.065 ;
        RECT 104.185 162.285 105.555 163.065 ;
        RECT 105.565 162.255 109.235 163.065 ;
        RECT 109.395 162.155 113.050 163.065 ;
        RECT 113.395 162.195 113.825 162.980 ;
        RECT 113.995 162.155 117.650 163.065 ;
        RECT 117.985 162.255 123.495 163.065 ;
        RECT 123.650 163.035 123.820 163.255 ;
        RECT 124.105 163.085 124.275 163.255 ;
        RECT 126.405 163.065 126.575 163.255 ;
        RECT 127.780 163.085 127.950 163.275 ;
        RECT 128.245 163.085 128.415 163.275 ;
        RECT 128.695 163.065 128.865 163.255 ;
        RECT 129.165 163.065 129.335 163.255 ;
        RECT 131.010 163.065 131.180 163.255 ;
        RECT 132.845 163.065 133.015 163.255 ;
        RECT 133.765 163.085 133.935 163.275 ;
        RECT 134.685 163.105 134.855 163.255 ;
        RECT 135.615 163.110 135.775 163.220 ;
        RECT 125.310 163.035 126.255 163.065 ;
        RECT 123.505 162.355 126.255 163.035 ;
        RECT 125.310 162.155 126.255 162.355 ;
        RECT 126.265 162.255 127.635 163.065 ;
        RECT 127.645 162.285 129.015 163.065 ;
        RECT 129.025 162.255 130.855 163.065 ;
        RECT 130.865 162.155 132.695 163.065 ;
        RECT 132.705 162.255 134.535 163.065 ;
        RECT 134.565 162.155 135.455 163.105 ;
        RECT 136.530 163.035 136.700 163.255 ;
        RECT 137.445 163.085 137.615 163.275 ;
        RECT 139.745 163.065 139.915 163.255 ;
        RECT 140.670 163.085 140.840 163.305 ;
        RECT 140.985 163.275 142.815 163.955 ;
        RECT 142.825 163.275 144.175 164.185 ;
        RECT 144.205 163.275 147.875 164.085 ;
        RECT 148.805 163.275 150.175 164.085 ;
        RECT 142.505 163.085 142.675 163.275 ;
        RECT 143.890 163.085 144.060 163.275 ;
        RECT 144.345 163.085 144.515 163.275 ;
        RECT 147.105 163.065 147.275 163.255 ;
        RECT 148.035 163.120 148.195 163.230 ;
        RECT 149.865 163.065 150.035 163.275 ;
        RECT 138.190 163.035 139.135 163.065 ;
        RECT 136.385 162.355 139.135 163.035 ;
        RECT 138.190 162.155 139.135 162.355 ;
        RECT 139.155 162.195 139.585 162.980 ;
        RECT 139.605 162.385 146.915 163.065 ;
        RECT 143.120 162.165 144.030 162.385 ;
        RECT 145.565 162.155 146.915 162.385 ;
        RECT 146.965 162.255 148.795 163.065 ;
        RECT 148.805 162.255 150.175 163.065 ;
      LAYER nwell ;
        RECT 35.910 159.035 150.370 161.865 ;
      LAYER pwell ;
        RECT 36.105 157.835 37.475 158.645 ;
        RECT 37.485 157.835 41.155 158.645 ;
        RECT 42.100 157.835 43.915 158.745 ;
        RECT 45.985 158.655 46.935 158.745 ;
        RECT 45.005 157.835 46.935 158.655 ;
        RECT 47.145 157.835 48.975 158.645 ;
        RECT 48.995 157.920 49.425 158.705 ;
        RECT 49.445 157.835 53.115 158.645 ;
        RECT 53.625 157.835 56.795 158.745 ;
        RECT 56.805 157.835 58.175 158.645 ;
        RECT 58.195 157.835 60.925 158.745 ;
        RECT 72.665 158.655 73.615 158.745 ;
        RECT 60.945 157.835 66.455 158.645 ;
        RECT 66.465 157.835 70.135 158.645 ;
        RECT 70.145 157.835 71.515 158.645 ;
        RECT 71.685 157.835 73.615 158.655 ;
        RECT 74.755 157.920 75.185 158.705 ;
        RECT 75.205 157.835 76.555 158.745 ;
        RECT 76.585 157.835 78.415 158.645 ;
        RECT 78.425 157.835 84.245 158.745 ;
        RECT 84.405 157.835 89.915 158.645 ;
        RECT 89.925 157.835 95.435 158.645 ;
        RECT 95.445 157.835 96.815 158.645 ;
        RECT 97.020 157.835 100.495 158.745 ;
        RECT 100.515 157.920 100.945 158.705 ;
        RECT 101.115 157.835 104.770 158.745 ;
        RECT 105.105 157.835 107.855 158.745 ;
        RECT 107.865 157.835 109.235 158.645 ;
        RECT 109.570 157.835 113.225 158.745 ;
        RECT 113.385 157.835 116.135 158.745 ;
        RECT 116.145 157.835 121.655 158.645 ;
        RECT 121.665 157.835 124.415 158.645 ;
        RECT 124.885 157.835 126.255 158.615 ;
        RECT 126.275 157.920 126.705 158.705 ;
        RECT 127.385 158.515 131.315 158.745 ;
        RECT 126.900 157.835 131.315 158.515 ;
        RECT 131.325 157.835 132.695 158.645 ;
        RECT 132.900 157.835 136.375 158.745 ;
        RECT 136.580 157.835 140.055 158.745 ;
        RECT 140.065 157.835 141.435 158.615 ;
        RECT 141.445 157.835 142.815 158.615 ;
        RECT 142.825 157.835 144.655 158.515 ;
        RECT 144.665 157.835 146.035 158.615 ;
        RECT 146.045 157.835 147.415 158.615 ;
        RECT 147.425 157.835 148.795 158.645 ;
        RECT 148.805 157.835 150.175 158.645 ;
        RECT 36.245 157.625 36.415 157.835 ;
        RECT 37.625 157.785 37.795 157.835 ;
        RECT 37.620 157.675 37.795 157.785 ;
        RECT 37.625 157.645 37.795 157.675 ;
        RECT 38.085 157.625 38.255 157.815 ;
        RECT 41.315 157.680 41.475 157.790 ;
        RECT 42.225 157.645 42.395 157.835 ;
        RECT 45.005 157.815 45.155 157.835 ;
        RECT 44.075 157.680 44.235 157.790 ;
        RECT 44.985 157.645 45.155 157.815 ;
        RECT 45.445 157.625 45.615 157.815 ;
        RECT 46.825 157.625 46.995 157.815 ;
        RECT 47.285 157.645 47.455 157.835 ;
        RECT 48.665 157.625 48.835 157.815 ;
        RECT 49.585 157.645 49.755 157.835 ;
        RECT 53.260 157.675 53.380 157.785 ;
        RECT 53.725 157.645 53.895 157.835 ;
        RECT 56.945 157.645 57.115 157.835 ;
        RECT 58.325 157.625 58.495 157.815 ;
        RECT 60.625 157.645 60.795 157.835 ;
        RECT 61.085 157.645 61.255 157.835 ;
        RECT 61.545 157.625 61.715 157.815 ;
        RECT 62.475 157.670 62.635 157.780 ;
        RECT 63.385 157.645 63.555 157.815 ;
        RECT 63.535 157.625 63.555 157.645 ;
        RECT 66.145 157.625 66.315 157.815 ;
        RECT 66.605 157.645 66.775 157.835 ;
        RECT 68.905 157.625 69.075 157.815 ;
        RECT 70.285 157.645 70.455 157.835 ;
        RECT 71.685 157.815 71.835 157.835 ;
        RECT 71.665 157.645 71.845 157.815 ;
        RECT 71.675 157.625 71.845 157.645 ;
        RECT 73.960 157.790 74.130 157.815 ;
        RECT 73.960 157.680 74.135 157.790 ;
        RECT 73.960 157.625 74.130 157.680 ;
        RECT 74.435 157.625 74.605 157.815 ;
        RECT 75.350 157.645 75.520 157.835 ;
        RECT 76.725 157.645 76.895 157.835 ;
        RECT 78.565 157.815 78.735 157.835 ;
        RECT 78.560 157.645 78.735 157.815 ;
        RECT 82.245 157.645 82.415 157.815 ;
        RECT 84.545 157.645 84.715 157.835 ;
        RECT 78.560 157.625 78.730 157.645 ;
        RECT 82.215 157.625 82.415 157.645 ;
        RECT 85.920 157.625 86.090 157.815 ;
        RECT 87.310 157.625 87.480 157.815 ;
        RECT 88.235 157.670 88.395 157.780 ;
        RECT 90.065 157.645 90.235 157.835 ;
        RECT 91.445 157.625 91.615 157.815 ;
        RECT 91.900 157.675 92.020 157.785 ;
        RECT 94.205 157.625 94.375 157.815 ;
        RECT 94.675 157.625 94.845 157.815 ;
        RECT 95.585 157.645 95.755 157.835 ;
        RECT 96.045 157.625 96.215 157.815 ;
        RECT 98.805 157.625 98.975 157.815 ;
        RECT 100.180 157.645 100.350 157.835 ;
        RECT 101.115 157.815 101.275 157.835 ;
        RECT 101.105 157.645 101.275 157.815 ;
        RECT 102.020 157.625 102.190 157.815 ;
        RECT 103.405 157.625 103.575 157.815 ;
        RECT 107.545 157.645 107.715 157.835 ;
        RECT 108.005 157.645 108.175 157.835 ;
        RECT 113.065 157.815 113.225 157.835 ;
        RECT 112.140 157.625 112.310 157.815 ;
        RECT 112.615 157.670 112.775 157.780 ;
        RECT 113.065 157.645 113.235 157.815 ;
        RECT 114.910 157.625 115.080 157.815 ;
        RECT 115.365 157.625 115.535 157.815 ;
        RECT 115.825 157.645 115.995 157.835 ;
        RECT 116.285 157.645 116.455 157.835 ;
        RECT 119.055 157.670 119.215 157.780 ;
        RECT 119.970 157.625 120.140 157.815 ;
        RECT 121.345 157.625 121.515 157.815 ;
        RECT 121.805 157.645 121.975 157.835 ;
        RECT 124.105 157.625 124.275 157.815 ;
        RECT 124.575 157.785 124.745 157.815 ;
        RECT 124.560 157.675 124.745 157.785 ;
        RECT 124.575 157.625 124.745 157.675 ;
        RECT 125.935 157.645 126.105 157.835 ;
        RECT 126.900 157.815 127.010 157.835 ;
        RECT 126.840 157.645 127.035 157.815 ;
        RECT 127.335 157.670 127.495 157.780 ;
        RECT 126.865 157.625 127.035 157.645 ;
        RECT 128.245 157.625 128.415 157.815 ;
        RECT 130.555 157.670 130.715 157.780 ;
        RECT 131.465 157.645 131.635 157.835 ;
        RECT 131.470 157.625 131.635 157.645 ;
        RECT 134.675 157.625 134.845 157.815 ;
        RECT 135.145 157.625 135.315 157.815 ;
        RECT 136.060 157.645 136.230 157.835 ;
        RECT 139.740 157.815 139.910 157.835 ;
        RECT 138.820 157.675 138.940 157.785 ;
        RECT 139.740 157.645 139.915 157.815 ;
        RECT 141.115 157.645 141.285 157.835 ;
        RECT 142.495 157.645 142.665 157.835 ;
        RECT 144.345 157.645 144.515 157.835 ;
        RECT 145.715 157.645 145.885 157.835 ;
        RECT 147.095 157.815 147.265 157.835 ;
        RECT 147.095 157.645 147.275 157.815 ;
        RECT 147.565 157.645 147.735 157.835 ;
        RECT 139.745 157.625 139.915 157.645 ;
        RECT 147.105 157.625 147.275 157.645 ;
        RECT 149.865 157.625 150.035 157.835 ;
        RECT 36.105 156.815 37.475 157.625 ;
        RECT 37.945 156.945 45.255 157.625 ;
        RECT 41.460 156.725 42.370 156.945 ;
        RECT 43.905 156.715 45.255 156.945 ;
        RECT 45.305 156.815 46.675 157.625 ;
        RECT 46.685 156.945 48.515 157.625 ;
        RECT 48.525 156.815 51.275 157.625 ;
        RECT 51.325 156.945 58.635 157.625 ;
        RECT 51.325 156.715 52.675 156.945 ;
        RECT 54.210 156.725 55.120 156.945 ;
        RECT 58.645 156.715 61.755 157.625 ;
        RECT 61.875 156.755 62.305 157.540 ;
        RECT 63.535 156.945 65.985 157.625 ;
        RECT 64.025 156.715 65.985 156.945 ;
        RECT 66.005 156.715 68.755 157.625 ;
        RECT 68.765 156.815 71.515 157.625 ;
        RECT 71.525 156.845 72.895 157.625 ;
        RECT 72.925 156.715 74.275 157.625 ;
        RECT 74.285 156.845 75.655 157.625 ;
        RECT 75.955 156.715 78.875 157.625 ;
        RECT 78.885 156.945 82.415 157.625 ;
        RECT 78.885 156.715 81.710 156.945 ;
        RECT 82.565 156.715 86.235 157.625 ;
        RECT 86.245 156.715 87.595 157.625 ;
        RECT 87.635 156.755 88.065 157.540 ;
        RECT 89.005 156.945 91.755 157.625 ;
        RECT 92.225 156.945 94.515 157.625 ;
        RECT 89.005 156.715 89.935 156.945 ;
        RECT 92.225 156.715 93.145 156.945 ;
        RECT 94.525 156.845 95.895 157.625 ;
        RECT 95.905 156.815 98.655 157.625 ;
        RECT 98.665 156.715 101.875 157.625 ;
        RECT 101.905 156.715 103.255 157.625 ;
        RECT 103.265 156.815 108.775 157.625 ;
        RECT 108.980 156.715 112.455 157.625 ;
        RECT 113.395 156.755 113.825 157.540 ;
        RECT 113.845 156.715 115.195 157.625 ;
        RECT 115.225 156.815 118.895 157.625 ;
        RECT 119.825 156.715 121.175 157.625 ;
        RECT 121.205 156.815 123.035 157.625 ;
        RECT 123.055 156.715 124.405 157.625 ;
        RECT 124.425 156.845 125.795 157.625 ;
        RECT 125.815 156.715 127.165 157.625 ;
        RECT 128.105 156.945 130.395 157.625 ;
        RECT 131.470 156.945 133.305 157.625 ;
        RECT 129.475 156.715 130.395 156.945 ;
        RECT 132.375 156.715 133.305 156.945 ;
        RECT 133.625 156.845 134.995 157.625 ;
        RECT 135.005 156.815 138.675 157.625 ;
        RECT 139.155 156.755 139.585 157.540 ;
        RECT 139.605 156.945 146.915 157.625 ;
        RECT 143.120 156.725 144.030 156.945 ;
        RECT 145.565 156.715 146.915 156.945 ;
        RECT 146.965 156.815 148.795 157.625 ;
        RECT 148.805 156.815 150.175 157.625 ;
      LAYER nwell ;
        RECT 35.910 153.595 150.370 156.425 ;
      LAYER pwell ;
        RECT 36.105 152.395 37.475 153.205 ;
        RECT 37.485 152.395 40.235 153.205 ;
        RECT 40.245 152.395 41.615 153.175 ;
        RECT 42.085 152.395 43.455 153.175 ;
        RECT 43.465 152.395 44.835 153.205 ;
        RECT 44.845 152.395 46.195 153.305 ;
        RECT 46.225 153.075 47.145 153.305 ;
        RECT 46.225 152.395 48.515 153.075 ;
        RECT 48.995 152.480 49.425 153.265 ;
        RECT 49.755 153.075 50.685 153.305 ;
        RECT 49.755 152.395 51.590 153.075 ;
        RECT 51.745 152.395 57.255 153.205 ;
        RECT 57.265 152.395 62.775 153.205 ;
        RECT 62.785 152.395 64.615 153.205 ;
        RECT 65.085 153.105 66.035 153.305 ;
        RECT 67.365 153.105 68.295 153.305 ;
        RECT 65.085 152.625 68.295 153.105 ;
        RECT 65.085 152.425 68.150 152.625 ;
        RECT 65.085 152.395 66.020 152.425 ;
        RECT 36.245 152.185 36.415 152.395 ;
        RECT 37.625 152.185 37.795 152.395 ;
        RECT 39.005 152.185 39.175 152.375 ;
        RECT 41.305 152.205 41.475 152.395 ;
        RECT 41.760 152.235 41.880 152.345 ;
        RECT 43.145 152.205 43.315 152.395 ;
        RECT 43.605 152.205 43.775 152.395 ;
        RECT 45.910 152.205 46.080 152.395 ;
        RECT 46.835 152.230 46.995 152.340 ;
        RECT 47.720 152.205 47.890 152.375 ;
        RECT 48.205 152.205 48.375 152.395 ;
        RECT 51.425 152.375 51.590 152.395 ;
        RECT 48.660 152.235 48.780 152.345 ;
        RECT 51.425 152.205 51.595 152.375 ;
        RECT 51.885 152.205 52.055 152.395 ;
        RECT 47.780 152.185 47.890 152.205 ;
        RECT 53.265 152.185 53.435 152.375 ;
        RECT 53.725 152.185 53.895 152.375 ;
        RECT 55.540 152.205 55.710 152.375 ;
        RECT 57.405 152.205 57.575 152.395 ;
        RECT 55.600 152.185 55.710 152.205 ;
        RECT 60.165 152.185 60.335 152.375 ;
        RECT 62.465 152.185 62.635 152.375 ;
        RECT 62.925 152.205 63.095 152.395 ;
        RECT 67.980 152.375 68.150 152.425 ;
        RECT 68.305 152.395 70.135 153.205 ;
        RECT 70.915 153.075 71.845 153.305 ;
        RECT 70.915 152.395 72.750 153.075 ;
        RECT 72.905 152.395 74.735 153.205 ;
        RECT 74.755 152.480 75.185 153.265 ;
        RECT 75.205 152.395 77.955 153.205 ;
        RECT 77.965 152.395 79.335 153.175 ;
        RECT 79.345 152.395 82.555 153.305 ;
        RECT 84.075 153.075 85.005 153.305 ;
        RECT 86.445 153.075 90.375 153.305 ;
        RECT 83.170 152.395 85.005 153.075 ;
        RECT 85.960 152.395 90.375 153.075 ;
        RECT 90.385 152.395 95.895 153.205 ;
        RECT 96.825 152.395 98.195 153.175 ;
        RECT 99.255 153.075 100.185 153.305 ;
        RECT 98.350 152.395 100.185 153.075 ;
        RECT 100.515 152.480 100.945 153.265 ;
        RECT 101.255 152.395 104.175 153.305 ;
        RECT 104.185 152.395 107.105 153.305 ;
        RECT 108.455 153.075 109.385 153.305 ;
        RECT 107.550 152.395 109.385 153.075 ;
        RECT 109.705 152.395 112.625 153.305 ;
        RECT 112.925 152.395 115.845 153.305 ;
        RECT 116.145 152.395 119.345 153.305 ;
        RECT 119.365 152.395 124.875 153.205 ;
        RECT 124.885 152.395 126.255 153.205 ;
        RECT 126.275 152.480 126.705 153.265 ;
        RECT 126.725 152.395 128.935 153.305 ;
        RECT 129.945 153.105 130.875 153.305 ;
        RECT 132.205 153.105 133.155 153.305 ;
        RECT 129.945 152.625 133.155 153.105 ;
        RECT 130.090 152.425 133.155 152.625 ;
        RECT 64.760 152.235 64.880 152.345 ;
        RECT 67.980 152.205 68.155 152.375 ;
        RECT 68.445 152.205 68.615 152.395 ;
        RECT 72.585 152.375 72.750 152.395 ;
        RECT 70.280 152.235 70.400 152.345 ;
        RECT 72.585 152.205 72.755 152.375 ;
        RECT 73.045 152.205 73.215 152.395 ;
        RECT 67.985 152.185 68.155 152.205 ;
        RECT 73.505 152.185 73.675 152.375 ;
        RECT 75.345 152.205 75.515 152.395 ;
        RECT 78.115 152.205 78.285 152.395 ;
        RECT 79.025 152.185 79.195 152.375 ;
        RECT 80.870 152.185 81.040 152.375 ;
        RECT 82.255 152.205 82.425 152.395 ;
        RECT 83.170 152.375 83.335 152.395 ;
        RECT 85.960 152.375 86.070 152.395 ;
        RECT 82.700 152.235 82.820 152.345 ;
        RECT 83.160 152.205 83.335 152.375 ;
        RECT 83.160 152.185 83.330 152.205 ;
        RECT 84.545 152.185 84.715 152.375 ;
        RECT 85.460 152.235 85.580 152.345 ;
        RECT 85.900 152.205 86.095 152.375 ;
        RECT 90.525 152.205 90.695 152.395 ;
        RECT 85.925 152.185 86.095 152.205 ;
        RECT 90.980 152.185 91.150 152.375 ;
        RECT 91.420 152.205 91.590 152.375 ;
        RECT 91.480 152.185 91.590 152.205 ;
        RECT 96.045 152.185 96.215 152.375 ;
        RECT 97.875 152.205 98.045 152.395 ;
        RECT 98.350 152.375 98.515 152.395 ;
        RECT 98.345 152.205 98.515 152.375 ;
        RECT 99.255 152.185 99.425 152.375 ;
        RECT 99.725 152.185 99.895 152.375 ;
        RECT 101.105 152.185 101.275 152.375 ;
        RECT 103.860 152.205 104.030 152.395 ;
        RECT 104.330 152.205 104.500 152.395 ;
        RECT 107.550 152.375 107.715 152.395 ;
        RECT 104.775 152.185 104.945 152.375 ;
        RECT 105.245 152.185 105.415 152.375 ;
        RECT 107.545 152.205 107.715 152.375 ;
        RECT 109.850 152.205 110.020 152.395 ;
        RECT 110.765 152.185 110.935 152.375 ;
        RECT 113.070 152.205 113.240 152.395 ;
        RECT 113.980 152.185 114.150 152.375 ;
        RECT 117.665 152.185 117.835 152.375 ;
        RECT 119.050 152.205 119.220 152.395 ;
        RECT 119.505 152.205 119.675 152.395 ;
        RECT 123.185 152.185 123.355 152.375 ;
        RECT 124.565 152.185 124.735 152.375 ;
        RECT 125.025 152.205 125.195 152.395 ;
        RECT 125.945 152.185 126.115 152.375 ;
        RECT 126.870 152.205 127.040 152.395 ;
        RECT 127.785 152.205 127.955 152.375 ;
        RECT 129.175 152.240 129.335 152.350 ;
        RECT 127.805 152.185 127.955 152.205 ;
        RECT 130.090 152.185 130.260 152.425 ;
        RECT 132.220 152.395 133.155 152.425 ;
        RECT 133.475 153.075 134.405 153.305 ;
        RECT 133.475 152.395 135.310 153.075 ;
        RECT 135.465 152.395 138.215 153.205 ;
        RECT 138.685 152.395 140.055 153.175 ;
        RECT 140.065 152.395 145.575 153.205 ;
        RECT 145.585 152.395 148.335 153.205 ;
        RECT 148.805 152.395 150.175 153.205 ;
        RECT 135.145 152.375 135.310 152.395 ;
        RECT 132.840 152.185 133.010 152.375 ;
        RECT 133.305 152.185 133.475 152.375 ;
        RECT 135.145 152.205 135.315 152.375 ;
        RECT 135.605 152.205 135.775 152.395 ;
        RECT 138.825 152.345 138.995 152.395 ;
        RECT 138.360 152.235 138.480 152.345 ;
        RECT 138.820 152.235 138.995 152.345 ;
        RECT 138.825 152.205 138.995 152.235 ;
        RECT 139.755 152.230 139.915 152.340 ;
        RECT 140.205 152.205 140.375 152.395 ;
        RECT 140.665 152.185 140.835 152.375 ;
        RECT 145.725 152.205 145.895 152.395 ;
        RECT 148.035 152.230 148.195 152.340 ;
        RECT 148.480 152.235 148.600 152.345 ;
        RECT 149.865 152.185 150.035 152.395 ;
        RECT 36.105 151.375 37.475 152.185 ;
        RECT 37.485 151.375 38.855 152.185 ;
        RECT 38.865 151.505 46.595 152.185 ;
        RECT 47.780 151.505 52.195 152.185 ;
        RECT 42.380 151.285 43.290 151.505 ;
        RECT 44.825 151.275 46.595 151.505 ;
        RECT 48.265 151.275 52.195 151.505 ;
        RECT 52.205 151.405 53.575 152.185 ;
        RECT 53.585 151.375 55.415 152.185 ;
        RECT 55.600 151.505 60.015 152.185 ;
        RECT 56.085 151.275 60.015 151.505 ;
        RECT 60.025 151.375 61.855 152.185 ;
        RECT 61.875 151.315 62.305 152.100 ;
        RECT 62.325 151.375 67.835 152.185 ;
        RECT 67.845 151.375 73.355 152.185 ;
        RECT 73.365 151.375 78.875 152.185 ;
        RECT 78.885 151.375 80.715 152.185 ;
        RECT 80.725 151.275 82.555 152.185 ;
        RECT 83.045 151.275 84.395 152.185 ;
        RECT 84.415 151.275 85.765 152.185 ;
        RECT 85.785 151.375 87.615 152.185 ;
        RECT 87.635 151.315 88.065 152.100 ;
        RECT 88.375 151.275 91.295 152.185 ;
        RECT 91.480 151.505 95.895 152.185 ;
        RECT 91.965 151.275 95.895 151.505 ;
        RECT 95.905 151.375 97.735 152.185 ;
        RECT 98.205 151.405 99.575 152.185 ;
        RECT 99.585 151.375 100.955 152.185 ;
        RECT 100.965 151.505 103.715 152.185 ;
        RECT 102.785 151.275 103.715 151.505 ;
        RECT 103.725 151.405 105.095 152.185 ;
        RECT 105.105 151.375 110.615 152.185 ;
        RECT 110.625 151.375 113.375 152.185 ;
        RECT 113.395 151.315 113.825 152.100 ;
        RECT 113.855 151.275 117.515 152.185 ;
        RECT 117.525 151.375 123.035 152.185 ;
        RECT 123.045 151.375 124.415 152.185 ;
        RECT 124.435 151.275 125.785 152.185 ;
        RECT 125.805 151.375 127.635 152.185 ;
        RECT 127.805 151.365 129.735 152.185 ;
        RECT 128.785 151.275 129.735 151.365 ;
        RECT 129.945 151.275 131.775 152.185 ;
        RECT 131.805 151.275 133.155 152.185 ;
        RECT 133.165 151.375 138.675 152.185 ;
        RECT 139.155 151.315 139.585 152.100 ;
        RECT 140.525 151.505 147.835 152.185 ;
        RECT 144.040 151.285 144.950 151.505 ;
        RECT 146.485 151.275 147.835 151.505 ;
        RECT 148.805 151.375 150.175 152.185 ;
      LAYER nwell ;
        RECT 35.910 148.155 150.370 150.985 ;
      LAYER pwell ;
        RECT 36.105 146.955 37.475 147.765 ;
        RECT 37.485 146.955 40.235 147.765 ;
        RECT 40.245 146.955 41.615 147.735 ;
        RECT 41.625 146.955 42.995 147.735 ;
        RECT 43.005 146.955 48.515 147.765 ;
        RECT 48.995 147.040 49.425 147.825 ;
        RECT 53.345 147.775 54.295 147.865 ;
        RECT 49.445 146.955 52.195 147.765 ;
        RECT 52.365 146.955 54.295 147.775 ;
        RECT 54.515 146.955 57.245 147.865 ;
        RECT 57.305 146.955 60.475 147.865 ;
        RECT 60.485 146.955 64.155 147.865 ;
        RECT 64.165 146.955 65.995 147.765 ;
        RECT 66.005 146.955 67.375 147.735 ;
        RECT 67.385 146.955 68.755 147.765 ;
        RECT 68.785 146.955 70.135 147.865 ;
        RECT 70.165 146.955 71.515 147.865 ;
        RECT 71.815 146.955 74.735 147.865 ;
        RECT 74.755 147.040 75.185 147.825 ;
        RECT 75.495 146.955 78.415 147.865 ;
        RECT 79.565 147.775 80.515 147.865 ;
        RECT 78.585 146.955 80.515 147.775 ;
        RECT 82.235 147.635 83.165 147.865 ;
        RECT 81.330 146.955 83.165 147.635 ;
        RECT 84.405 146.955 87.325 147.865 ;
        RECT 87.625 146.955 91.100 147.865 ;
        RECT 91.305 146.955 94.055 147.765 ;
        RECT 94.545 146.955 95.895 147.865 ;
        RECT 95.905 146.955 98.655 147.765 ;
        RECT 98.665 146.955 100.495 147.635 ;
        RECT 100.515 147.040 100.945 147.825 ;
        RECT 100.965 146.955 102.795 147.635 ;
        RECT 102.805 146.955 105.555 147.765 ;
        RECT 105.565 146.955 107.395 147.635 ;
        RECT 107.405 146.955 110.155 147.765 ;
        RECT 110.165 146.955 113.640 147.865 ;
        RECT 114.135 146.955 117.055 147.865 ;
        RECT 118.295 147.635 119.225 147.865 ;
        RECT 118.295 146.955 120.130 147.635 ;
        RECT 120.285 146.955 121.635 147.865 ;
        RECT 122.595 146.955 125.795 147.865 ;
        RECT 126.275 147.040 126.705 147.825 ;
        RECT 126.725 147.665 127.670 147.865 ;
        RECT 126.725 146.985 129.475 147.665 ;
        RECT 126.725 146.955 127.670 146.985 ;
        RECT 36.245 146.745 36.415 146.955 ;
        RECT 37.625 146.765 37.795 146.955 ;
        RECT 39.925 146.745 40.095 146.935 ;
        RECT 40.395 146.790 40.555 146.900 ;
        RECT 41.305 146.765 41.475 146.955 ;
        RECT 42.685 146.765 42.855 146.955 ;
        RECT 43.145 146.765 43.315 146.955 ;
        RECT 43.605 146.745 43.775 146.935 ;
        RECT 44.060 146.795 44.180 146.905 ;
        RECT 44.525 146.745 44.695 146.935 ;
        RECT 48.660 146.795 48.780 146.905 ;
        RECT 49.585 146.765 49.755 146.955 ;
        RECT 52.365 146.935 52.515 146.955 ;
        RECT 51.885 146.745 52.055 146.935 ;
        RECT 52.345 146.765 52.515 146.935 ;
        RECT 55.115 146.745 55.285 146.935 ;
        RECT 56.495 146.790 56.655 146.900 ;
        RECT 56.945 146.765 57.115 146.955 ;
        RECT 57.405 146.745 57.575 146.955 ;
        RECT 60.625 146.745 60.795 146.935 ;
        RECT 62.465 146.745 62.635 146.935 ;
        RECT 63.840 146.765 64.010 146.955 ;
        RECT 64.305 146.905 64.475 146.955 ;
        RECT 64.300 146.795 64.475 146.905 ;
        RECT 64.305 146.765 64.475 146.795 ;
        RECT 64.765 146.765 64.935 146.935 ;
        RECT 66.155 146.765 66.325 146.955 ;
        RECT 67.075 146.790 67.235 146.900 ;
        RECT 67.525 146.765 67.695 146.955 ;
        RECT 64.785 146.745 64.935 146.765 ;
        RECT 68.900 146.745 69.070 146.955 ;
        RECT 70.280 146.745 70.450 146.955 ;
        RECT 70.745 146.745 70.915 146.935 ;
        RECT 72.125 146.745 72.295 146.935 ;
        RECT 74.420 146.765 74.590 146.955 ;
        RECT 75.345 146.745 75.515 146.935 ;
        RECT 78.100 146.765 78.270 146.955 ;
        RECT 78.585 146.935 78.735 146.955 ;
        RECT 81.330 146.935 81.495 146.955 ;
        RECT 78.565 146.745 78.735 146.935 ;
        RECT 80.860 146.795 80.980 146.905 ;
        RECT 81.325 146.765 81.495 146.935 ;
        RECT 82.245 146.745 82.415 146.935 ;
        RECT 83.635 146.800 83.795 146.910 ;
        RECT 84.550 146.765 84.720 146.955 ;
        RECT 87.305 146.745 87.475 146.935 ;
        RECT 87.770 146.765 87.940 146.955 ;
        RECT 88.220 146.795 88.340 146.905 ;
        RECT 88.690 146.745 88.860 146.935 ;
        RECT 91.445 146.765 91.615 146.955 ;
        RECT 92.365 146.745 92.535 146.935 ;
        RECT 94.200 146.795 94.320 146.905 ;
        RECT 94.660 146.765 94.830 146.955 ;
        RECT 96.045 146.765 96.215 146.955 ;
        RECT 96.505 146.745 96.675 146.935 ;
        RECT 96.965 146.745 97.135 146.935 ;
        RECT 98.345 146.745 98.515 146.935 ;
        RECT 100.185 146.765 100.355 146.955 ;
        RECT 101.105 146.745 101.275 146.935 ;
        RECT 102.485 146.765 102.655 146.955 ;
        RECT 102.945 146.765 103.115 146.955 ;
        RECT 104.775 146.745 104.945 146.935 ;
        RECT 105.245 146.745 105.415 146.935 ;
        RECT 105.705 146.765 105.875 146.955 ;
        RECT 107.545 146.765 107.715 146.955 ;
        RECT 108.005 146.745 108.175 146.935 ;
        RECT 109.395 146.745 109.565 146.935 ;
        RECT 110.310 146.765 110.480 146.955 ;
        RECT 113.065 146.745 113.235 146.935 ;
        RECT 116.285 146.745 116.455 146.935 ;
        RECT 116.740 146.765 116.910 146.955 ;
        RECT 119.965 146.935 120.130 146.955 ;
        RECT 117.215 146.800 117.375 146.910 ;
        RECT 119.045 146.745 119.215 146.935 ;
        RECT 119.505 146.745 119.675 146.935 ;
        RECT 119.965 146.765 120.135 146.935 ;
        RECT 121.350 146.765 121.520 146.955 ;
        RECT 121.815 146.800 121.975 146.910 ;
        RECT 122.720 146.765 122.890 146.955 ;
        RECT 129.160 146.935 129.330 146.985 ;
        RECT 129.485 146.955 134.995 147.765 ;
        RECT 135.005 146.955 136.835 147.765 ;
        RECT 136.855 146.955 139.585 147.865 ;
        RECT 139.805 147.775 140.755 147.865 ;
        RECT 139.805 146.955 141.735 147.775 ;
        RECT 141.905 146.955 143.275 147.735 ;
        RECT 143.295 146.955 144.645 147.865 ;
        RECT 144.665 146.955 148.335 147.765 ;
        RECT 148.805 146.955 150.175 147.765 ;
        RECT 123.185 146.745 123.355 146.935 ;
        RECT 125.940 146.795 126.060 146.905 ;
        RECT 129.160 146.765 129.335 146.935 ;
        RECT 129.165 146.745 129.335 146.765 ;
        RECT 129.625 146.745 129.795 146.955 ;
        RECT 131.460 146.795 131.580 146.905 ;
        RECT 131.925 146.745 132.095 146.935 ;
        RECT 135.145 146.765 135.315 146.955 ;
        RECT 136.985 146.765 137.155 146.955 ;
        RECT 141.585 146.935 141.735 146.955 ;
        RECT 139.745 146.745 139.915 146.935 ;
        RECT 141.585 146.765 141.755 146.935 ;
        RECT 142.955 146.765 143.125 146.955 ;
        RECT 144.345 146.765 144.515 146.955 ;
        RECT 144.805 146.765 144.975 146.955 ;
        RECT 145.725 146.745 145.895 146.935 ;
        RECT 147.565 146.745 147.735 146.935 ;
        RECT 148.480 146.795 148.600 146.905 ;
        RECT 149.865 146.745 150.035 146.955 ;
        RECT 36.105 145.935 37.475 146.745 ;
        RECT 37.495 146.065 40.235 146.745 ;
        RECT 41.175 146.065 43.915 146.745 ;
        RECT 44.385 146.065 51.695 146.745 ;
        RECT 47.900 145.845 48.810 146.065 ;
        RECT 50.345 145.835 51.695 146.065 ;
        RECT 51.785 145.835 54.955 146.745 ;
        RECT 54.965 145.965 56.335 146.745 ;
        RECT 57.365 145.835 60.475 146.745 ;
        RECT 60.485 145.935 61.855 146.745 ;
        RECT 61.875 145.875 62.305 146.660 ;
        RECT 62.325 145.935 64.155 146.745 ;
        RECT 64.785 145.925 66.715 146.745 ;
        RECT 65.765 145.835 66.715 145.925 ;
        RECT 67.865 145.835 69.215 146.745 ;
        RECT 69.245 145.835 70.595 146.745 ;
        RECT 70.605 145.935 71.975 146.745 ;
        RECT 72.065 145.835 75.065 146.745 ;
        RECT 75.205 145.835 77.955 146.745 ;
        RECT 78.425 145.835 81.175 146.745 ;
        RECT 82.105 145.835 84.855 146.745 ;
        RECT 84.865 145.835 87.615 146.745 ;
        RECT 87.635 145.875 88.065 146.660 ;
        RECT 88.545 145.835 92.020 146.745 ;
        RECT 92.225 145.935 94.055 146.745 ;
        RECT 94.065 145.835 96.815 146.745 ;
        RECT 96.825 145.935 98.195 146.745 ;
        RECT 98.205 145.835 100.955 146.745 ;
        RECT 100.965 145.835 103.715 146.745 ;
        RECT 103.725 145.965 105.095 146.745 ;
        RECT 105.105 145.835 107.855 146.745 ;
        RECT 107.865 145.965 109.235 146.745 ;
        RECT 109.245 145.965 110.615 146.745 ;
        RECT 110.625 145.835 113.375 146.745 ;
        RECT 113.395 145.875 113.825 146.660 ;
        RECT 113.845 145.835 116.595 146.745 ;
        RECT 116.605 145.835 119.355 146.745 ;
        RECT 119.365 145.965 120.735 146.745 ;
        RECT 120.745 145.835 123.495 146.745 ;
        RECT 123.655 145.835 129.475 146.745 ;
        RECT 129.485 145.935 131.315 146.745 ;
        RECT 131.785 146.065 139.095 146.745 ;
        RECT 135.300 145.845 136.210 146.065 ;
        RECT 137.745 145.835 139.095 146.065 ;
        RECT 139.155 145.875 139.585 146.660 ;
        RECT 139.605 145.835 145.425 146.745 ;
        RECT 145.585 146.065 147.415 146.745 ;
        RECT 146.070 145.835 147.415 146.065 ;
        RECT 147.425 145.935 148.795 146.745 ;
        RECT 148.805 145.935 150.175 146.745 ;
      LAYER nwell ;
        RECT 35.910 142.715 150.370 145.545 ;
      LAYER pwell ;
        RECT 36.105 141.515 37.475 142.325 ;
        RECT 37.945 142.195 39.290 142.425 ;
        RECT 43.760 142.195 44.670 142.415 ;
        RECT 46.205 142.195 47.555 142.425 ;
        RECT 37.945 141.515 39.775 142.195 ;
        RECT 40.245 141.515 47.555 142.195 ;
        RECT 47.605 141.515 48.975 142.325 ;
        RECT 48.995 141.600 49.425 142.385 ;
        RECT 49.445 142.195 50.790 142.425 ;
        RECT 54.505 142.195 55.850 142.425 ;
        RECT 49.445 141.515 51.275 142.195 ;
        RECT 51.295 141.515 54.035 142.195 ;
        RECT 54.505 141.515 56.335 142.195 ;
        RECT 56.345 141.515 58.175 142.325 ;
        RECT 58.645 142.195 59.990 142.425 ;
        RECT 58.645 141.515 60.475 142.195 ;
        RECT 60.485 141.515 61.855 142.325 ;
        RECT 61.875 141.600 62.305 142.385 ;
        RECT 62.785 142.195 64.130 142.425 ;
        RECT 62.785 141.515 64.615 142.195 ;
        RECT 64.625 141.515 70.135 142.325 ;
        RECT 70.145 141.515 73.815 142.325 ;
        RECT 74.755 141.600 75.185 142.385 ;
        RECT 75.205 142.195 76.550 142.425 ;
        RECT 75.205 141.515 77.035 142.195 ;
        RECT 77.505 141.515 78.875 142.295 ;
        RECT 79.830 142.195 81.175 142.425 ;
        RECT 79.345 141.515 81.175 142.195 ;
        RECT 81.185 141.515 82.555 142.295 ;
        RECT 83.970 142.195 85.315 142.425 ;
        RECT 83.485 141.515 85.315 142.195 ;
        RECT 85.325 141.515 87.155 142.325 ;
        RECT 87.635 141.600 88.065 142.385 ;
        RECT 88.085 141.515 90.825 142.195 ;
        RECT 91.305 141.515 94.055 142.425 ;
        RECT 94.550 142.195 95.895 142.425 ;
        RECT 94.065 141.515 95.895 142.195 ;
        RECT 95.905 142.195 97.250 142.425 ;
        RECT 95.905 141.515 97.735 142.195 ;
        RECT 97.745 141.515 100.495 142.325 ;
        RECT 100.515 141.600 100.945 142.385 ;
        RECT 101.450 142.195 102.795 142.425 ;
        RECT 100.965 141.515 102.795 142.195 ;
        RECT 102.805 141.515 104.175 142.325 ;
        RECT 104.185 142.195 105.530 142.425 ;
        RECT 104.185 141.515 106.015 142.195 ;
        RECT 106.025 141.515 111.535 142.325 ;
        RECT 111.545 141.515 113.375 142.325 ;
        RECT 113.395 141.600 113.825 142.385 ;
        RECT 113.845 141.515 116.595 142.425 ;
        RECT 117.090 142.195 118.435 142.425 ;
        RECT 116.605 141.515 118.435 142.195 ;
        RECT 118.445 141.515 120.275 142.325 ;
        RECT 121.230 142.195 122.575 142.425 ;
        RECT 120.745 141.515 122.575 142.195 ;
        RECT 122.585 141.515 124.415 142.325 ;
        RECT 124.910 142.195 126.255 142.425 ;
        RECT 124.425 141.515 126.255 142.195 ;
        RECT 126.275 141.600 126.705 142.385 ;
        RECT 126.725 141.515 129.475 142.425 ;
        RECT 133.650 142.195 134.995 142.425 ;
        RECT 129.485 141.515 132.225 142.195 ;
        RECT 133.165 141.515 134.995 142.195 ;
        RECT 135.005 141.515 136.835 142.325 ;
        RECT 137.790 142.195 139.135 142.425 ;
        RECT 137.305 141.515 139.135 142.195 ;
        RECT 139.155 141.600 139.585 142.385 ;
        RECT 140.195 141.515 146.035 142.425 ;
        RECT 146.530 142.195 147.875 142.425 ;
        RECT 146.045 141.515 147.875 142.195 ;
        RECT 148.805 141.515 150.175 142.325 ;
        RECT 36.245 141.325 36.415 141.515 ;
        RECT 37.620 141.355 37.740 141.465 ;
        RECT 39.465 141.325 39.635 141.515 ;
        RECT 39.920 141.355 40.040 141.465 ;
        RECT 40.385 141.325 40.555 141.515 ;
        RECT 47.745 141.325 47.915 141.515 ;
        RECT 50.965 141.325 51.135 141.515 ;
        RECT 53.725 141.325 53.895 141.515 ;
        RECT 54.180 141.355 54.300 141.465 ;
        RECT 56.025 141.325 56.195 141.515 ;
        RECT 56.485 141.325 56.655 141.515 ;
        RECT 58.320 141.355 58.440 141.465 ;
        RECT 60.165 141.325 60.335 141.515 ;
        RECT 60.625 141.325 60.795 141.515 ;
        RECT 62.460 141.355 62.580 141.465 ;
        RECT 64.305 141.325 64.475 141.515 ;
        RECT 64.765 141.325 64.935 141.515 ;
        RECT 70.285 141.325 70.455 141.515 ;
        RECT 73.975 141.360 74.135 141.470 ;
        RECT 76.725 141.325 76.895 141.515 ;
        RECT 77.180 141.355 77.300 141.465 ;
        RECT 77.645 141.325 77.815 141.515 ;
        RECT 79.020 141.355 79.140 141.465 ;
        RECT 79.485 141.325 79.655 141.515 ;
        RECT 82.245 141.325 82.415 141.515 ;
        RECT 82.715 141.360 82.875 141.470 ;
        RECT 83.625 141.325 83.795 141.515 ;
        RECT 85.465 141.325 85.635 141.515 ;
        RECT 87.300 141.355 87.420 141.465 ;
        RECT 88.225 141.325 88.395 141.515 ;
        RECT 90.980 141.355 91.100 141.465 ;
        RECT 93.745 141.325 93.915 141.515 ;
        RECT 94.205 141.325 94.375 141.515 ;
        RECT 97.425 141.325 97.595 141.515 ;
        RECT 97.885 141.325 98.055 141.515 ;
        RECT 101.105 141.325 101.275 141.515 ;
        RECT 102.945 141.325 103.115 141.515 ;
        RECT 105.705 141.325 105.875 141.515 ;
        RECT 106.165 141.325 106.335 141.515 ;
        RECT 111.685 141.325 111.855 141.515 ;
        RECT 116.285 141.325 116.455 141.515 ;
        RECT 116.745 141.325 116.915 141.515 ;
        RECT 118.585 141.325 118.755 141.515 ;
        RECT 120.420 141.355 120.540 141.465 ;
        RECT 120.885 141.325 121.055 141.515 ;
        RECT 122.725 141.325 122.895 141.515 ;
        RECT 124.565 141.325 124.735 141.515 ;
        RECT 129.165 141.325 129.335 141.515 ;
        RECT 129.625 141.325 129.795 141.515 ;
        RECT 132.395 141.360 132.555 141.470 ;
        RECT 133.305 141.325 133.475 141.515 ;
        RECT 135.145 141.325 135.315 141.515 ;
        RECT 136.980 141.355 137.100 141.465 ;
        RECT 137.445 141.325 137.615 141.515 ;
        RECT 139.740 141.355 139.860 141.465 ;
        RECT 145.725 141.325 145.895 141.515 ;
        RECT 146.185 141.325 146.355 141.515 ;
        RECT 148.035 141.360 148.195 141.470 ;
        RECT 149.865 141.325 150.035 141.515 ;
        RECT 33.930 83.110 36.280 128.830 ;
        RECT 37.930 83.110 40.280 128.830 ;
        RECT 41.930 83.110 44.280 128.830 ;
        RECT 45.930 83.110 48.280 128.830 ;
        RECT 49.930 83.110 52.280 128.830 ;
        RECT 53.930 83.110 56.280 128.830 ;
        RECT 57.930 83.110 60.280 128.830 ;
        RECT 61.930 83.110 64.280 128.830 ;
        RECT 74.930 83.110 77.280 128.830 ;
        RECT 78.930 83.110 81.280 128.830 ;
        RECT 82.930 83.110 85.280 128.830 ;
        RECT 86.930 83.110 89.280 128.830 ;
        RECT 90.930 83.110 93.280 128.830 ;
        RECT 94.930 83.110 97.280 128.830 ;
        RECT 98.930 83.110 101.280 128.830 ;
        RECT 102.930 83.110 105.280 128.830 ;
        RECT 115.930 83.110 118.280 128.830 ;
        RECT 119.930 83.110 122.280 128.830 ;
        RECT 123.930 83.110 126.280 128.830 ;
        RECT 127.930 83.110 130.280 128.830 ;
        RECT 131.930 83.110 134.280 128.830 ;
        RECT 135.930 83.110 138.280 128.830 ;
        RECT 139.930 83.110 142.280 128.830 ;
        RECT 143.930 83.110 146.280 128.830 ;
        RECT 33.930 55.460 36.280 80.830 ;
        RECT 37.930 55.460 40.280 80.830 ;
        RECT 41.930 55.460 44.280 80.830 ;
        RECT 45.930 55.460 48.280 80.830 ;
        RECT 49.930 55.460 52.280 80.830 ;
        RECT 53.930 55.460 56.280 80.830 ;
        RECT 57.930 55.460 60.280 80.830 ;
        RECT 61.930 55.460 64.280 80.830 ;
        RECT 74.930 55.460 77.280 80.830 ;
        RECT 78.930 55.460 81.280 80.830 ;
        RECT 82.930 55.460 85.280 80.830 ;
        RECT 86.930 55.460 89.280 80.830 ;
        RECT 90.930 55.460 93.280 80.830 ;
        RECT 94.930 55.460 97.280 80.830 ;
        RECT 98.930 55.460 101.280 80.830 ;
        RECT 102.930 55.460 105.280 80.830 ;
        RECT 115.930 55.460 118.280 80.830 ;
        RECT 119.930 55.460 122.280 80.830 ;
        RECT 123.930 55.460 126.280 80.830 ;
        RECT 127.930 55.460 130.280 80.830 ;
        RECT 131.930 55.460 134.280 80.830 ;
        RECT 135.930 55.460 138.280 80.830 ;
        RECT 139.930 55.460 142.280 80.830 ;
        RECT 143.930 55.460 146.280 80.830 ;
      LAYER nwell ;
        RECT 26.685 10.800 28.795 20.990 ;
      LAYER pwell ;
        RECT 29.500 12.865 31.610 18.965 ;
      LAYER li1 ;
        RECT 36.100 214.765 150.180 214.935 ;
        RECT 36.185 213.675 37.395 214.765 ;
        RECT 37.565 214.330 42.910 214.765 ;
        RECT 36.185 212.965 36.705 213.505 ;
        RECT 36.875 213.135 37.395 213.675 ;
        RECT 36.185 212.215 37.395 212.965 ;
        RECT 39.150 212.760 39.490 213.590 ;
        RECT 40.970 213.080 41.320 214.330 ;
        RECT 43.085 213.675 44.755 214.765 ;
        RECT 45.040 214.135 45.325 214.595 ;
        RECT 45.495 214.305 45.765 214.765 ;
        RECT 45.040 213.915 45.995 214.135 ;
        RECT 43.085 212.985 43.835 213.505 ;
        RECT 44.005 213.155 44.755 213.675 ;
        RECT 44.925 213.185 45.615 213.745 ;
        RECT 45.785 213.015 45.995 213.915 ;
        RECT 37.565 212.215 42.910 212.760 ;
        RECT 43.085 212.215 44.755 212.985 ;
        RECT 45.040 212.845 45.995 213.015 ;
        RECT 46.165 213.745 46.565 214.595 ;
        RECT 46.755 214.135 47.035 214.595 ;
        RECT 47.555 214.305 47.880 214.765 ;
        RECT 46.755 213.915 47.880 214.135 ;
        RECT 46.165 213.185 47.260 213.745 ;
        RECT 47.430 213.455 47.880 213.915 ;
        RECT 48.050 213.625 48.435 214.595 ;
        RECT 45.040 212.385 45.325 212.845 ;
        RECT 45.495 212.215 45.765 212.675 ;
        RECT 46.165 212.385 46.565 213.185 ;
        RECT 47.430 213.125 47.985 213.455 ;
        RECT 47.430 213.015 47.880 213.125 ;
        RECT 46.755 212.845 47.880 213.015 ;
        RECT 48.155 212.955 48.435 213.625 ;
        RECT 49.065 213.600 49.355 214.765 ;
        RECT 49.525 214.330 54.870 214.765 ;
        RECT 46.755 212.385 47.035 212.845 ;
        RECT 47.555 212.215 47.880 212.675 ;
        RECT 48.050 212.385 48.435 212.955 ;
        RECT 49.065 212.215 49.355 212.940 ;
        RECT 51.110 212.760 51.450 213.590 ;
        RECT 52.930 213.080 53.280 214.330 ;
        RECT 55.970 213.615 56.230 214.765 ;
        RECT 56.405 213.690 56.660 214.595 ;
        RECT 56.830 214.005 57.160 214.765 ;
        RECT 57.375 213.835 57.545 214.595 ;
        RECT 58.780 213.895 59.065 214.765 ;
        RECT 59.235 214.135 59.495 214.595 ;
        RECT 59.670 214.305 59.925 214.765 ;
        RECT 60.095 214.135 60.355 214.595 ;
        RECT 59.235 213.965 60.355 214.135 ;
        RECT 60.525 213.965 60.835 214.765 ;
        RECT 49.525 212.215 54.870 212.760 ;
        RECT 55.970 212.215 56.230 213.055 ;
        RECT 56.405 212.960 56.575 213.690 ;
        RECT 56.830 213.665 57.545 213.835 ;
        RECT 59.235 213.715 59.495 213.965 ;
        RECT 61.005 213.795 61.315 214.595 ;
        RECT 56.830 213.455 57.000 213.665 ;
        RECT 58.740 213.545 59.495 213.715 ;
        RECT 60.285 213.625 61.315 213.795 ;
        RECT 56.745 213.125 57.000 213.455 ;
        RECT 56.405 212.385 56.660 212.960 ;
        RECT 56.830 212.935 57.000 213.125 ;
        RECT 57.280 213.115 57.635 213.485 ;
        RECT 58.740 213.035 59.145 213.545 ;
        RECT 60.285 213.375 60.455 213.625 ;
        RECT 59.315 213.205 60.455 213.375 ;
        RECT 56.830 212.765 57.545 212.935 ;
        RECT 58.740 212.865 60.390 213.035 ;
        RECT 60.625 212.885 60.975 213.455 ;
        RECT 56.830 212.215 57.160 212.595 ;
        RECT 57.375 212.385 57.545 212.765 ;
        RECT 58.785 212.215 59.065 212.695 ;
        RECT 59.235 212.475 59.495 212.865 ;
        RECT 59.670 212.215 59.925 212.695 ;
        RECT 60.095 212.475 60.390 212.865 ;
        RECT 61.145 212.715 61.315 213.625 ;
        RECT 61.945 213.600 62.235 214.765 ;
        RECT 63.415 213.835 63.585 214.595 ;
        RECT 63.800 214.005 64.130 214.765 ;
        RECT 63.415 213.665 64.130 213.835 ;
        RECT 64.300 213.690 64.555 214.595 ;
        RECT 63.325 213.115 63.680 213.485 ;
        RECT 63.960 213.455 64.130 213.665 ;
        RECT 63.960 213.125 64.215 213.455 ;
        RECT 60.570 212.215 60.845 212.695 ;
        RECT 61.015 212.385 61.315 212.715 ;
        RECT 61.945 212.215 62.235 212.940 ;
        RECT 63.960 212.935 64.130 213.125 ;
        RECT 64.385 212.960 64.555 213.690 ;
        RECT 64.730 213.615 64.990 214.765 ;
        RECT 66.140 213.895 66.425 214.765 ;
        RECT 66.595 214.135 66.855 214.595 ;
        RECT 67.030 214.305 67.285 214.765 ;
        RECT 67.455 214.135 67.715 214.595 ;
        RECT 66.595 213.965 67.715 214.135 ;
        RECT 67.885 213.965 68.195 214.765 ;
        RECT 66.595 213.715 66.855 213.965 ;
        RECT 68.365 213.795 68.675 214.595 ;
        RECT 66.100 213.545 66.855 213.715 ;
        RECT 67.645 213.625 68.675 213.795 ;
        RECT 68.845 213.675 70.515 214.765 ;
        RECT 63.415 212.765 64.130 212.935 ;
        RECT 63.415 212.385 63.585 212.765 ;
        RECT 63.800 212.215 64.130 212.595 ;
        RECT 64.300 212.385 64.555 212.960 ;
        RECT 64.730 212.215 64.990 213.055 ;
        RECT 66.100 213.035 66.505 213.545 ;
        RECT 67.645 213.375 67.815 213.625 ;
        RECT 66.675 213.205 67.815 213.375 ;
        RECT 66.100 212.865 67.750 213.035 ;
        RECT 67.985 212.885 68.335 213.455 ;
        RECT 66.145 212.215 66.425 212.695 ;
        RECT 66.595 212.475 66.855 212.865 ;
        RECT 67.030 212.215 67.285 212.695 ;
        RECT 67.455 212.475 67.750 212.865 ;
        RECT 68.505 212.715 68.675 213.625 ;
        RECT 67.930 212.215 68.205 212.695 ;
        RECT 68.375 212.385 68.675 212.715 ;
        RECT 68.845 212.985 69.595 213.505 ;
        RECT 69.765 213.155 70.515 213.675 ;
        RECT 70.690 213.615 70.950 214.765 ;
        RECT 71.125 213.690 71.380 214.595 ;
        RECT 71.550 214.005 71.880 214.765 ;
        RECT 72.095 213.835 72.265 214.595 ;
        RECT 68.845 212.215 70.515 212.985 ;
        RECT 70.690 212.215 70.950 213.055 ;
        RECT 71.125 212.960 71.295 213.690 ;
        RECT 71.550 213.665 72.265 213.835 ;
        RECT 72.535 213.795 72.865 214.580 ;
        RECT 71.550 213.455 71.720 213.665 ;
        RECT 72.535 213.625 73.215 213.795 ;
        RECT 73.395 213.625 73.725 214.765 ;
        RECT 71.465 213.125 71.720 213.455 ;
        RECT 71.125 212.385 71.380 212.960 ;
        RECT 71.550 212.935 71.720 213.125 ;
        RECT 72.000 213.115 72.355 213.485 ;
        RECT 72.525 213.205 72.875 213.455 ;
        RECT 73.045 213.025 73.215 213.625 ;
        RECT 74.825 213.600 75.115 214.765 ;
        RECT 75.340 213.895 75.625 214.765 ;
        RECT 75.795 214.135 76.055 214.595 ;
        RECT 76.230 214.305 76.485 214.765 ;
        RECT 76.655 214.135 76.915 214.595 ;
        RECT 75.795 213.965 76.915 214.135 ;
        RECT 77.085 213.965 77.395 214.765 ;
        RECT 75.795 213.715 76.055 213.965 ;
        RECT 77.565 213.795 77.875 214.595 ;
        RECT 75.300 213.545 76.055 213.715 ;
        RECT 76.845 213.625 77.875 213.795 ;
        RECT 78.135 213.835 78.305 214.595 ;
        RECT 78.520 214.005 78.850 214.765 ;
        RECT 78.135 213.665 78.850 213.835 ;
        RECT 79.020 213.690 79.275 214.595 ;
        RECT 73.385 213.205 73.735 213.455 ;
        RECT 75.300 213.035 75.705 213.545 ;
        RECT 76.845 213.375 77.015 213.625 ;
        RECT 75.875 213.205 77.015 213.375 ;
        RECT 71.550 212.765 72.265 212.935 ;
        RECT 71.550 212.215 71.880 212.595 ;
        RECT 72.095 212.385 72.265 212.765 ;
        RECT 72.545 212.215 72.785 213.025 ;
        RECT 72.955 212.385 73.285 213.025 ;
        RECT 73.455 212.215 73.725 213.025 ;
        RECT 74.825 212.215 75.115 212.940 ;
        RECT 75.300 212.865 76.950 213.035 ;
        RECT 77.185 212.885 77.535 213.455 ;
        RECT 75.345 212.215 75.625 212.695 ;
        RECT 75.795 212.475 76.055 212.865 ;
        RECT 76.230 212.215 76.485 212.695 ;
        RECT 76.655 212.475 76.950 212.865 ;
        RECT 77.705 212.715 77.875 213.625 ;
        RECT 78.045 213.115 78.400 213.485 ;
        RECT 78.680 213.455 78.850 213.665 ;
        RECT 78.680 213.125 78.935 213.455 ;
        RECT 78.680 212.935 78.850 213.125 ;
        RECT 79.105 212.960 79.275 213.690 ;
        RECT 79.450 213.615 79.710 214.765 ;
        RECT 80.860 213.895 81.145 214.765 ;
        RECT 81.315 214.135 81.575 214.595 ;
        RECT 81.750 214.305 82.005 214.765 ;
        RECT 82.175 214.135 82.435 214.595 ;
        RECT 81.315 213.965 82.435 214.135 ;
        RECT 82.605 213.965 82.915 214.765 ;
        RECT 81.315 213.715 81.575 213.965 ;
        RECT 83.085 213.795 83.395 214.595 ;
        RECT 80.820 213.545 81.575 213.715 ;
        RECT 82.365 213.625 83.395 213.795 ;
        RECT 83.565 213.675 85.235 214.765 ;
        RECT 77.130 212.215 77.405 212.695 ;
        RECT 77.575 212.385 77.875 212.715 ;
        RECT 78.135 212.765 78.850 212.935 ;
        RECT 78.135 212.385 78.305 212.765 ;
        RECT 78.520 212.215 78.850 212.595 ;
        RECT 79.020 212.385 79.275 212.960 ;
        RECT 79.450 212.215 79.710 213.055 ;
        RECT 80.820 213.035 81.225 213.545 ;
        RECT 82.365 213.375 82.535 213.625 ;
        RECT 81.395 213.205 82.535 213.375 ;
        RECT 80.820 212.865 82.470 213.035 ;
        RECT 82.705 212.885 83.055 213.455 ;
        RECT 80.865 212.215 81.145 212.695 ;
        RECT 81.315 212.475 81.575 212.865 ;
        RECT 81.750 212.215 82.005 212.695 ;
        RECT 82.175 212.475 82.470 212.865 ;
        RECT 83.225 212.715 83.395 213.625 ;
        RECT 82.650 212.215 82.925 212.695 ;
        RECT 83.095 212.385 83.395 212.715 ;
        RECT 83.565 212.985 84.315 213.505 ;
        RECT 84.485 213.155 85.235 213.675 ;
        RECT 85.410 213.615 85.670 214.765 ;
        RECT 85.845 213.690 86.100 214.595 ;
        RECT 86.270 214.005 86.600 214.765 ;
        RECT 86.815 213.835 86.985 214.595 ;
        RECT 83.565 212.215 85.235 212.985 ;
        RECT 85.410 212.215 85.670 213.055 ;
        RECT 85.845 212.960 86.015 213.690 ;
        RECT 86.270 213.665 86.985 213.835 ;
        RECT 86.270 213.455 86.440 213.665 ;
        RECT 87.705 213.600 87.995 214.765 ;
        RECT 88.220 213.895 88.505 214.765 ;
        RECT 88.675 214.135 88.935 214.595 ;
        RECT 89.110 214.305 89.365 214.765 ;
        RECT 89.535 214.135 89.795 214.595 ;
        RECT 88.675 213.965 89.795 214.135 ;
        RECT 89.965 213.965 90.275 214.765 ;
        RECT 88.675 213.715 88.935 213.965 ;
        RECT 90.445 213.795 90.755 214.595 ;
        RECT 90.925 214.330 96.270 214.765 ;
        RECT 88.180 213.545 88.935 213.715 ;
        RECT 89.725 213.625 90.755 213.795 ;
        RECT 86.185 213.125 86.440 213.455 ;
        RECT 85.845 212.385 86.100 212.960 ;
        RECT 86.270 212.935 86.440 213.125 ;
        RECT 86.720 213.115 87.075 213.485 ;
        RECT 88.180 213.035 88.585 213.545 ;
        RECT 89.725 213.375 89.895 213.625 ;
        RECT 88.755 213.205 89.895 213.375 ;
        RECT 86.270 212.765 86.985 212.935 ;
        RECT 86.270 212.215 86.600 212.595 ;
        RECT 86.815 212.385 86.985 212.765 ;
        RECT 87.705 212.215 87.995 212.940 ;
        RECT 88.180 212.865 89.830 213.035 ;
        RECT 90.065 212.885 90.415 213.455 ;
        RECT 88.225 212.215 88.505 212.695 ;
        RECT 88.675 212.475 88.935 212.865 ;
        RECT 89.110 212.215 89.365 212.695 ;
        RECT 89.535 212.475 89.830 212.865 ;
        RECT 90.585 212.715 90.755 213.625 ;
        RECT 92.510 212.760 92.850 213.590 ;
        RECT 94.330 213.080 94.680 214.330 ;
        RECT 96.445 213.675 98.115 214.765 ;
        RECT 96.445 212.985 97.195 213.505 ;
        RECT 97.365 213.155 98.115 213.675 ;
        RECT 98.345 213.625 98.555 214.765 ;
        RECT 98.725 213.615 99.055 214.595 ;
        RECT 99.225 213.625 99.455 214.765 ;
        RECT 90.010 212.215 90.285 212.695 ;
        RECT 90.455 212.385 90.755 212.715 ;
        RECT 90.925 212.215 96.270 212.760 ;
        RECT 96.445 212.215 98.115 212.985 ;
        RECT 98.345 212.215 98.555 213.035 ;
        RECT 98.725 213.015 98.975 213.615 ;
        RECT 100.585 213.600 100.875 214.765 ;
        RECT 101.045 214.170 101.480 214.595 ;
        RECT 101.650 214.340 102.035 214.765 ;
        RECT 101.045 214.000 102.035 214.170 ;
        RECT 99.145 213.205 99.475 213.455 ;
        RECT 101.045 213.125 101.530 213.830 ;
        RECT 101.700 213.455 102.035 214.000 ;
        RECT 102.205 213.805 102.630 214.595 ;
        RECT 102.800 214.170 103.075 214.595 ;
        RECT 103.245 214.340 103.630 214.765 ;
        RECT 102.800 213.975 103.630 214.170 ;
        RECT 102.205 213.625 103.110 213.805 ;
        RECT 101.700 213.125 102.110 213.455 ;
        RECT 102.280 213.125 103.110 213.625 ;
        RECT 103.280 213.455 103.630 213.975 ;
        RECT 103.800 213.805 104.045 214.595 ;
        RECT 104.235 214.170 104.490 214.595 ;
        RECT 104.660 214.340 105.045 214.765 ;
        RECT 104.235 213.975 105.045 214.170 ;
        RECT 103.800 213.625 104.525 213.805 ;
        RECT 103.280 213.125 103.705 213.455 ;
        RECT 103.875 213.125 104.525 213.625 ;
        RECT 104.695 213.455 105.045 213.975 ;
        RECT 105.215 213.625 105.475 214.595 ;
        RECT 105.645 214.330 110.990 214.765 ;
        RECT 104.695 213.125 105.120 213.455 ;
        RECT 98.725 212.385 99.055 213.015 ;
        RECT 99.225 212.215 99.455 213.035 ;
        RECT 101.700 212.955 102.035 213.125 ;
        RECT 102.280 212.955 102.630 213.125 ;
        RECT 103.280 212.955 103.630 213.125 ;
        RECT 103.875 212.955 104.045 213.125 ;
        RECT 104.695 212.955 105.045 213.125 ;
        RECT 105.290 212.955 105.475 213.625 ;
        RECT 100.585 212.215 100.875 212.940 ;
        RECT 101.045 212.785 102.035 212.955 ;
        RECT 101.045 212.385 101.480 212.785 ;
        RECT 101.650 212.215 102.035 212.615 ;
        RECT 102.205 212.385 102.630 212.955 ;
        RECT 102.820 212.785 103.630 212.955 ;
        RECT 102.820 212.385 103.075 212.785 ;
        RECT 103.245 212.215 103.630 212.615 ;
        RECT 103.800 212.385 104.045 212.955 ;
        RECT 104.235 212.785 105.045 212.955 ;
        RECT 104.235 212.385 104.490 212.785 ;
        RECT 104.660 212.215 105.045 212.615 ;
        RECT 105.215 212.385 105.475 212.955 ;
        RECT 107.230 212.760 107.570 213.590 ;
        RECT 109.050 213.080 109.400 214.330 ;
        RECT 111.165 213.675 112.835 214.765 ;
        RECT 111.165 212.985 111.915 213.505 ;
        RECT 112.085 213.155 112.835 213.675 ;
        RECT 113.465 213.600 113.755 214.765 ;
        RECT 113.930 213.625 114.265 214.595 ;
        RECT 114.435 213.625 114.605 214.765 ;
        RECT 114.775 214.425 116.805 214.595 ;
        RECT 105.645 212.215 110.990 212.760 ;
        RECT 111.165 212.215 112.835 212.985 ;
        RECT 113.930 212.955 114.100 213.625 ;
        RECT 114.775 213.455 114.945 214.425 ;
        RECT 114.270 213.125 114.525 213.455 ;
        RECT 114.750 213.125 114.945 213.455 ;
        RECT 115.115 214.085 116.240 214.255 ;
        RECT 114.355 212.955 114.525 213.125 ;
        RECT 115.115 212.955 115.285 214.085 ;
        RECT 113.465 212.215 113.755 212.940 ;
        RECT 113.930 212.385 114.185 212.955 ;
        RECT 114.355 212.785 115.285 212.955 ;
        RECT 115.455 213.745 116.465 213.915 ;
        RECT 115.455 212.945 115.625 213.745 ;
        RECT 115.830 213.065 116.105 213.545 ;
        RECT 115.825 212.895 116.105 213.065 ;
        RECT 115.110 212.750 115.285 212.785 ;
        RECT 114.355 212.215 114.685 212.615 ;
        RECT 115.110 212.385 115.640 212.750 ;
        RECT 115.830 212.385 116.105 212.895 ;
        RECT 116.275 212.385 116.465 213.745 ;
        RECT 116.635 213.760 116.805 214.425 ;
        RECT 116.975 214.005 117.145 214.765 ;
        RECT 117.380 214.005 117.895 214.415 ;
        RECT 116.635 213.570 117.385 213.760 ;
        RECT 117.555 213.195 117.895 214.005 ;
        RECT 118.065 213.675 121.575 214.765 ;
        RECT 116.665 213.025 117.895 213.195 ;
        RECT 116.645 212.215 117.155 212.750 ;
        RECT 117.375 212.420 117.620 213.025 ;
        RECT 118.065 212.985 119.715 213.505 ;
        RECT 119.885 213.155 121.575 213.675 ;
        RECT 122.295 213.835 122.465 214.595 ;
        RECT 122.645 214.005 122.975 214.765 ;
        RECT 122.295 213.665 122.960 213.835 ;
        RECT 123.145 213.690 123.415 214.595 ;
        RECT 122.790 213.520 122.960 213.665 ;
        RECT 122.225 213.115 122.555 213.485 ;
        RECT 122.790 213.190 123.075 213.520 ;
        RECT 118.065 212.215 121.575 212.985 ;
        RECT 122.790 212.935 122.960 213.190 ;
        RECT 122.295 212.765 122.960 212.935 ;
        RECT 123.245 212.890 123.415 213.690 ;
        RECT 123.585 213.675 126.175 214.765 ;
        RECT 122.295 212.385 122.465 212.765 ;
        RECT 122.645 212.215 122.975 212.595 ;
        RECT 123.155 212.385 123.415 212.890 ;
        RECT 123.585 212.985 124.795 213.505 ;
        RECT 124.965 213.155 126.175 213.675 ;
        RECT 126.345 213.600 126.635 214.765 ;
        RECT 126.895 213.835 127.065 214.595 ;
        RECT 127.245 214.005 127.575 214.765 ;
        RECT 126.895 213.665 127.560 213.835 ;
        RECT 127.745 213.690 128.015 214.595 ;
        RECT 127.390 213.520 127.560 213.665 ;
        RECT 126.825 213.115 127.155 213.485 ;
        RECT 127.390 213.190 127.675 213.520 ;
        RECT 123.585 212.215 126.175 212.985 ;
        RECT 126.345 212.215 126.635 212.940 ;
        RECT 127.390 212.935 127.560 213.190 ;
        RECT 126.895 212.765 127.560 212.935 ;
        RECT 127.845 212.890 128.015 213.690 ;
        RECT 128.185 213.675 129.395 214.765 ;
        RECT 126.895 212.385 127.065 212.765 ;
        RECT 127.245 212.215 127.575 212.595 ;
        RECT 127.755 212.385 128.015 212.890 ;
        RECT 128.185 212.965 128.705 213.505 ;
        RECT 128.875 213.135 129.395 213.675 ;
        RECT 129.565 213.690 129.835 214.595 ;
        RECT 130.005 214.005 130.335 214.765 ;
        RECT 130.515 213.835 130.685 214.595 ;
        RECT 128.185 212.215 129.395 212.965 ;
        RECT 129.565 212.890 129.735 213.690 ;
        RECT 130.020 213.665 130.685 213.835 ;
        RECT 130.945 213.675 132.615 214.765 ;
        RECT 130.020 213.520 130.190 213.665 ;
        RECT 129.905 213.190 130.190 213.520 ;
        RECT 130.020 212.935 130.190 213.190 ;
        RECT 130.425 213.115 130.755 213.485 ;
        RECT 130.945 212.985 131.695 213.505 ;
        RECT 131.865 213.155 132.615 213.675 ;
        RECT 132.785 213.690 133.055 214.595 ;
        RECT 133.225 214.005 133.555 214.765 ;
        RECT 133.735 213.835 133.905 214.595 ;
        RECT 129.565 212.385 129.825 212.890 ;
        RECT 130.020 212.765 130.685 212.935 ;
        RECT 130.005 212.215 130.335 212.595 ;
        RECT 130.515 212.385 130.685 212.765 ;
        RECT 130.945 212.215 132.615 212.985 ;
        RECT 132.785 212.890 132.955 213.690 ;
        RECT 133.240 213.665 133.905 213.835 ;
        RECT 134.165 213.690 134.435 214.595 ;
        RECT 134.605 214.005 134.935 214.765 ;
        RECT 135.115 213.835 135.285 214.595 ;
        RECT 133.240 213.520 133.410 213.665 ;
        RECT 133.125 213.190 133.410 213.520 ;
        RECT 133.240 212.935 133.410 213.190 ;
        RECT 133.645 213.115 133.975 213.485 ;
        RECT 132.785 212.385 133.045 212.890 ;
        RECT 133.240 212.765 133.905 212.935 ;
        RECT 133.225 212.215 133.555 212.595 ;
        RECT 133.735 212.385 133.905 212.765 ;
        RECT 134.165 212.890 134.335 213.690 ;
        RECT 134.620 213.665 135.285 213.835 ;
        RECT 135.545 213.675 136.755 214.765 ;
        RECT 134.620 213.520 134.790 213.665 ;
        RECT 134.505 213.190 134.790 213.520 ;
        RECT 134.620 212.935 134.790 213.190 ;
        RECT 135.025 213.115 135.355 213.485 ;
        RECT 135.545 212.965 136.065 213.505 ;
        RECT 136.235 213.135 136.755 213.675 ;
        RECT 136.925 213.690 137.195 214.595 ;
        RECT 137.365 214.005 137.695 214.765 ;
        RECT 137.875 213.835 138.055 214.595 ;
        RECT 134.165 212.385 134.425 212.890 ;
        RECT 134.620 212.765 135.285 212.935 ;
        RECT 134.605 212.215 134.935 212.595 ;
        RECT 135.115 212.385 135.285 212.765 ;
        RECT 135.545 212.215 136.755 212.965 ;
        RECT 136.925 212.890 137.105 213.690 ;
        RECT 137.380 213.665 138.055 213.835 ;
        RECT 137.380 213.520 137.550 213.665 ;
        RECT 139.225 213.600 139.515 214.765 ;
        RECT 139.685 213.625 139.955 214.595 ;
        RECT 140.165 213.965 140.445 214.765 ;
        RECT 140.625 214.215 141.820 214.545 ;
        RECT 140.950 213.795 141.370 214.045 ;
        RECT 140.125 213.625 141.370 213.795 ;
        RECT 137.275 213.190 137.550 213.520 ;
        RECT 137.380 212.935 137.550 213.190 ;
        RECT 137.775 213.115 138.115 213.485 ;
        RECT 136.925 212.385 137.185 212.890 ;
        RECT 137.380 212.765 138.045 212.935 ;
        RECT 137.365 212.215 137.695 212.595 ;
        RECT 137.875 212.385 138.045 212.765 ;
        RECT 139.225 212.215 139.515 212.940 ;
        RECT 139.685 212.890 139.855 213.625 ;
        RECT 140.125 213.455 140.295 213.625 ;
        RECT 141.595 213.455 141.765 214.015 ;
        RECT 142.015 213.625 142.270 214.765 ;
        RECT 142.445 213.690 142.715 214.595 ;
        RECT 142.885 214.005 143.215 214.765 ;
        RECT 143.395 213.835 143.575 214.595 ;
        RECT 140.065 213.125 140.295 213.455 ;
        RECT 141.025 213.125 141.765 213.455 ;
        RECT 141.935 213.205 142.270 213.455 ;
        RECT 140.125 212.955 140.295 213.125 ;
        RECT 141.515 213.035 141.765 213.125 ;
        RECT 139.685 212.545 139.955 212.890 ;
        RECT 140.125 212.785 140.865 212.955 ;
        RECT 141.515 212.865 142.250 213.035 ;
        RECT 140.145 212.215 140.525 212.615 ;
        RECT 140.695 212.435 140.865 212.785 ;
        RECT 141.035 212.215 141.770 212.695 ;
        RECT 141.940 212.395 142.250 212.865 ;
        RECT 142.445 212.890 142.625 213.690 ;
        RECT 142.900 213.665 143.575 213.835 ;
        RECT 144.285 213.690 144.555 214.595 ;
        RECT 144.725 214.005 145.055 214.765 ;
        RECT 145.235 213.835 145.415 214.595 ;
        RECT 142.900 213.520 143.070 213.665 ;
        RECT 142.795 213.190 143.070 213.520 ;
        RECT 142.900 212.935 143.070 213.190 ;
        RECT 143.295 213.115 143.635 213.485 ;
        RECT 142.445 212.385 142.705 212.890 ;
        RECT 142.900 212.765 143.565 212.935 ;
        RECT 142.885 212.215 143.215 212.595 ;
        RECT 143.395 212.385 143.565 212.765 ;
        RECT 144.285 212.890 144.465 213.690 ;
        RECT 144.740 213.665 145.415 213.835 ;
        RECT 145.665 213.675 147.335 214.765 ;
        RECT 144.740 213.520 144.910 213.665 ;
        RECT 144.635 213.190 144.910 213.520 ;
        RECT 144.740 212.935 144.910 213.190 ;
        RECT 145.135 213.115 145.475 213.485 ;
        RECT 145.665 212.985 146.415 213.505 ;
        RECT 146.585 213.155 147.335 213.675 ;
        RECT 147.505 213.690 147.775 214.595 ;
        RECT 147.945 214.005 148.275 214.765 ;
        RECT 148.455 213.835 148.635 214.595 ;
        RECT 144.285 212.385 144.545 212.890 ;
        RECT 144.740 212.765 145.405 212.935 ;
        RECT 144.725 212.215 145.055 212.595 ;
        RECT 145.235 212.385 145.405 212.765 ;
        RECT 145.665 212.215 147.335 212.985 ;
        RECT 147.505 212.890 147.685 213.690 ;
        RECT 147.960 213.665 148.635 213.835 ;
        RECT 148.885 213.675 150.095 214.765 ;
        RECT 147.960 213.520 148.130 213.665 ;
        RECT 147.855 213.190 148.130 213.520 ;
        RECT 147.960 212.935 148.130 213.190 ;
        RECT 148.355 213.115 148.695 213.485 ;
        RECT 148.885 213.135 149.405 213.675 ;
        RECT 149.575 212.965 150.095 213.505 ;
        RECT 147.505 212.385 147.765 212.890 ;
        RECT 147.960 212.765 148.625 212.935 ;
        RECT 147.945 212.215 148.275 212.595 ;
        RECT 148.455 212.385 148.625 212.765 ;
        RECT 148.885 212.215 150.095 212.965 ;
        RECT 36.100 212.045 150.180 212.215 ;
        RECT 36.185 211.295 37.395 212.045 ;
        RECT 37.655 211.495 37.825 211.785 ;
        RECT 37.995 211.665 38.325 212.045 ;
        RECT 37.655 211.325 38.320 211.495 ;
        RECT 36.185 210.755 36.705 211.295 ;
        RECT 36.875 210.585 37.395 211.125 ;
        RECT 36.185 209.495 37.395 210.585 ;
        RECT 37.570 210.505 37.920 211.155 ;
        RECT 38.090 210.335 38.320 211.325 ;
        RECT 37.655 210.165 38.320 210.335 ;
        RECT 37.655 209.665 37.825 210.165 ;
        RECT 37.995 209.495 38.325 209.995 ;
        RECT 38.495 209.665 38.680 211.785 ;
        RECT 38.935 211.585 39.185 212.045 ;
        RECT 39.355 211.595 39.690 211.765 ;
        RECT 39.885 211.595 40.560 211.765 ;
        RECT 39.355 211.455 39.525 211.595 ;
        RECT 38.850 210.465 39.130 211.415 ;
        RECT 39.300 211.325 39.525 211.455 ;
        RECT 39.300 210.220 39.470 211.325 ;
        RECT 39.695 211.175 40.220 211.395 ;
        RECT 39.640 210.410 39.880 211.005 ;
        RECT 40.050 210.475 40.220 211.175 ;
        RECT 40.390 210.815 40.560 211.595 ;
        RECT 40.880 211.545 41.250 212.045 ;
        RECT 41.430 211.595 41.835 211.765 ;
        RECT 42.005 211.595 42.790 211.765 ;
        RECT 41.430 211.365 41.600 211.595 ;
        RECT 40.770 211.065 41.600 211.365 ;
        RECT 41.985 211.095 42.450 211.425 ;
        RECT 40.770 211.035 40.970 211.065 ;
        RECT 41.090 210.815 41.260 210.885 ;
        RECT 40.390 210.645 41.260 210.815 ;
        RECT 40.750 210.555 41.260 210.645 ;
        RECT 39.300 210.090 39.605 210.220 ;
        RECT 40.050 210.110 40.580 210.475 ;
        RECT 38.920 209.495 39.185 209.955 ;
        RECT 39.355 209.665 39.605 210.090 ;
        RECT 40.750 209.940 40.920 210.555 ;
        RECT 39.815 209.770 40.920 209.940 ;
        RECT 41.090 209.495 41.260 210.295 ;
        RECT 41.430 209.995 41.600 211.065 ;
        RECT 41.770 210.165 41.960 210.885 ;
        RECT 42.130 210.135 42.450 211.095 ;
        RECT 42.620 211.135 42.790 211.595 ;
        RECT 43.065 211.515 43.275 212.045 ;
        RECT 43.535 211.305 43.865 211.830 ;
        RECT 44.035 211.435 44.205 212.045 ;
        RECT 44.375 211.390 44.705 211.825 ;
        RECT 44.375 211.305 44.755 211.390 ;
        RECT 43.665 211.135 43.865 211.305 ;
        RECT 44.530 211.265 44.755 211.305 ;
        RECT 42.620 210.805 43.495 211.135 ;
        RECT 43.665 210.805 44.415 211.135 ;
        RECT 41.430 209.665 41.680 209.995 ;
        RECT 42.620 209.965 42.790 210.805 ;
        RECT 43.665 210.600 43.855 210.805 ;
        RECT 44.585 210.685 44.755 211.265 ;
        RECT 44.985 211.225 45.195 212.045 ;
        RECT 45.365 211.245 45.695 211.875 ;
        RECT 44.540 210.635 44.755 210.685 ;
        RECT 45.365 210.645 45.615 211.245 ;
        RECT 45.865 211.225 46.095 212.045 ;
        RECT 46.395 211.495 46.565 211.785 ;
        RECT 46.735 211.665 47.065 212.045 ;
        RECT 46.395 211.325 47.060 211.495 ;
        RECT 45.785 210.805 46.115 211.055 ;
        RECT 42.960 210.225 43.855 210.600 ;
        RECT 44.365 210.555 44.755 210.635 ;
        RECT 41.905 209.795 42.790 209.965 ;
        RECT 42.970 209.495 43.285 209.995 ;
        RECT 43.515 209.665 43.855 210.225 ;
        RECT 44.025 209.495 44.195 210.505 ;
        RECT 44.365 209.710 44.695 210.555 ;
        RECT 44.985 209.495 45.195 210.635 ;
        RECT 45.365 209.665 45.695 210.645 ;
        RECT 45.865 209.495 46.095 210.635 ;
        RECT 46.310 210.505 46.660 211.155 ;
        RECT 46.830 210.335 47.060 211.325 ;
        RECT 46.395 210.165 47.060 210.335 ;
        RECT 46.395 209.665 46.565 210.165 ;
        RECT 46.735 209.495 47.065 209.995 ;
        RECT 47.235 209.665 47.420 211.785 ;
        RECT 47.675 211.585 47.925 212.045 ;
        RECT 48.095 211.595 48.430 211.765 ;
        RECT 48.625 211.595 49.300 211.765 ;
        RECT 48.095 211.455 48.265 211.595 ;
        RECT 47.590 210.465 47.870 211.415 ;
        RECT 48.040 211.325 48.265 211.455 ;
        RECT 48.040 210.220 48.210 211.325 ;
        RECT 48.435 211.175 48.960 211.395 ;
        RECT 48.380 210.410 48.620 211.005 ;
        RECT 48.790 210.475 48.960 211.175 ;
        RECT 49.130 210.815 49.300 211.595 ;
        RECT 49.620 211.545 49.990 212.045 ;
        RECT 50.170 211.595 50.575 211.765 ;
        RECT 50.745 211.595 51.530 211.765 ;
        RECT 50.170 211.365 50.340 211.595 ;
        RECT 49.510 211.065 50.340 211.365 ;
        RECT 50.725 211.095 51.190 211.425 ;
        RECT 49.510 211.035 49.710 211.065 ;
        RECT 49.830 210.815 50.000 210.885 ;
        RECT 49.130 210.645 50.000 210.815 ;
        RECT 49.490 210.555 50.000 210.645 ;
        RECT 48.040 210.090 48.345 210.220 ;
        RECT 48.790 210.110 49.320 210.475 ;
        RECT 47.660 209.495 47.925 209.955 ;
        RECT 48.095 209.665 48.345 210.090 ;
        RECT 49.490 209.940 49.660 210.555 ;
        RECT 48.555 209.770 49.660 209.940 ;
        RECT 49.830 209.495 50.000 210.295 ;
        RECT 50.170 209.995 50.340 211.065 ;
        RECT 50.510 210.165 50.700 210.885 ;
        RECT 50.870 210.135 51.190 211.095 ;
        RECT 51.360 211.135 51.530 211.595 ;
        RECT 51.805 211.515 52.015 212.045 ;
        RECT 52.275 211.305 52.605 211.830 ;
        RECT 52.775 211.435 52.945 212.045 ;
        RECT 53.115 211.390 53.445 211.825 ;
        RECT 54.675 211.495 54.845 211.785 ;
        RECT 55.015 211.665 55.345 212.045 ;
        RECT 53.115 211.305 53.495 211.390 ;
        RECT 54.675 211.325 55.340 211.495 ;
        RECT 52.405 211.135 52.605 211.305 ;
        RECT 53.270 211.265 53.495 211.305 ;
        RECT 51.360 210.805 52.235 211.135 ;
        RECT 52.405 210.805 53.155 211.135 ;
        RECT 50.170 209.665 50.420 209.995 ;
        RECT 51.360 209.965 51.530 210.805 ;
        RECT 52.405 210.600 52.595 210.805 ;
        RECT 53.325 210.685 53.495 211.265 ;
        RECT 53.280 210.635 53.495 210.685 ;
        RECT 51.700 210.225 52.595 210.600 ;
        RECT 53.105 210.555 53.495 210.635 ;
        RECT 50.645 209.795 51.530 209.965 ;
        RECT 51.710 209.495 52.025 209.995 ;
        RECT 52.255 209.665 52.595 210.225 ;
        RECT 52.765 209.495 52.935 210.505 ;
        RECT 53.105 209.710 53.435 210.555 ;
        RECT 54.590 210.505 54.940 211.155 ;
        RECT 55.110 210.335 55.340 211.325 ;
        RECT 54.675 210.165 55.340 210.335 ;
        RECT 54.675 209.665 54.845 210.165 ;
        RECT 55.015 209.495 55.345 209.995 ;
        RECT 55.515 209.665 55.700 211.785 ;
        RECT 55.955 211.585 56.205 212.045 ;
        RECT 56.375 211.595 56.710 211.765 ;
        RECT 56.905 211.595 57.580 211.765 ;
        RECT 56.375 211.455 56.545 211.595 ;
        RECT 55.870 210.465 56.150 211.415 ;
        RECT 56.320 211.325 56.545 211.455 ;
        RECT 56.320 210.220 56.490 211.325 ;
        RECT 56.715 211.175 57.240 211.395 ;
        RECT 56.660 210.410 56.900 211.005 ;
        RECT 57.070 210.475 57.240 211.175 ;
        RECT 57.410 210.815 57.580 211.595 ;
        RECT 57.900 211.545 58.270 212.045 ;
        RECT 58.450 211.595 58.855 211.765 ;
        RECT 59.025 211.595 59.810 211.765 ;
        RECT 58.450 211.365 58.620 211.595 ;
        RECT 57.790 211.065 58.620 211.365 ;
        RECT 59.005 211.095 59.470 211.425 ;
        RECT 57.790 211.035 57.990 211.065 ;
        RECT 58.110 210.815 58.280 210.885 ;
        RECT 57.410 210.645 58.280 210.815 ;
        RECT 57.770 210.555 58.280 210.645 ;
        RECT 56.320 210.090 56.625 210.220 ;
        RECT 57.070 210.110 57.600 210.475 ;
        RECT 55.940 209.495 56.205 209.955 ;
        RECT 56.375 209.665 56.625 210.090 ;
        RECT 57.770 209.940 57.940 210.555 ;
        RECT 56.835 209.770 57.940 209.940 ;
        RECT 58.110 209.495 58.280 210.295 ;
        RECT 58.450 209.995 58.620 211.065 ;
        RECT 58.790 210.165 58.980 210.885 ;
        RECT 59.150 210.135 59.470 211.095 ;
        RECT 59.640 211.135 59.810 211.595 ;
        RECT 60.085 211.515 60.295 212.045 ;
        RECT 60.555 211.305 60.885 211.830 ;
        RECT 61.055 211.435 61.225 212.045 ;
        RECT 61.395 211.390 61.725 211.825 ;
        RECT 61.395 211.305 61.775 211.390 ;
        RECT 61.945 211.320 62.235 212.045 ;
        RECT 63.325 211.545 63.585 211.875 ;
        RECT 63.795 211.565 64.070 212.045 ;
        RECT 60.685 211.135 60.885 211.305 ;
        RECT 61.550 211.265 61.775 211.305 ;
        RECT 59.640 210.805 60.515 211.135 ;
        RECT 60.685 210.805 61.435 211.135 ;
        RECT 58.450 209.665 58.700 209.995 ;
        RECT 59.640 209.965 59.810 210.805 ;
        RECT 60.685 210.600 60.875 210.805 ;
        RECT 61.605 210.685 61.775 211.265 ;
        RECT 61.560 210.635 61.775 210.685 ;
        RECT 59.980 210.225 60.875 210.600 ;
        RECT 61.385 210.555 61.775 210.635 ;
        RECT 58.925 209.795 59.810 209.965 ;
        RECT 59.990 209.495 60.305 209.995 ;
        RECT 60.535 209.665 60.875 210.225 ;
        RECT 61.045 209.495 61.215 210.505 ;
        RECT 61.385 209.710 61.715 210.555 ;
        RECT 61.945 209.495 62.235 210.660 ;
        RECT 63.325 210.635 63.495 211.545 ;
        RECT 64.280 211.475 64.485 211.875 ;
        RECT 64.655 211.645 64.990 212.045 ;
        RECT 63.665 210.805 64.025 211.385 ;
        RECT 64.280 211.305 64.965 211.475 ;
        RECT 64.205 210.635 64.455 211.135 ;
        RECT 63.325 210.465 64.455 210.635 ;
        RECT 63.325 209.695 63.595 210.465 ;
        RECT 64.625 210.275 64.965 211.305 ;
        RECT 63.765 209.495 64.095 210.275 ;
        RECT 64.300 210.100 64.965 210.275 ;
        RECT 65.165 211.370 65.425 211.875 ;
        RECT 65.605 211.665 65.935 212.045 ;
        RECT 66.115 211.495 66.285 211.875 ;
        RECT 65.165 210.570 65.335 211.370 ;
        RECT 65.620 211.325 66.285 211.495 ;
        RECT 65.620 211.070 65.790 211.325 ;
        RECT 66.565 211.235 66.805 212.045 ;
        RECT 66.975 211.235 67.305 211.875 ;
        RECT 67.475 211.235 67.745 212.045 ;
        RECT 67.925 211.370 68.185 211.875 ;
        RECT 68.365 211.665 68.695 212.045 ;
        RECT 68.875 211.495 69.045 211.875 ;
        RECT 65.505 210.740 65.790 211.070 ;
        RECT 66.025 210.775 66.355 211.145 ;
        RECT 66.545 210.805 66.895 211.055 ;
        RECT 65.620 210.595 65.790 210.740 ;
        RECT 67.065 210.635 67.235 211.235 ;
        RECT 67.405 210.805 67.755 211.055 ;
        RECT 64.300 209.695 64.485 210.100 ;
        RECT 64.655 209.495 64.990 209.920 ;
        RECT 65.165 209.665 65.435 210.570 ;
        RECT 65.620 210.425 66.285 210.595 ;
        RECT 65.605 209.495 65.935 210.255 ;
        RECT 66.115 209.665 66.285 210.425 ;
        RECT 66.555 210.465 67.235 210.635 ;
        RECT 66.555 209.680 66.885 210.465 ;
        RECT 67.415 209.495 67.745 210.635 ;
        RECT 67.925 210.570 68.095 211.370 ;
        RECT 68.380 211.325 69.045 211.495 ;
        RECT 68.380 211.070 68.550 211.325 ;
        RECT 70.225 211.305 70.690 211.850 ;
        RECT 68.265 210.740 68.550 211.070 ;
        RECT 68.785 210.775 69.115 211.145 ;
        RECT 68.380 210.595 68.550 210.740 ;
        RECT 67.925 209.665 68.195 210.570 ;
        RECT 68.380 210.425 69.045 210.595 ;
        RECT 68.365 209.495 68.695 210.255 ;
        RECT 68.875 209.665 69.045 210.425 ;
        RECT 70.225 210.345 70.395 211.305 ;
        RECT 71.195 211.225 71.365 212.045 ;
        RECT 71.535 211.395 71.865 211.875 ;
        RECT 72.035 211.655 72.385 212.045 ;
        RECT 72.555 211.475 72.785 211.875 ;
        RECT 72.275 211.395 72.785 211.475 ;
        RECT 71.535 211.305 72.785 211.395 ;
        RECT 72.955 211.305 73.275 211.785 ;
        RECT 71.535 211.225 72.445 211.305 ;
        RECT 70.565 210.685 70.810 211.135 ;
        RECT 71.070 210.855 71.765 211.055 ;
        RECT 71.935 210.885 72.535 211.055 ;
        RECT 71.935 210.685 72.105 210.885 ;
        RECT 72.765 210.715 72.935 211.135 ;
        RECT 70.565 210.515 72.105 210.685 ;
        RECT 72.275 210.545 72.935 210.715 ;
        RECT 72.275 210.345 72.445 210.545 ;
        RECT 73.105 210.375 73.275 211.305 ;
        RECT 70.225 210.175 72.445 210.345 ;
        RECT 72.615 210.175 73.275 210.375 ;
        RECT 73.445 211.305 73.910 211.850 ;
        RECT 73.445 210.345 73.615 211.305 ;
        RECT 74.415 211.225 74.585 212.045 ;
        RECT 74.755 211.395 75.085 211.875 ;
        RECT 75.255 211.655 75.605 212.045 ;
        RECT 75.775 211.475 76.005 211.875 ;
        RECT 75.495 211.395 76.005 211.475 ;
        RECT 74.755 211.305 76.005 211.395 ;
        RECT 76.175 211.305 76.495 211.785 ;
        RECT 74.755 211.225 75.665 211.305 ;
        RECT 73.785 210.685 74.030 211.135 ;
        RECT 74.290 210.855 74.985 211.055 ;
        RECT 75.155 210.885 75.755 211.055 ;
        RECT 75.155 210.685 75.325 210.885 ;
        RECT 75.985 210.715 76.155 211.135 ;
        RECT 73.785 210.515 75.325 210.685 ;
        RECT 75.495 210.545 76.155 210.715 ;
        RECT 75.495 210.345 75.665 210.545 ;
        RECT 76.325 210.375 76.495 211.305 ;
        RECT 76.665 211.275 79.255 212.045 ;
        RECT 80.085 211.415 80.415 211.775 ;
        RECT 81.035 211.585 81.285 212.045 ;
        RECT 81.455 211.585 82.015 211.875 ;
        RECT 76.665 210.755 77.875 211.275 ;
        RECT 80.085 211.225 81.475 211.415 ;
        RECT 81.305 211.135 81.475 211.225 ;
        RECT 78.045 210.585 79.255 211.105 ;
        RECT 73.445 210.175 75.665 210.345 ;
        RECT 75.835 210.175 76.495 210.375 ;
        RECT 70.225 209.495 70.525 210.005 ;
        RECT 70.695 209.665 71.025 210.175 ;
        RECT 72.615 210.005 72.785 210.175 ;
        RECT 71.195 209.495 71.825 210.005 ;
        RECT 72.405 209.835 72.785 210.005 ;
        RECT 72.955 209.495 73.255 210.005 ;
        RECT 73.445 209.495 73.745 210.005 ;
        RECT 73.915 209.665 74.245 210.175 ;
        RECT 75.835 210.005 76.005 210.175 ;
        RECT 74.415 209.495 75.045 210.005 ;
        RECT 75.625 209.835 76.005 210.005 ;
        RECT 76.175 209.495 76.475 210.005 ;
        RECT 76.665 209.495 79.255 210.585 ;
        RECT 79.900 210.805 80.575 211.055 ;
        RECT 80.795 210.805 81.135 211.055 ;
        RECT 81.305 210.805 81.595 211.135 ;
        RECT 79.900 210.445 80.165 210.805 ;
        RECT 81.305 210.555 81.475 210.805 ;
        RECT 80.535 210.385 81.475 210.555 ;
        RECT 80.085 209.495 80.365 210.165 ;
        RECT 80.535 209.835 80.835 210.385 ;
        RECT 81.765 210.215 82.015 211.585 ;
        RECT 82.190 211.540 82.525 212.045 ;
        RECT 82.695 211.475 82.935 211.850 ;
        RECT 83.215 211.715 83.385 211.860 ;
        RECT 83.215 211.520 83.590 211.715 ;
        RECT 83.950 211.550 84.345 212.045 ;
        RECT 82.245 210.515 82.545 211.365 ;
        RECT 82.715 211.325 82.935 211.475 ;
        RECT 82.715 210.995 83.250 211.325 ;
        RECT 83.420 211.185 83.590 211.520 ;
        RECT 84.515 211.355 84.755 211.875 ;
        RECT 82.715 210.345 82.950 210.995 ;
        RECT 83.420 210.825 84.405 211.185 ;
        RECT 81.035 209.495 81.365 210.215 ;
        RECT 81.555 209.665 82.015 210.215 ;
        RECT 82.275 210.115 82.950 210.345 ;
        RECT 83.120 210.805 84.405 210.825 ;
        RECT 83.120 210.655 83.980 210.805 ;
        RECT 82.275 209.685 82.445 210.115 ;
        RECT 82.615 209.495 82.945 209.945 ;
        RECT 83.120 209.710 83.405 210.655 ;
        RECT 84.580 210.550 84.755 211.355 ;
        RECT 84.965 211.315 85.255 212.045 ;
        RECT 84.955 210.805 85.255 211.135 ;
        RECT 85.435 211.115 85.665 211.755 ;
        RECT 85.845 211.495 86.155 211.865 ;
        RECT 86.335 211.675 87.005 212.045 ;
        RECT 85.845 211.295 87.075 211.495 ;
        RECT 85.435 210.805 85.960 211.115 ;
        RECT 86.140 210.805 86.605 211.115 ;
        RECT 86.785 210.625 87.075 211.295 ;
        RECT 83.580 210.175 84.275 210.485 ;
        RECT 83.585 209.495 84.270 209.965 ;
        RECT 84.450 209.765 84.755 210.550 ;
        RECT 84.965 210.385 86.125 210.625 ;
        RECT 84.965 209.675 85.225 210.385 ;
        RECT 85.395 209.495 85.725 210.205 ;
        RECT 85.895 209.675 86.125 210.385 ;
        RECT 86.305 210.405 87.075 210.625 ;
        RECT 86.305 209.675 86.575 210.405 ;
        RECT 86.755 209.495 87.095 210.225 ;
        RECT 87.265 209.675 87.525 211.865 ;
        RECT 87.705 211.320 87.995 212.045 ;
        RECT 88.165 211.535 88.505 212.045 ;
        RECT 88.175 210.805 88.515 211.365 ;
        RECT 88.685 211.135 88.935 211.865 ;
        RECT 89.260 211.505 89.445 211.865 ;
        RECT 89.625 211.675 89.955 212.045 ;
        RECT 90.135 211.505 90.360 211.865 ;
        RECT 89.260 211.315 90.740 211.505 ;
        RECT 88.685 210.805 89.325 211.135 ;
        RECT 89.505 210.805 89.835 211.135 ;
        RECT 87.705 209.495 87.995 210.660 ;
        RECT 88.330 210.405 89.435 210.605 ;
        RECT 88.330 209.675 88.580 210.405 ;
        RECT 88.750 209.495 89.080 210.225 ;
        RECT 89.250 209.675 89.435 210.405 ;
        RECT 89.605 209.675 89.835 210.805 ;
        RECT 90.015 210.515 90.315 211.135 ;
        RECT 90.525 210.345 90.740 211.315 ;
        RECT 90.925 211.275 93.515 212.045 ;
        RECT 93.775 211.495 93.945 211.875 ;
        RECT 94.125 211.665 94.455 212.045 ;
        RECT 93.775 211.325 94.440 211.495 ;
        RECT 94.635 211.370 94.895 211.875 ;
        RECT 90.925 210.755 92.135 211.275 ;
        RECT 92.305 210.585 93.515 211.105 ;
        RECT 93.705 210.775 94.035 211.145 ;
        RECT 94.270 211.070 94.440 211.325 ;
        RECT 94.270 210.740 94.555 211.070 ;
        RECT 94.270 210.595 94.440 210.740 ;
        RECT 90.015 209.675 90.740 210.345 ;
        RECT 90.925 209.495 93.515 210.585 ;
        RECT 93.775 210.425 94.440 210.595 ;
        RECT 94.725 210.570 94.895 211.370 ;
        RECT 95.155 211.495 95.325 211.785 ;
        RECT 95.495 211.665 95.825 212.045 ;
        RECT 95.155 211.325 95.820 211.495 ;
        RECT 93.775 209.665 93.945 210.425 ;
        RECT 94.125 209.495 94.455 210.255 ;
        RECT 94.625 209.665 94.895 210.570 ;
        RECT 95.070 210.505 95.420 211.155 ;
        RECT 95.590 210.335 95.820 211.325 ;
        RECT 95.155 210.165 95.820 210.335 ;
        RECT 95.155 209.665 95.325 210.165 ;
        RECT 95.495 209.495 95.825 209.995 ;
        RECT 95.995 209.665 96.180 211.785 ;
        RECT 96.435 211.585 96.685 212.045 ;
        RECT 96.855 211.595 97.190 211.765 ;
        RECT 97.385 211.595 98.060 211.765 ;
        RECT 96.855 211.455 97.025 211.595 ;
        RECT 96.350 210.465 96.630 211.415 ;
        RECT 96.800 211.325 97.025 211.455 ;
        RECT 96.800 210.220 96.970 211.325 ;
        RECT 97.195 211.175 97.720 211.395 ;
        RECT 97.140 210.410 97.380 211.005 ;
        RECT 97.550 210.475 97.720 211.175 ;
        RECT 97.890 210.815 98.060 211.595 ;
        RECT 98.380 211.545 98.750 212.045 ;
        RECT 98.930 211.595 99.335 211.765 ;
        RECT 99.505 211.595 100.290 211.765 ;
        RECT 98.930 211.365 99.100 211.595 ;
        RECT 98.270 211.065 99.100 211.365 ;
        RECT 99.485 211.095 99.950 211.425 ;
        RECT 98.270 211.035 98.470 211.065 ;
        RECT 98.590 210.815 98.760 210.885 ;
        RECT 97.890 210.645 98.760 210.815 ;
        RECT 98.250 210.555 98.760 210.645 ;
        RECT 96.800 210.090 97.105 210.220 ;
        RECT 97.550 210.110 98.080 210.475 ;
        RECT 96.420 209.495 96.685 209.955 ;
        RECT 96.855 209.665 97.105 210.090 ;
        RECT 98.250 209.940 98.420 210.555 ;
        RECT 97.315 209.770 98.420 209.940 ;
        RECT 98.590 209.495 98.760 210.295 ;
        RECT 98.930 209.995 99.100 211.065 ;
        RECT 99.270 210.165 99.460 210.885 ;
        RECT 99.630 210.135 99.950 211.095 ;
        RECT 100.120 211.135 100.290 211.595 ;
        RECT 100.565 211.515 100.775 212.045 ;
        RECT 101.035 211.305 101.365 211.830 ;
        RECT 101.535 211.435 101.705 212.045 ;
        RECT 101.875 211.390 102.205 211.825 ;
        RECT 102.515 211.495 102.685 211.785 ;
        RECT 102.855 211.665 103.185 212.045 ;
        RECT 101.875 211.305 102.255 211.390 ;
        RECT 102.515 211.325 103.180 211.495 ;
        RECT 101.165 211.135 101.365 211.305 ;
        RECT 102.030 211.265 102.255 211.305 ;
        RECT 100.120 210.805 100.995 211.135 ;
        RECT 101.165 210.805 101.915 211.135 ;
        RECT 98.930 209.665 99.180 209.995 ;
        RECT 100.120 209.965 100.290 210.805 ;
        RECT 101.165 210.600 101.355 210.805 ;
        RECT 102.085 210.685 102.255 211.265 ;
        RECT 102.040 210.635 102.255 210.685 ;
        RECT 100.460 210.225 101.355 210.600 ;
        RECT 101.865 210.555 102.255 210.635 ;
        RECT 99.405 209.795 100.290 209.965 ;
        RECT 100.470 209.495 100.785 209.995 ;
        RECT 101.015 209.665 101.355 210.225 ;
        RECT 101.525 209.495 101.695 210.505 ;
        RECT 101.865 209.710 102.195 210.555 ;
        RECT 102.430 210.505 102.780 211.155 ;
        RECT 102.950 210.335 103.180 211.325 ;
        RECT 102.515 210.165 103.180 210.335 ;
        RECT 102.515 209.665 102.685 210.165 ;
        RECT 102.855 209.495 103.185 209.995 ;
        RECT 103.355 209.665 103.540 211.785 ;
        RECT 103.795 211.585 104.045 212.045 ;
        RECT 104.215 211.595 104.550 211.765 ;
        RECT 104.745 211.595 105.420 211.765 ;
        RECT 104.215 211.455 104.385 211.595 ;
        RECT 103.710 210.465 103.990 211.415 ;
        RECT 104.160 211.325 104.385 211.455 ;
        RECT 104.160 210.220 104.330 211.325 ;
        RECT 104.555 211.175 105.080 211.395 ;
        RECT 104.500 210.410 104.740 211.005 ;
        RECT 104.910 210.475 105.080 211.175 ;
        RECT 105.250 210.815 105.420 211.595 ;
        RECT 105.740 211.545 106.110 212.045 ;
        RECT 106.290 211.595 106.695 211.765 ;
        RECT 106.865 211.595 107.650 211.765 ;
        RECT 106.290 211.365 106.460 211.595 ;
        RECT 105.630 211.065 106.460 211.365 ;
        RECT 106.845 211.095 107.310 211.425 ;
        RECT 105.630 211.035 105.830 211.065 ;
        RECT 105.950 210.815 106.120 210.885 ;
        RECT 105.250 210.645 106.120 210.815 ;
        RECT 105.610 210.555 106.120 210.645 ;
        RECT 104.160 210.090 104.465 210.220 ;
        RECT 104.910 210.110 105.440 210.475 ;
        RECT 103.780 209.495 104.045 209.955 ;
        RECT 104.215 209.665 104.465 210.090 ;
        RECT 105.610 209.940 105.780 210.555 ;
        RECT 104.675 209.770 105.780 209.940 ;
        RECT 105.950 209.495 106.120 210.295 ;
        RECT 106.290 209.995 106.460 211.065 ;
        RECT 106.630 210.165 106.820 210.885 ;
        RECT 106.990 210.135 107.310 211.095 ;
        RECT 107.480 211.135 107.650 211.595 ;
        RECT 107.925 211.515 108.135 212.045 ;
        RECT 108.395 211.305 108.725 211.830 ;
        RECT 108.895 211.435 109.065 212.045 ;
        RECT 109.235 211.390 109.565 211.825 ;
        RECT 109.235 211.305 109.615 211.390 ;
        RECT 108.525 211.135 108.725 211.305 ;
        RECT 109.390 211.265 109.615 211.305 ;
        RECT 107.480 210.805 108.355 211.135 ;
        RECT 108.525 210.805 109.275 211.135 ;
        RECT 106.290 209.665 106.540 209.995 ;
        RECT 107.480 209.965 107.650 210.805 ;
        RECT 108.525 210.600 108.715 210.805 ;
        RECT 109.445 210.685 109.615 211.265 ;
        RECT 109.400 210.635 109.615 210.685 ;
        RECT 107.820 210.225 108.715 210.600 ;
        RECT 109.225 210.555 109.615 210.635 ;
        RECT 110.705 211.100 111.045 211.875 ;
        RECT 111.215 211.585 111.385 212.045 ;
        RECT 111.625 211.610 111.985 211.875 ;
        RECT 111.625 211.605 111.980 211.610 ;
        RECT 111.625 211.595 111.975 211.605 ;
        RECT 111.625 211.590 111.970 211.595 ;
        RECT 111.625 211.580 111.965 211.590 ;
        RECT 112.615 211.585 112.785 212.045 ;
        RECT 111.625 211.575 111.960 211.580 ;
        RECT 111.625 211.565 111.950 211.575 ;
        RECT 111.625 211.555 111.940 211.565 ;
        RECT 111.625 211.415 111.925 211.555 ;
        RECT 111.215 211.225 111.925 211.415 ;
        RECT 112.115 211.415 112.445 211.495 ;
        RECT 112.955 211.415 113.295 211.875 ;
        RECT 112.115 211.225 113.295 211.415 ;
        RECT 113.465 211.320 113.755 212.045 ;
        RECT 113.930 211.305 114.185 211.875 ;
        RECT 114.355 211.645 114.685 212.045 ;
        RECT 115.110 211.510 115.640 211.875 ;
        RECT 115.110 211.475 115.285 211.510 ;
        RECT 114.355 211.305 115.285 211.475 ;
        RECT 106.765 209.795 107.650 209.965 ;
        RECT 107.830 209.495 108.145 209.995 ;
        RECT 108.375 209.665 108.715 210.225 ;
        RECT 108.885 209.495 109.055 210.505 ;
        RECT 109.225 209.710 109.555 210.555 ;
        RECT 110.705 209.665 110.985 211.100 ;
        RECT 111.215 210.655 111.500 211.225 ;
        RECT 111.685 210.825 112.155 211.055 ;
        RECT 112.325 211.035 112.655 211.055 ;
        RECT 112.325 210.855 112.775 211.035 ;
        RECT 112.965 210.855 113.295 211.055 ;
        RECT 111.215 210.440 112.365 210.655 ;
        RECT 111.155 209.495 111.865 210.270 ;
        RECT 112.035 209.665 112.365 210.440 ;
        RECT 112.560 209.740 112.775 210.855 ;
        RECT 113.065 210.515 113.295 210.855 ;
        RECT 112.955 209.495 113.285 210.215 ;
        RECT 113.465 209.495 113.755 210.660 ;
        RECT 113.930 210.635 114.100 211.305 ;
        RECT 114.355 211.135 114.525 211.305 ;
        RECT 114.270 210.805 114.525 211.135 ;
        RECT 114.750 210.805 114.945 211.135 ;
        RECT 113.930 209.665 114.265 210.635 ;
        RECT 114.435 209.495 114.605 210.635 ;
        RECT 114.775 209.835 114.945 210.805 ;
        RECT 115.115 210.175 115.285 211.305 ;
        RECT 115.455 210.515 115.625 211.315 ;
        RECT 115.830 211.025 116.105 211.875 ;
        RECT 115.825 210.855 116.105 211.025 ;
        RECT 115.830 210.715 116.105 210.855 ;
        RECT 116.275 210.515 116.465 211.875 ;
        RECT 116.645 211.510 117.155 212.045 ;
        RECT 117.375 211.235 117.620 211.840 ;
        RECT 116.665 211.065 117.895 211.235 ;
        RECT 115.455 210.345 116.465 210.515 ;
        RECT 116.635 210.500 117.385 210.690 ;
        RECT 115.115 210.005 116.240 210.175 ;
        RECT 116.635 209.835 116.805 210.500 ;
        RECT 117.555 210.255 117.895 211.065 ;
        RECT 114.775 209.665 116.805 209.835 ;
        RECT 116.975 209.495 117.145 210.255 ;
        RECT 117.380 209.845 117.895 210.255 ;
        RECT 118.065 211.100 118.405 211.875 ;
        RECT 118.575 211.585 118.745 212.045 ;
        RECT 118.985 211.610 119.345 211.875 ;
        RECT 118.985 211.605 119.340 211.610 ;
        RECT 118.985 211.595 119.335 211.605 ;
        RECT 118.985 211.590 119.330 211.595 ;
        RECT 118.985 211.580 119.325 211.590 ;
        RECT 119.975 211.585 120.145 212.045 ;
        RECT 118.985 211.575 119.320 211.580 ;
        RECT 118.985 211.565 119.310 211.575 ;
        RECT 118.985 211.555 119.300 211.565 ;
        RECT 118.985 211.415 119.285 211.555 ;
        RECT 118.575 211.225 119.285 211.415 ;
        RECT 119.475 211.415 119.805 211.495 ;
        RECT 120.315 211.415 120.655 211.875 ;
        RECT 119.475 211.225 120.655 211.415 ;
        RECT 118.065 209.665 118.345 211.100 ;
        RECT 118.575 210.655 118.860 211.225 ;
        RECT 120.825 211.100 121.165 211.875 ;
        RECT 121.335 211.585 121.505 212.045 ;
        RECT 121.745 211.610 122.105 211.875 ;
        RECT 121.745 211.605 122.100 211.610 ;
        RECT 121.745 211.595 122.095 211.605 ;
        RECT 121.745 211.590 122.090 211.595 ;
        RECT 121.745 211.580 122.085 211.590 ;
        RECT 122.735 211.585 122.905 212.045 ;
        RECT 121.745 211.575 122.080 211.580 ;
        RECT 121.745 211.565 122.070 211.575 ;
        RECT 121.745 211.555 122.060 211.565 ;
        RECT 121.745 211.415 122.045 211.555 ;
        RECT 121.335 211.225 122.045 211.415 ;
        RECT 122.235 211.415 122.565 211.495 ;
        RECT 123.075 211.415 123.415 211.875 ;
        RECT 122.235 211.225 123.415 211.415 ;
        RECT 123.590 211.305 123.845 211.875 ;
        RECT 124.015 211.645 124.345 212.045 ;
        RECT 124.770 211.510 125.300 211.875 ;
        RECT 125.490 211.705 125.765 211.875 ;
        RECT 125.485 211.535 125.765 211.705 ;
        RECT 124.770 211.475 124.945 211.510 ;
        RECT 124.015 211.305 124.945 211.475 ;
        RECT 119.045 210.825 119.515 211.055 ;
        RECT 119.685 211.035 120.015 211.055 ;
        RECT 119.685 210.855 120.135 211.035 ;
        RECT 120.325 210.855 120.655 211.055 ;
        RECT 118.575 210.440 119.725 210.655 ;
        RECT 118.515 209.495 119.225 210.270 ;
        RECT 119.395 209.665 119.725 210.440 ;
        RECT 119.920 209.740 120.135 210.855 ;
        RECT 120.425 210.515 120.655 210.855 ;
        RECT 120.315 209.495 120.645 210.215 ;
        RECT 120.825 209.665 121.105 211.100 ;
        RECT 121.335 210.655 121.620 211.225 ;
        RECT 121.805 210.825 122.275 211.055 ;
        RECT 122.445 211.035 122.775 211.055 ;
        RECT 122.445 210.855 122.895 211.035 ;
        RECT 123.085 210.855 123.415 211.055 ;
        RECT 121.335 210.440 122.485 210.655 ;
        RECT 121.275 209.495 121.985 210.270 ;
        RECT 122.155 209.665 122.485 210.440 ;
        RECT 122.680 209.740 122.895 210.855 ;
        RECT 123.185 210.515 123.415 210.855 ;
        RECT 123.590 210.635 123.760 211.305 ;
        RECT 124.015 211.135 124.185 211.305 ;
        RECT 123.930 210.805 124.185 211.135 ;
        RECT 124.410 210.805 124.605 211.135 ;
        RECT 123.075 209.495 123.405 210.215 ;
        RECT 123.590 209.665 123.925 210.635 ;
        RECT 124.095 209.495 124.265 210.635 ;
        RECT 124.435 209.835 124.605 210.805 ;
        RECT 124.775 210.175 124.945 211.305 ;
        RECT 125.115 210.515 125.285 211.315 ;
        RECT 125.490 210.715 125.765 211.535 ;
        RECT 125.935 210.515 126.125 211.875 ;
        RECT 126.305 211.510 126.815 212.045 ;
        RECT 127.035 211.235 127.280 211.840 ;
        RECT 128.000 211.235 128.245 211.840 ;
        RECT 128.465 211.510 128.975 212.045 ;
        RECT 126.325 211.065 127.555 211.235 ;
        RECT 125.115 210.345 126.125 210.515 ;
        RECT 126.295 210.500 127.045 210.690 ;
        RECT 124.775 210.005 125.900 210.175 ;
        RECT 126.295 209.835 126.465 210.500 ;
        RECT 127.215 210.255 127.555 211.065 ;
        RECT 124.435 209.665 126.465 209.835 ;
        RECT 126.635 209.495 126.805 210.255 ;
        RECT 127.040 209.845 127.555 210.255 ;
        RECT 127.725 211.065 128.955 211.235 ;
        RECT 127.725 210.255 128.065 211.065 ;
        RECT 128.235 210.500 128.985 210.690 ;
        RECT 127.725 209.845 128.240 210.255 ;
        RECT 128.475 209.495 128.645 210.255 ;
        RECT 128.815 209.835 128.985 210.500 ;
        RECT 129.155 210.515 129.345 211.875 ;
        RECT 129.515 211.025 129.790 211.875 ;
        RECT 129.980 211.510 130.510 211.875 ;
        RECT 130.935 211.645 131.265 212.045 ;
        RECT 130.335 211.475 130.510 211.510 ;
        RECT 129.515 210.855 129.795 211.025 ;
        RECT 129.515 210.715 129.790 210.855 ;
        RECT 129.995 210.515 130.165 211.315 ;
        RECT 129.155 210.345 130.165 210.515 ;
        RECT 130.335 211.305 131.265 211.475 ;
        RECT 131.435 211.305 131.690 211.875 ;
        RECT 131.955 211.495 132.125 211.785 ;
        RECT 132.295 211.665 132.625 212.045 ;
        RECT 131.955 211.325 132.620 211.495 ;
        RECT 130.335 210.175 130.505 211.305 ;
        RECT 131.095 211.135 131.265 211.305 ;
        RECT 129.380 210.005 130.505 210.175 ;
        RECT 130.675 210.805 130.870 211.135 ;
        RECT 131.095 210.805 131.350 211.135 ;
        RECT 130.675 209.835 130.845 210.805 ;
        RECT 131.520 210.635 131.690 211.305 ;
        RECT 128.815 209.665 130.845 209.835 ;
        RECT 131.015 209.495 131.185 210.635 ;
        RECT 131.355 209.665 131.690 210.635 ;
        RECT 131.870 210.505 132.220 211.155 ;
        RECT 132.390 210.335 132.620 211.325 ;
        RECT 131.955 210.165 132.620 210.335 ;
        RECT 131.955 209.665 132.125 210.165 ;
        RECT 132.295 209.495 132.625 209.995 ;
        RECT 132.795 209.665 132.980 211.785 ;
        RECT 133.235 211.585 133.485 212.045 ;
        RECT 133.655 211.595 133.990 211.765 ;
        RECT 134.185 211.595 134.860 211.765 ;
        RECT 133.655 211.455 133.825 211.595 ;
        RECT 133.150 210.465 133.430 211.415 ;
        RECT 133.600 211.325 133.825 211.455 ;
        RECT 133.600 210.220 133.770 211.325 ;
        RECT 133.995 211.175 134.520 211.395 ;
        RECT 133.940 210.410 134.180 211.005 ;
        RECT 134.350 210.475 134.520 211.175 ;
        RECT 134.690 210.815 134.860 211.595 ;
        RECT 135.180 211.545 135.550 212.045 ;
        RECT 135.730 211.595 136.135 211.765 ;
        RECT 136.305 211.595 137.090 211.765 ;
        RECT 135.730 211.365 135.900 211.595 ;
        RECT 135.070 211.065 135.900 211.365 ;
        RECT 136.285 211.095 136.750 211.425 ;
        RECT 135.070 211.035 135.270 211.065 ;
        RECT 135.390 210.815 135.560 210.885 ;
        RECT 134.690 210.645 135.560 210.815 ;
        RECT 135.050 210.555 135.560 210.645 ;
        RECT 133.600 210.090 133.905 210.220 ;
        RECT 134.350 210.110 134.880 210.475 ;
        RECT 133.220 209.495 133.485 209.955 ;
        RECT 133.655 209.665 133.905 210.090 ;
        RECT 135.050 209.940 135.220 210.555 ;
        RECT 134.115 209.770 135.220 209.940 ;
        RECT 135.390 209.495 135.560 210.295 ;
        RECT 135.730 209.995 135.900 211.065 ;
        RECT 136.070 210.165 136.260 210.885 ;
        RECT 136.430 210.135 136.750 211.095 ;
        RECT 136.920 211.135 137.090 211.595 ;
        RECT 137.365 211.515 137.575 212.045 ;
        RECT 137.835 211.305 138.165 211.830 ;
        RECT 138.335 211.435 138.505 212.045 ;
        RECT 138.675 211.390 139.005 211.825 ;
        RECT 138.675 211.305 139.055 211.390 ;
        RECT 139.225 211.320 139.515 212.045 ;
        RECT 140.235 211.495 140.405 211.875 ;
        RECT 140.585 211.665 140.915 212.045 ;
        RECT 140.235 211.325 140.900 211.495 ;
        RECT 141.095 211.370 141.355 211.875 ;
        RECT 137.965 211.135 138.165 211.305 ;
        RECT 138.830 211.265 139.055 211.305 ;
        RECT 136.920 210.805 137.795 211.135 ;
        RECT 137.965 210.805 138.715 211.135 ;
        RECT 135.730 209.665 135.980 209.995 ;
        RECT 136.920 209.965 137.090 210.805 ;
        RECT 137.965 210.600 138.155 210.805 ;
        RECT 138.885 210.685 139.055 211.265 ;
        RECT 140.165 210.775 140.495 211.145 ;
        RECT 140.730 211.070 140.900 211.325 ;
        RECT 138.840 210.635 139.055 210.685 ;
        RECT 140.730 210.740 141.015 211.070 ;
        RECT 137.260 210.225 138.155 210.600 ;
        RECT 138.665 210.555 139.055 210.635 ;
        RECT 136.205 209.795 137.090 209.965 ;
        RECT 137.270 209.495 137.585 209.995 ;
        RECT 137.815 209.665 138.155 210.225 ;
        RECT 138.325 209.495 138.495 210.505 ;
        RECT 138.665 209.710 138.995 210.555 ;
        RECT 139.225 209.495 139.515 210.660 ;
        RECT 140.730 210.595 140.900 210.740 ;
        RECT 140.235 210.425 140.900 210.595 ;
        RECT 141.185 210.570 141.355 211.370 ;
        RECT 141.615 211.495 141.785 211.785 ;
        RECT 141.955 211.665 142.285 212.045 ;
        RECT 141.615 211.325 142.280 211.495 ;
        RECT 140.235 209.665 140.405 210.425 ;
        RECT 140.585 209.495 140.915 210.255 ;
        RECT 141.085 209.665 141.355 210.570 ;
        RECT 141.530 210.505 141.880 211.155 ;
        RECT 142.050 210.335 142.280 211.325 ;
        RECT 141.615 210.165 142.280 210.335 ;
        RECT 141.615 209.665 141.785 210.165 ;
        RECT 141.955 209.495 142.285 209.995 ;
        RECT 142.455 209.665 142.640 211.785 ;
        RECT 142.895 211.585 143.145 212.045 ;
        RECT 143.315 211.595 143.650 211.765 ;
        RECT 143.845 211.595 144.520 211.765 ;
        RECT 143.315 211.455 143.485 211.595 ;
        RECT 142.810 210.465 143.090 211.415 ;
        RECT 143.260 211.325 143.485 211.455 ;
        RECT 143.260 210.220 143.430 211.325 ;
        RECT 143.655 211.175 144.180 211.395 ;
        RECT 143.600 210.410 143.840 211.005 ;
        RECT 144.010 210.475 144.180 211.175 ;
        RECT 144.350 210.815 144.520 211.595 ;
        RECT 144.840 211.545 145.210 212.045 ;
        RECT 145.390 211.595 145.795 211.765 ;
        RECT 145.965 211.595 146.750 211.765 ;
        RECT 145.390 211.365 145.560 211.595 ;
        RECT 144.730 211.065 145.560 211.365 ;
        RECT 145.945 211.095 146.410 211.425 ;
        RECT 144.730 211.035 144.930 211.065 ;
        RECT 145.050 210.815 145.220 210.885 ;
        RECT 144.350 210.645 145.220 210.815 ;
        RECT 144.710 210.555 145.220 210.645 ;
        RECT 143.260 210.090 143.565 210.220 ;
        RECT 144.010 210.110 144.540 210.475 ;
        RECT 142.880 209.495 143.145 209.955 ;
        RECT 143.315 209.665 143.565 210.090 ;
        RECT 144.710 209.940 144.880 210.555 ;
        RECT 143.775 209.770 144.880 209.940 ;
        RECT 145.050 209.495 145.220 210.295 ;
        RECT 145.390 209.995 145.560 211.065 ;
        RECT 145.730 210.165 145.920 210.885 ;
        RECT 146.090 210.135 146.410 211.095 ;
        RECT 146.580 211.135 146.750 211.595 ;
        RECT 147.025 211.515 147.235 212.045 ;
        RECT 147.495 211.305 147.825 211.830 ;
        RECT 147.995 211.435 148.165 212.045 ;
        RECT 148.335 211.390 148.665 211.825 ;
        RECT 148.335 211.305 148.715 211.390 ;
        RECT 147.625 211.135 147.825 211.305 ;
        RECT 148.490 211.265 148.715 211.305 ;
        RECT 148.885 211.295 150.095 212.045 ;
        RECT 146.580 210.805 147.455 211.135 ;
        RECT 147.625 210.805 148.375 211.135 ;
        RECT 145.390 209.665 145.640 209.995 ;
        RECT 146.580 209.965 146.750 210.805 ;
        RECT 147.625 210.600 147.815 210.805 ;
        RECT 148.545 210.685 148.715 211.265 ;
        RECT 148.500 210.635 148.715 210.685 ;
        RECT 146.920 210.225 147.815 210.600 ;
        RECT 148.325 210.555 148.715 210.635 ;
        RECT 148.885 210.585 149.405 211.125 ;
        RECT 149.575 210.755 150.095 211.295 ;
        RECT 145.865 209.795 146.750 209.965 ;
        RECT 146.930 209.495 147.245 209.995 ;
        RECT 147.475 209.665 147.815 210.225 ;
        RECT 147.985 209.495 148.155 210.505 ;
        RECT 148.325 209.710 148.655 210.555 ;
        RECT 148.885 209.495 150.095 210.585 ;
        RECT 36.100 209.325 150.180 209.495 ;
        RECT 36.185 208.235 37.395 209.325 ;
        RECT 37.565 208.235 41.075 209.325 ;
        RECT 41.245 208.235 42.455 209.325 ;
        RECT 36.185 207.525 36.705 208.065 ;
        RECT 36.875 207.695 37.395 208.235 ;
        RECT 37.565 207.545 39.215 208.065 ;
        RECT 39.385 207.715 41.075 208.235 ;
        RECT 36.185 206.775 37.395 207.525 ;
        RECT 37.565 206.775 41.075 207.545 ;
        RECT 41.245 207.525 41.765 208.065 ;
        RECT 41.935 207.695 42.455 208.235 ;
        RECT 42.635 208.375 42.910 209.145 ;
        RECT 43.080 208.715 43.410 209.145 ;
        RECT 43.580 208.885 43.775 209.325 ;
        RECT 43.955 208.715 44.285 209.145 ;
        RECT 43.080 208.545 44.285 208.715 ;
        RECT 42.635 208.185 43.220 208.375 ;
        RECT 43.390 208.215 44.285 208.545 ;
        RECT 45.015 208.395 45.185 209.155 ;
        RECT 45.365 208.565 45.695 209.325 ;
        RECT 45.015 208.225 45.680 208.395 ;
        RECT 45.865 208.250 46.135 209.155 ;
        RECT 41.245 206.775 42.455 207.525 ;
        RECT 42.635 207.365 42.875 208.015 ;
        RECT 43.045 207.515 43.220 208.185 ;
        RECT 45.510 208.080 45.680 208.225 ;
        RECT 43.390 207.685 43.805 208.015 ;
        RECT 43.985 207.685 44.280 208.015 ;
        RECT 43.045 207.335 43.375 207.515 ;
        RECT 42.650 206.775 42.980 207.165 ;
        RECT 43.150 206.955 43.375 207.335 ;
        RECT 43.575 207.065 43.805 207.685 ;
        RECT 44.945 207.675 45.275 208.045 ;
        RECT 45.510 207.750 45.795 208.080 ;
        RECT 43.985 206.775 44.285 207.505 ;
        RECT 45.510 207.495 45.680 207.750 ;
        RECT 45.015 207.325 45.680 207.495 ;
        RECT 45.965 207.450 46.135 208.250 ;
        RECT 46.855 208.395 47.025 209.155 ;
        RECT 47.205 208.565 47.535 209.325 ;
        RECT 46.855 208.225 47.520 208.395 ;
        RECT 47.705 208.250 47.975 209.155 ;
        RECT 47.350 208.080 47.520 208.225 ;
        RECT 46.785 207.675 47.115 208.045 ;
        RECT 47.350 207.750 47.635 208.080 ;
        RECT 47.350 207.495 47.520 207.750 ;
        RECT 45.015 206.945 45.185 207.325 ;
        RECT 45.365 206.775 45.695 207.155 ;
        RECT 45.875 206.945 46.135 207.450 ;
        RECT 46.855 207.325 47.520 207.495 ;
        RECT 47.805 207.450 47.975 208.250 ;
        RECT 49.065 208.160 49.355 209.325 ;
        RECT 49.525 208.890 54.870 209.325 ;
        RECT 46.855 206.945 47.025 207.325 ;
        RECT 47.205 206.775 47.535 207.155 ;
        RECT 47.715 206.945 47.975 207.450 ;
        RECT 49.065 206.775 49.355 207.500 ;
        RECT 51.110 207.320 51.450 208.150 ;
        RECT 52.930 207.640 53.280 208.890 ;
        RECT 55.045 208.235 57.635 209.325 ;
        RECT 57.865 208.265 58.195 209.110 ;
        RECT 58.365 208.315 58.535 209.325 ;
        RECT 58.705 208.595 59.045 209.155 ;
        RECT 59.275 208.825 59.590 209.325 ;
        RECT 59.770 208.855 60.655 209.025 ;
        RECT 55.045 207.545 56.255 208.065 ;
        RECT 56.425 207.715 57.635 208.235 ;
        RECT 57.805 208.185 58.195 208.265 ;
        RECT 58.705 208.220 59.600 208.595 ;
        RECT 57.805 208.135 58.020 208.185 ;
        RECT 57.805 207.555 57.975 208.135 ;
        RECT 58.705 208.015 58.895 208.220 ;
        RECT 59.770 208.015 59.940 208.855 ;
        RECT 60.880 208.825 61.130 209.155 ;
        RECT 58.145 207.685 58.895 208.015 ;
        RECT 59.065 207.685 59.940 208.015 ;
        RECT 49.525 206.775 54.870 207.320 ;
        RECT 55.045 206.775 57.635 207.545 ;
        RECT 57.805 207.515 58.030 207.555 ;
        RECT 58.695 207.515 58.895 207.685 ;
        RECT 57.805 207.430 58.185 207.515 ;
        RECT 57.855 206.995 58.185 207.430 ;
        RECT 58.355 206.775 58.525 207.385 ;
        RECT 58.695 206.990 59.025 207.515 ;
        RECT 59.285 206.775 59.495 207.305 ;
        RECT 59.770 207.225 59.940 207.685 ;
        RECT 60.110 207.725 60.430 208.685 ;
        RECT 60.600 207.935 60.790 208.655 ;
        RECT 60.960 207.755 61.130 208.825 ;
        RECT 61.300 208.525 61.470 209.325 ;
        RECT 61.640 208.880 62.745 209.050 ;
        RECT 61.640 208.265 61.810 208.880 ;
        RECT 62.955 208.730 63.205 209.155 ;
        RECT 63.375 208.865 63.640 209.325 ;
        RECT 61.980 208.345 62.510 208.710 ;
        RECT 62.955 208.600 63.260 208.730 ;
        RECT 61.300 208.175 61.810 208.265 ;
        RECT 61.300 208.005 62.170 208.175 ;
        RECT 61.300 207.935 61.470 208.005 ;
        RECT 61.590 207.755 61.790 207.785 ;
        RECT 60.110 207.395 60.575 207.725 ;
        RECT 60.960 207.455 61.790 207.755 ;
        RECT 60.960 207.225 61.130 207.455 ;
        RECT 59.770 207.055 60.555 207.225 ;
        RECT 60.725 207.055 61.130 207.225 ;
        RECT 61.310 206.775 61.680 207.275 ;
        RECT 62.000 207.225 62.170 208.005 ;
        RECT 62.340 207.645 62.510 208.345 ;
        RECT 62.680 207.815 62.920 208.410 ;
        RECT 62.340 207.425 62.865 207.645 ;
        RECT 63.090 207.495 63.260 208.600 ;
        RECT 63.035 207.365 63.260 207.495 ;
        RECT 63.430 207.405 63.710 208.355 ;
        RECT 63.035 207.225 63.205 207.365 ;
        RECT 62.000 207.055 62.675 207.225 ;
        RECT 62.870 207.055 63.205 207.225 ;
        RECT 63.375 206.775 63.625 207.235 ;
        RECT 63.880 207.035 64.065 209.155 ;
        RECT 64.235 208.825 64.565 209.325 ;
        RECT 64.735 208.655 64.905 209.155 ;
        RECT 65.170 208.900 65.505 209.325 ;
        RECT 65.675 208.720 65.860 209.125 ;
        RECT 64.240 208.485 64.905 208.655 ;
        RECT 65.195 208.545 65.860 208.720 ;
        RECT 66.065 208.545 66.395 209.325 ;
        RECT 64.240 207.495 64.470 208.485 ;
        RECT 64.640 207.665 64.990 208.315 ;
        RECT 65.195 207.515 65.535 208.545 ;
        RECT 66.565 208.355 66.835 209.125 ;
        RECT 67.005 208.890 72.350 209.325 ;
        RECT 65.705 208.185 66.835 208.355 ;
        RECT 65.705 207.685 65.955 208.185 ;
        RECT 64.240 207.325 64.905 207.495 ;
        RECT 65.195 207.345 65.880 207.515 ;
        RECT 66.135 207.435 66.495 208.015 ;
        RECT 64.235 206.775 64.565 207.155 ;
        RECT 64.735 207.035 64.905 207.325 ;
        RECT 65.170 206.775 65.505 207.175 ;
        RECT 65.675 206.945 65.880 207.345 ;
        RECT 66.665 207.275 66.835 208.185 ;
        RECT 68.590 207.320 68.930 208.150 ;
        RECT 70.410 207.640 70.760 208.890 ;
        RECT 72.535 208.355 72.865 209.140 ;
        RECT 72.535 208.185 73.215 208.355 ;
        RECT 73.395 208.185 73.725 209.325 ;
        RECT 72.525 207.765 72.875 208.015 ;
        RECT 73.045 207.585 73.215 208.185 ;
        RECT 74.825 208.160 75.115 209.325 ;
        RECT 75.295 208.605 75.625 209.325 ;
        RECT 73.385 207.765 73.735 208.015 ;
        RECT 75.285 207.965 75.515 208.305 ;
        RECT 75.805 207.965 76.020 209.080 ;
        RECT 76.215 208.380 76.545 209.155 ;
        RECT 76.715 208.550 77.425 209.325 ;
        RECT 76.215 208.165 77.365 208.380 ;
        RECT 75.285 207.765 75.615 207.965 ;
        RECT 75.805 207.785 76.255 207.965 ;
        RECT 75.925 207.765 76.255 207.785 ;
        RECT 76.425 207.765 76.895 207.995 ;
        RECT 77.080 207.595 77.365 208.165 ;
        RECT 77.595 207.720 77.875 209.155 ;
        RECT 78.085 208.185 78.315 209.325 ;
        RECT 78.485 208.175 78.815 209.155 ;
        RECT 78.985 208.185 79.195 209.325 ;
        RECT 80.530 208.355 80.920 208.530 ;
        RECT 81.405 208.525 81.735 209.325 ;
        RECT 81.905 208.535 82.440 209.155 ;
        RECT 83.565 208.815 83.865 209.325 ;
        RECT 84.035 208.645 84.365 209.155 ;
        RECT 84.535 208.815 85.165 209.325 ;
        RECT 85.745 208.815 86.125 208.985 ;
        RECT 86.295 208.815 86.595 209.325 ;
        RECT 85.955 208.645 86.125 208.815 ;
        RECT 80.530 208.185 81.955 208.355 ;
        RECT 78.065 207.765 78.395 208.015 ;
        RECT 66.090 206.775 66.365 207.255 ;
        RECT 66.575 206.945 66.835 207.275 ;
        RECT 67.005 206.775 72.350 207.320 ;
        RECT 72.545 206.775 72.785 207.585 ;
        RECT 72.955 206.945 73.285 207.585 ;
        RECT 73.455 206.775 73.725 207.585 ;
        RECT 74.825 206.775 75.115 207.500 ;
        RECT 75.285 207.405 76.465 207.595 ;
        RECT 75.285 206.945 75.625 207.405 ;
        RECT 76.135 207.325 76.465 207.405 ;
        RECT 76.655 207.405 77.365 207.595 ;
        RECT 76.655 207.265 76.955 207.405 ;
        RECT 76.640 207.255 76.955 207.265 ;
        RECT 76.630 207.245 76.955 207.255 ;
        RECT 76.620 207.240 76.955 207.245 ;
        RECT 75.795 206.775 75.965 207.235 ;
        RECT 76.615 207.230 76.955 207.240 ;
        RECT 76.610 207.225 76.955 207.230 ;
        RECT 76.605 207.215 76.955 207.225 ;
        RECT 76.600 207.210 76.955 207.215 ;
        RECT 76.595 206.945 76.955 207.210 ;
        RECT 77.195 206.775 77.365 207.235 ;
        RECT 77.535 206.945 77.875 207.720 ;
        RECT 78.085 206.775 78.315 207.595 ;
        RECT 78.565 207.575 78.815 208.175 ;
        RECT 78.485 206.945 78.815 207.575 ;
        RECT 78.985 206.775 79.195 207.595 ;
        RECT 80.405 207.455 80.760 208.015 ;
        RECT 80.930 207.285 81.100 208.185 ;
        RECT 81.270 207.455 81.535 208.015 ;
        RECT 81.785 207.685 81.955 208.185 ;
        RECT 82.125 207.515 82.440 208.535 ;
        RECT 80.510 206.775 80.750 207.285 ;
        RECT 80.930 206.955 81.210 207.285 ;
        RECT 81.440 206.775 81.655 207.285 ;
        RECT 81.825 206.945 82.440 207.515 ;
        RECT 83.565 208.475 85.785 208.645 ;
        RECT 83.565 207.515 83.735 208.475 ;
        RECT 83.905 208.135 85.445 208.305 ;
        RECT 83.905 207.685 84.150 208.135 ;
        RECT 84.410 207.765 85.105 207.965 ;
        RECT 85.275 207.935 85.445 208.135 ;
        RECT 85.615 208.275 85.785 208.475 ;
        RECT 85.955 208.445 86.615 208.645 ;
        RECT 85.615 208.105 86.275 208.275 ;
        RECT 85.275 207.765 85.875 207.935 ;
        RECT 86.105 207.685 86.275 208.105 ;
        RECT 83.565 206.970 84.030 207.515 ;
        RECT 84.535 206.775 84.705 207.595 ;
        RECT 84.875 207.515 85.785 207.595 ;
        RECT 86.445 207.515 86.615 208.445 ;
        RECT 86.850 208.355 87.120 209.150 ;
        RECT 87.300 208.525 87.515 209.325 ;
        RECT 87.695 208.355 87.980 209.150 ;
        RECT 86.850 208.185 87.980 208.355 ;
        RECT 86.830 207.715 87.330 207.980 ;
        RECT 87.550 207.685 87.935 208.015 ;
        RECT 88.160 207.685 88.440 209.155 ;
        RECT 88.620 207.740 88.950 209.155 ;
        RECT 89.120 207.980 89.325 209.155 ;
        RECT 89.495 208.335 89.705 209.150 ;
        RECT 89.945 208.505 90.275 209.325 ;
        RECT 89.495 208.155 90.145 208.335 ;
        RECT 90.450 208.310 90.705 209.150 ;
        RECT 89.120 207.740 89.550 207.980 ;
        RECT 87.550 207.535 87.855 207.685 ;
        RECT 84.875 207.425 86.125 207.515 ;
        RECT 84.875 206.945 85.205 207.425 ;
        RECT 85.615 207.345 86.125 207.425 ;
        RECT 85.375 206.775 85.725 207.165 ;
        RECT 85.895 206.945 86.125 207.345 ;
        RECT 86.295 207.035 86.615 207.515 ;
        RECT 86.885 206.775 87.125 207.450 ;
        RECT 87.300 206.975 87.855 207.535 ;
        RECT 89.925 207.515 90.145 208.155 ;
        RECT 88.035 207.345 90.145 207.515 ;
        RECT 88.035 206.950 88.240 207.345 ;
        RECT 88.925 207.340 90.145 207.345 ;
        RECT 88.410 206.775 88.755 207.175 ;
        RECT 88.925 206.950 89.255 207.340 ;
        RECT 89.530 206.775 90.205 207.160 ;
        RECT 90.375 206.945 90.705 208.310 ;
        RECT 90.935 208.355 91.265 209.140 ;
        RECT 90.935 208.185 91.615 208.355 ;
        RECT 91.795 208.185 92.125 209.325 ;
        RECT 92.305 208.890 97.650 209.325 ;
        RECT 90.925 207.765 91.275 208.015 ;
        RECT 91.445 207.585 91.615 208.185 ;
        RECT 91.785 207.765 92.135 208.015 ;
        RECT 90.945 206.775 91.185 207.585 ;
        RECT 91.355 206.945 91.685 207.585 ;
        RECT 91.855 206.775 92.125 207.585 ;
        RECT 93.890 207.320 94.230 208.150 ;
        RECT 95.710 207.640 96.060 208.890 ;
        RECT 98.755 208.355 99.085 209.140 ;
        RECT 98.755 208.185 99.435 208.355 ;
        RECT 99.615 208.185 99.945 209.325 ;
        RECT 98.745 207.765 99.095 208.015 ;
        RECT 99.265 207.585 99.435 208.185 ;
        RECT 100.585 208.160 100.875 209.325 ;
        RECT 101.545 208.985 102.685 209.155 ;
        RECT 101.545 208.525 101.845 208.985 ;
        RECT 102.015 208.355 102.345 208.815 ;
        RECT 101.585 208.135 102.345 208.355 ;
        RECT 102.515 208.355 102.685 208.985 ;
        RECT 102.855 208.525 103.185 209.325 ;
        RECT 103.355 208.355 103.630 209.155 ;
        RECT 102.515 208.145 103.630 208.355 ;
        RECT 103.805 208.235 105.475 209.325 ;
        RECT 99.605 207.765 99.955 208.015 ;
        RECT 101.585 207.595 101.800 208.135 ;
        RECT 101.970 207.765 102.740 207.965 ;
        RECT 102.910 207.765 103.630 207.965 ;
        RECT 92.305 206.775 97.650 207.320 ;
        RECT 98.765 206.775 99.005 207.585 ;
        RECT 99.175 206.945 99.505 207.585 ;
        RECT 99.675 206.775 99.945 207.585 ;
        RECT 100.585 206.775 100.875 207.500 ;
        RECT 101.585 207.425 103.185 207.595 ;
        RECT 102.015 207.415 103.185 207.425 ;
        RECT 101.555 206.775 101.845 207.245 ;
        RECT 102.015 206.945 102.345 207.415 ;
        RECT 102.515 206.775 102.685 207.245 ;
        RECT 102.855 206.945 103.185 207.415 ;
        RECT 103.355 206.775 103.630 207.595 ;
        RECT 103.805 207.545 104.555 208.065 ;
        RECT 104.725 207.715 105.475 208.235 ;
        RECT 106.105 208.250 106.375 209.155 ;
        RECT 106.545 208.565 106.875 209.325 ;
        RECT 107.055 208.395 107.225 209.155 ;
        RECT 103.805 206.775 105.475 207.545 ;
        RECT 106.105 207.450 106.275 208.250 ;
        RECT 106.560 208.225 107.225 208.395 ;
        RECT 107.485 208.235 110.075 209.325 ;
        RECT 110.245 208.730 110.680 209.155 ;
        RECT 110.850 208.900 111.235 209.325 ;
        RECT 110.245 208.560 111.235 208.730 ;
        RECT 106.560 208.080 106.730 208.225 ;
        RECT 106.445 207.750 106.730 208.080 ;
        RECT 106.560 207.495 106.730 207.750 ;
        RECT 106.965 207.675 107.295 208.045 ;
        RECT 107.485 207.545 108.695 208.065 ;
        RECT 108.865 207.715 110.075 208.235 ;
        RECT 110.245 207.685 110.730 208.390 ;
        RECT 110.900 208.015 111.235 208.560 ;
        RECT 111.405 208.365 111.830 209.155 ;
        RECT 112.000 208.730 112.275 209.155 ;
        RECT 112.445 208.900 112.830 209.325 ;
        RECT 112.000 208.535 112.830 208.730 ;
        RECT 111.405 208.185 112.310 208.365 ;
        RECT 110.900 207.685 111.310 208.015 ;
        RECT 111.480 207.685 112.310 208.185 ;
        RECT 112.480 208.015 112.830 208.535 ;
        RECT 113.000 208.365 113.245 209.155 ;
        RECT 113.435 208.730 113.690 209.155 ;
        RECT 113.860 208.900 114.245 209.325 ;
        RECT 113.435 208.535 114.245 208.730 ;
        RECT 113.000 208.185 113.725 208.365 ;
        RECT 112.480 207.685 112.905 208.015 ;
        RECT 113.075 207.685 113.725 208.185 ;
        RECT 113.895 208.015 114.245 208.535 ;
        RECT 114.415 208.185 114.675 209.155 ;
        RECT 113.895 207.685 114.320 208.015 ;
        RECT 106.105 206.945 106.365 207.450 ;
        RECT 106.560 207.325 107.225 207.495 ;
        RECT 106.545 206.775 106.875 207.155 ;
        RECT 107.055 206.945 107.225 207.325 ;
        RECT 107.485 206.775 110.075 207.545 ;
        RECT 110.900 207.515 111.235 207.685 ;
        RECT 111.480 207.515 111.830 207.685 ;
        RECT 112.480 207.515 112.830 207.685 ;
        RECT 113.075 207.515 113.245 207.685 ;
        RECT 113.895 207.515 114.245 207.685 ;
        RECT 114.490 207.515 114.675 208.185 ;
        RECT 110.245 207.345 111.235 207.515 ;
        RECT 110.245 206.945 110.680 207.345 ;
        RECT 110.850 206.775 111.235 207.175 ;
        RECT 111.405 206.945 111.830 207.515 ;
        RECT 112.020 207.345 112.830 207.515 ;
        RECT 112.020 206.945 112.275 207.345 ;
        RECT 112.445 206.775 112.830 207.175 ;
        RECT 113.000 206.945 113.245 207.515 ;
        RECT 113.435 207.345 114.245 207.515 ;
        RECT 113.435 206.945 113.690 207.345 ;
        RECT 113.860 206.775 114.245 207.175 ;
        RECT 114.415 206.945 114.675 207.515 ;
        RECT 114.850 208.185 115.185 209.155 ;
        RECT 115.355 208.185 115.525 209.325 ;
        RECT 115.695 208.985 117.725 209.155 ;
        RECT 114.850 207.515 115.020 208.185 ;
        RECT 115.695 208.015 115.865 208.985 ;
        RECT 115.190 207.685 115.445 208.015 ;
        RECT 115.670 207.685 115.865 208.015 ;
        RECT 116.035 208.645 117.160 208.815 ;
        RECT 115.275 207.515 115.445 207.685 ;
        RECT 116.035 207.515 116.205 208.645 ;
        RECT 114.850 206.945 115.105 207.515 ;
        RECT 115.275 207.345 116.205 207.515 ;
        RECT 116.375 208.305 117.385 208.475 ;
        RECT 116.375 207.505 116.545 208.305 ;
        RECT 116.030 207.310 116.205 207.345 ;
        RECT 115.275 206.775 115.605 207.175 ;
        RECT 116.030 206.945 116.560 207.310 ;
        RECT 116.750 207.285 117.025 208.105 ;
        RECT 116.745 207.115 117.025 207.285 ;
        RECT 116.750 206.945 117.025 207.115 ;
        RECT 117.195 206.945 117.385 208.305 ;
        RECT 117.555 208.320 117.725 208.985 ;
        RECT 117.895 208.565 118.065 209.325 ;
        RECT 118.300 208.565 118.815 208.975 ;
        RECT 117.555 208.130 118.305 208.320 ;
        RECT 118.475 207.755 118.815 208.565 ;
        RECT 117.585 207.585 118.815 207.755 ;
        RECT 118.985 208.250 119.255 209.155 ;
        RECT 119.425 208.565 119.755 209.325 ;
        RECT 119.935 208.395 120.115 209.155 ;
        RECT 117.565 206.775 118.075 207.310 ;
        RECT 118.295 206.980 118.540 207.585 ;
        RECT 118.985 207.450 119.165 208.250 ;
        RECT 119.440 208.225 120.115 208.395 ;
        RECT 120.445 208.395 120.625 209.155 ;
        RECT 120.805 208.565 121.135 209.325 ;
        RECT 120.445 208.225 121.120 208.395 ;
        RECT 121.305 208.250 121.575 209.155 ;
        RECT 119.440 208.080 119.610 208.225 ;
        RECT 119.335 207.750 119.610 208.080 ;
        RECT 120.950 208.080 121.120 208.225 ;
        RECT 119.440 207.495 119.610 207.750 ;
        RECT 119.835 207.675 120.175 208.045 ;
        RECT 120.385 207.675 120.725 208.045 ;
        RECT 120.950 207.750 121.225 208.080 ;
        RECT 120.950 207.495 121.120 207.750 ;
        RECT 118.985 206.945 119.245 207.450 ;
        RECT 119.440 207.325 120.105 207.495 ;
        RECT 119.425 206.775 119.755 207.155 ;
        RECT 119.935 206.945 120.105 207.325 ;
        RECT 120.455 207.325 121.120 207.495 ;
        RECT 121.395 207.450 121.575 208.250 ;
        RECT 120.455 206.945 120.625 207.325 ;
        RECT 120.805 206.775 121.135 207.155 ;
        RECT 121.315 206.945 121.575 207.450 ;
        RECT 122.665 207.720 122.945 209.155 ;
        RECT 123.115 208.550 123.825 209.325 ;
        RECT 123.995 208.380 124.325 209.155 ;
        RECT 123.175 208.165 124.325 208.380 ;
        RECT 122.665 206.945 123.005 207.720 ;
        RECT 123.175 207.595 123.460 208.165 ;
        RECT 123.645 207.765 124.115 207.995 ;
        RECT 124.520 207.965 124.735 209.080 ;
        RECT 124.915 208.605 125.245 209.325 ;
        RECT 125.025 207.965 125.255 208.305 ;
        RECT 126.345 208.160 126.635 209.325 ;
        RECT 126.810 208.185 127.085 209.155 ;
        RECT 127.295 208.525 127.575 209.325 ;
        RECT 127.745 208.815 128.935 209.105 ;
        RECT 127.745 208.475 128.915 208.645 ;
        RECT 127.745 208.355 127.915 208.475 ;
        RECT 127.255 208.185 127.915 208.355 ;
        RECT 124.285 207.785 124.735 207.965 ;
        RECT 124.285 207.765 124.615 207.785 ;
        RECT 124.925 207.765 125.255 207.965 ;
        RECT 123.175 207.405 123.885 207.595 ;
        RECT 123.585 207.265 123.885 207.405 ;
        RECT 124.075 207.405 125.255 207.595 ;
        RECT 124.075 207.325 124.405 207.405 ;
        RECT 123.585 207.255 123.900 207.265 ;
        RECT 123.585 207.245 123.910 207.255 ;
        RECT 123.585 207.240 123.920 207.245 ;
        RECT 123.175 206.775 123.345 207.235 ;
        RECT 123.585 207.230 123.925 207.240 ;
        RECT 123.585 207.225 123.930 207.230 ;
        RECT 123.585 207.215 123.935 207.225 ;
        RECT 123.585 207.210 123.940 207.215 ;
        RECT 123.585 206.945 123.945 207.210 ;
        RECT 124.575 206.775 124.745 207.235 ;
        RECT 124.915 206.945 125.255 207.405 ;
        RECT 126.345 206.775 126.635 207.500 ;
        RECT 126.810 207.450 126.980 208.185 ;
        RECT 127.255 208.015 127.425 208.185 ;
        RECT 128.225 208.015 128.420 208.305 ;
        RECT 128.590 208.185 128.915 208.475 ;
        RECT 130.025 208.565 130.540 208.975 ;
        RECT 130.775 208.565 130.945 209.325 ;
        RECT 131.115 208.985 133.145 209.155 ;
        RECT 127.150 207.685 127.425 208.015 ;
        RECT 127.595 207.685 128.420 208.015 ;
        RECT 128.590 207.685 128.935 208.015 ;
        RECT 130.025 207.755 130.365 208.565 ;
        RECT 131.115 208.320 131.285 208.985 ;
        RECT 131.680 208.645 132.805 208.815 ;
        RECT 130.535 208.130 131.285 208.320 ;
        RECT 131.455 208.305 132.465 208.475 ;
        RECT 127.255 207.515 127.425 207.685 ;
        RECT 130.025 207.585 131.255 207.755 ;
        RECT 126.810 207.105 127.085 207.450 ;
        RECT 127.255 207.345 128.920 207.515 ;
        RECT 127.275 206.775 127.655 207.175 ;
        RECT 127.825 206.995 127.995 207.345 ;
        RECT 128.165 206.775 128.495 207.175 ;
        RECT 128.665 206.995 128.920 207.345 ;
        RECT 130.300 206.980 130.545 207.585 ;
        RECT 130.765 206.775 131.275 207.310 ;
        RECT 131.455 206.945 131.645 208.305 ;
        RECT 131.815 207.965 132.090 208.105 ;
        RECT 131.815 207.795 132.095 207.965 ;
        RECT 131.815 206.945 132.090 207.795 ;
        RECT 132.295 207.505 132.465 208.305 ;
        RECT 132.635 207.515 132.805 208.645 ;
        RECT 132.975 208.015 133.145 208.985 ;
        RECT 133.315 208.185 133.485 209.325 ;
        RECT 133.655 208.185 133.990 209.155 ;
        RECT 134.165 208.235 135.835 209.325 ;
        RECT 136.470 208.900 136.805 209.325 ;
        RECT 136.975 208.720 137.160 209.125 ;
        RECT 132.975 207.685 133.170 208.015 ;
        RECT 133.395 207.685 133.650 208.015 ;
        RECT 133.395 207.515 133.565 207.685 ;
        RECT 133.820 207.515 133.990 208.185 ;
        RECT 132.635 207.345 133.565 207.515 ;
        RECT 132.635 207.310 132.810 207.345 ;
        RECT 132.280 206.945 132.810 207.310 ;
        RECT 133.235 206.775 133.565 207.175 ;
        RECT 133.735 206.945 133.990 207.515 ;
        RECT 134.165 207.545 134.915 208.065 ;
        RECT 135.085 207.715 135.835 208.235 ;
        RECT 136.495 208.545 137.160 208.720 ;
        RECT 137.365 208.545 137.695 209.325 ;
        RECT 134.165 206.775 135.835 207.545 ;
        RECT 136.495 207.515 136.835 208.545 ;
        RECT 137.865 208.355 138.135 209.125 ;
        RECT 138.305 208.890 143.650 209.325 ;
        RECT 137.005 208.185 138.135 208.355 ;
        RECT 137.005 207.685 137.255 208.185 ;
        RECT 136.495 207.345 137.180 207.515 ;
        RECT 137.435 207.435 137.795 208.015 ;
        RECT 136.470 206.775 136.805 207.175 ;
        RECT 136.975 206.945 137.180 207.345 ;
        RECT 137.965 207.275 138.135 208.185 ;
        RECT 139.890 207.320 140.230 208.150 ;
        RECT 141.710 207.640 142.060 208.890 ;
        RECT 143.825 208.235 147.335 209.325 ;
        RECT 147.505 208.235 148.715 209.325 ;
        RECT 143.825 207.545 145.475 208.065 ;
        RECT 145.645 207.715 147.335 208.235 ;
        RECT 137.390 206.775 137.665 207.255 ;
        RECT 137.875 206.945 138.135 207.275 ;
        RECT 138.305 206.775 143.650 207.320 ;
        RECT 143.825 206.775 147.335 207.545 ;
        RECT 147.505 207.525 148.025 208.065 ;
        RECT 148.195 207.695 148.715 208.235 ;
        RECT 148.885 208.235 150.095 209.325 ;
        RECT 148.885 207.695 149.405 208.235 ;
        RECT 149.575 207.525 150.095 208.065 ;
        RECT 147.505 206.775 148.715 207.525 ;
        RECT 148.885 206.775 150.095 207.525 ;
        RECT 36.100 206.605 150.180 206.775 ;
        RECT 36.185 205.855 37.395 206.605 ;
        RECT 36.185 205.315 36.705 205.855 ;
        RECT 37.565 205.835 41.075 206.605 ;
        RECT 41.245 205.855 42.455 206.605 ;
        RECT 42.625 206.225 43.515 206.395 ;
        RECT 36.875 205.145 37.395 205.685 ;
        RECT 37.565 205.315 39.215 205.835 ;
        RECT 39.385 205.145 41.075 205.665 ;
        RECT 41.245 205.315 41.765 205.855 ;
        RECT 41.935 205.145 42.455 205.685 ;
        RECT 42.625 205.670 43.175 206.055 ;
        RECT 43.345 205.500 43.515 206.225 ;
        RECT 36.185 204.055 37.395 205.145 ;
        RECT 37.565 204.055 41.075 205.145 ;
        RECT 41.245 204.055 42.455 205.145 ;
        RECT 42.625 205.430 43.515 205.500 ;
        RECT 43.685 205.925 43.905 206.385 ;
        RECT 44.075 206.065 44.325 206.605 ;
        RECT 44.495 205.955 44.755 206.435 ;
        RECT 43.685 205.900 43.935 205.925 ;
        RECT 43.685 205.475 44.015 205.900 ;
        RECT 42.625 205.405 43.520 205.430 ;
        RECT 42.625 205.390 43.530 205.405 ;
        RECT 42.625 205.375 43.535 205.390 ;
        RECT 42.625 205.370 43.545 205.375 ;
        RECT 42.625 205.360 43.550 205.370 ;
        RECT 42.625 205.350 43.555 205.360 ;
        RECT 42.625 205.345 43.565 205.350 ;
        RECT 42.625 205.335 43.575 205.345 ;
        RECT 42.625 205.330 43.585 205.335 ;
        RECT 42.625 204.880 42.885 205.330 ;
        RECT 43.250 205.325 43.585 205.330 ;
        RECT 43.250 205.320 43.600 205.325 ;
        RECT 43.250 205.310 43.615 205.320 ;
        RECT 43.250 205.305 43.640 205.310 ;
        RECT 44.185 205.305 44.415 205.700 ;
        RECT 43.250 205.300 44.415 205.305 ;
        RECT 43.280 205.265 44.415 205.300 ;
        RECT 43.315 205.240 44.415 205.265 ;
        RECT 43.345 205.210 44.415 205.240 ;
        RECT 43.365 205.180 44.415 205.210 ;
        RECT 43.385 205.150 44.415 205.180 ;
        RECT 43.455 205.140 44.415 205.150 ;
        RECT 43.480 205.130 44.415 205.140 ;
        RECT 43.500 205.115 44.415 205.130 ;
        RECT 43.520 205.100 44.415 205.115 ;
        RECT 43.525 205.090 44.310 205.100 ;
        RECT 43.540 205.055 44.310 205.090 ;
        RECT 43.055 204.735 43.385 204.980 ;
        RECT 43.555 204.805 44.310 205.055 ;
        RECT 44.585 204.925 44.755 205.955 ;
        RECT 45.015 206.055 45.185 206.345 ;
        RECT 45.355 206.225 45.685 206.605 ;
        RECT 45.015 205.885 45.680 206.055 ;
        RECT 44.930 205.065 45.280 205.715 ;
        RECT 43.055 204.710 43.240 204.735 ;
        RECT 42.625 204.610 43.240 204.710 ;
        RECT 42.625 204.055 43.230 204.610 ;
        RECT 43.405 204.225 43.885 204.565 ;
        RECT 44.055 204.055 44.310 204.600 ;
        RECT 44.480 204.225 44.755 204.925 ;
        RECT 45.450 204.895 45.680 205.885 ;
        RECT 45.015 204.725 45.680 204.895 ;
        RECT 45.015 204.225 45.185 204.725 ;
        RECT 45.355 204.055 45.685 204.555 ;
        RECT 45.855 204.225 46.040 206.345 ;
        RECT 46.295 206.145 46.545 206.605 ;
        RECT 46.715 206.155 47.050 206.325 ;
        RECT 47.245 206.155 47.920 206.325 ;
        RECT 46.715 206.015 46.885 206.155 ;
        RECT 46.210 205.025 46.490 205.975 ;
        RECT 46.660 205.885 46.885 206.015 ;
        RECT 46.660 204.780 46.830 205.885 ;
        RECT 47.055 205.735 47.580 205.955 ;
        RECT 47.000 204.970 47.240 205.565 ;
        RECT 47.410 205.035 47.580 205.735 ;
        RECT 47.750 205.375 47.920 206.155 ;
        RECT 48.240 206.105 48.610 206.605 ;
        RECT 48.790 206.155 49.195 206.325 ;
        RECT 49.365 206.155 50.150 206.325 ;
        RECT 48.790 205.925 48.960 206.155 ;
        RECT 48.130 205.625 48.960 205.925 ;
        RECT 49.345 205.655 49.810 205.985 ;
        RECT 48.130 205.595 48.330 205.625 ;
        RECT 48.450 205.375 48.620 205.445 ;
        RECT 47.750 205.205 48.620 205.375 ;
        RECT 48.110 205.115 48.620 205.205 ;
        RECT 46.660 204.650 46.965 204.780 ;
        RECT 47.410 204.670 47.940 205.035 ;
        RECT 46.280 204.055 46.545 204.515 ;
        RECT 46.715 204.225 46.965 204.650 ;
        RECT 48.110 204.500 48.280 205.115 ;
        RECT 47.175 204.330 48.280 204.500 ;
        RECT 48.450 204.055 48.620 204.855 ;
        RECT 48.790 204.555 48.960 205.625 ;
        RECT 49.130 204.725 49.320 205.445 ;
        RECT 49.490 204.695 49.810 205.655 ;
        RECT 49.980 205.695 50.150 206.155 ;
        RECT 50.425 206.075 50.635 206.605 ;
        RECT 50.895 205.865 51.225 206.390 ;
        RECT 51.395 205.995 51.565 206.605 ;
        RECT 51.735 205.950 52.065 206.385 ;
        RECT 52.285 206.060 57.630 206.605 ;
        RECT 51.735 205.865 52.115 205.950 ;
        RECT 51.025 205.695 51.225 205.865 ;
        RECT 51.890 205.825 52.115 205.865 ;
        RECT 49.980 205.365 50.855 205.695 ;
        RECT 51.025 205.365 51.775 205.695 ;
        RECT 48.790 204.225 49.040 204.555 ;
        RECT 49.980 204.525 50.150 205.365 ;
        RECT 51.025 205.160 51.215 205.365 ;
        RECT 51.945 205.245 52.115 205.825 ;
        RECT 51.900 205.195 52.115 205.245 ;
        RECT 53.870 205.230 54.210 206.060 ;
        RECT 57.805 205.835 61.315 206.605 ;
        RECT 61.945 205.880 62.235 206.605 ;
        RECT 50.320 204.785 51.215 205.160 ;
        RECT 51.725 205.115 52.115 205.195 ;
        RECT 49.265 204.355 50.150 204.525 ;
        RECT 50.330 204.055 50.645 204.555 ;
        RECT 50.875 204.225 51.215 204.785 ;
        RECT 51.385 204.055 51.555 205.065 ;
        RECT 51.725 204.270 52.055 205.115 ;
        RECT 55.690 204.490 56.040 205.740 ;
        RECT 57.805 205.315 59.455 205.835 ;
        RECT 63.330 205.765 63.590 206.605 ;
        RECT 63.765 205.860 64.020 206.435 ;
        RECT 64.190 206.225 64.520 206.605 ;
        RECT 64.735 206.055 64.905 206.435 ;
        RECT 64.190 205.885 64.905 206.055 ;
        RECT 59.625 205.145 61.315 205.665 ;
        RECT 52.285 204.055 57.630 204.490 ;
        RECT 57.805 204.055 61.315 205.145 ;
        RECT 61.945 204.055 62.235 205.220 ;
        RECT 63.330 204.055 63.590 205.205 ;
        RECT 63.765 205.130 63.935 205.860 ;
        RECT 64.190 205.695 64.360 205.885 ;
        RECT 65.205 205.785 65.435 206.605 ;
        RECT 65.605 205.805 65.935 206.435 ;
        RECT 64.105 205.365 64.360 205.695 ;
        RECT 64.190 205.155 64.360 205.365 ;
        RECT 64.640 205.335 64.995 205.705 ;
        RECT 65.185 205.365 65.515 205.615 ;
        RECT 65.685 205.205 65.935 205.805 ;
        RECT 66.105 205.785 66.315 206.605 ;
        RECT 66.545 205.835 70.055 206.605 ;
        RECT 70.225 205.855 71.435 206.605 ;
        RECT 66.545 205.315 68.195 205.835 ;
        RECT 63.765 204.225 64.020 205.130 ;
        RECT 64.190 204.985 64.905 205.155 ;
        RECT 64.190 204.055 64.520 204.815 ;
        RECT 64.735 204.225 64.905 204.985 ;
        RECT 65.205 204.055 65.435 205.195 ;
        RECT 65.605 204.225 65.935 205.205 ;
        RECT 66.105 204.055 66.315 205.195 ;
        RECT 68.365 205.145 70.055 205.665 ;
        RECT 70.225 205.315 70.745 205.855 ;
        RECT 71.605 205.805 71.915 206.605 ;
        RECT 72.120 205.805 72.815 206.435 ;
        RECT 72.985 205.835 76.495 206.605 ;
        RECT 77.215 206.055 77.385 206.435 ;
        RECT 77.565 206.225 77.895 206.605 ;
        RECT 77.215 205.885 77.880 206.055 ;
        RECT 78.075 205.930 78.335 206.435 ;
        RECT 78.505 206.060 83.850 206.605 ;
        RECT 70.915 205.145 71.435 205.685 ;
        RECT 71.615 205.365 71.950 205.635 ;
        RECT 72.120 205.205 72.290 205.805 ;
        RECT 72.460 205.365 72.795 205.615 ;
        RECT 72.985 205.315 74.635 205.835 ;
        RECT 66.545 204.055 70.055 205.145 ;
        RECT 70.225 204.055 71.435 205.145 ;
        RECT 71.605 204.055 71.885 205.195 ;
        RECT 72.055 204.225 72.385 205.205 ;
        RECT 72.555 204.055 72.815 205.195 ;
        RECT 74.805 205.145 76.495 205.665 ;
        RECT 77.145 205.335 77.485 205.705 ;
        RECT 77.710 205.630 77.880 205.885 ;
        RECT 77.710 205.300 77.985 205.630 ;
        RECT 77.710 205.155 77.880 205.300 ;
        RECT 72.985 204.055 76.495 205.145 ;
        RECT 77.205 204.985 77.880 205.155 ;
        RECT 78.155 205.130 78.335 205.930 ;
        RECT 80.090 205.230 80.430 206.060 ;
        RECT 84.025 205.805 84.720 206.435 ;
        RECT 84.925 205.805 85.235 206.605 ;
        RECT 85.570 206.095 85.810 206.605 ;
        RECT 85.990 206.095 86.270 206.425 ;
        RECT 86.500 206.095 86.715 206.605 ;
        RECT 77.205 204.225 77.385 204.985 ;
        RECT 77.565 204.055 77.895 204.815 ;
        RECT 78.065 204.225 78.335 205.130 ;
        RECT 81.910 204.490 82.260 205.740 ;
        RECT 84.045 205.365 84.380 205.615 ;
        RECT 84.550 205.205 84.720 205.805 ;
        RECT 84.890 205.365 85.225 205.635 ;
        RECT 85.465 205.365 85.820 205.925 ;
        RECT 78.505 204.055 83.850 204.490 ;
        RECT 84.025 204.055 84.285 205.195 ;
        RECT 84.455 204.225 84.785 205.205 ;
        RECT 85.990 205.195 86.160 206.095 ;
        RECT 86.330 205.365 86.595 205.925 ;
        RECT 86.885 205.865 87.500 206.435 ;
        RECT 87.705 205.880 87.995 206.605 ;
        RECT 86.845 205.195 87.015 205.695 ;
        RECT 84.955 204.055 85.235 205.195 ;
        RECT 85.590 205.025 87.015 205.195 ;
        RECT 85.590 204.850 85.980 205.025 ;
        RECT 86.465 204.055 86.795 204.855 ;
        RECT 87.185 204.845 87.500 205.865 ;
        RECT 88.290 205.825 88.585 206.605 ;
        RECT 89.160 206.075 89.490 206.435 ;
        RECT 89.950 206.245 90.280 206.605 ;
        RECT 90.500 206.075 90.700 206.435 ;
        RECT 89.160 205.905 90.700 206.075 ;
        RECT 88.425 205.395 88.835 205.655 ;
        RECT 88.545 205.245 88.835 205.395 ;
        RECT 89.005 205.365 89.615 205.695 ;
        RECT 89.795 205.445 90.125 205.615 ;
        RECT 86.965 204.225 87.500 204.845 ;
        RECT 87.705 204.055 87.995 205.220 ;
        RECT 88.545 205.195 88.855 205.245 ;
        RECT 89.795 205.195 90.120 205.445 ;
        RECT 88.545 205.015 90.120 205.195 ;
        RECT 88.300 204.665 90.335 204.835 ;
        RECT 88.300 204.585 89.410 204.665 ;
        RECT 88.300 204.225 88.560 204.585 ;
        RECT 88.730 204.055 89.060 204.415 ;
        RECT 89.240 204.225 89.410 204.585 ;
        RECT 89.665 204.055 89.835 204.495 ;
        RECT 90.005 204.405 90.335 204.665 ;
        RECT 90.505 204.575 90.700 205.905 ;
        RECT 90.995 205.805 91.235 206.605 ;
        RECT 91.425 206.160 91.955 206.330 ;
        RECT 91.425 205.620 91.625 206.160 ;
        RECT 92.305 206.060 97.650 206.605 ;
        RECT 97.825 206.060 103.170 206.605 ;
        RECT 103.345 206.060 108.690 206.605 ;
        RECT 90.895 205.405 91.625 205.620 ;
        RECT 90.870 204.405 91.175 204.895 ;
        RECT 91.365 204.425 91.625 205.405 ;
        RECT 91.795 204.885 92.100 205.925 ;
        RECT 93.890 205.230 94.230 206.060 ;
        RECT 90.005 204.225 91.175 204.405 ;
        RECT 91.795 204.055 92.125 204.610 ;
        RECT 95.710 204.490 96.060 205.740 ;
        RECT 99.410 205.230 99.750 206.060 ;
        RECT 101.230 204.490 101.580 205.740 ;
        RECT 104.930 205.230 105.270 206.060 ;
        RECT 108.865 205.835 112.375 206.605 ;
        RECT 113.465 205.880 113.755 206.605 ;
        RECT 106.750 204.490 107.100 205.740 ;
        RECT 108.865 205.315 110.515 205.835 ;
        RECT 110.685 205.145 112.375 205.665 ;
        RECT 113.925 205.660 114.265 206.435 ;
        RECT 114.435 206.145 114.605 206.605 ;
        RECT 114.845 206.170 115.205 206.435 ;
        RECT 114.845 206.165 115.200 206.170 ;
        RECT 114.845 206.155 115.195 206.165 ;
        RECT 114.845 206.150 115.190 206.155 ;
        RECT 114.845 206.140 115.185 206.150 ;
        RECT 115.835 206.145 116.005 206.605 ;
        RECT 114.845 206.135 115.180 206.140 ;
        RECT 114.845 206.125 115.170 206.135 ;
        RECT 114.845 206.115 115.160 206.125 ;
        RECT 114.845 205.975 115.145 206.115 ;
        RECT 114.435 205.785 115.145 205.975 ;
        RECT 115.335 205.975 115.665 206.055 ;
        RECT 116.175 205.975 116.515 206.435 ;
        RECT 115.335 205.785 116.515 205.975 ;
        RECT 92.305 204.055 97.650 204.490 ;
        RECT 97.825 204.055 103.170 204.490 ;
        RECT 103.345 204.055 108.690 204.490 ;
        RECT 108.865 204.055 112.375 205.145 ;
        RECT 113.465 204.055 113.755 205.220 ;
        RECT 113.925 204.225 114.205 205.660 ;
        RECT 114.435 205.215 114.720 205.785 ;
        RECT 116.685 205.660 117.025 206.435 ;
        RECT 117.195 206.145 117.365 206.605 ;
        RECT 117.605 206.170 117.965 206.435 ;
        RECT 117.605 206.165 117.960 206.170 ;
        RECT 117.605 206.155 117.955 206.165 ;
        RECT 117.605 206.150 117.950 206.155 ;
        RECT 117.605 206.140 117.945 206.150 ;
        RECT 118.595 206.145 118.765 206.605 ;
        RECT 117.605 206.135 117.940 206.140 ;
        RECT 117.605 206.125 117.930 206.135 ;
        RECT 117.605 206.115 117.920 206.125 ;
        RECT 117.605 205.975 117.905 206.115 ;
        RECT 117.195 205.785 117.905 205.975 ;
        RECT 118.095 205.975 118.425 206.055 ;
        RECT 118.935 205.975 119.275 206.435 ;
        RECT 118.095 205.785 119.275 205.975 ;
        RECT 119.445 205.835 121.115 206.605 ;
        RECT 121.285 205.930 121.545 206.435 ;
        RECT 121.725 206.225 122.055 206.605 ;
        RECT 122.235 206.055 122.405 206.435 ;
        RECT 114.905 205.385 115.375 205.615 ;
        RECT 115.545 205.595 115.875 205.615 ;
        RECT 115.545 205.415 115.995 205.595 ;
        RECT 116.185 205.415 116.515 205.615 ;
        RECT 114.435 205.000 115.585 205.215 ;
        RECT 114.375 204.055 115.085 204.830 ;
        RECT 115.255 204.225 115.585 205.000 ;
        RECT 115.780 204.300 115.995 205.415 ;
        RECT 116.285 205.075 116.515 205.415 ;
        RECT 116.175 204.055 116.505 204.775 ;
        RECT 116.685 204.225 116.965 205.660 ;
        RECT 117.195 205.215 117.480 205.785 ;
        RECT 117.665 205.385 118.135 205.615 ;
        RECT 118.305 205.595 118.635 205.615 ;
        RECT 118.305 205.415 118.755 205.595 ;
        RECT 118.945 205.415 119.275 205.615 ;
        RECT 117.195 205.000 118.345 205.215 ;
        RECT 117.135 204.055 117.845 204.830 ;
        RECT 118.015 204.225 118.345 205.000 ;
        RECT 118.540 204.300 118.755 205.415 ;
        RECT 119.045 205.075 119.275 205.415 ;
        RECT 119.445 205.315 120.195 205.835 ;
        RECT 120.365 205.145 121.115 205.665 ;
        RECT 118.935 204.055 119.265 204.775 ;
        RECT 119.445 204.055 121.115 205.145 ;
        RECT 121.285 205.130 121.465 205.930 ;
        RECT 121.740 205.885 122.405 206.055 ;
        RECT 122.665 205.930 122.925 206.435 ;
        RECT 123.105 206.225 123.435 206.605 ;
        RECT 123.615 206.055 123.785 206.435 ;
        RECT 121.740 205.630 121.910 205.885 ;
        RECT 121.635 205.300 121.910 205.630 ;
        RECT 122.135 205.335 122.475 205.705 ;
        RECT 121.740 205.155 121.910 205.300 ;
        RECT 121.285 204.225 121.555 205.130 ;
        RECT 121.740 204.985 122.415 205.155 ;
        RECT 121.725 204.055 122.055 204.815 ;
        RECT 122.235 204.225 122.415 204.985 ;
        RECT 122.665 205.130 122.845 205.930 ;
        RECT 123.120 205.885 123.785 206.055 ;
        RECT 123.120 205.630 123.290 205.885 ;
        RECT 124.320 205.795 124.565 206.400 ;
        RECT 124.785 206.070 125.295 206.605 ;
        RECT 123.015 205.300 123.290 205.630 ;
        RECT 123.515 205.335 123.855 205.705 ;
        RECT 124.045 205.625 125.275 205.795 ;
        RECT 123.120 205.155 123.290 205.300 ;
        RECT 122.665 204.225 122.935 205.130 ;
        RECT 123.120 204.985 123.795 205.155 ;
        RECT 123.105 204.055 123.435 204.815 ;
        RECT 123.615 204.225 123.795 204.985 ;
        RECT 124.045 204.815 124.385 205.625 ;
        RECT 124.555 205.060 125.305 205.250 ;
        RECT 124.045 204.405 124.560 204.815 ;
        RECT 124.795 204.055 124.965 204.815 ;
        RECT 125.135 204.395 125.305 205.060 ;
        RECT 125.475 205.075 125.665 206.435 ;
        RECT 125.835 206.265 126.110 206.435 ;
        RECT 125.835 206.095 126.115 206.265 ;
        RECT 125.835 205.275 126.110 206.095 ;
        RECT 126.300 206.070 126.830 206.435 ;
        RECT 127.255 206.205 127.585 206.605 ;
        RECT 126.655 206.035 126.830 206.070 ;
        RECT 126.315 205.075 126.485 205.875 ;
        RECT 125.475 204.905 126.485 205.075 ;
        RECT 126.655 205.865 127.585 206.035 ;
        RECT 127.755 205.865 128.010 206.435 ;
        RECT 128.650 206.205 128.985 206.605 ;
        RECT 129.155 206.035 129.360 206.435 ;
        RECT 129.570 206.125 129.845 206.605 ;
        RECT 130.055 206.105 130.315 206.435 ;
        RECT 126.655 204.735 126.825 205.865 ;
        RECT 127.415 205.695 127.585 205.865 ;
        RECT 125.700 204.565 126.825 204.735 ;
        RECT 126.995 205.365 127.190 205.695 ;
        RECT 127.415 205.365 127.670 205.695 ;
        RECT 126.995 204.395 127.165 205.365 ;
        RECT 127.840 205.195 128.010 205.865 ;
        RECT 125.135 204.225 127.165 204.395 ;
        RECT 127.335 204.055 127.505 205.195 ;
        RECT 127.675 204.225 128.010 205.195 ;
        RECT 128.675 205.865 129.360 206.035 ;
        RECT 128.675 204.835 129.015 205.865 ;
        RECT 129.185 205.195 129.435 205.695 ;
        RECT 129.615 205.365 129.975 205.945 ;
        RECT 130.145 205.195 130.315 206.105 ;
        RECT 130.485 205.835 133.075 206.605 ;
        RECT 133.335 206.055 133.505 206.435 ;
        RECT 133.685 206.225 134.015 206.605 ;
        RECT 133.335 205.885 134.000 206.055 ;
        RECT 134.195 205.930 134.455 206.435 ;
        RECT 130.485 205.315 131.695 205.835 ;
        RECT 129.185 205.025 130.315 205.195 ;
        RECT 131.865 205.145 133.075 205.665 ;
        RECT 133.265 205.335 133.595 205.705 ;
        RECT 133.830 205.630 134.000 205.885 ;
        RECT 133.830 205.300 134.115 205.630 ;
        RECT 133.830 205.155 134.000 205.300 ;
        RECT 128.675 204.660 129.340 204.835 ;
        RECT 128.650 204.055 128.985 204.480 ;
        RECT 129.155 204.255 129.340 204.660 ;
        RECT 129.545 204.055 129.875 204.835 ;
        RECT 130.045 204.255 130.315 205.025 ;
        RECT 130.485 204.055 133.075 205.145 ;
        RECT 133.335 204.985 134.000 205.155 ;
        RECT 134.285 205.130 134.455 205.930 ;
        RECT 134.625 205.835 138.135 206.605 ;
        RECT 139.225 205.880 139.515 206.605 ;
        RECT 140.235 206.055 140.405 206.435 ;
        RECT 140.585 206.225 140.915 206.605 ;
        RECT 140.235 205.885 140.900 206.055 ;
        RECT 141.095 205.930 141.355 206.435 ;
        RECT 134.625 205.315 136.275 205.835 ;
        RECT 136.445 205.145 138.135 205.665 ;
        RECT 140.165 205.335 140.495 205.705 ;
        RECT 140.730 205.630 140.900 205.885 ;
        RECT 140.730 205.300 141.015 205.630 ;
        RECT 133.335 204.225 133.505 204.985 ;
        RECT 133.685 204.055 134.015 204.815 ;
        RECT 134.185 204.225 134.455 205.130 ;
        RECT 134.625 204.055 138.135 205.145 ;
        RECT 139.225 204.055 139.515 205.220 ;
        RECT 140.730 205.155 140.900 205.300 ;
        RECT 140.235 204.985 140.900 205.155 ;
        RECT 141.185 205.130 141.355 205.930 ;
        RECT 141.615 206.055 141.785 206.345 ;
        RECT 141.955 206.225 142.285 206.605 ;
        RECT 141.615 205.885 142.280 206.055 ;
        RECT 140.235 204.225 140.405 204.985 ;
        RECT 140.585 204.055 140.915 204.815 ;
        RECT 141.085 204.225 141.355 205.130 ;
        RECT 141.530 205.065 141.880 205.715 ;
        RECT 142.050 204.895 142.280 205.885 ;
        RECT 141.615 204.725 142.280 204.895 ;
        RECT 141.615 204.225 141.785 204.725 ;
        RECT 141.955 204.055 142.285 204.555 ;
        RECT 142.455 204.225 142.640 206.345 ;
        RECT 142.895 206.145 143.145 206.605 ;
        RECT 143.315 206.155 143.650 206.325 ;
        RECT 143.845 206.155 144.520 206.325 ;
        RECT 143.315 206.015 143.485 206.155 ;
        RECT 142.810 205.025 143.090 205.975 ;
        RECT 143.260 205.885 143.485 206.015 ;
        RECT 143.260 204.780 143.430 205.885 ;
        RECT 143.655 205.735 144.180 205.955 ;
        RECT 143.600 204.970 143.840 205.565 ;
        RECT 144.010 205.035 144.180 205.735 ;
        RECT 144.350 205.375 144.520 206.155 ;
        RECT 144.840 206.105 145.210 206.605 ;
        RECT 145.390 206.155 145.795 206.325 ;
        RECT 145.965 206.155 146.750 206.325 ;
        RECT 145.390 205.925 145.560 206.155 ;
        RECT 144.730 205.625 145.560 205.925 ;
        RECT 145.945 205.655 146.410 205.985 ;
        RECT 144.730 205.595 144.930 205.625 ;
        RECT 145.050 205.375 145.220 205.445 ;
        RECT 144.350 205.205 145.220 205.375 ;
        RECT 144.710 205.115 145.220 205.205 ;
        RECT 143.260 204.650 143.565 204.780 ;
        RECT 144.010 204.670 144.540 205.035 ;
        RECT 142.880 204.055 143.145 204.515 ;
        RECT 143.315 204.225 143.565 204.650 ;
        RECT 144.710 204.500 144.880 205.115 ;
        RECT 143.775 204.330 144.880 204.500 ;
        RECT 145.050 204.055 145.220 204.855 ;
        RECT 145.390 204.555 145.560 205.625 ;
        RECT 145.730 204.725 145.920 205.445 ;
        RECT 146.090 204.695 146.410 205.655 ;
        RECT 146.580 205.695 146.750 206.155 ;
        RECT 147.025 206.075 147.235 206.605 ;
        RECT 147.495 205.865 147.825 206.390 ;
        RECT 147.995 205.995 148.165 206.605 ;
        RECT 148.335 205.950 148.665 206.385 ;
        RECT 148.335 205.865 148.715 205.950 ;
        RECT 147.625 205.695 147.825 205.865 ;
        RECT 148.490 205.825 148.715 205.865 ;
        RECT 148.885 205.855 150.095 206.605 ;
        RECT 146.580 205.365 147.455 205.695 ;
        RECT 147.625 205.365 148.375 205.695 ;
        RECT 145.390 204.225 145.640 204.555 ;
        RECT 146.580 204.525 146.750 205.365 ;
        RECT 147.625 205.160 147.815 205.365 ;
        RECT 148.545 205.245 148.715 205.825 ;
        RECT 148.500 205.195 148.715 205.245 ;
        RECT 146.920 204.785 147.815 205.160 ;
        RECT 148.325 205.115 148.715 205.195 ;
        RECT 148.885 205.145 149.405 205.685 ;
        RECT 149.575 205.315 150.095 205.855 ;
        RECT 145.865 204.355 146.750 204.525 ;
        RECT 146.930 204.055 147.245 204.555 ;
        RECT 147.475 204.225 147.815 204.785 ;
        RECT 147.985 204.055 148.155 205.065 ;
        RECT 148.325 204.270 148.655 205.115 ;
        RECT 148.885 204.055 150.095 205.145 ;
        RECT 36.100 203.885 150.180 204.055 ;
        RECT 36.185 202.795 37.395 203.885 ;
        RECT 37.565 202.795 39.235 203.885 ;
        RECT 36.185 202.085 36.705 202.625 ;
        RECT 36.875 202.255 37.395 202.795 ;
        RECT 37.565 202.105 38.315 202.625 ;
        RECT 38.485 202.275 39.235 202.795 ;
        RECT 39.405 202.745 39.685 203.885 ;
        RECT 39.855 202.735 40.185 203.715 ;
        RECT 40.355 202.745 40.615 203.885 ;
        RECT 40.785 203.330 41.390 203.885 ;
        RECT 41.565 203.375 42.045 203.715 ;
        RECT 42.215 203.340 42.470 203.885 ;
        RECT 40.785 203.230 41.400 203.330 ;
        RECT 41.215 203.205 41.400 203.230 ;
        RECT 39.415 202.305 39.750 202.575 ;
        RECT 39.920 202.135 40.090 202.735 ;
        RECT 40.785 202.610 41.045 203.060 ;
        RECT 41.215 202.960 41.545 203.205 ;
        RECT 41.715 202.885 42.470 203.135 ;
        RECT 42.640 203.015 42.915 203.715 ;
        RECT 41.700 202.850 42.470 202.885 ;
        RECT 41.685 202.840 42.470 202.850 ;
        RECT 41.680 202.825 42.575 202.840 ;
        RECT 41.660 202.810 42.575 202.825 ;
        RECT 41.640 202.800 42.575 202.810 ;
        RECT 41.615 202.790 42.575 202.800 ;
        RECT 41.545 202.760 42.575 202.790 ;
        RECT 41.525 202.730 42.575 202.760 ;
        RECT 41.505 202.700 42.575 202.730 ;
        RECT 41.475 202.675 42.575 202.700 ;
        RECT 41.440 202.640 42.575 202.675 ;
        RECT 41.410 202.635 42.575 202.640 ;
        RECT 41.410 202.630 41.800 202.635 ;
        RECT 41.410 202.620 41.775 202.630 ;
        RECT 41.410 202.615 41.760 202.620 ;
        RECT 41.410 202.610 41.745 202.615 ;
        RECT 40.785 202.605 41.745 202.610 ;
        RECT 40.785 202.595 41.735 202.605 ;
        RECT 40.785 202.590 41.725 202.595 ;
        RECT 40.785 202.580 41.715 202.590 ;
        RECT 40.260 202.325 40.595 202.575 ;
        RECT 40.785 202.570 41.710 202.580 ;
        RECT 40.785 202.565 41.705 202.570 ;
        RECT 40.785 202.550 41.695 202.565 ;
        RECT 40.785 202.535 41.690 202.550 ;
        RECT 40.785 202.510 41.680 202.535 ;
        RECT 40.785 202.440 41.675 202.510 ;
        RECT 36.185 201.335 37.395 202.085 ;
        RECT 37.565 201.335 39.235 202.105 ;
        RECT 39.405 201.335 39.715 202.135 ;
        RECT 39.920 201.505 40.615 202.135 ;
        RECT 40.785 201.885 41.335 202.270 ;
        RECT 41.505 201.715 41.675 202.440 ;
        RECT 40.785 201.545 41.675 201.715 ;
        RECT 41.845 202.040 42.175 202.465 ;
        RECT 42.345 202.240 42.575 202.635 ;
        RECT 41.845 201.555 42.065 202.040 ;
        RECT 42.745 201.985 42.915 203.015 ;
        RECT 43.270 202.915 43.660 203.090 ;
        RECT 44.145 203.085 44.475 203.885 ;
        RECT 44.645 203.095 45.180 203.715 ;
        RECT 43.270 202.745 44.695 202.915 ;
        RECT 43.145 202.015 43.500 202.575 ;
        RECT 42.235 201.335 42.485 201.875 ;
        RECT 42.655 201.505 42.915 201.985 ;
        RECT 43.670 201.845 43.840 202.745 ;
        RECT 44.010 202.015 44.275 202.575 ;
        RECT 44.525 202.245 44.695 202.745 ;
        RECT 44.865 202.075 45.180 203.095 ;
        RECT 45.590 202.915 45.920 203.715 ;
        RECT 46.090 203.085 46.420 203.885 ;
        RECT 46.720 202.915 47.050 203.715 ;
        RECT 47.695 203.085 47.945 203.885 ;
        RECT 45.590 202.745 48.025 202.915 ;
        RECT 48.215 202.745 48.385 203.885 ;
        RECT 48.555 202.745 48.895 203.715 ;
        RECT 45.385 202.325 45.735 202.575 ;
        RECT 45.920 202.115 46.090 202.745 ;
        RECT 46.260 202.325 46.590 202.525 ;
        RECT 46.760 202.325 47.090 202.525 ;
        RECT 47.260 202.355 47.685 202.525 ;
        RECT 47.855 202.495 48.025 202.745 ;
        RECT 47.260 202.325 47.680 202.355 ;
        RECT 47.855 202.325 48.550 202.495 ;
        RECT 43.250 201.335 43.490 201.845 ;
        RECT 43.670 201.515 43.950 201.845 ;
        RECT 44.180 201.335 44.395 201.845 ;
        RECT 44.565 201.505 45.180 202.075 ;
        RECT 45.590 201.505 46.090 202.115 ;
        RECT 46.720 201.985 47.945 202.155 ;
        RECT 48.720 202.135 48.895 202.745 ;
        RECT 49.065 202.720 49.355 203.885 ;
        RECT 49.525 202.745 49.805 203.885 ;
        RECT 49.975 202.735 50.305 203.715 ;
        RECT 50.475 202.745 50.735 203.885 ;
        RECT 50.995 203.215 51.165 203.715 ;
        RECT 51.335 203.385 51.665 203.885 ;
        RECT 50.995 203.045 51.660 203.215 ;
        RECT 49.535 202.305 49.870 202.575 ;
        RECT 50.040 202.135 50.210 202.735 ;
        RECT 50.380 202.325 50.715 202.575 ;
        RECT 50.910 202.225 51.260 202.875 ;
        RECT 46.720 201.505 47.050 201.985 ;
        RECT 47.220 201.335 47.445 201.795 ;
        RECT 47.615 201.505 47.945 201.985 ;
        RECT 48.135 201.335 48.385 202.135 ;
        RECT 48.555 201.505 48.895 202.135 ;
        RECT 49.065 201.335 49.355 202.060 ;
        RECT 49.525 201.335 49.835 202.135 ;
        RECT 50.040 201.505 50.735 202.135 ;
        RECT 51.430 202.055 51.660 203.045 ;
        RECT 50.995 201.885 51.660 202.055 ;
        RECT 50.995 201.595 51.165 201.885 ;
        RECT 51.335 201.335 51.665 201.715 ;
        RECT 51.835 201.595 52.020 203.715 ;
        RECT 52.260 203.425 52.525 203.885 ;
        RECT 52.695 203.290 52.945 203.715 ;
        RECT 53.155 203.440 54.260 203.610 ;
        RECT 52.640 203.160 52.945 203.290 ;
        RECT 52.190 201.965 52.470 202.915 ;
        RECT 52.640 202.055 52.810 203.160 ;
        RECT 52.980 202.375 53.220 202.970 ;
        RECT 53.390 202.905 53.920 203.270 ;
        RECT 53.390 202.205 53.560 202.905 ;
        RECT 54.090 202.825 54.260 203.440 ;
        RECT 54.430 203.085 54.600 203.885 ;
        RECT 54.770 203.385 55.020 203.715 ;
        RECT 55.245 203.415 56.130 203.585 ;
        RECT 54.090 202.735 54.600 202.825 ;
        RECT 52.640 201.925 52.865 202.055 ;
        RECT 53.035 201.985 53.560 202.205 ;
        RECT 53.730 202.565 54.600 202.735 ;
        RECT 52.275 201.335 52.525 201.795 ;
        RECT 52.695 201.785 52.865 201.925 ;
        RECT 53.730 201.785 53.900 202.565 ;
        RECT 54.430 202.495 54.600 202.565 ;
        RECT 54.110 202.315 54.310 202.345 ;
        RECT 54.770 202.315 54.940 203.385 ;
        RECT 55.110 202.495 55.300 203.215 ;
        RECT 54.110 202.015 54.940 202.315 ;
        RECT 55.470 202.285 55.790 203.245 ;
        RECT 52.695 201.615 53.030 201.785 ;
        RECT 53.225 201.615 53.900 201.785 ;
        RECT 54.220 201.335 54.590 201.835 ;
        RECT 54.770 201.785 54.940 202.015 ;
        RECT 55.325 201.955 55.790 202.285 ;
        RECT 55.960 202.575 56.130 203.415 ;
        RECT 56.310 203.385 56.625 203.885 ;
        RECT 56.855 203.155 57.195 203.715 ;
        RECT 56.300 202.780 57.195 203.155 ;
        RECT 57.365 202.875 57.535 203.885 ;
        RECT 57.005 202.575 57.195 202.780 ;
        RECT 57.705 202.825 58.035 203.670 ;
        RECT 58.725 203.125 59.240 203.535 ;
        RECT 59.475 203.125 59.645 203.885 ;
        RECT 59.815 203.545 61.845 203.715 ;
        RECT 57.705 202.745 58.095 202.825 ;
        RECT 57.880 202.695 58.095 202.745 ;
        RECT 55.960 202.245 56.835 202.575 ;
        RECT 57.005 202.245 57.755 202.575 ;
        RECT 55.960 201.785 56.130 202.245 ;
        RECT 57.005 202.075 57.205 202.245 ;
        RECT 57.925 202.115 58.095 202.695 ;
        RECT 58.725 202.315 59.065 203.125 ;
        RECT 59.815 202.880 59.985 203.545 ;
        RECT 60.380 203.205 61.505 203.375 ;
        RECT 59.235 202.690 59.985 202.880 ;
        RECT 60.155 202.865 61.165 203.035 ;
        RECT 58.725 202.145 59.955 202.315 ;
        RECT 57.870 202.075 58.095 202.115 ;
        RECT 54.770 201.615 55.175 201.785 ;
        RECT 55.345 201.615 56.130 201.785 ;
        RECT 56.405 201.335 56.615 201.865 ;
        RECT 56.875 201.550 57.205 202.075 ;
        RECT 57.715 201.990 58.095 202.075 ;
        RECT 57.375 201.335 57.545 201.945 ;
        RECT 57.715 201.555 58.045 201.990 ;
        RECT 59.000 201.540 59.245 202.145 ;
        RECT 59.465 201.335 59.975 201.870 ;
        RECT 60.155 201.505 60.345 202.865 ;
        RECT 60.515 202.525 60.790 202.665 ;
        RECT 60.515 202.355 60.795 202.525 ;
        RECT 60.515 201.505 60.790 202.355 ;
        RECT 60.995 202.065 61.165 202.865 ;
        RECT 61.335 202.075 61.505 203.205 ;
        RECT 61.675 202.575 61.845 203.545 ;
        RECT 62.015 202.745 62.185 203.885 ;
        RECT 62.355 202.745 62.690 203.715 ;
        RECT 61.675 202.245 61.870 202.575 ;
        RECT 62.095 202.245 62.350 202.575 ;
        RECT 62.095 202.075 62.265 202.245 ;
        RECT 62.520 202.075 62.690 202.745 ;
        RECT 61.335 201.905 62.265 202.075 ;
        RECT 61.335 201.870 61.510 201.905 ;
        RECT 60.980 201.505 61.510 201.870 ;
        RECT 61.935 201.335 62.265 201.735 ;
        RECT 62.435 201.505 62.690 202.075 ;
        RECT 62.865 203.085 63.305 203.715 ;
        RECT 62.865 202.075 63.175 203.085 ;
        RECT 63.480 203.035 63.795 203.885 ;
        RECT 63.965 203.545 65.395 203.715 ;
        RECT 63.965 202.865 64.135 203.545 ;
        RECT 63.345 202.695 64.135 202.865 ;
        RECT 63.345 202.245 63.515 202.695 ;
        RECT 64.305 202.575 64.505 203.375 ;
        RECT 63.685 202.245 64.075 202.525 ;
        RECT 64.260 202.245 64.505 202.575 ;
        RECT 64.705 202.245 64.955 203.375 ;
        RECT 65.145 202.915 65.395 203.545 ;
        RECT 65.575 203.085 65.905 203.885 ;
        RECT 65.145 202.745 65.915 202.915 ;
        RECT 66.085 202.745 66.345 203.885 ;
        RECT 65.170 202.245 65.575 202.575 ;
        RECT 65.745 202.075 65.915 202.745 ;
        RECT 66.515 202.735 66.845 203.715 ;
        RECT 67.015 202.745 67.295 203.885 ;
        RECT 67.555 203.215 67.725 203.715 ;
        RECT 67.895 203.385 68.225 203.885 ;
        RECT 67.555 203.045 68.220 203.215 ;
        RECT 66.105 202.325 66.440 202.575 ;
        RECT 66.610 202.185 66.780 202.735 ;
        RECT 66.950 202.305 67.285 202.575 ;
        RECT 67.470 202.225 67.820 202.875 ;
        RECT 66.605 202.135 66.780 202.185 ;
        RECT 62.865 201.515 63.305 202.075 ;
        RECT 63.475 201.335 63.925 202.075 ;
        RECT 64.095 201.905 65.255 202.075 ;
        RECT 64.095 201.505 64.265 201.905 ;
        RECT 64.435 201.335 64.855 201.735 ;
        RECT 65.025 201.505 65.255 201.905 ;
        RECT 65.425 201.505 65.915 202.075 ;
        RECT 66.085 201.505 66.780 202.135 ;
        RECT 66.985 201.335 67.295 202.135 ;
        RECT 67.990 202.055 68.220 203.045 ;
        RECT 67.555 201.885 68.220 202.055 ;
        RECT 67.555 201.595 67.725 201.885 ;
        RECT 67.895 201.335 68.225 201.715 ;
        RECT 68.395 201.595 68.580 203.715 ;
        RECT 68.820 203.425 69.085 203.885 ;
        RECT 69.255 203.290 69.505 203.715 ;
        RECT 69.715 203.440 70.820 203.610 ;
        RECT 69.200 203.160 69.505 203.290 ;
        RECT 68.750 201.965 69.030 202.915 ;
        RECT 69.200 202.055 69.370 203.160 ;
        RECT 69.540 202.375 69.780 202.970 ;
        RECT 69.950 202.905 70.480 203.270 ;
        RECT 69.950 202.205 70.120 202.905 ;
        RECT 70.650 202.825 70.820 203.440 ;
        RECT 70.990 203.085 71.160 203.885 ;
        RECT 71.330 203.385 71.580 203.715 ;
        RECT 71.805 203.415 72.690 203.585 ;
        RECT 70.650 202.735 71.160 202.825 ;
        RECT 69.200 201.925 69.425 202.055 ;
        RECT 69.595 201.985 70.120 202.205 ;
        RECT 70.290 202.565 71.160 202.735 ;
        RECT 68.835 201.335 69.085 201.795 ;
        RECT 69.255 201.785 69.425 201.925 ;
        RECT 70.290 201.785 70.460 202.565 ;
        RECT 70.990 202.495 71.160 202.565 ;
        RECT 70.670 202.315 70.870 202.345 ;
        RECT 71.330 202.315 71.500 203.385 ;
        RECT 71.670 202.495 71.860 203.215 ;
        RECT 70.670 202.015 71.500 202.315 ;
        RECT 72.030 202.285 72.350 203.245 ;
        RECT 69.255 201.615 69.590 201.785 ;
        RECT 69.785 201.615 70.460 201.785 ;
        RECT 70.780 201.335 71.150 201.835 ;
        RECT 71.330 201.785 71.500 202.015 ;
        RECT 71.885 201.955 72.350 202.285 ;
        RECT 72.520 202.575 72.690 203.415 ;
        RECT 72.870 203.385 73.185 203.885 ;
        RECT 73.415 203.155 73.755 203.715 ;
        RECT 72.860 202.780 73.755 203.155 ;
        RECT 73.925 202.875 74.095 203.885 ;
        RECT 73.565 202.575 73.755 202.780 ;
        RECT 74.265 202.825 74.595 203.670 ;
        RECT 74.265 202.745 74.655 202.825 ;
        RECT 74.440 202.695 74.655 202.745 ;
        RECT 74.825 202.720 75.115 203.885 ;
        RECT 75.285 202.795 78.795 203.885 ;
        RECT 72.520 202.245 73.395 202.575 ;
        RECT 73.565 202.245 74.315 202.575 ;
        RECT 72.520 201.785 72.690 202.245 ;
        RECT 73.565 202.075 73.765 202.245 ;
        RECT 74.485 202.115 74.655 202.695 ;
        RECT 74.430 202.075 74.655 202.115 ;
        RECT 71.330 201.615 71.735 201.785 ;
        RECT 71.905 201.615 72.690 201.785 ;
        RECT 72.965 201.335 73.175 201.865 ;
        RECT 73.435 201.550 73.765 202.075 ;
        RECT 74.275 201.990 74.655 202.075 ;
        RECT 75.285 202.105 76.935 202.625 ;
        RECT 77.105 202.275 78.795 202.795 ;
        RECT 79.425 202.280 79.705 203.715 ;
        RECT 79.875 203.110 80.585 203.885 ;
        RECT 80.755 202.940 81.085 203.715 ;
        RECT 79.935 202.725 81.085 202.940 ;
        RECT 73.935 201.335 74.105 201.945 ;
        RECT 74.275 201.555 74.605 201.990 ;
        RECT 74.825 201.335 75.115 202.060 ;
        RECT 75.285 201.335 78.795 202.105 ;
        RECT 79.425 201.505 79.765 202.280 ;
        RECT 79.935 202.155 80.220 202.725 ;
        RECT 80.405 202.325 80.875 202.555 ;
        RECT 81.280 202.525 81.495 203.640 ;
        RECT 81.675 203.165 82.005 203.885 ;
        RECT 81.785 202.525 82.015 202.865 ;
        RECT 82.185 202.795 85.695 203.885 ;
        RECT 81.045 202.345 81.495 202.525 ;
        RECT 81.045 202.325 81.375 202.345 ;
        RECT 81.685 202.325 82.015 202.525 ;
        RECT 79.935 201.965 80.645 202.155 ;
        RECT 80.345 201.825 80.645 201.965 ;
        RECT 80.835 201.965 82.015 202.155 ;
        RECT 80.835 201.885 81.165 201.965 ;
        RECT 80.345 201.815 80.660 201.825 ;
        RECT 80.345 201.805 80.670 201.815 ;
        RECT 80.345 201.800 80.680 201.805 ;
        RECT 79.935 201.335 80.105 201.795 ;
        RECT 80.345 201.790 80.685 201.800 ;
        RECT 80.345 201.785 80.690 201.790 ;
        RECT 80.345 201.775 80.695 201.785 ;
        RECT 80.345 201.770 80.700 201.775 ;
        RECT 80.345 201.505 80.705 201.770 ;
        RECT 81.335 201.335 81.505 201.795 ;
        RECT 81.675 201.505 82.015 201.965 ;
        RECT 82.185 202.105 83.835 202.625 ;
        RECT 84.005 202.275 85.695 202.795 ;
        RECT 86.335 202.825 86.665 203.675 ;
        RECT 86.335 202.695 86.555 202.825 ;
        RECT 86.835 202.745 87.085 203.885 ;
        RECT 87.275 203.245 87.525 203.665 ;
        RECT 87.755 203.415 88.085 203.885 ;
        RECT 88.315 203.245 88.565 203.665 ;
        RECT 87.275 203.075 88.565 203.245 ;
        RECT 88.745 203.245 89.075 203.675 ;
        RECT 88.745 203.075 89.200 203.245 ;
        RECT 82.185 201.335 85.695 202.105 ;
        RECT 86.335 202.060 86.525 202.695 ;
        RECT 87.265 202.575 87.480 202.905 ;
        RECT 86.695 202.245 87.005 202.575 ;
        RECT 87.175 202.245 87.480 202.575 ;
        RECT 87.655 202.245 87.940 202.905 ;
        RECT 88.135 202.245 88.400 202.905 ;
        RECT 88.615 202.245 88.860 202.905 ;
        RECT 86.835 202.075 87.005 202.245 ;
        RECT 89.030 202.075 89.200 203.075 ;
        RECT 86.335 201.550 86.665 202.060 ;
        RECT 86.835 201.905 89.200 202.075 ;
        RECT 89.545 202.280 89.825 203.715 ;
        RECT 89.995 203.110 90.705 203.885 ;
        RECT 90.875 202.940 91.205 203.715 ;
        RECT 90.055 202.725 91.205 202.940 ;
        RECT 86.835 201.335 87.165 201.735 ;
        RECT 88.215 201.565 88.545 201.905 ;
        RECT 88.715 201.335 89.045 201.735 ;
        RECT 89.545 201.505 89.885 202.280 ;
        RECT 90.055 202.155 90.340 202.725 ;
        RECT 90.525 202.325 90.995 202.555 ;
        RECT 91.400 202.525 91.615 203.640 ;
        RECT 91.795 203.165 92.125 203.885 ;
        RECT 92.305 203.450 97.650 203.885 ;
        RECT 91.905 202.525 92.135 202.865 ;
        RECT 91.165 202.345 91.615 202.525 ;
        RECT 91.165 202.325 91.495 202.345 ;
        RECT 91.805 202.325 92.135 202.525 ;
        RECT 90.055 201.965 90.765 202.155 ;
        RECT 90.465 201.825 90.765 201.965 ;
        RECT 90.955 201.965 92.135 202.155 ;
        RECT 90.955 201.885 91.285 201.965 ;
        RECT 90.465 201.815 90.780 201.825 ;
        RECT 90.465 201.805 90.790 201.815 ;
        RECT 90.465 201.800 90.800 201.805 ;
        RECT 90.055 201.335 90.225 201.795 ;
        RECT 90.465 201.790 90.805 201.800 ;
        RECT 90.465 201.785 90.810 201.790 ;
        RECT 90.465 201.775 90.815 201.785 ;
        RECT 90.465 201.770 90.820 201.775 ;
        RECT 90.465 201.505 90.825 201.770 ;
        RECT 91.455 201.335 91.625 201.795 ;
        RECT 91.795 201.505 92.135 201.965 ;
        RECT 93.890 201.880 94.230 202.710 ;
        RECT 95.710 202.200 96.060 203.450 ;
        RECT 97.825 202.280 98.105 203.715 ;
        RECT 98.275 203.110 98.985 203.885 ;
        RECT 99.155 202.940 99.485 203.715 ;
        RECT 98.335 202.725 99.485 202.940 ;
        RECT 92.305 201.335 97.650 201.880 ;
        RECT 97.825 201.505 98.165 202.280 ;
        RECT 98.335 202.155 98.620 202.725 ;
        RECT 98.805 202.325 99.275 202.555 ;
        RECT 99.680 202.525 99.895 203.640 ;
        RECT 100.075 203.165 100.405 203.885 ;
        RECT 100.185 202.525 100.415 202.865 ;
        RECT 100.585 202.720 100.875 203.885 ;
        RECT 101.065 203.375 101.365 203.885 ;
        RECT 101.535 203.375 101.915 203.545 ;
        RECT 102.495 203.375 103.125 203.885 ;
        RECT 101.535 203.205 101.705 203.375 ;
        RECT 103.295 203.205 103.625 203.715 ;
        RECT 103.795 203.375 104.095 203.885 ;
        RECT 101.045 203.005 101.705 203.205 ;
        RECT 101.875 203.035 104.095 203.205 ;
        RECT 104.275 203.165 104.605 203.885 ;
        RECT 99.445 202.345 99.895 202.525 ;
        RECT 99.445 202.325 99.775 202.345 ;
        RECT 100.085 202.325 100.415 202.525 ;
        RECT 98.335 201.965 99.045 202.155 ;
        RECT 98.745 201.825 99.045 201.965 ;
        RECT 99.235 201.965 100.415 202.155 ;
        RECT 101.045 202.075 101.215 203.005 ;
        RECT 101.875 202.835 102.045 203.035 ;
        RECT 101.385 202.665 102.045 202.835 ;
        RECT 102.215 202.695 103.755 202.865 ;
        RECT 101.385 202.245 101.555 202.665 ;
        RECT 102.215 202.495 102.385 202.695 ;
        RECT 101.785 202.325 102.385 202.495 ;
        RECT 102.555 202.325 103.250 202.525 ;
        RECT 103.510 202.245 103.755 202.695 ;
        RECT 101.875 202.075 102.785 202.155 ;
        RECT 99.235 201.885 99.565 201.965 ;
        RECT 98.745 201.815 99.060 201.825 ;
        RECT 98.745 201.805 99.070 201.815 ;
        RECT 98.745 201.800 99.080 201.805 ;
        RECT 98.335 201.335 98.505 201.795 ;
        RECT 98.745 201.790 99.085 201.800 ;
        RECT 98.745 201.785 99.090 201.790 ;
        RECT 98.745 201.775 99.095 201.785 ;
        RECT 98.745 201.770 99.100 201.775 ;
        RECT 98.745 201.505 99.105 201.770 ;
        RECT 99.735 201.335 99.905 201.795 ;
        RECT 100.075 201.505 100.415 201.965 ;
        RECT 100.585 201.335 100.875 202.060 ;
        RECT 101.045 201.595 101.365 202.075 ;
        RECT 101.535 201.985 102.785 202.075 ;
        RECT 101.535 201.905 102.045 201.985 ;
        RECT 101.535 201.505 101.765 201.905 ;
        RECT 101.935 201.335 102.285 201.725 ;
        RECT 102.455 201.505 102.785 201.985 ;
        RECT 102.955 201.335 103.125 202.155 ;
        RECT 103.925 202.075 104.095 203.035 ;
        RECT 104.265 202.525 104.495 202.865 ;
        RECT 104.785 202.525 105.000 203.640 ;
        RECT 105.195 202.940 105.525 203.715 ;
        RECT 105.695 203.110 106.405 203.885 ;
        RECT 105.195 202.725 106.345 202.940 ;
        RECT 104.265 202.325 104.595 202.525 ;
        RECT 104.785 202.345 105.235 202.525 ;
        RECT 104.905 202.325 105.235 202.345 ;
        RECT 105.405 202.325 105.875 202.555 ;
        RECT 106.060 202.155 106.345 202.725 ;
        RECT 106.575 202.280 106.855 203.715 ;
        RECT 107.025 203.450 112.370 203.885 ;
        RECT 103.630 201.530 104.095 202.075 ;
        RECT 104.265 201.965 105.445 202.155 ;
        RECT 104.265 201.505 104.605 201.965 ;
        RECT 105.115 201.885 105.445 201.965 ;
        RECT 105.635 201.965 106.345 202.155 ;
        RECT 105.635 201.825 105.935 201.965 ;
        RECT 105.620 201.815 105.935 201.825 ;
        RECT 105.610 201.805 105.935 201.815 ;
        RECT 105.600 201.800 105.935 201.805 ;
        RECT 104.775 201.335 104.945 201.795 ;
        RECT 105.595 201.790 105.935 201.800 ;
        RECT 105.590 201.785 105.935 201.790 ;
        RECT 105.585 201.775 105.935 201.785 ;
        RECT 105.580 201.770 105.935 201.775 ;
        RECT 105.575 201.505 105.935 201.770 ;
        RECT 106.175 201.335 106.345 201.795 ;
        RECT 106.515 201.505 106.855 202.280 ;
        RECT 108.610 201.880 108.950 202.710 ;
        RECT 110.430 202.200 110.780 203.450 ;
        RECT 112.545 202.795 114.215 203.885 ;
        RECT 112.545 202.105 113.295 202.625 ;
        RECT 113.465 202.275 114.215 202.795 ;
        RECT 114.385 202.280 114.665 203.715 ;
        RECT 114.835 203.110 115.545 203.885 ;
        RECT 115.715 202.940 116.045 203.715 ;
        RECT 114.895 202.725 116.045 202.940 ;
        RECT 107.025 201.335 112.370 201.880 ;
        RECT 112.545 201.335 114.215 202.105 ;
        RECT 114.385 201.505 114.725 202.280 ;
        RECT 114.895 202.155 115.180 202.725 ;
        RECT 115.365 202.325 115.835 202.555 ;
        RECT 116.240 202.525 116.455 203.640 ;
        RECT 116.635 203.165 116.965 203.885 ;
        RECT 117.145 203.450 122.490 203.885 ;
        RECT 116.745 202.525 116.975 202.865 ;
        RECT 116.005 202.345 116.455 202.525 ;
        RECT 116.005 202.325 116.335 202.345 ;
        RECT 116.645 202.325 116.975 202.525 ;
        RECT 114.895 201.965 115.605 202.155 ;
        RECT 115.305 201.825 115.605 201.965 ;
        RECT 115.795 201.965 116.975 202.155 ;
        RECT 115.795 201.885 116.125 201.965 ;
        RECT 115.305 201.815 115.620 201.825 ;
        RECT 115.305 201.805 115.630 201.815 ;
        RECT 115.305 201.800 115.640 201.805 ;
        RECT 114.895 201.335 115.065 201.795 ;
        RECT 115.305 201.790 115.645 201.800 ;
        RECT 115.305 201.785 115.650 201.790 ;
        RECT 115.305 201.775 115.655 201.785 ;
        RECT 115.305 201.770 115.660 201.775 ;
        RECT 115.305 201.505 115.665 201.770 ;
        RECT 116.295 201.335 116.465 201.795 ;
        RECT 116.635 201.505 116.975 201.965 ;
        RECT 118.730 201.880 119.070 202.710 ;
        RECT 120.550 202.200 120.900 203.450 ;
        RECT 123.585 202.280 123.865 203.715 ;
        RECT 124.035 203.110 124.745 203.885 ;
        RECT 124.915 202.940 125.245 203.715 ;
        RECT 124.095 202.725 125.245 202.940 ;
        RECT 117.145 201.335 122.490 201.880 ;
        RECT 123.585 201.505 123.925 202.280 ;
        RECT 124.095 202.155 124.380 202.725 ;
        RECT 124.565 202.325 125.035 202.555 ;
        RECT 125.440 202.525 125.655 203.640 ;
        RECT 125.835 203.165 126.165 203.885 ;
        RECT 125.945 202.525 126.175 202.865 ;
        RECT 126.345 202.720 126.635 203.885 ;
        RECT 126.805 202.745 127.065 203.715 ;
        RECT 127.235 203.460 127.620 203.885 ;
        RECT 127.790 203.290 128.045 203.715 ;
        RECT 127.235 203.095 128.045 203.290 ;
        RECT 125.205 202.345 125.655 202.525 ;
        RECT 125.205 202.325 125.535 202.345 ;
        RECT 125.845 202.325 126.175 202.525 ;
        RECT 124.095 201.965 124.805 202.155 ;
        RECT 124.505 201.825 124.805 201.965 ;
        RECT 124.995 201.965 126.175 202.155 ;
        RECT 126.805 202.075 126.990 202.745 ;
        RECT 127.235 202.575 127.585 203.095 ;
        RECT 128.235 202.925 128.480 203.715 ;
        RECT 128.650 203.460 129.035 203.885 ;
        RECT 129.205 203.290 129.480 203.715 ;
        RECT 127.160 202.245 127.585 202.575 ;
        RECT 127.755 202.745 128.480 202.925 ;
        RECT 128.650 203.095 129.480 203.290 ;
        RECT 127.755 202.245 128.405 202.745 ;
        RECT 128.650 202.575 129.000 203.095 ;
        RECT 129.650 202.925 130.075 203.715 ;
        RECT 130.245 203.460 130.630 203.885 ;
        RECT 130.800 203.290 131.235 203.715 ;
        RECT 128.575 202.245 129.000 202.575 ;
        RECT 129.170 202.745 130.075 202.925 ;
        RECT 130.245 203.120 131.235 203.290 ;
        RECT 129.170 202.245 130.000 202.745 ;
        RECT 130.245 202.575 130.580 203.120 ;
        RECT 130.170 202.245 130.580 202.575 ;
        RECT 130.750 202.245 131.235 202.950 ;
        RECT 131.405 202.810 131.675 203.715 ;
        RECT 131.845 203.125 132.175 203.885 ;
        RECT 132.355 202.955 132.535 203.715 ;
        RECT 127.235 202.075 127.585 202.245 ;
        RECT 128.235 202.075 128.405 202.245 ;
        RECT 128.650 202.075 129.000 202.245 ;
        RECT 129.650 202.075 130.000 202.245 ;
        RECT 130.245 202.075 130.580 202.245 ;
        RECT 124.995 201.885 125.325 201.965 ;
        RECT 124.505 201.815 124.820 201.825 ;
        RECT 124.505 201.805 124.830 201.815 ;
        RECT 124.505 201.800 124.840 201.805 ;
        RECT 124.095 201.335 124.265 201.795 ;
        RECT 124.505 201.790 124.845 201.800 ;
        RECT 124.505 201.785 124.850 201.790 ;
        RECT 124.505 201.775 124.855 201.785 ;
        RECT 124.505 201.770 124.860 201.775 ;
        RECT 124.505 201.505 124.865 201.770 ;
        RECT 125.495 201.335 125.665 201.795 ;
        RECT 125.835 201.505 126.175 201.965 ;
        RECT 126.345 201.335 126.635 202.060 ;
        RECT 126.805 201.505 127.065 202.075 ;
        RECT 127.235 201.905 128.045 202.075 ;
        RECT 127.235 201.335 127.620 201.735 ;
        RECT 127.790 201.505 128.045 201.905 ;
        RECT 128.235 201.505 128.480 202.075 ;
        RECT 128.650 201.905 129.460 202.075 ;
        RECT 128.650 201.335 129.035 201.735 ;
        RECT 129.205 201.505 129.460 201.905 ;
        RECT 129.650 201.505 130.075 202.075 ;
        RECT 130.245 201.905 131.235 202.075 ;
        RECT 130.245 201.335 130.630 201.735 ;
        RECT 130.800 201.505 131.235 201.905 ;
        RECT 131.405 202.010 131.585 202.810 ;
        RECT 131.860 202.785 132.535 202.955 ;
        RECT 132.785 202.795 133.995 203.885 ;
        RECT 134.255 203.215 134.425 203.715 ;
        RECT 134.595 203.385 134.925 203.885 ;
        RECT 134.255 203.045 134.920 203.215 ;
        RECT 131.860 202.640 132.030 202.785 ;
        RECT 131.755 202.310 132.030 202.640 ;
        RECT 131.860 202.055 132.030 202.310 ;
        RECT 132.255 202.235 132.595 202.605 ;
        RECT 132.785 202.085 133.305 202.625 ;
        RECT 133.475 202.255 133.995 202.795 ;
        RECT 134.170 202.225 134.520 202.875 ;
        RECT 131.405 201.505 131.665 202.010 ;
        RECT 131.860 201.885 132.525 202.055 ;
        RECT 131.845 201.335 132.175 201.715 ;
        RECT 132.355 201.505 132.525 201.885 ;
        RECT 132.785 201.335 133.995 202.085 ;
        RECT 134.690 202.055 134.920 203.045 ;
        RECT 134.255 201.885 134.920 202.055 ;
        RECT 134.255 201.595 134.425 201.885 ;
        RECT 134.595 201.335 134.925 201.715 ;
        RECT 135.095 201.595 135.280 203.715 ;
        RECT 135.520 203.425 135.785 203.885 ;
        RECT 135.955 203.290 136.205 203.715 ;
        RECT 136.415 203.440 137.520 203.610 ;
        RECT 135.900 203.160 136.205 203.290 ;
        RECT 135.450 201.965 135.730 202.915 ;
        RECT 135.900 202.055 136.070 203.160 ;
        RECT 136.240 202.375 136.480 202.970 ;
        RECT 136.650 202.905 137.180 203.270 ;
        RECT 136.650 202.205 136.820 202.905 ;
        RECT 137.350 202.825 137.520 203.440 ;
        RECT 137.690 203.085 137.860 203.885 ;
        RECT 138.030 203.385 138.280 203.715 ;
        RECT 138.505 203.415 139.390 203.585 ;
        RECT 137.350 202.735 137.860 202.825 ;
        RECT 135.900 201.925 136.125 202.055 ;
        RECT 136.295 201.985 136.820 202.205 ;
        RECT 136.990 202.565 137.860 202.735 ;
        RECT 135.535 201.335 135.785 201.795 ;
        RECT 135.955 201.785 136.125 201.925 ;
        RECT 136.990 201.785 137.160 202.565 ;
        RECT 137.690 202.495 137.860 202.565 ;
        RECT 137.370 202.315 137.570 202.345 ;
        RECT 138.030 202.315 138.200 203.385 ;
        RECT 138.370 202.495 138.560 203.215 ;
        RECT 137.370 202.015 138.200 202.315 ;
        RECT 138.730 202.285 139.050 203.245 ;
        RECT 135.955 201.615 136.290 201.785 ;
        RECT 136.485 201.615 137.160 201.785 ;
        RECT 137.480 201.335 137.850 201.835 ;
        RECT 138.030 201.785 138.200 202.015 ;
        RECT 138.585 201.955 139.050 202.285 ;
        RECT 139.220 202.575 139.390 203.415 ;
        RECT 139.570 203.385 139.885 203.885 ;
        RECT 140.115 203.155 140.455 203.715 ;
        RECT 139.560 202.780 140.455 203.155 ;
        RECT 140.625 202.875 140.795 203.885 ;
        RECT 140.265 202.575 140.455 202.780 ;
        RECT 140.965 202.825 141.295 203.670 ;
        RECT 140.965 202.745 141.355 202.825 ;
        RECT 141.140 202.695 141.355 202.745 ;
        RECT 139.220 202.245 140.095 202.575 ;
        RECT 140.265 202.245 141.015 202.575 ;
        RECT 139.220 201.785 139.390 202.245 ;
        RECT 140.265 202.075 140.465 202.245 ;
        RECT 141.185 202.115 141.355 202.695 ;
        RECT 141.130 202.075 141.355 202.115 ;
        RECT 138.030 201.615 138.435 201.785 ;
        RECT 138.605 201.615 139.390 201.785 ;
        RECT 139.665 201.335 139.875 201.865 ;
        RECT 140.135 201.550 140.465 202.075 ;
        RECT 140.975 201.990 141.355 202.075 ;
        RECT 141.530 202.745 141.865 203.715 ;
        RECT 142.035 202.745 142.205 203.885 ;
        RECT 142.375 203.545 144.405 203.715 ;
        RECT 141.530 202.075 141.700 202.745 ;
        RECT 142.375 202.575 142.545 203.545 ;
        RECT 141.870 202.245 142.125 202.575 ;
        RECT 142.350 202.245 142.545 202.575 ;
        RECT 142.715 203.205 143.840 203.375 ;
        RECT 141.955 202.075 142.125 202.245 ;
        RECT 142.715 202.075 142.885 203.205 ;
        RECT 140.635 201.335 140.805 201.945 ;
        RECT 140.975 201.555 141.305 201.990 ;
        RECT 141.530 201.505 141.785 202.075 ;
        RECT 141.955 201.905 142.885 202.075 ;
        RECT 143.055 202.865 144.065 203.035 ;
        RECT 143.055 202.065 143.225 202.865 ;
        RECT 143.430 202.185 143.705 202.665 ;
        RECT 143.425 202.015 143.705 202.185 ;
        RECT 142.710 201.870 142.885 201.905 ;
        RECT 141.955 201.335 142.285 201.735 ;
        RECT 142.710 201.505 143.240 201.870 ;
        RECT 143.430 201.505 143.705 202.015 ;
        RECT 143.875 201.505 144.065 202.865 ;
        RECT 144.235 202.880 144.405 203.545 ;
        RECT 144.575 203.125 144.745 203.885 ;
        RECT 144.980 203.125 145.495 203.535 ;
        RECT 144.235 202.690 144.985 202.880 ;
        RECT 145.155 202.315 145.495 203.125 ;
        RECT 145.665 202.795 147.335 203.885 ;
        RECT 144.265 202.145 145.495 202.315 ;
        RECT 144.245 201.335 144.755 201.870 ;
        RECT 144.975 201.540 145.220 202.145 ;
        RECT 145.665 202.105 146.415 202.625 ;
        RECT 146.585 202.275 147.335 202.795 ;
        RECT 147.505 202.810 147.775 203.715 ;
        RECT 147.945 203.125 148.275 203.885 ;
        RECT 148.455 202.955 148.635 203.715 ;
        RECT 145.665 201.335 147.335 202.105 ;
        RECT 147.505 202.010 147.685 202.810 ;
        RECT 147.960 202.785 148.635 202.955 ;
        RECT 148.885 202.795 150.095 203.885 ;
        RECT 147.960 202.640 148.130 202.785 ;
        RECT 147.855 202.310 148.130 202.640 ;
        RECT 147.960 202.055 148.130 202.310 ;
        RECT 148.355 202.235 148.695 202.605 ;
        RECT 148.885 202.255 149.405 202.795 ;
        RECT 149.575 202.085 150.095 202.625 ;
        RECT 147.505 201.505 147.765 202.010 ;
        RECT 147.960 201.885 148.625 202.055 ;
        RECT 147.945 201.335 148.275 201.715 ;
        RECT 148.455 201.505 148.625 201.885 ;
        RECT 148.885 201.335 150.095 202.085 ;
        RECT 36.100 201.165 150.180 201.335 ;
        RECT 36.185 200.415 37.395 201.165 ;
        RECT 36.185 199.875 36.705 200.415 ;
        RECT 37.565 200.395 41.075 201.165 ;
        RECT 41.710 200.675 41.965 201.165 ;
        RECT 42.135 200.655 43.365 200.995 ;
        RECT 36.875 199.705 37.395 200.245 ;
        RECT 37.565 199.875 39.215 200.395 ;
        RECT 39.385 199.705 41.075 200.225 ;
        RECT 41.730 199.925 41.950 200.505 ;
        RECT 42.135 199.755 42.315 200.655 ;
        RECT 42.485 199.925 42.860 200.485 ;
        RECT 43.035 200.425 43.365 200.655 ;
        RECT 43.555 200.440 43.885 200.950 ;
        RECT 44.055 200.765 44.385 201.165 ;
        RECT 45.435 200.595 45.765 200.935 ;
        RECT 45.935 200.765 46.265 201.165 ;
        RECT 46.765 200.665 47.025 200.995 ;
        RECT 47.235 200.685 47.510 201.165 ;
        RECT 43.065 199.925 43.375 200.255 ;
        RECT 36.185 198.615 37.395 199.705 ;
        RECT 37.565 198.615 41.075 199.705 ;
        RECT 41.710 198.615 41.965 199.755 ;
        RECT 42.135 199.585 43.365 199.755 ;
        RECT 42.135 198.785 42.465 199.585 ;
        RECT 42.635 198.615 42.865 199.415 ;
        RECT 43.035 198.785 43.365 199.585 ;
        RECT 43.555 199.675 43.745 200.440 ;
        RECT 44.055 200.425 46.420 200.595 ;
        RECT 44.055 200.255 44.225 200.425 ;
        RECT 43.915 199.925 44.225 200.255 ;
        RECT 44.395 199.925 44.700 200.255 ;
        RECT 43.555 198.825 43.885 199.675 ;
        RECT 44.055 198.615 44.305 199.755 ;
        RECT 44.485 199.595 44.700 199.925 ;
        RECT 44.875 199.595 45.160 200.255 ;
        RECT 45.355 199.595 45.620 200.255 ;
        RECT 45.835 199.595 46.080 200.255 ;
        RECT 46.250 199.425 46.420 200.425 ;
        RECT 44.495 199.255 45.785 199.425 ;
        RECT 44.495 198.835 44.745 199.255 ;
        RECT 44.975 198.615 45.305 199.085 ;
        RECT 45.535 198.835 45.785 199.255 ;
        RECT 45.965 199.255 46.420 199.425 ;
        RECT 46.765 199.755 46.935 200.665 ;
        RECT 47.720 200.595 47.925 200.995 ;
        RECT 48.095 200.765 48.430 201.165 ;
        RECT 48.605 200.595 49.040 200.995 ;
        RECT 49.210 200.765 49.595 201.165 ;
        RECT 47.105 199.925 47.465 200.505 ;
        RECT 47.720 200.425 48.405 200.595 ;
        RECT 48.605 200.425 49.595 200.595 ;
        RECT 49.765 200.425 50.190 200.995 ;
        RECT 50.380 200.595 50.635 200.995 ;
        RECT 50.805 200.765 51.190 201.165 ;
        RECT 50.380 200.425 51.190 200.595 ;
        RECT 51.360 200.425 51.605 200.995 ;
        RECT 51.795 200.595 52.050 200.995 ;
        RECT 52.220 200.765 52.605 201.165 ;
        RECT 51.795 200.425 52.605 200.595 ;
        RECT 52.775 200.425 53.035 200.995 ;
        RECT 47.645 199.755 47.895 200.255 ;
        RECT 46.765 199.585 47.895 199.755 ;
        RECT 45.965 198.825 46.295 199.255 ;
        RECT 46.765 198.815 47.035 199.585 ;
        RECT 48.065 199.395 48.405 200.425 ;
        RECT 49.260 200.255 49.595 200.425 ;
        RECT 49.840 200.255 50.190 200.425 ;
        RECT 50.840 200.255 51.190 200.425 ;
        RECT 51.435 200.255 51.605 200.425 ;
        RECT 52.255 200.255 52.605 200.425 ;
        RECT 48.605 199.550 49.090 200.255 ;
        RECT 49.260 199.925 49.670 200.255 ;
        RECT 47.205 198.615 47.535 199.395 ;
        RECT 47.740 199.220 48.405 199.395 ;
        RECT 49.260 199.380 49.595 199.925 ;
        RECT 49.840 199.755 50.670 200.255 ;
        RECT 47.740 198.815 47.925 199.220 ;
        RECT 48.605 199.210 49.595 199.380 ;
        RECT 49.765 199.575 50.670 199.755 ;
        RECT 50.840 199.925 51.265 200.255 ;
        RECT 48.095 198.615 48.430 199.040 ;
        RECT 48.605 198.785 49.040 199.210 ;
        RECT 49.210 198.615 49.595 199.040 ;
        RECT 49.765 198.785 50.190 199.575 ;
        RECT 50.840 199.405 51.190 199.925 ;
        RECT 51.435 199.755 52.085 200.255 ;
        RECT 50.360 199.210 51.190 199.405 ;
        RECT 51.360 199.575 52.085 199.755 ;
        RECT 52.255 199.925 52.680 200.255 ;
        RECT 50.360 198.785 50.635 199.210 ;
        RECT 50.805 198.615 51.190 199.040 ;
        RECT 51.360 198.785 51.605 199.575 ;
        RECT 52.255 199.405 52.605 199.925 ;
        RECT 52.850 199.755 53.035 200.425 ;
        RECT 53.205 200.395 54.875 201.165 ;
        RECT 55.595 200.615 55.765 200.995 ;
        RECT 55.945 200.785 56.275 201.165 ;
        RECT 55.595 200.445 56.260 200.615 ;
        RECT 56.455 200.490 56.715 200.995 ;
        RECT 53.205 199.875 53.955 200.395 ;
        RECT 51.795 199.210 52.605 199.405 ;
        RECT 51.795 198.785 52.050 199.210 ;
        RECT 52.220 198.615 52.605 199.040 ;
        RECT 52.775 198.785 53.035 199.755 ;
        RECT 54.125 199.705 54.875 200.225 ;
        RECT 55.525 199.895 55.865 200.265 ;
        RECT 56.090 200.190 56.260 200.445 ;
        RECT 56.090 199.860 56.365 200.190 ;
        RECT 56.090 199.715 56.260 199.860 ;
        RECT 53.205 198.615 54.875 199.705 ;
        RECT 55.585 199.545 56.260 199.715 ;
        RECT 56.535 199.690 56.715 200.490 ;
        RECT 57.435 200.615 57.605 200.995 ;
        RECT 57.785 200.785 58.115 201.165 ;
        RECT 57.435 200.445 58.100 200.615 ;
        RECT 58.295 200.490 58.555 200.995 ;
        RECT 57.365 199.895 57.705 200.265 ;
        RECT 57.930 200.190 58.100 200.445 ;
        RECT 57.930 199.860 58.205 200.190 ;
        RECT 57.930 199.715 58.100 199.860 ;
        RECT 55.585 198.785 55.765 199.545 ;
        RECT 55.945 198.615 56.275 199.375 ;
        RECT 56.445 198.785 56.715 199.690 ;
        RECT 57.425 199.545 58.100 199.715 ;
        RECT 58.375 199.690 58.555 200.490 ;
        RECT 57.425 198.785 57.605 199.545 ;
        RECT 57.785 198.615 58.115 199.375 ;
        RECT 58.285 198.785 58.555 199.690 ;
        RECT 58.725 200.425 59.215 200.995 ;
        RECT 59.385 200.595 59.615 200.995 ;
        RECT 59.785 200.765 60.205 201.165 ;
        RECT 60.375 200.595 60.545 200.995 ;
        RECT 59.385 200.425 60.545 200.595 ;
        RECT 60.715 200.425 61.165 201.165 ;
        RECT 61.335 200.425 61.775 200.985 ;
        RECT 61.945 200.440 62.235 201.165 ;
        RECT 62.405 200.595 62.840 200.995 ;
        RECT 63.010 200.765 63.395 201.165 ;
        RECT 62.405 200.425 63.395 200.595 ;
        RECT 63.565 200.425 63.990 200.995 ;
        RECT 64.180 200.595 64.435 200.995 ;
        RECT 64.605 200.765 64.990 201.165 ;
        RECT 64.180 200.425 64.990 200.595 ;
        RECT 65.160 200.425 65.405 200.995 ;
        RECT 65.595 200.595 65.850 200.995 ;
        RECT 66.020 200.765 66.405 201.165 ;
        RECT 65.595 200.425 66.405 200.595 ;
        RECT 66.575 200.425 66.835 200.995 ;
        RECT 58.725 199.755 58.895 200.425 ;
        RECT 59.065 199.925 59.470 200.255 ;
        RECT 58.725 199.585 59.495 199.755 ;
        RECT 58.735 198.615 59.065 199.415 ;
        RECT 59.245 198.955 59.495 199.585 ;
        RECT 59.685 199.125 59.935 200.255 ;
        RECT 60.135 199.925 60.380 200.255 ;
        RECT 60.565 199.975 60.955 200.255 ;
        RECT 60.135 199.125 60.335 199.925 ;
        RECT 61.125 199.805 61.295 200.255 ;
        RECT 60.505 199.635 61.295 199.805 ;
        RECT 60.505 198.955 60.675 199.635 ;
        RECT 59.245 198.785 60.675 198.955 ;
        RECT 60.845 198.615 61.160 199.465 ;
        RECT 61.465 199.415 61.775 200.425 ;
        RECT 63.060 200.255 63.395 200.425 ;
        RECT 63.640 200.255 63.990 200.425 ;
        RECT 64.640 200.255 64.990 200.425 ;
        RECT 65.235 200.255 65.405 200.425 ;
        RECT 66.055 200.255 66.405 200.425 ;
        RECT 61.335 198.785 61.775 199.415 ;
        RECT 61.945 198.615 62.235 199.780 ;
        RECT 62.405 199.550 62.890 200.255 ;
        RECT 63.060 199.925 63.470 200.255 ;
        RECT 63.060 199.380 63.395 199.925 ;
        RECT 63.640 199.755 64.470 200.255 ;
        RECT 62.405 199.210 63.395 199.380 ;
        RECT 63.565 199.575 64.470 199.755 ;
        RECT 64.640 199.925 65.065 200.255 ;
        RECT 62.405 198.785 62.840 199.210 ;
        RECT 63.010 198.615 63.395 199.040 ;
        RECT 63.565 198.785 63.990 199.575 ;
        RECT 64.640 199.405 64.990 199.925 ;
        RECT 65.235 199.755 65.885 200.255 ;
        RECT 64.160 199.210 64.990 199.405 ;
        RECT 65.160 199.575 65.885 199.755 ;
        RECT 66.055 199.925 66.480 200.255 ;
        RECT 64.160 198.785 64.435 199.210 ;
        RECT 64.605 198.615 64.990 199.040 ;
        RECT 65.160 198.785 65.405 199.575 ;
        RECT 66.055 199.405 66.405 199.925 ;
        RECT 66.650 199.755 66.835 200.425 ;
        RECT 67.005 200.395 70.515 201.165 ;
        RECT 70.685 200.490 70.945 200.995 ;
        RECT 71.125 200.785 71.455 201.165 ;
        RECT 71.635 200.615 71.805 200.995 ;
        RECT 67.005 199.875 68.655 200.395 ;
        RECT 65.595 199.210 66.405 199.405 ;
        RECT 65.595 198.785 65.850 199.210 ;
        RECT 66.020 198.615 66.405 199.040 ;
        RECT 66.575 198.785 66.835 199.755 ;
        RECT 68.825 199.705 70.515 200.225 ;
        RECT 67.005 198.615 70.515 199.705 ;
        RECT 70.685 199.690 70.855 200.490 ;
        RECT 71.140 200.445 71.805 200.615 ;
        RECT 72.155 200.615 72.325 200.905 ;
        RECT 72.495 200.785 72.825 201.165 ;
        RECT 72.155 200.445 72.820 200.615 ;
        RECT 71.140 200.190 71.310 200.445 ;
        RECT 71.025 199.860 71.310 200.190 ;
        RECT 71.545 199.895 71.875 200.265 ;
        RECT 71.140 199.715 71.310 199.860 ;
        RECT 70.685 198.785 70.955 199.690 ;
        RECT 71.140 199.545 71.805 199.715 ;
        RECT 72.070 199.625 72.420 200.275 ;
        RECT 71.125 198.615 71.455 199.375 ;
        RECT 71.635 198.785 71.805 199.545 ;
        RECT 72.590 199.455 72.820 200.445 ;
        RECT 72.155 199.285 72.820 199.455 ;
        RECT 72.155 198.785 72.325 199.285 ;
        RECT 72.495 198.615 72.825 199.115 ;
        RECT 72.995 198.785 73.180 200.905 ;
        RECT 73.435 200.705 73.685 201.165 ;
        RECT 73.855 200.715 74.190 200.885 ;
        RECT 74.385 200.715 75.060 200.885 ;
        RECT 73.855 200.575 74.025 200.715 ;
        RECT 73.350 199.585 73.630 200.535 ;
        RECT 73.800 200.445 74.025 200.575 ;
        RECT 73.800 199.340 73.970 200.445 ;
        RECT 74.195 200.295 74.720 200.515 ;
        RECT 74.140 199.530 74.380 200.125 ;
        RECT 74.550 199.595 74.720 200.295 ;
        RECT 74.890 199.935 75.060 200.715 ;
        RECT 75.380 200.665 75.750 201.165 ;
        RECT 75.930 200.715 76.335 200.885 ;
        RECT 76.505 200.715 77.290 200.885 ;
        RECT 75.930 200.485 76.100 200.715 ;
        RECT 75.270 200.185 76.100 200.485 ;
        RECT 76.485 200.215 76.950 200.545 ;
        RECT 75.270 200.155 75.470 200.185 ;
        RECT 75.590 199.935 75.760 200.005 ;
        RECT 74.890 199.765 75.760 199.935 ;
        RECT 75.250 199.675 75.760 199.765 ;
        RECT 73.800 199.210 74.105 199.340 ;
        RECT 74.550 199.230 75.080 199.595 ;
        RECT 73.420 198.615 73.685 199.075 ;
        RECT 73.855 198.785 74.105 199.210 ;
        RECT 75.250 199.060 75.420 199.675 ;
        RECT 74.315 198.890 75.420 199.060 ;
        RECT 75.590 198.615 75.760 199.415 ;
        RECT 75.930 199.115 76.100 200.185 ;
        RECT 76.270 199.285 76.460 200.005 ;
        RECT 76.630 199.255 76.950 200.215 ;
        RECT 77.120 200.255 77.290 200.715 ;
        RECT 77.565 200.635 77.775 201.165 ;
        RECT 78.035 200.425 78.365 200.950 ;
        RECT 78.535 200.555 78.705 201.165 ;
        RECT 78.875 200.510 79.205 200.945 ;
        RECT 78.875 200.425 79.255 200.510 ;
        RECT 78.165 200.255 78.365 200.425 ;
        RECT 79.030 200.385 79.255 200.425 ;
        RECT 77.120 199.925 77.995 200.255 ;
        RECT 78.165 199.925 78.915 200.255 ;
        RECT 75.930 198.785 76.180 199.115 ;
        RECT 77.120 199.085 77.290 199.925 ;
        RECT 78.165 199.720 78.355 199.925 ;
        RECT 79.085 199.805 79.255 200.385 ;
        RECT 79.425 200.415 80.635 201.165 ;
        RECT 79.425 199.875 79.945 200.415 ;
        RECT 79.040 199.755 79.255 199.805 ;
        RECT 77.460 199.345 78.355 199.720 ;
        RECT 78.865 199.675 79.255 199.755 ;
        RECT 80.115 199.705 80.635 200.245 ;
        RECT 76.405 198.915 77.290 199.085 ;
        RECT 77.470 198.615 77.785 199.115 ;
        RECT 78.015 198.785 78.355 199.345 ;
        RECT 78.525 198.615 78.695 199.625 ;
        RECT 78.865 198.830 79.195 199.675 ;
        RECT 79.425 198.615 80.635 199.705 ;
        RECT 80.805 200.220 81.145 200.995 ;
        RECT 81.315 200.705 81.485 201.165 ;
        RECT 81.725 200.730 82.085 200.995 ;
        RECT 81.725 200.725 82.080 200.730 ;
        RECT 81.725 200.715 82.075 200.725 ;
        RECT 81.725 200.710 82.070 200.715 ;
        RECT 81.725 200.700 82.065 200.710 ;
        RECT 82.715 200.705 82.885 201.165 ;
        RECT 81.725 200.695 82.060 200.700 ;
        RECT 81.725 200.685 82.050 200.695 ;
        RECT 81.725 200.675 82.040 200.685 ;
        RECT 81.725 200.535 82.025 200.675 ;
        RECT 81.315 200.345 82.025 200.535 ;
        RECT 82.215 200.535 82.545 200.615 ;
        RECT 83.055 200.535 83.395 200.995 ;
        RECT 82.215 200.345 83.395 200.535 ;
        RECT 83.565 200.395 86.155 201.165 ;
        RECT 80.805 198.785 81.085 200.220 ;
        RECT 81.315 199.775 81.600 200.345 ;
        RECT 81.785 199.945 82.255 200.175 ;
        RECT 82.425 200.155 82.755 200.175 ;
        RECT 82.425 199.975 82.875 200.155 ;
        RECT 83.065 199.975 83.395 200.175 ;
        RECT 81.315 199.560 82.465 199.775 ;
        RECT 81.255 198.615 81.965 199.390 ;
        RECT 82.135 198.785 82.465 199.560 ;
        RECT 82.660 198.860 82.875 199.975 ;
        RECT 83.165 199.635 83.395 199.975 ;
        RECT 83.565 199.875 84.775 200.395 ;
        RECT 86.325 200.365 86.635 201.165 ;
        RECT 86.840 200.365 87.535 200.995 ;
        RECT 87.705 200.440 87.995 201.165 ;
        RECT 88.255 200.615 88.425 200.995 ;
        RECT 88.605 200.785 88.935 201.165 ;
        RECT 88.255 200.445 88.920 200.615 ;
        RECT 89.115 200.490 89.375 200.995 ;
        RECT 89.550 200.765 89.885 201.165 ;
        RECT 90.055 200.595 90.260 200.995 ;
        RECT 90.470 200.685 90.745 201.165 ;
        RECT 90.955 200.665 91.215 200.995 ;
        RECT 84.945 199.705 86.155 200.225 ;
        RECT 86.335 199.925 86.670 200.195 ;
        RECT 86.840 199.765 87.010 200.365 ;
        RECT 87.180 199.925 87.515 200.175 ;
        RECT 88.185 199.895 88.525 200.265 ;
        RECT 88.750 200.190 88.920 200.445 ;
        RECT 88.750 199.860 89.025 200.190 ;
        RECT 83.055 198.615 83.385 199.335 ;
        RECT 83.565 198.615 86.155 199.705 ;
        RECT 86.325 198.615 86.605 199.755 ;
        RECT 86.775 198.785 87.105 199.765 ;
        RECT 87.275 198.615 87.535 199.755 ;
        RECT 87.705 198.615 87.995 199.780 ;
        RECT 88.750 199.715 88.920 199.860 ;
        RECT 88.245 199.545 88.920 199.715 ;
        RECT 89.195 199.690 89.375 200.490 ;
        RECT 88.245 198.785 88.425 199.545 ;
        RECT 88.605 198.615 88.935 199.375 ;
        RECT 89.105 198.785 89.375 199.690 ;
        RECT 89.575 200.425 90.260 200.595 ;
        RECT 89.575 199.395 89.915 200.425 ;
        RECT 90.085 199.755 90.335 200.255 ;
        RECT 90.515 199.925 90.875 200.505 ;
        RECT 91.045 199.755 91.215 200.665 ;
        RECT 91.385 200.395 93.975 201.165 ;
        RECT 94.155 200.440 94.485 200.950 ;
        RECT 94.655 200.765 94.985 201.165 ;
        RECT 96.035 200.595 96.365 200.935 ;
        RECT 96.535 200.765 96.865 201.165 ;
        RECT 97.415 200.775 97.745 201.165 ;
        RECT 97.915 200.595 98.085 200.915 ;
        RECT 98.255 200.775 98.585 201.165 ;
        RECT 99.000 200.765 99.955 200.935 ;
        RECT 91.385 199.875 92.595 200.395 ;
        RECT 90.085 199.585 91.215 199.755 ;
        RECT 92.765 199.705 93.975 200.225 ;
        RECT 89.575 199.220 90.240 199.395 ;
        RECT 89.550 198.615 89.885 199.040 ;
        RECT 90.055 198.815 90.240 199.220 ;
        RECT 90.445 198.615 90.775 199.395 ;
        RECT 90.945 198.815 91.215 199.585 ;
        RECT 91.385 198.615 93.975 199.705 ;
        RECT 94.155 199.675 94.345 200.440 ;
        RECT 94.655 200.425 97.020 200.595 ;
        RECT 94.655 200.255 94.825 200.425 ;
        RECT 94.515 199.925 94.825 200.255 ;
        RECT 94.995 199.925 95.300 200.255 ;
        RECT 94.155 198.825 94.485 199.675 ;
        RECT 94.655 198.615 94.905 199.755 ;
        RECT 95.085 199.595 95.300 199.925 ;
        RECT 95.475 199.595 95.760 200.255 ;
        RECT 95.955 199.595 96.220 200.255 ;
        RECT 96.435 199.595 96.680 200.255 ;
        RECT 96.850 199.425 97.020 200.425 ;
        RECT 95.095 199.255 96.385 199.425 ;
        RECT 95.095 198.835 95.345 199.255 ;
        RECT 95.575 198.615 95.905 199.085 ;
        RECT 96.135 198.835 96.385 199.255 ;
        RECT 96.565 199.255 97.020 199.425 ;
        RECT 97.365 200.425 99.615 200.595 ;
        RECT 97.365 199.465 97.535 200.425 ;
        RECT 97.705 199.805 97.950 200.255 ;
        RECT 98.120 199.975 98.670 200.175 ;
        RECT 98.840 200.005 99.215 200.175 ;
        RECT 98.840 199.805 99.010 200.005 ;
        RECT 99.385 199.925 99.615 200.425 ;
        RECT 97.705 199.635 99.010 199.805 ;
        RECT 99.785 199.885 99.955 200.765 ;
        RECT 100.125 200.330 100.415 201.165 ;
        RECT 100.590 200.400 101.045 201.165 ;
        RECT 101.320 200.785 102.620 200.995 ;
        RECT 102.875 200.805 103.205 201.165 ;
        RECT 102.450 200.635 102.620 200.785 ;
        RECT 103.375 200.665 103.635 200.995 ;
        RECT 103.405 200.655 103.635 200.665 ;
        RECT 101.520 200.175 101.740 200.575 ;
        RECT 100.585 199.975 101.075 200.175 ;
        RECT 101.265 199.965 101.740 200.175 ;
        RECT 101.985 200.175 102.195 200.575 ;
        RECT 102.450 200.510 103.205 200.635 ;
        RECT 102.450 200.465 103.295 200.510 ;
        RECT 103.025 200.345 103.295 200.465 ;
        RECT 101.985 199.965 102.315 200.175 ;
        RECT 102.485 199.905 102.895 200.210 ;
        RECT 99.785 199.715 100.415 199.885 ;
        RECT 96.565 198.825 96.895 199.255 ;
        RECT 97.365 198.785 97.745 199.465 ;
        RECT 98.335 198.615 98.505 199.465 ;
        RECT 98.675 199.295 99.915 199.465 ;
        RECT 98.675 198.785 99.005 199.295 ;
        RECT 99.175 198.615 99.345 199.125 ;
        RECT 99.515 198.785 99.915 199.295 ;
        RECT 100.095 198.785 100.415 199.715 ;
        RECT 100.590 199.735 101.765 199.795 ;
        RECT 103.125 199.770 103.295 200.345 ;
        RECT 103.095 199.735 103.295 199.770 ;
        RECT 100.590 199.625 103.295 199.735 ;
        RECT 100.590 199.005 100.845 199.625 ;
        RECT 101.435 199.565 103.235 199.625 ;
        RECT 101.435 199.535 101.765 199.565 ;
        RECT 103.465 199.465 103.635 200.655 ;
        RECT 103.805 200.620 109.150 201.165 ;
        RECT 105.390 199.790 105.730 200.620 ;
        RECT 109.325 200.395 111.915 201.165 ;
        RECT 112.175 200.615 112.345 200.995 ;
        RECT 112.525 200.785 112.855 201.165 ;
        RECT 112.175 200.445 112.840 200.615 ;
        RECT 113.035 200.490 113.295 200.995 ;
        RECT 101.095 199.365 101.280 199.455 ;
        RECT 101.870 199.365 102.705 199.375 ;
        RECT 101.095 199.165 102.705 199.365 ;
        RECT 101.095 199.125 101.325 199.165 ;
        RECT 100.590 198.785 100.925 199.005 ;
        RECT 101.930 198.615 102.285 198.995 ;
        RECT 102.455 198.785 102.705 199.165 ;
        RECT 102.955 198.615 103.205 199.395 ;
        RECT 103.375 198.785 103.635 199.465 ;
        RECT 107.210 199.050 107.560 200.300 ;
        RECT 109.325 199.875 110.535 200.395 ;
        RECT 110.705 199.705 111.915 200.225 ;
        RECT 112.105 199.895 112.435 200.265 ;
        RECT 112.670 200.190 112.840 200.445 ;
        RECT 112.670 199.860 112.955 200.190 ;
        RECT 112.670 199.715 112.840 199.860 ;
        RECT 103.805 198.615 109.150 199.050 ;
        RECT 109.325 198.615 111.915 199.705 ;
        RECT 112.175 199.545 112.840 199.715 ;
        RECT 113.125 199.690 113.295 200.490 ;
        RECT 113.465 200.440 113.755 201.165 ;
        RECT 113.975 200.510 114.305 200.945 ;
        RECT 114.475 200.555 114.645 201.165 ;
        RECT 113.925 200.425 114.305 200.510 ;
        RECT 114.815 200.425 115.145 200.950 ;
        RECT 115.405 200.635 115.615 201.165 ;
        RECT 115.890 200.715 116.675 200.885 ;
        RECT 116.845 200.715 117.250 200.885 ;
        RECT 113.925 200.385 114.150 200.425 ;
        RECT 113.925 199.805 114.095 200.385 ;
        RECT 114.815 200.255 115.015 200.425 ;
        RECT 115.890 200.255 116.060 200.715 ;
        RECT 114.265 199.925 115.015 200.255 ;
        RECT 115.185 199.925 116.060 200.255 ;
        RECT 112.175 198.785 112.345 199.545 ;
        RECT 112.525 198.615 112.855 199.375 ;
        RECT 113.025 198.785 113.295 199.690 ;
        RECT 113.465 198.615 113.755 199.780 ;
        RECT 113.925 199.755 114.140 199.805 ;
        RECT 113.925 199.675 114.315 199.755 ;
        RECT 113.985 198.830 114.315 199.675 ;
        RECT 114.825 199.720 115.015 199.925 ;
        RECT 114.485 198.615 114.655 199.625 ;
        RECT 114.825 199.345 115.720 199.720 ;
        RECT 114.825 198.785 115.165 199.345 ;
        RECT 115.395 198.615 115.710 199.115 ;
        RECT 115.890 199.085 116.060 199.925 ;
        RECT 116.230 200.215 116.695 200.545 ;
        RECT 117.080 200.485 117.250 200.715 ;
        RECT 117.430 200.665 117.800 201.165 ;
        RECT 118.120 200.715 118.795 200.885 ;
        RECT 118.990 200.715 119.325 200.885 ;
        RECT 116.230 199.255 116.550 200.215 ;
        RECT 117.080 200.185 117.910 200.485 ;
        RECT 116.720 199.285 116.910 200.005 ;
        RECT 117.080 199.115 117.250 200.185 ;
        RECT 117.710 200.155 117.910 200.185 ;
        RECT 117.420 199.935 117.590 200.005 ;
        RECT 118.120 199.935 118.290 200.715 ;
        RECT 119.155 200.575 119.325 200.715 ;
        RECT 119.495 200.705 119.745 201.165 ;
        RECT 117.420 199.765 118.290 199.935 ;
        RECT 118.460 200.295 118.985 200.515 ;
        RECT 119.155 200.445 119.380 200.575 ;
        RECT 117.420 199.675 117.930 199.765 ;
        RECT 115.890 198.915 116.775 199.085 ;
        RECT 117.000 198.785 117.250 199.115 ;
        RECT 117.420 198.615 117.590 199.415 ;
        RECT 117.760 199.060 117.930 199.675 ;
        RECT 118.460 199.595 118.630 200.295 ;
        RECT 118.100 199.230 118.630 199.595 ;
        RECT 118.800 199.530 119.040 200.125 ;
        RECT 119.210 199.340 119.380 200.445 ;
        RECT 119.550 199.585 119.830 200.535 ;
        RECT 119.075 199.210 119.380 199.340 ;
        RECT 117.760 198.890 118.865 199.060 ;
        RECT 119.075 198.785 119.325 199.210 ;
        RECT 119.495 198.615 119.760 199.075 ;
        RECT 120.000 198.785 120.185 200.905 ;
        RECT 120.355 200.785 120.685 201.165 ;
        RECT 120.855 200.615 121.025 200.905 ;
        RECT 120.360 200.445 121.025 200.615 ;
        RECT 120.360 199.455 120.590 200.445 ;
        RECT 121.285 200.395 124.795 201.165 ;
        RECT 120.760 199.625 121.110 200.275 ;
        RECT 121.285 199.875 122.935 200.395 ;
        RECT 125.425 200.365 125.735 201.165 ;
        RECT 125.940 200.365 126.635 200.995 ;
        RECT 126.855 200.510 127.185 200.945 ;
        RECT 127.355 200.555 127.525 201.165 ;
        RECT 126.805 200.425 127.185 200.510 ;
        RECT 127.695 200.425 128.025 200.950 ;
        RECT 128.285 200.635 128.495 201.165 ;
        RECT 128.770 200.715 129.555 200.885 ;
        RECT 129.725 200.715 130.130 200.885 ;
        RECT 126.805 200.385 127.030 200.425 ;
        RECT 123.105 199.705 124.795 200.225 ;
        RECT 125.435 199.925 125.770 200.195 ;
        RECT 125.940 199.765 126.110 200.365 ;
        RECT 126.280 199.925 126.615 200.175 ;
        RECT 126.805 199.805 126.975 200.385 ;
        RECT 127.695 200.255 127.895 200.425 ;
        RECT 128.770 200.255 128.940 200.715 ;
        RECT 127.145 199.925 127.895 200.255 ;
        RECT 128.065 199.925 128.940 200.255 ;
        RECT 120.360 199.285 121.025 199.455 ;
        RECT 120.355 198.615 120.685 199.115 ;
        RECT 120.855 198.785 121.025 199.285 ;
        RECT 121.285 198.615 124.795 199.705 ;
        RECT 125.425 198.615 125.705 199.755 ;
        RECT 125.875 198.785 126.205 199.765 ;
        RECT 126.805 199.755 127.020 199.805 ;
        RECT 126.375 198.615 126.635 199.755 ;
        RECT 126.805 199.675 127.195 199.755 ;
        RECT 126.865 198.830 127.195 199.675 ;
        RECT 127.705 199.720 127.895 199.925 ;
        RECT 127.365 198.615 127.535 199.625 ;
        RECT 127.705 199.345 128.600 199.720 ;
        RECT 127.705 198.785 128.045 199.345 ;
        RECT 128.275 198.615 128.590 199.115 ;
        RECT 128.770 199.085 128.940 199.925 ;
        RECT 129.110 200.215 129.575 200.545 ;
        RECT 129.960 200.485 130.130 200.715 ;
        RECT 130.310 200.665 130.680 201.165 ;
        RECT 131.000 200.715 131.675 200.885 ;
        RECT 131.870 200.715 132.205 200.885 ;
        RECT 129.110 199.255 129.430 200.215 ;
        RECT 129.960 200.185 130.790 200.485 ;
        RECT 129.600 199.285 129.790 200.005 ;
        RECT 129.960 199.115 130.130 200.185 ;
        RECT 130.590 200.155 130.790 200.185 ;
        RECT 130.300 199.935 130.470 200.005 ;
        RECT 131.000 199.935 131.170 200.715 ;
        RECT 132.035 200.575 132.205 200.715 ;
        RECT 132.375 200.705 132.625 201.165 ;
        RECT 130.300 199.765 131.170 199.935 ;
        RECT 131.340 200.295 131.865 200.515 ;
        RECT 132.035 200.445 132.260 200.575 ;
        RECT 130.300 199.675 130.810 199.765 ;
        RECT 128.770 198.915 129.655 199.085 ;
        RECT 129.880 198.785 130.130 199.115 ;
        RECT 130.300 198.615 130.470 199.415 ;
        RECT 130.640 199.060 130.810 199.675 ;
        RECT 131.340 199.595 131.510 200.295 ;
        RECT 130.980 199.230 131.510 199.595 ;
        RECT 131.680 199.530 131.920 200.125 ;
        RECT 132.090 199.340 132.260 200.445 ;
        RECT 132.430 199.585 132.710 200.535 ;
        RECT 131.955 199.210 132.260 199.340 ;
        RECT 130.640 198.890 131.745 199.060 ;
        RECT 131.955 198.785 132.205 199.210 ;
        RECT 132.375 198.615 132.640 199.075 ;
        RECT 132.880 198.785 133.065 200.905 ;
        RECT 133.235 200.785 133.565 201.165 ;
        RECT 133.735 200.615 133.905 200.905 ;
        RECT 133.240 200.445 133.905 200.615 ;
        RECT 133.240 199.455 133.470 200.445 ;
        RECT 134.165 200.395 137.675 201.165 ;
        RECT 137.845 200.415 139.055 201.165 ;
        RECT 139.225 200.440 139.515 201.165 ;
        RECT 139.685 200.620 145.030 201.165 ;
        RECT 133.640 199.625 133.990 200.275 ;
        RECT 134.165 199.875 135.815 200.395 ;
        RECT 135.985 199.705 137.675 200.225 ;
        RECT 137.845 199.875 138.365 200.415 ;
        RECT 138.535 199.705 139.055 200.245 ;
        RECT 141.270 199.790 141.610 200.620 ;
        RECT 145.205 200.395 148.715 201.165 ;
        RECT 148.885 200.415 150.095 201.165 ;
        RECT 133.240 199.285 133.905 199.455 ;
        RECT 133.235 198.615 133.565 199.115 ;
        RECT 133.735 198.785 133.905 199.285 ;
        RECT 134.165 198.615 137.675 199.705 ;
        RECT 137.845 198.615 139.055 199.705 ;
        RECT 139.225 198.615 139.515 199.780 ;
        RECT 143.090 199.050 143.440 200.300 ;
        RECT 145.205 199.875 146.855 200.395 ;
        RECT 147.025 199.705 148.715 200.225 ;
        RECT 139.685 198.615 145.030 199.050 ;
        RECT 145.205 198.615 148.715 199.705 ;
        RECT 148.885 199.705 149.405 200.245 ;
        RECT 149.575 199.875 150.095 200.415 ;
        RECT 148.885 198.615 150.095 199.705 ;
        RECT 36.100 198.445 150.180 198.615 ;
        RECT 36.185 197.355 37.395 198.445 ;
        RECT 37.565 197.355 41.075 198.445 ;
        RECT 36.185 196.645 36.705 197.185 ;
        RECT 36.875 196.815 37.395 197.355 ;
        RECT 37.565 196.665 39.215 197.185 ;
        RECT 39.385 196.835 41.075 197.355 ;
        RECT 41.255 197.305 41.585 198.445 ;
        RECT 42.115 197.475 42.445 198.260 ;
        RECT 41.765 197.305 42.445 197.475 ;
        RECT 42.625 197.355 43.835 198.445 ;
        RECT 41.245 196.885 41.595 197.135 ;
        RECT 41.765 196.705 41.935 197.305 ;
        RECT 42.105 196.885 42.455 197.135 ;
        RECT 36.185 195.895 37.395 196.645 ;
        RECT 37.565 195.895 41.075 196.665 ;
        RECT 41.255 195.895 41.525 196.705 ;
        RECT 41.695 196.065 42.025 196.705 ;
        RECT 42.195 195.895 42.435 196.705 ;
        RECT 42.625 196.645 43.145 197.185 ;
        RECT 43.315 196.815 43.835 197.355 ;
        RECT 44.005 197.725 44.465 198.275 ;
        RECT 44.655 197.725 44.985 198.445 ;
        RECT 42.625 195.895 43.835 196.645 ;
        RECT 44.005 196.355 44.255 197.725 ;
        RECT 45.185 197.555 45.485 198.105 ;
        RECT 45.655 197.775 45.935 198.445 ;
        RECT 44.545 197.385 45.485 197.555 ;
        RECT 44.545 197.135 44.715 197.385 ;
        RECT 45.855 197.135 46.120 197.495 ;
        RECT 46.305 197.355 48.895 198.445 ;
        RECT 44.425 196.805 44.715 197.135 ;
        RECT 44.885 196.885 45.225 197.135 ;
        RECT 45.445 196.885 46.120 197.135 ;
        RECT 44.545 196.715 44.715 196.805 ;
        RECT 44.545 196.525 45.935 196.715 ;
        RECT 44.005 196.065 44.565 196.355 ;
        RECT 44.735 195.895 44.985 196.355 ;
        RECT 45.605 196.165 45.935 196.525 ;
        RECT 46.305 196.665 47.515 197.185 ;
        RECT 47.685 196.835 48.895 197.355 ;
        RECT 49.065 197.280 49.355 198.445 ;
        RECT 49.525 197.850 49.960 198.275 ;
        RECT 50.130 198.020 50.515 198.445 ;
        RECT 49.525 197.680 50.515 197.850 ;
        RECT 49.525 196.805 50.010 197.510 ;
        RECT 50.180 197.135 50.515 197.680 ;
        RECT 50.685 197.485 51.110 198.275 ;
        RECT 51.280 197.850 51.555 198.275 ;
        RECT 51.725 198.020 52.110 198.445 ;
        RECT 51.280 197.655 52.110 197.850 ;
        RECT 50.685 197.305 51.590 197.485 ;
        RECT 50.180 196.805 50.590 197.135 ;
        RECT 50.760 196.805 51.590 197.305 ;
        RECT 51.760 197.135 52.110 197.655 ;
        RECT 52.280 197.485 52.525 198.275 ;
        RECT 52.715 197.850 52.970 198.275 ;
        RECT 53.140 198.020 53.525 198.445 ;
        RECT 52.715 197.655 53.525 197.850 ;
        RECT 52.280 197.305 53.005 197.485 ;
        RECT 51.760 196.805 52.185 197.135 ;
        RECT 52.355 196.805 53.005 197.305 ;
        RECT 53.175 197.135 53.525 197.655 ;
        RECT 53.695 197.305 53.955 198.275 ;
        RECT 55.125 197.515 55.305 198.275 ;
        RECT 55.485 197.685 55.815 198.445 ;
        RECT 55.125 197.345 55.800 197.515 ;
        RECT 55.985 197.370 56.255 198.275 ;
        RECT 53.175 196.805 53.600 197.135 ;
        RECT 46.305 195.895 48.895 196.665 ;
        RECT 50.180 196.635 50.515 196.805 ;
        RECT 50.760 196.635 51.110 196.805 ;
        RECT 51.760 196.635 52.110 196.805 ;
        RECT 52.355 196.635 52.525 196.805 ;
        RECT 53.175 196.635 53.525 196.805 ;
        RECT 53.770 196.635 53.955 197.305 ;
        RECT 55.630 197.200 55.800 197.345 ;
        RECT 55.065 196.795 55.405 197.165 ;
        RECT 55.630 196.870 55.905 197.200 ;
        RECT 49.065 195.895 49.355 196.620 ;
        RECT 49.525 196.465 50.515 196.635 ;
        RECT 49.525 196.065 49.960 196.465 ;
        RECT 50.130 195.895 50.515 196.295 ;
        RECT 50.685 196.065 51.110 196.635 ;
        RECT 51.300 196.465 52.110 196.635 ;
        RECT 51.300 196.065 51.555 196.465 ;
        RECT 51.725 195.895 52.110 196.295 ;
        RECT 52.280 196.065 52.525 196.635 ;
        RECT 52.715 196.465 53.525 196.635 ;
        RECT 52.715 196.065 52.970 196.465 ;
        RECT 53.140 195.895 53.525 196.295 ;
        RECT 53.695 196.065 53.955 196.635 ;
        RECT 55.630 196.615 55.800 196.870 ;
        RECT 55.135 196.445 55.800 196.615 ;
        RECT 56.075 196.570 56.255 197.370 ;
        RECT 55.135 196.065 55.305 196.445 ;
        RECT 55.485 195.895 55.815 196.275 ;
        RECT 55.995 196.065 56.255 196.570 ;
        RECT 56.425 197.370 56.695 198.275 ;
        RECT 56.865 197.685 57.195 198.445 ;
        RECT 57.375 197.515 57.555 198.275 ;
        RECT 56.425 196.570 56.605 197.370 ;
        RECT 56.880 197.345 57.555 197.515 ;
        RECT 57.805 197.370 58.075 198.275 ;
        RECT 58.245 197.685 58.575 198.445 ;
        RECT 58.755 197.515 58.935 198.275 ;
        RECT 56.880 197.200 57.050 197.345 ;
        RECT 56.775 196.870 57.050 197.200 ;
        RECT 56.880 196.615 57.050 196.870 ;
        RECT 57.275 196.795 57.615 197.165 ;
        RECT 56.425 196.065 56.685 196.570 ;
        RECT 56.880 196.445 57.545 196.615 ;
        RECT 56.865 195.895 57.195 196.275 ;
        RECT 57.375 196.065 57.545 196.445 ;
        RECT 57.805 196.570 57.985 197.370 ;
        RECT 58.260 197.345 58.935 197.515 ;
        RECT 59.655 197.385 59.985 198.235 ;
        RECT 58.260 197.200 58.430 197.345 ;
        RECT 58.155 196.870 58.430 197.200 ;
        RECT 58.260 196.615 58.430 196.870 ;
        RECT 58.655 196.795 58.995 197.165 ;
        RECT 59.655 196.620 59.845 197.385 ;
        RECT 60.155 197.305 60.405 198.445 ;
        RECT 60.595 197.805 60.845 198.225 ;
        RECT 61.075 197.975 61.405 198.445 ;
        RECT 61.635 197.805 61.885 198.225 ;
        RECT 60.595 197.635 61.885 197.805 ;
        RECT 62.065 197.805 62.395 198.235 ;
        RECT 63.330 198.020 63.665 198.445 ;
        RECT 63.835 197.840 64.020 198.245 ;
        RECT 62.065 197.635 62.520 197.805 ;
        RECT 60.585 197.135 60.800 197.465 ;
        RECT 60.015 196.805 60.325 197.135 ;
        RECT 60.495 196.805 60.800 197.135 ;
        RECT 60.975 196.805 61.260 197.465 ;
        RECT 61.455 196.805 61.720 197.465 ;
        RECT 61.935 196.805 62.180 197.465 ;
        RECT 60.155 196.635 60.325 196.805 ;
        RECT 62.350 196.635 62.520 197.635 ;
        RECT 57.805 196.065 58.065 196.570 ;
        RECT 58.260 196.445 58.925 196.615 ;
        RECT 58.245 195.895 58.575 196.275 ;
        RECT 58.755 196.065 58.925 196.445 ;
        RECT 59.655 196.110 59.985 196.620 ;
        RECT 60.155 196.465 62.520 196.635 ;
        RECT 63.355 197.665 64.020 197.840 ;
        RECT 64.225 197.665 64.555 198.445 ;
        RECT 63.355 196.635 63.695 197.665 ;
        RECT 64.725 197.475 64.995 198.245 ;
        RECT 63.865 197.305 64.995 197.475 ;
        RECT 63.865 196.805 64.115 197.305 ;
        RECT 63.355 196.465 64.040 196.635 ;
        RECT 64.295 196.555 64.655 197.135 ;
        RECT 60.155 195.895 60.485 196.295 ;
        RECT 61.535 196.125 61.865 196.465 ;
        RECT 62.035 195.895 62.365 196.295 ;
        RECT 63.330 195.895 63.665 196.295 ;
        RECT 63.835 196.065 64.040 196.465 ;
        RECT 64.825 196.395 64.995 197.305 ;
        RECT 64.250 195.895 64.525 196.375 ;
        RECT 64.735 196.065 64.995 196.395 ;
        RECT 66.085 197.475 66.355 198.245 ;
        RECT 66.525 197.665 66.855 198.445 ;
        RECT 67.060 197.840 67.245 198.245 ;
        RECT 67.415 198.020 67.750 198.445 ;
        RECT 67.925 198.010 73.270 198.445 ;
        RECT 67.060 197.665 67.725 197.840 ;
        RECT 66.085 197.305 67.215 197.475 ;
        RECT 66.085 196.395 66.255 197.305 ;
        RECT 66.425 196.555 66.785 197.135 ;
        RECT 66.965 196.805 67.215 197.305 ;
        RECT 67.385 196.635 67.725 197.665 ;
        RECT 67.040 196.465 67.725 196.635 ;
        RECT 66.085 196.065 66.345 196.395 ;
        RECT 66.555 195.895 66.830 196.375 ;
        RECT 67.040 196.065 67.245 196.465 ;
        RECT 69.510 196.440 69.850 197.270 ;
        RECT 71.330 196.760 71.680 198.010 ;
        RECT 73.445 197.355 74.655 198.445 ;
        RECT 73.445 196.645 73.965 197.185 ;
        RECT 74.135 196.815 74.655 197.355 ;
        RECT 74.825 197.280 75.115 198.445 ;
        RECT 75.285 198.010 80.630 198.445 ;
        RECT 67.415 195.895 67.750 196.295 ;
        RECT 67.925 195.895 73.270 196.440 ;
        RECT 73.445 195.895 74.655 196.645 ;
        RECT 74.825 195.895 75.115 196.620 ;
        RECT 76.870 196.440 77.210 197.270 ;
        RECT 78.690 196.760 79.040 198.010 ;
        RECT 80.805 197.355 83.395 198.445 ;
        RECT 80.805 196.665 82.015 197.185 ;
        RECT 82.185 196.835 83.395 197.355 ;
        RECT 84.210 197.475 84.600 197.650 ;
        RECT 85.085 197.645 85.415 198.445 ;
        RECT 85.585 197.655 86.120 198.275 ;
        RECT 84.210 197.305 85.635 197.475 ;
        RECT 75.285 195.895 80.630 196.440 ;
        RECT 80.805 195.895 83.395 196.665 ;
        RECT 84.085 196.575 84.440 197.135 ;
        RECT 84.610 196.405 84.780 197.305 ;
        RECT 84.950 196.575 85.215 197.135 ;
        RECT 85.465 196.805 85.635 197.305 ;
        RECT 85.805 196.635 86.120 197.655 ;
        RECT 84.190 195.895 84.430 196.405 ;
        RECT 84.610 196.075 84.890 196.405 ;
        RECT 85.120 195.895 85.335 196.405 ;
        RECT 85.505 196.065 86.120 196.635 ;
        RECT 86.335 197.385 86.665 198.235 ;
        RECT 86.335 196.620 86.525 197.385 ;
        RECT 86.835 197.305 87.085 198.445 ;
        RECT 87.275 197.805 87.525 198.225 ;
        RECT 87.755 197.975 88.085 198.445 ;
        RECT 88.315 197.805 88.565 198.225 ;
        RECT 87.275 197.635 88.565 197.805 ;
        RECT 88.745 197.805 89.075 198.235 ;
        RECT 88.745 197.635 89.200 197.805 ;
        RECT 87.265 197.135 87.480 197.465 ;
        RECT 86.695 196.805 87.005 197.135 ;
        RECT 87.175 196.805 87.480 197.135 ;
        RECT 87.655 196.805 87.940 197.465 ;
        RECT 88.135 196.805 88.400 197.465 ;
        RECT 88.615 196.805 88.860 197.465 ;
        RECT 86.835 196.635 87.005 196.805 ;
        RECT 89.030 196.635 89.200 197.635 ;
        RECT 86.335 196.110 86.665 196.620 ;
        RECT 86.835 196.465 89.200 196.635 ;
        RECT 89.555 197.385 89.885 198.235 ;
        RECT 89.555 196.620 89.745 197.385 ;
        RECT 90.055 197.305 90.305 198.445 ;
        RECT 90.495 197.805 90.745 198.225 ;
        RECT 90.975 197.975 91.305 198.445 ;
        RECT 91.535 197.805 91.785 198.225 ;
        RECT 90.495 197.635 91.785 197.805 ;
        RECT 91.965 197.805 92.295 198.235 ;
        RECT 92.765 198.010 98.110 198.445 ;
        RECT 91.965 197.635 92.420 197.805 ;
        RECT 90.485 197.135 90.700 197.465 ;
        RECT 89.915 196.805 90.225 197.135 ;
        RECT 90.395 196.805 90.700 197.135 ;
        RECT 90.875 196.805 91.160 197.465 ;
        RECT 91.355 196.805 91.620 197.465 ;
        RECT 91.835 196.805 92.080 197.465 ;
        RECT 90.055 196.635 90.225 196.805 ;
        RECT 92.250 196.635 92.420 197.635 ;
        RECT 86.835 195.895 87.165 196.295 ;
        RECT 88.215 196.125 88.545 196.465 ;
        RECT 88.715 195.895 89.045 196.295 ;
        RECT 89.555 196.110 89.885 196.620 ;
        RECT 90.055 196.465 92.420 196.635 ;
        RECT 90.055 195.895 90.385 196.295 ;
        RECT 91.435 196.125 91.765 196.465 ;
        RECT 94.350 196.440 94.690 197.270 ;
        RECT 96.170 196.760 96.520 198.010 ;
        RECT 98.285 197.355 99.955 198.445 ;
        RECT 98.285 196.665 99.035 197.185 ;
        RECT 99.205 196.835 99.955 197.355 ;
        RECT 100.585 197.280 100.875 198.445 ;
        RECT 101.045 197.595 101.385 198.235 ;
        RECT 101.555 197.985 101.800 198.445 ;
        RECT 101.975 197.815 102.225 198.275 ;
        RECT 102.415 198.065 103.085 198.445 ;
        RECT 103.285 197.815 103.535 198.275 ;
        RECT 101.975 197.645 103.535 197.815 ;
        RECT 91.935 195.895 92.265 196.295 ;
        RECT 92.765 195.895 98.110 196.440 ;
        RECT 98.285 195.895 99.955 196.665 ;
        RECT 100.585 195.895 100.875 196.620 ;
        RECT 101.045 196.480 101.215 197.595 ;
        RECT 104.295 197.475 104.465 198.275 ;
        RECT 101.525 197.305 104.465 197.475 ;
        RECT 104.725 197.575 105.000 198.275 ;
        RECT 105.170 197.900 105.425 198.445 ;
        RECT 105.595 197.935 106.075 198.275 ;
        RECT 106.250 197.890 106.855 198.445 ;
        RECT 106.240 197.790 106.855 197.890 ;
        RECT 106.240 197.765 106.425 197.790 ;
        RECT 101.525 197.135 101.695 197.305 ;
        RECT 101.385 196.805 101.695 197.135 ;
        RECT 101.865 196.805 102.200 197.135 ;
        RECT 101.525 196.635 101.695 196.805 ;
        RECT 101.045 196.065 101.355 196.480 ;
        RECT 101.525 196.465 102.220 196.635 ;
        RECT 102.470 196.560 102.665 197.135 ;
        RECT 102.925 196.805 103.270 197.135 ;
        RECT 103.580 196.805 104.055 197.135 ;
        RECT 104.310 196.805 104.495 197.135 ;
        RECT 102.925 196.575 103.115 196.805 ;
        RECT 101.550 195.895 101.880 196.275 ;
        RECT 102.050 196.235 102.220 196.465 ;
        RECT 103.285 196.465 104.465 196.635 ;
        RECT 103.285 196.235 103.455 196.465 ;
        RECT 102.050 196.065 103.455 196.235 ;
        RECT 103.725 195.895 104.055 196.295 ;
        RECT 104.295 196.065 104.465 196.465 ;
        RECT 104.725 196.545 104.895 197.575 ;
        RECT 105.170 197.445 105.925 197.695 ;
        RECT 106.095 197.520 106.425 197.765 ;
        RECT 105.170 197.410 105.940 197.445 ;
        RECT 105.170 197.400 105.955 197.410 ;
        RECT 105.065 197.385 105.960 197.400 ;
        RECT 105.065 197.370 105.980 197.385 ;
        RECT 105.065 197.360 106.000 197.370 ;
        RECT 105.065 197.350 106.025 197.360 ;
        RECT 105.065 197.320 106.095 197.350 ;
        RECT 105.065 197.290 106.115 197.320 ;
        RECT 105.065 197.260 106.135 197.290 ;
        RECT 105.065 197.235 106.165 197.260 ;
        RECT 105.065 197.200 106.200 197.235 ;
        RECT 105.065 197.195 106.230 197.200 ;
        RECT 105.065 196.800 105.295 197.195 ;
        RECT 105.840 197.190 106.230 197.195 ;
        RECT 105.865 197.180 106.230 197.190 ;
        RECT 105.880 197.175 106.230 197.180 ;
        RECT 105.895 197.170 106.230 197.175 ;
        RECT 106.595 197.170 106.855 197.620 ;
        RECT 107.945 197.305 108.205 198.445 ;
        RECT 108.375 197.295 108.705 198.275 ;
        RECT 108.875 197.305 109.155 198.445 ;
        RECT 109.385 197.305 109.595 198.445 ;
        RECT 109.765 197.295 110.095 198.275 ;
        RECT 110.265 197.305 110.495 198.445 ;
        RECT 110.705 197.355 112.375 198.445 ;
        RECT 105.895 197.165 106.855 197.170 ;
        RECT 105.905 197.155 106.855 197.165 ;
        RECT 105.915 197.150 106.855 197.155 ;
        RECT 105.925 197.140 106.855 197.150 ;
        RECT 105.930 197.130 106.855 197.140 ;
        RECT 105.935 197.125 106.855 197.130 ;
        RECT 105.945 197.110 106.855 197.125 ;
        RECT 105.950 197.095 106.855 197.110 ;
        RECT 105.960 197.070 106.855 197.095 ;
        RECT 105.465 196.600 105.795 197.025 ;
        RECT 104.725 196.065 104.985 196.545 ;
        RECT 105.155 195.895 105.405 196.435 ;
        RECT 105.575 196.115 105.795 196.600 ;
        RECT 105.965 197.000 106.855 197.070 ;
        RECT 105.965 196.275 106.135 197.000 ;
        RECT 107.965 196.885 108.300 197.135 ;
        RECT 106.305 196.445 106.855 196.830 ;
        RECT 108.470 196.695 108.640 197.295 ;
        RECT 108.810 196.865 109.145 197.135 ;
        RECT 105.965 196.105 106.855 196.275 ;
        RECT 107.945 196.065 108.640 196.695 ;
        RECT 108.845 195.895 109.155 196.695 ;
        RECT 109.385 195.895 109.595 196.715 ;
        RECT 109.765 196.695 110.015 197.295 ;
        RECT 110.185 196.885 110.515 197.135 ;
        RECT 109.765 196.065 110.095 196.695 ;
        RECT 110.265 195.895 110.495 196.715 ;
        RECT 110.705 196.665 111.455 197.185 ;
        RECT 111.625 196.835 112.375 197.355 ;
        RECT 113.085 197.515 113.265 198.275 ;
        RECT 113.445 197.685 113.775 198.445 ;
        RECT 113.085 197.345 113.760 197.515 ;
        RECT 113.945 197.370 114.215 198.275 ;
        RECT 113.590 197.200 113.760 197.345 ;
        RECT 113.025 196.795 113.365 197.165 ;
        RECT 113.590 196.870 113.865 197.200 ;
        RECT 110.705 195.895 112.375 196.665 ;
        RECT 113.590 196.615 113.760 196.870 ;
        RECT 113.095 196.445 113.760 196.615 ;
        RECT 114.035 196.570 114.215 197.370 ;
        RECT 113.095 196.065 113.265 196.445 ;
        RECT 113.445 195.895 113.775 196.275 ;
        RECT 113.955 196.065 114.215 196.570 ;
        RECT 114.390 197.305 114.725 198.275 ;
        RECT 114.895 197.305 115.065 198.445 ;
        RECT 115.235 198.105 117.265 198.275 ;
        RECT 114.390 196.635 114.560 197.305 ;
        RECT 115.235 197.135 115.405 198.105 ;
        RECT 114.730 196.805 114.985 197.135 ;
        RECT 115.210 196.805 115.405 197.135 ;
        RECT 115.575 197.765 116.700 197.935 ;
        RECT 114.815 196.635 114.985 196.805 ;
        RECT 115.575 196.635 115.745 197.765 ;
        RECT 114.390 196.065 114.645 196.635 ;
        RECT 114.815 196.465 115.745 196.635 ;
        RECT 115.915 197.425 116.925 197.595 ;
        RECT 115.915 196.625 116.085 197.425 ;
        RECT 116.290 197.085 116.565 197.225 ;
        RECT 116.285 196.915 116.565 197.085 ;
        RECT 115.570 196.430 115.745 196.465 ;
        RECT 114.815 195.895 115.145 196.295 ;
        RECT 115.570 196.065 116.100 196.430 ;
        RECT 116.290 196.065 116.565 196.915 ;
        RECT 116.735 196.065 116.925 197.425 ;
        RECT 117.095 197.440 117.265 198.105 ;
        RECT 117.435 197.685 117.605 198.445 ;
        RECT 117.840 197.685 118.355 198.095 ;
        RECT 117.095 197.250 117.845 197.440 ;
        RECT 118.015 196.875 118.355 197.685 ;
        RECT 117.125 196.705 118.355 196.875 ;
        RECT 119.445 197.475 119.715 198.245 ;
        RECT 119.885 197.665 120.215 198.445 ;
        RECT 120.420 197.840 120.605 198.245 ;
        RECT 120.775 198.020 121.110 198.445 ;
        RECT 120.420 197.665 121.085 197.840 ;
        RECT 119.445 197.305 120.575 197.475 ;
        RECT 117.105 195.895 117.615 196.430 ;
        RECT 117.835 196.100 118.080 196.705 ;
        RECT 119.445 196.395 119.615 197.305 ;
        RECT 119.785 196.555 120.145 197.135 ;
        RECT 120.325 196.805 120.575 197.305 ;
        RECT 120.745 196.635 121.085 197.665 ;
        RECT 121.285 197.355 123.875 198.445 ;
        RECT 120.400 196.465 121.085 196.635 ;
        RECT 121.285 196.665 122.495 197.185 ;
        RECT 122.665 196.835 123.875 197.355 ;
        RECT 124.125 197.515 124.305 198.275 ;
        RECT 124.485 197.685 124.815 198.445 ;
        RECT 124.125 197.345 124.800 197.515 ;
        RECT 124.985 197.370 125.255 198.275 ;
        RECT 124.630 197.200 124.800 197.345 ;
        RECT 124.065 196.795 124.405 197.165 ;
        RECT 124.630 196.870 124.905 197.200 ;
        RECT 119.445 196.065 119.705 196.395 ;
        RECT 119.915 195.895 120.190 196.375 ;
        RECT 120.400 196.065 120.605 196.465 ;
        RECT 120.775 195.895 121.110 196.295 ;
        RECT 121.285 195.895 123.875 196.665 ;
        RECT 124.630 196.615 124.800 196.870 ;
        RECT 124.135 196.445 124.800 196.615 ;
        RECT 125.075 196.570 125.255 197.370 ;
        RECT 126.345 197.280 126.635 198.445 ;
        RECT 126.805 197.305 127.145 198.275 ;
        RECT 127.315 197.305 127.485 198.445 ;
        RECT 127.755 197.645 128.005 198.445 ;
        RECT 128.650 197.475 128.980 198.275 ;
        RECT 129.280 197.645 129.610 198.445 ;
        RECT 129.780 197.475 130.110 198.275 ;
        RECT 130.485 198.010 135.830 198.445 ;
        RECT 127.675 197.305 130.110 197.475 ;
        RECT 126.805 196.695 126.980 197.305 ;
        RECT 127.675 197.055 127.845 197.305 ;
        RECT 127.150 196.885 127.845 197.055 ;
        RECT 128.020 196.885 128.440 197.085 ;
        RECT 128.610 196.885 128.940 197.085 ;
        RECT 129.110 196.885 129.440 197.085 ;
        RECT 124.135 196.065 124.305 196.445 ;
        RECT 124.485 195.895 124.815 196.275 ;
        RECT 124.995 196.065 125.255 196.570 ;
        RECT 126.345 195.895 126.635 196.620 ;
        RECT 126.805 196.065 127.145 196.695 ;
        RECT 127.315 195.895 127.565 196.695 ;
        RECT 127.755 196.545 128.980 196.715 ;
        RECT 127.755 196.065 128.085 196.545 ;
        RECT 128.255 195.895 128.480 196.355 ;
        RECT 128.650 196.065 128.980 196.545 ;
        RECT 129.610 196.675 129.780 197.305 ;
        RECT 129.965 196.885 130.315 197.135 ;
        RECT 129.610 196.065 130.110 196.675 ;
        RECT 132.070 196.440 132.410 197.270 ;
        RECT 133.890 196.760 134.240 198.010 ;
        RECT 136.005 197.355 137.215 198.445 ;
        RECT 136.005 196.645 136.525 197.185 ;
        RECT 136.695 196.815 137.215 197.355 ;
        RECT 137.475 197.515 137.645 198.275 ;
        RECT 137.825 197.685 138.155 198.445 ;
        RECT 137.475 197.345 138.140 197.515 ;
        RECT 138.325 197.370 138.595 198.275 ;
        RECT 139.315 197.775 139.485 198.275 ;
        RECT 139.655 197.945 139.985 198.445 ;
        RECT 139.315 197.605 139.980 197.775 ;
        RECT 137.970 197.200 138.140 197.345 ;
        RECT 137.405 196.795 137.735 197.165 ;
        RECT 137.970 196.870 138.255 197.200 ;
        RECT 130.485 195.895 135.830 196.440 ;
        RECT 136.005 195.895 137.215 196.645 ;
        RECT 137.970 196.615 138.140 196.870 ;
        RECT 137.475 196.445 138.140 196.615 ;
        RECT 138.425 196.570 138.595 197.370 ;
        RECT 139.230 196.785 139.580 197.435 ;
        RECT 139.750 196.615 139.980 197.605 ;
        RECT 137.475 196.065 137.645 196.445 ;
        RECT 137.825 195.895 138.155 196.275 ;
        RECT 138.335 196.065 138.595 196.570 ;
        RECT 139.315 196.445 139.980 196.615 ;
        RECT 139.315 196.155 139.485 196.445 ;
        RECT 139.655 195.895 139.985 196.275 ;
        RECT 140.155 196.155 140.340 198.275 ;
        RECT 140.580 197.985 140.845 198.445 ;
        RECT 141.015 197.850 141.265 198.275 ;
        RECT 141.475 198.000 142.580 198.170 ;
        RECT 140.960 197.720 141.265 197.850 ;
        RECT 140.510 196.525 140.790 197.475 ;
        RECT 140.960 196.615 141.130 197.720 ;
        RECT 141.300 196.935 141.540 197.530 ;
        RECT 141.710 197.465 142.240 197.830 ;
        RECT 141.710 196.765 141.880 197.465 ;
        RECT 142.410 197.385 142.580 198.000 ;
        RECT 142.750 197.645 142.920 198.445 ;
        RECT 143.090 197.945 143.340 198.275 ;
        RECT 143.565 197.975 144.450 198.145 ;
        RECT 142.410 197.295 142.920 197.385 ;
        RECT 140.960 196.485 141.185 196.615 ;
        RECT 141.355 196.545 141.880 196.765 ;
        RECT 142.050 197.125 142.920 197.295 ;
        RECT 140.595 195.895 140.845 196.355 ;
        RECT 141.015 196.345 141.185 196.485 ;
        RECT 142.050 196.345 142.220 197.125 ;
        RECT 142.750 197.055 142.920 197.125 ;
        RECT 142.430 196.875 142.630 196.905 ;
        RECT 143.090 196.875 143.260 197.945 ;
        RECT 143.430 197.055 143.620 197.775 ;
        RECT 142.430 196.575 143.260 196.875 ;
        RECT 143.790 196.845 144.110 197.805 ;
        RECT 141.015 196.175 141.350 196.345 ;
        RECT 141.545 196.175 142.220 196.345 ;
        RECT 142.540 195.895 142.910 196.395 ;
        RECT 143.090 196.345 143.260 196.575 ;
        RECT 143.645 196.515 144.110 196.845 ;
        RECT 144.280 197.135 144.450 197.975 ;
        RECT 144.630 197.945 144.945 198.445 ;
        RECT 145.175 197.715 145.515 198.275 ;
        RECT 144.620 197.340 145.515 197.715 ;
        RECT 145.685 197.435 145.855 198.445 ;
        RECT 145.325 197.135 145.515 197.340 ;
        RECT 146.025 197.385 146.355 198.230 ;
        RECT 146.025 197.305 146.415 197.385 ;
        RECT 146.585 197.355 148.255 198.445 ;
        RECT 146.200 197.255 146.415 197.305 ;
        RECT 144.280 196.805 145.155 197.135 ;
        RECT 145.325 196.805 146.075 197.135 ;
        RECT 144.280 196.345 144.450 196.805 ;
        RECT 145.325 196.635 145.525 196.805 ;
        RECT 146.245 196.675 146.415 197.255 ;
        RECT 146.190 196.635 146.415 196.675 ;
        RECT 143.090 196.175 143.495 196.345 ;
        RECT 143.665 196.175 144.450 196.345 ;
        RECT 144.725 195.895 144.935 196.425 ;
        RECT 145.195 196.110 145.525 196.635 ;
        RECT 146.035 196.550 146.415 196.635 ;
        RECT 146.585 196.665 147.335 197.185 ;
        RECT 147.505 196.835 148.255 197.355 ;
        RECT 148.885 197.355 150.095 198.445 ;
        RECT 148.885 196.815 149.405 197.355 ;
        RECT 145.695 195.895 145.865 196.505 ;
        RECT 146.035 196.115 146.365 196.550 ;
        RECT 146.585 195.895 148.255 196.665 ;
        RECT 149.575 196.645 150.095 197.185 ;
        RECT 148.885 195.895 150.095 196.645 ;
        RECT 36.100 195.725 150.180 195.895 ;
        RECT 36.185 194.975 37.395 195.725 ;
        RECT 36.185 194.435 36.705 194.975 ;
        RECT 37.565 194.955 39.235 195.725 ;
        RECT 39.495 195.175 39.665 195.465 ;
        RECT 39.835 195.345 40.165 195.725 ;
        RECT 39.495 195.005 40.160 195.175 ;
        RECT 36.875 194.265 37.395 194.805 ;
        RECT 37.565 194.435 38.315 194.955 ;
        RECT 38.485 194.265 39.235 194.785 ;
        RECT 36.185 193.175 37.395 194.265 ;
        RECT 37.565 193.175 39.235 194.265 ;
        RECT 39.410 194.185 39.760 194.835 ;
        RECT 39.930 194.015 40.160 195.005 ;
        RECT 39.495 193.845 40.160 194.015 ;
        RECT 39.495 193.345 39.665 193.845 ;
        RECT 39.835 193.175 40.165 193.675 ;
        RECT 40.335 193.345 40.520 195.465 ;
        RECT 40.775 195.265 41.025 195.725 ;
        RECT 41.195 195.275 41.530 195.445 ;
        RECT 41.725 195.275 42.400 195.445 ;
        RECT 41.195 195.135 41.365 195.275 ;
        RECT 40.690 194.145 40.970 195.095 ;
        RECT 41.140 195.005 41.365 195.135 ;
        RECT 41.140 193.900 41.310 195.005 ;
        RECT 41.535 194.855 42.060 195.075 ;
        RECT 41.480 194.090 41.720 194.685 ;
        RECT 41.890 194.155 42.060 194.855 ;
        RECT 42.230 194.495 42.400 195.275 ;
        RECT 42.720 195.225 43.090 195.725 ;
        RECT 43.270 195.275 43.675 195.445 ;
        RECT 43.845 195.275 44.630 195.445 ;
        RECT 43.270 195.045 43.440 195.275 ;
        RECT 42.610 194.745 43.440 195.045 ;
        RECT 43.825 194.775 44.290 195.105 ;
        RECT 42.610 194.715 42.810 194.745 ;
        RECT 42.930 194.495 43.100 194.565 ;
        RECT 42.230 194.325 43.100 194.495 ;
        RECT 42.590 194.235 43.100 194.325 ;
        RECT 41.140 193.770 41.445 193.900 ;
        RECT 41.890 193.790 42.420 194.155 ;
        RECT 40.760 193.175 41.025 193.635 ;
        RECT 41.195 193.345 41.445 193.770 ;
        RECT 42.590 193.620 42.760 194.235 ;
        RECT 41.655 193.450 42.760 193.620 ;
        RECT 42.930 193.175 43.100 193.975 ;
        RECT 43.270 193.675 43.440 194.745 ;
        RECT 43.610 193.845 43.800 194.565 ;
        RECT 43.970 193.815 44.290 194.775 ;
        RECT 44.460 194.815 44.630 195.275 ;
        RECT 44.905 195.195 45.115 195.725 ;
        RECT 45.375 194.985 45.705 195.510 ;
        RECT 45.875 195.115 46.045 195.725 ;
        RECT 46.215 195.070 46.545 195.505 ;
        RECT 46.215 194.985 46.595 195.070 ;
        RECT 45.505 194.815 45.705 194.985 ;
        RECT 46.370 194.945 46.595 194.985 ;
        RECT 44.460 194.485 45.335 194.815 ;
        RECT 45.505 194.485 46.255 194.815 ;
        RECT 43.270 193.345 43.520 193.675 ;
        RECT 44.460 193.645 44.630 194.485 ;
        RECT 45.505 194.280 45.695 194.485 ;
        RECT 46.425 194.365 46.595 194.945 ;
        RECT 46.765 194.955 49.355 195.725 ;
        RECT 49.525 195.050 49.785 195.555 ;
        RECT 49.965 195.345 50.295 195.725 ;
        RECT 50.475 195.175 50.645 195.555 ;
        RECT 46.765 194.435 47.975 194.955 ;
        RECT 46.380 194.315 46.595 194.365 ;
        RECT 44.800 193.905 45.695 194.280 ;
        RECT 46.205 194.235 46.595 194.315 ;
        RECT 48.145 194.265 49.355 194.785 ;
        RECT 43.745 193.475 44.630 193.645 ;
        RECT 44.810 193.175 45.125 193.675 ;
        RECT 45.355 193.345 45.695 193.905 ;
        RECT 45.865 193.175 46.035 194.185 ;
        RECT 46.205 193.390 46.535 194.235 ;
        RECT 46.765 193.175 49.355 194.265 ;
        RECT 49.525 194.250 49.705 195.050 ;
        RECT 49.980 195.005 50.645 195.175 ;
        RECT 49.980 194.750 50.150 195.005 ;
        RECT 50.905 194.975 52.115 195.725 ;
        RECT 49.875 194.420 50.150 194.750 ;
        RECT 50.375 194.455 50.715 194.825 ;
        RECT 50.905 194.435 51.425 194.975 ;
        RECT 52.345 194.905 52.555 195.725 ;
        RECT 52.725 194.925 53.055 195.555 ;
        RECT 49.980 194.275 50.150 194.420 ;
        RECT 49.525 193.345 49.795 194.250 ;
        RECT 49.980 194.105 50.655 194.275 ;
        RECT 51.595 194.265 52.115 194.805 ;
        RECT 52.725 194.325 52.975 194.925 ;
        RECT 53.225 194.905 53.455 195.725 ;
        RECT 53.665 194.925 54.005 195.555 ;
        RECT 54.295 195.265 54.465 195.725 ;
        RECT 54.735 195.095 55.065 195.540 ;
        RECT 53.145 194.485 53.475 194.735 ;
        RECT 53.665 194.355 53.935 194.925 ;
        RECT 54.315 194.905 55.065 195.095 ;
        RECT 55.235 195.075 55.405 195.395 ;
        RECT 55.630 195.265 55.960 195.725 ;
        RECT 56.160 195.075 56.490 195.555 ;
        RECT 56.705 195.265 57.035 195.725 ;
        RECT 57.205 195.075 57.535 195.555 ;
        RECT 55.235 194.905 57.535 195.075 ;
        RECT 58.785 194.905 58.995 195.725 ;
        RECT 59.165 194.925 59.495 195.555 ;
        RECT 54.315 194.735 54.685 194.905 ;
        RECT 54.105 194.525 54.685 194.735 ;
        RECT 54.855 194.525 55.275 194.735 ;
        RECT 54.425 194.355 54.685 194.525 ;
        RECT 49.965 193.175 50.295 193.935 ;
        RECT 50.475 193.345 50.655 194.105 ;
        RECT 50.905 193.175 52.115 194.265 ;
        RECT 52.345 193.175 52.555 194.315 ;
        RECT 52.725 193.345 53.055 194.325 ;
        RECT 53.225 193.175 53.455 194.315 ;
        RECT 53.665 193.345 54.190 194.355 ;
        RECT 54.425 194.065 55.175 194.355 ;
        RECT 54.425 193.175 54.755 193.895 ;
        RECT 54.925 193.345 55.175 194.065 ;
        RECT 55.445 193.420 55.775 194.735 ;
        RECT 55.985 193.420 56.315 194.735 ;
        RECT 56.485 193.420 56.855 194.735 ;
        RECT 57.065 194.485 57.575 194.735 ;
        RECT 59.165 194.325 59.415 194.925 ;
        RECT 59.665 194.905 59.895 195.725 ;
        RECT 60.195 195.175 60.365 195.555 ;
        RECT 60.545 195.345 60.875 195.725 ;
        RECT 60.195 195.005 60.860 195.175 ;
        RECT 61.055 195.050 61.315 195.555 ;
        RECT 59.585 194.485 59.915 194.735 ;
        RECT 60.125 194.455 60.465 194.825 ;
        RECT 60.690 194.750 60.860 195.005 ;
        RECT 60.690 194.420 60.965 194.750 ;
        RECT 57.185 193.175 57.515 194.295 ;
        RECT 58.785 193.175 58.995 194.315 ;
        RECT 59.165 193.345 59.495 194.325 ;
        RECT 59.665 193.175 59.895 194.315 ;
        RECT 60.690 194.275 60.860 194.420 ;
        RECT 60.185 194.105 60.860 194.275 ;
        RECT 61.135 194.250 61.315 195.050 ;
        RECT 61.945 195.000 62.235 195.725 ;
        RECT 62.490 195.175 62.665 195.465 ;
        RECT 62.835 195.345 63.165 195.725 ;
        RECT 62.490 195.005 62.985 195.175 ;
        RECT 63.340 195.045 63.555 195.415 ;
        RECT 63.790 195.275 64.390 195.445 ;
        RECT 60.185 193.345 60.365 194.105 ;
        RECT 60.545 193.175 60.875 193.935 ;
        RECT 61.045 193.345 61.315 194.250 ;
        RECT 61.945 193.175 62.235 194.340 ;
        RECT 62.465 194.065 62.645 194.835 ;
        RECT 62.815 194.025 62.985 195.005 ;
        RECT 63.155 194.715 63.555 195.045 ;
        RECT 63.725 194.775 64.050 195.105 ;
        RECT 63.540 194.365 63.710 194.525 ;
        RECT 63.325 194.195 63.710 194.365 ;
        RECT 63.880 194.235 64.050 194.775 ;
        RECT 64.220 194.575 64.390 195.275 ;
        RECT 64.770 195.265 65.100 195.725 ;
        RECT 65.305 195.345 65.735 195.515 ;
        RECT 64.560 194.795 64.935 195.095 ;
        RECT 64.220 194.405 64.560 194.575 ;
        RECT 64.730 194.490 64.935 194.795 ;
        RECT 65.105 194.490 65.395 195.095 ;
        RECT 65.565 194.750 65.735 195.345 ;
        RECT 65.905 195.135 66.140 195.465 ;
        RECT 63.880 194.025 64.220 194.235 ;
        RECT 62.815 193.895 64.220 194.025 ;
        RECT 62.495 193.855 64.220 193.895 ;
        RECT 62.495 193.725 62.985 193.855 ;
        RECT 62.495 193.435 62.665 193.725 ;
        RECT 64.390 193.685 64.560 194.405 ;
        RECT 65.565 194.420 65.800 194.750 ;
        RECT 65.565 194.320 65.735 194.420 ;
        RECT 65.465 194.150 65.735 194.320 ;
        RECT 65.465 194.025 65.635 194.150 ;
        RECT 65.290 193.855 65.635 194.025 ;
        RECT 65.970 194.000 66.140 195.135 ;
        RECT 62.835 193.175 63.165 193.555 ;
        RECT 63.730 193.515 64.560 193.685 ;
        RECT 64.915 193.175 65.145 193.755 ;
        RECT 65.885 193.685 66.140 194.000 ;
        RECT 65.625 193.515 66.140 193.685 ;
        RECT 66.310 193.685 66.500 195.465 ;
        RECT 66.715 195.225 66.920 195.555 ;
        RECT 67.115 195.265 67.445 195.725 ;
        RECT 67.645 195.345 68.540 195.515 ;
        RECT 66.715 194.245 66.885 195.225 ;
        RECT 67.065 194.415 67.435 195.095 ;
        RECT 67.645 194.245 67.815 195.345 ;
        RECT 66.715 194.075 67.815 194.245 ;
        RECT 66.715 193.915 66.905 194.075 ;
        RECT 66.310 193.515 66.835 193.685 ;
        RECT 67.075 193.175 67.420 193.805 ;
        RECT 67.645 193.655 67.815 194.075 ;
        RECT 67.985 194.775 68.605 195.105 ;
        RECT 68.855 194.815 69.165 195.435 ;
        RECT 69.335 194.995 69.585 195.725 ;
        RECT 69.755 195.085 70.085 195.545 ;
        RECT 67.985 193.825 68.275 194.775 ;
        RECT 68.855 194.735 69.265 194.815 ;
        RECT 68.445 194.165 68.785 194.565 ;
        RECT 68.955 194.485 69.265 194.735 ;
        RECT 69.435 194.485 69.745 194.815 ;
        RECT 69.435 194.315 69.605 194.485 ;
        RECT 69.915 194.315 70.085 195.085 ;
        RECT 70.255 194.925 70.510 195.725 ;
        RECT 70.685 194.955 72.355 195.725 ;
        RECT 72.985 195.075 73.245 195.555 ;
        RECT 73.415 195.265 73.745 195.725 ;
        RECT 73.935 195.085 74.135 195.505 ;
        RECT 70.685 194.435 71.435 194.955 ;
        RECT 68.995 194.145 69.605 194.315 ;
        RECT 68.995 193.685 69.165 194.145 ;
        RECT 69.775 193.975 70.085 194.315 ;
        RECT 67.645 193.485 68.595 193.655 ;
        RECT 68.845 193.515 69.165 193.685 ;
        RECT 69.335 193.175 69.505 193.975 ;
        RECT 69.675 193.355 70.085 193.975 ;
        RECT 70.255 193.175 70.505 194.315 ;
        RECT 71.605 194.265 72.355 194.785 ;
        RECT 70.685 193.175 72.355 194.265 ;
        RECT 72.985 194.045 73.155 195.075 ;
        RECT 73.325 194.385 73.555 194.815 ;
        RECT 73.725 194.565 74.135 195.085 ;
        RECT 74.305 195.240 75.095 195.505 ;
        RECT 74.305 194.385 74.560 195.240 ;
        RECT 75.275 194.905 75.605 195.325 ;
        RECT 75.775 194.905 76.035 195.725 ;
        RECT 76.215 194.995 76.515 195.725 ;
        RECT 75.275 194.815 75.525 194.905 ;
        RECT 76.695 194.815 76.925 195.435 ;
        RECT 77.125 195.165 77.350 195.545 ;
        RECT 77.520 195.335 77.850 195.725 ;
        RECT 77.125 194.985 77.455 195.165 ;
        RECT 74.730 194.565 75.525 194.815 ;
        RECT 73.325 194.215 75.115 194.385 ;
        RECT 72.985 193.345 73.260 194.045 ;
        RECT 73.430 193.920 74.145 194.215 ;
        RECT 74.365 193.855 74.695 194.045 ;
        RECT 73.470 193.175 73.685 193.720 ;
        RECT 73.855 193.345 74.330 193.685 ;
        RECT 74.500 193.680 74.695 193.855 ;
        RECT 74.865 193.850 75.115 194.215 ;
        RECT 74.500 193.175 75.115 193.680 ;
        RECT 75.355 193.345 75.525 194.565 ;
        RECT 75.695 193.855 76.035 194.735 ;
        RECT 76.220 194.485 76.515 194.815 ;
        RECT 76.695 194.485 77.110 194.815 ;
        RECT 77.280 194.315 77.455 194.985 ;
        RECT 77.625 194.485 77.865 195.135 ;
        RECT 78.045 194.955 79.715 195.725 ;
        RECT 79.885 195.050 80.145 195.555 ;
        RECT 80.325 195.345 80.655 195.725 ;
        RECT 80.835 195.175 81.005 195.555 ;
        RECT 78.045 194.435 78.795 194.955 ;
        RECT 76.215 193.955 77.110 194.285 ;
        RECT 77.280 194.125 77.865 194.315 ;
        RECT 78.965 194.265 79.715 194.785 ;
        RECT 76.215 193.785 77.420 193.955 ;
        RECT 75.775 193.175 76.035 193.685 ;
        RECT 76.215 193.355 76.545 193.785 ;
        RECT 76.725 193.175 76.920 193.615 ;
        RECT 77.090 193.355 77.420 193.785 ;
        RECT 77.590 193.355 77.865 194.125 ;
        RECT 78.045 193.175 79.715 194.265 ;
        RECT 79.885 194.250 80.065 195.050 ;
        RECT 80.340 195.005 81.005 195.175 ;
        RECT 80.340 194.750 80.510 195.005 ;
        RECT 81.265 194.955 84.775 195.725 ;
        RECT 85.495 195.175 85.665 195.555 ;
        RECT 85.845 195.345 86.175 195.725 ;
        RECT 85.495 195.005 86.160 195.175 ;
        RECT 86.355 195.050 86.615 195.555 ;
        RECT 80.235 194.420 80.510 194.750 ;
        RECT 80.735 194.455 81.075 194.825 ;
        RECT 81.265 194.435 82.915 194.955 ;
        RECT 80.340 194.275 80.510 194.420 ;
        RECT 79.885 193.345 80.155 194.250 ;
        RECT 80.340 194.105 81.015 194.275 ;
        RECT 83.085 194.265 84.775 194.785 ;
        RECT 85.425 194.455 85.765 194.825 ;
        RECT 85.990 194.750 86.160 195.005 ;
        RECT 85.990 194.420 86.265 194.750 ;
        RECT 85.990 194.275 86.160 194.420 ;
        RECT 80.325 193.175 80.655 193.935 ;
        RECT 80.835 193.345 81.015 194.105 ;
        RECT 81.265 193.175 84.775 194.265 ;
        RECT 85.485 194.105 86.160 194.275 ;
        RECT 86.435 194.250 86.615 195.050 ;
        RECT 87.705 195.000 87.995 195.725 ;
        RECT 88.625 194.780 88.965 195.555 ;
        RECT 89.135 195.265 89.305 195.725 ;
        RECT 89.545 195.290 89.905 195.555 ;
        RECT 89.545 195.285 89.900 195.290 ;
        RECT 89.545 195.275 89.895 195.285 ;
        RECT 89.545 195.270 89.890 195.275 ;
        RECT 89.545 195.260 89.885 195.270 ;
        RECT 90.535 195.265 90.705 195.725 ;
        RECT 89.545 195.255 89.880 195.260 ;
        RECT 89.545 195.245 89.870 195.255 ;
        RECT 89.545 195.235 89.860 195.245 ;
        RECT 89.545 195.095 89.845 195.235 ;
        RECT 89.135 194.905 89.845 195.095 ;
        RECT 90.035 195.095 90.365 195.175 ;
        RECT 90.875 195.095 91.215 195.555 ;
        RECT 90.035 194.905 91.215 195.095 ;
        RECT 91.385 195.155 91.820 195.555 ;
        RECT 91.990 195.325 92.375 195.725 ;
        RECT 91.385 194.985 92.375 195.155 ;
        RECT 92.545 194.985 92.970 195.555 ;
        RECT 93.160 195.155 93.415 195.555 ;
        RECT 93.585 195.325 93.970 195.725 ;
        RECT 93.160 194.985 93.970 195.155 ;
        RECT 94.140 194.985 94.385 195.555 ;
        RECT 94.575 195.155 94.830 195.555 ;
        RECT 95.000 195.325 95.385 195.725 ;
        RECT 94.575 194.985 95.385 195.155 ;
        RECT 95.555 194.985 95.815 195.555 ;
        RECT 85.485 193.345 85.665 194.105 ;
        RECT 85.845 193.175 86.175 193.935 ;
        RECT 86.345 193.345 86.615 194.250 ;
        RECT 87.705 193.175 87.995 194.340 ;
        RECT 88.625 193.345 88.905 194.780 ;
        RECT 89.135 194.335 89.420 194.905 ;
        RECT 92.040 194.815 92.375 194.985 ;
        RECT 92.620 194.815 92.970 194.985 ;
        RECT 93.620 194.815 93.970 194.985 ;
        RECT 94.215 194.815 94.385 194.985 ;
        RECT 95.035 194.815 95.385 194.985 ;
        RECT 89.605 194.505 90.075 194.735 ;
        RECT 90.245 194.715 90.575 194.735 ;
        RECT 90.245 194.535 90.695 194.715 ;
        RECT 90.885 194.535 91.215 194.735 ;
        RECT 89.135 194.120 90.285 194.335 ;
        RECT 89.075 193.175 89.785 193.950 ;
        RECT 89.955 193.345 90.285 194.120 ;
        RECT 90.480 193.420 90.695 194.535 ;
        RECT 90.985 194.195 91.215 194.535 ;
        RECT 91.385 194.110 91.870 194.815 ;
        RECT 92.040 194.485 92.450 194.815 ;
        RECT 92.040 193.940 92.375 194.485 ;
        RECT 92.620 194.315 93.450 194.815 ;
        RECT 90.875 193.175 91.205 193.895 ;
        RECT 91.385 193.770 92.375 193.940 ;
        RECT 92.545 194.135 93.450 194.315 ;
        RECT 93.620 194.485 94.045 194.815 ;
        RECT 91.385 193.345 91.820 193.770 ;
        RECT 91.990 193.175 92.375 193.600 ;
        RECT 92.545 193.345 92.970 194.135 ;
        RECT 93.620 193.965 93.970 194.485 ;
        RECT 94.215 194.315 94.865 194.815 ;
        RECT 93.140 193.770 93.970 193.965 ;
        RECT 94.140 194.135 94.865 194.315 ;
        RECT 95.035 194.485 95.460 194.815 ;
        RECT 93.140 193.345 93.415 193.770 ;
        RECT 93.585 193.175 93.970 193.600 ;
        RECT 94.140 193.345 94.385 194.135 ;
        RECT 95.035 193.965 95.385 194.485 ;
        RECT 95.630 194.315 95.815 194.985 ;
        RECT 95.985 194.955 98.575 195.725 ;
        RECT 98.745 195.155 99.180 195.555 ;
        RECT 99.350 195.325 99.735 195.725 ;
        RECT 98.745 194.985 99.735 195.155 ;
        RECT 99.905 194.985 100.330 195.555 ;
        RECT 100.520 195.155 100.775 195.555 ;
        RECT 100.945 195.325 101.330 195.725 ;
        RECT 100.520 194.985 101.330 195.155 ;
        RECT 101.500 194.985 101.745 195.555 ;
        RECT 101.935 195.155 102.190 195.555 ;
        RECT 102.360 195.325 102.745 195.725 ;
        RECT 101.935 194.985 102.745 195.155 ;
        RECT 102.915 194.985 103.175 195.555 ;
        RECT 95.985 194.435 97.195 194.955 ;
        RECT 99.400 194.815 99.735 194.985 ;
        RECT 99.980 194.815 100.330 194.985 ;
        RECT 100.980 194.815 101.330 194.985 ;
        RECT 101.575 194.815 101.745 194.985 ;
        RECT 102.395 194.815 102.745 194.985 ;
        RECT 94.575 193.770 95.385 193.965 ;
        RECT 94.575 193.345 94.830 193.770 ;
        RECT 95.000 193.175 95.385 193.600 ;
        RECT 95.555 193.345 95.815 194.315 ;
        RECT 97.365 194.265 98.575 194.785 ;
        RECT 95.985 193.175 98.575 194.265 ;
        RECT 98.745 194.110 99.230 194.815 ;
        RECT 99.400 194.485 99.810 194.815 ;
        RECT 99.400 193.940 99.735 194.485 ;
        RECT 99.980 194.315 100.810 194.815 ;
        RECT 98.745 193.770 99.735 193.940 ;
        RECT 99.905 194.135 100.810 194.315 ;
        RECT 100.980 194.485 101.405 194.815 ;
        RECT 98.745 193.345 99.180 193.770 ;
        RECT 99.350 193.175 99.735 193.600 ;
        RECT 99.905 193.345 100.330 194.135 ;
        RECT 100.980 193.965 101.330 194.485 ;
        RECT 101.575 194.315 102.225 194.815 ;
        RECT 100.500 193.770 101.330 193.965 ;
        RECT 101.500 194.135 102.225 194.315 ;
        RECT 102.395 194.485 102.820 194.815 ;
        RECT 100.500 193.345 100.775 193.770 ;
        RECT 100.945 193.175 101.330 193.600 ;
        RECT 101.500 193.345 101.745 194.135 ;
        RECT 102.395 193.965 102.745 194.485 ;
        RECT 102.990 194.315 103.175 194.985 ;
        RECT 103.365 194.915 103.605 195.725 ;
        RECT 103.775 194.915 104.105 195.555 ;
        RECT 104.275 194.915 104.545 195.725 ;
        RECT 104.725 195.050 104.985 195.555 ;
        RECT 105.165 195.345 105.495 195.725 ;
        RECT 105.675 195.175 105.845 195.555 ;
        RECT 103.345 194.485 103.695 194.735 ;
        RECT 103.865 194.315 104.035 194.915 ;
        RECT 104.205 194.485 104.555 194.735 ;
        RECT 101.935 193.770 102.745 193.965 ;
        RECT 101.935 193.345 102.190 193.770 ;
        RECT 102.360 193.175 102.745 193.600 ;
        RECT 102.915 193.345 103.175 194.315 ;
        RECT 103.355 194.145 104.035 194.315 ;
        RECT 103.355 193.360 103.685 194.145 ;
        RECT 104.215 193.175 104.545 194.315 ;
        RECT 104.725 194.250 104.905 195.050 ;
        RECT 105.180 195.005 105.845 195.175 ;
        RECT 105.180 194.750 105.350 195.005 ;
        RECT 106.105 194.985 106.365 195.555 ;
        RECT 106.535 195.325 106.920 195.725 ;
        RECT 107.090 195.155 107.345 195.555 ;
        RECT 106.535 194.985 107.345 195.155 ;
        RECT 107.535 194.985 107.780 195.555 ;
        RECT 107.950 195.325 108.335 195.725 ;
        RECT 108.505 195.155 108.760 195.555 ;
        RECT 107.950 194.985 108.760 195.155 ;
        RECT 108.950 194.985 109.375 195.555 ;
        RECT 109.545 195.325 109.930 195.725 ;
        RECT 110.100 195.155 110.535 195.555 ;
        RECT 109.545 194.985 110.535 195.155 ;
        RECT 110.740 194.985 111.355 195.555 ;
        RECT 111.525 195.215 111.740 195.725 ;
        RECT 111.970 195.215 112.250 195.545 ;
        RECT 112.430 195.215 112.670 195.725 ;
        RECT 105.075 194.420 105.350 194.750 ;
        RECT 105.575 194.455 105.915 194.825 ;
        RECT 105.180 194.275 105.350 194.420 ;
        RECT 106.105 194.315 106.290 194.985 ;
        RECT 106.535 194.815 106.885 194.985 ;
        RECT 107.535 194.815 107.705 194.985 ;
        RECT 107.950 194.815 108.300 194.985 ;
        RECT 108.950 194.815 109.300 194.985 ;
        RECT 109.545 194.815 109.880 194.985 ;
        RECT 106.460 194.485 106.885 194.815 ;
        RECT 104.725 193.345 104.995 194.250 ;
        RECT 105.180 194.105 105.855 194.275 ;
        RECT 105.165 193.175 105.495 193.935 ;
        RECT 105.675 193.345 105.855 194.105 ;
        RECT 106.105 193.345 106.365 194.315 ;
        RECT 106.535 193.965 106.885 194.485 ;
        RECT 107.055 194.315 107.705 194.815 ;
        RECT 107.875 194.485 108.300 194.815 ;
        RECT 107.055 194.135 107.780 194.315 ;
        RECT 106.535 193.770 107.345 193.965 ;
        RECT 106.535 193.175 106.920 193.600 ;
        RECT 107.090 193.345 107.345 193.770 ;
        RECT 107.535 193.345 107.780 194.135 ;
        RECT 107.950 193.965 108.300 194.485 ;
        RECT 108.470 194.315 109.300 194.815 ;
        RECT 109.470 194.485 109.880 194.815 ;
        RECT 108.470 194.135 109.375 194.315 ;
        RECT 107.950 193.770 108.780 193.965 ;
        RECT 107.950 193.175 108.335 193.600 ;
        RECT 108.505 193.345 108.780 193.770 ;
        RECT 108.950 193.345 109.375 194.135 ;
        RECT 109.545 193.940 109.880 194.485 ;
        RECT 110.050 194.110 110.535 194.815 ;
        RECT 110.740 193.965 111.055 194.985 ;
        RECT 111.225 194.315 111.395 194.815 ;
        RECT 111.645 194.485 111.910 195.045 ;
        RECT 112.080 194.315 112.250 195.215 ;
        RECT 112.420 194.485 112.775 195.045 ;
        RECT 113.465 195.000 113.755 195.725 ;
        RECT 113.965 194.905 114.195 195.725 ;
        RECT 114.365 194.925 114.695 195.555 ;
        RECT 113.945 194.485 114.275 194.735 ;
        RECT 111.225 194.145 112.650 194.315 ;
        RECT 109.545 193.770 110.535 193.940 ;
        RECT 109.545 193.175 109.930 193.600 ;
        RECT 110.100 193.345 110.535 193.770 ;
        RECT 110.740 193.345 111.275 193.965 ;
        RECT 111.445 193.175 111.775 193.975 ;
        RECT 112.260 193.970 112.650 194.145 ;
        RECT 113.465 193.175 113.755 194.340 ;
        RECT 114.445 194.325 114.695 194.925 ;
        RECT 114.865 194.905 115.075 195.725 ;
        RECT 115.305 194.955 116.975 195.725 ;
        RECT 117.145 194.985 117.405 195.555 ;
        RECT 117.575 195.325 117.960 195.725 ;
        RECT 118.130 195.155 118.385 195.555 ;
        RECT 117.575 194.985 118.385 195.155 ;
        RECT 118.575 194.985 118.820 195.555 ;
        RECT 118.990 195.325 119.375 195.725 ;
        RECT 119.545 195.155 119.800 195.555 ;
        RECT 118.990 194.985 119.800 195.155 ;
        RECT 119.990 194.985 120.415 195.555 ;
        RECT 120.585 195.325 120.970 195.725 ;
        RECT 121.140 195.155 121.575 195.555 ;
        RECT 122.535 195.325 122.865 195.725 ;
        RECT 123.035 195.155 123.365 195.495 ;
        RECT 124.415 195.325 124.745 195.725 ;
        RECT 120.585 194.985 121.575 195.155 ;
        RECT 122.380 194.985 124.745 195.155 ;
        RECT 124.915 195.000 125.245 195.510 ;
        RECT 115.305 194.435 116.055 194.955 ;
        RECT 113.965 193.175 114.195 194.315 ;
        RECT 114.365 193.345 114.695 194.325 ;
        RECT 114.865 193.175 115.075 194.315 ;
        RECT 116.225 194.265 116.975 194.785 ;
        RECT 115.305 193.175 116.975 194.265 ;
        RECT 117.145 194.315 117.330 194.985 ;
        RECT 117.575 194.815 117.925 194.985 ;
        RECT 118.575 194.815 118.745 194.985 ;
        RECT 118.990 194.815 119.340 194.985 ;
        RECT 119.990 194.815 120.340 194.985 ;
        RECT 120.585 194.815 120.920 194.985 ;
        RECT 117.500 194.485 117.925 194.815 ;
        RECT 117.145 193.345 117.405 194.315 ;
        RECT 117.575 193.965 117.925 194.485 ;
        RECT 118.095 194.315 118.745 194.815 ;
        RECT 118.915 194.485 119.340 194.815 ;
        RECT 118.095 194.135 118.820 194.315 ;
        RECT 117.575 193.770 118.385 193.965 ;
        RECT 117.575 193.175 117.960 193.600 ;
        RECT 118.130 193.345 118.385 193.770 ;
        RECT 118.575 193.345 118.820 194.135 ;
        RECT 118.990 193.965 119.340 194.485 ;
        RECT 119.510 194.315 120.340 194.815 ;
        RECT 120.510 194.485 120.920 194.815 ;
        RECT 119.510 194.135 120.415 194.315 ;
        RECT 118.990 193.770 119.820 193.965 ;
        RECT 118.990 193.175 119.375 193.600 ;
        RECT 119.545 193.345 119.820 193.770 ;
        RECT 119.990 193.345 120.415 194.135 ;
        RECT 120.585 193.940 120.920 194.485 ;
        RECT 121.090 194.110 121.575 194.815 ;
        RECT 122.380 193.985 122.550 194.985 ;
        RECT 124.575 194.815 124.745 194.985 ;
        RECT 122.720 194.155 122.965 194.815 ;
        RECT 123.180 194.155 123.445 194.815 ;
        RECT 123.640 194.155 123.925 194.815 ;
        RECT 124.100 194.485 124.405 194.815 ;
        RECT 124.575 194.485 124.885 194.815 ;
        RECT 124.100 194.155 124.315 194.485 ;
        RECT 125.055 194.365 125.245 195.000 ;
        RECT 125.445 194.995 125.735 195.725 ;
        RECT 125.435 194.485 125.735 194.815 ;
        RECT 125.915 194.795 126.145 195.435 ;
        RECT 126.325 195.175 126.635 195.545 ;
        RECT 126.815 195.355 127.485 195.725 ;
        RECT 126.325 194.975 127.555 195.175 ;
        RECT 125.915 194.485 126.440 194.795 ;
        RECT 126.620 194.485 127.085 194.795 ;
        RECT 120.585 193.770 121.575 193.940 ;
        RECT 122.380 193.815 122.835 193.985 ;
        RECT 120.585 193.175 120.970 193.600 ;
        RECT 121.140 193.345 121.575 193.770 ;
        RECT 122.505 193.385 122.835 193.815 ;
        RECT 123.015 193.815 124.305 193.985 ;
        RECT 123.015 193.395 123.265 193.815 ;
        RECT 123.495 193.175 123.825 193.645 ;
        RECT 124.055 193.395 124.305 193.815 ;
        RECT 124.495 193.175 124.745 194.315 ;
        RECT 125.025 194.235 125.245 194.365 ;
        RECT 127.265 194.305 127.555 194.975 ;
        RECT 124.915 193.385 125.245 194.235 ;
        RECT 125.445 194.065 126.605 194.305 ;
        RECT 125.445 193.355 125.705 194.065 ;
        RECT 125.875 193.175 126.205 193.885 ;
        RECT 126.375 193.355 126.605 194.065 ;
        RECT 126.785 194.085 127.555 194.305 ;
        RECT 126.785 193.355 127.055 194.085 ;
        RECT 127.235 193.175 127.575 193.905 ;
        RECT 127.745 193.355 128.005 195.545 ;
        RECT 128.185 194.955 131.695 195.725 ;
        RECT 128.185 194.435 129.835 194.955 ;
        RECT 133.060 194.915 133.305 195.520 ;
        RECT 133.525 195.190 134.035 195.725 ;
        RECT 130.005 194.265 131.695 194.785 ;
        RECT 128.185 193.175 131.695 194.265 ;
        RECT 132.785 194.745 134.015 194.915 ;
        RECT 132.785 193.935 133.125 194.745 ;
        RECT 133.295 194.180 134.045 194.370 ;
        RECT 132.785 193.525 133.300 193.935 ;
        RECT 133.535 193.175 133.705 193.935 ;
        RECT 133.875 193.515 134.045 194.180 ;
        RECT 134.215 194.195 134.405 195.555 ;
        RECT 134.575 195.385 134.850 195.555 ;
        RECT 134.575 195.215 134.855 195.385 ;
        RECT 134.575 194.395 134.850 195.215 ;
        RECT 135.040 195.190 135.570 195.555 ;
        RECT 135.995 195.325 136.325 195.725 ;
        RECT 135.395 195.155 135.570 195.190 ;
        RECT 135.055 194.195 135.225 194.995 ;
        RECT 134.215 194.025 135.225 194.195 ;
        RECT 135.395 194.985 136.325 195.155 ;
        RECT 136.495 194.985 136.750 195.555 ;
        RECT 135.395 193.855 135.565 194.985 ;
        RECT 136.155 194.815 136.325 194.985 ;
        RECT 134.440 193.685 135.565 193.855 ;
        RECT 135.735 194.485 135.930 194.815 ;
        RECT 136.155 194.485 136.410 194.815 ;
        RECT 135.735 193.515 135.905 194.485 ;
        RECT 136.580 194.315 136.750 194.985 ;
        RECT 137.125 195.095 137.455 195.455 ;
        RECT 138.075 195.265 138.325 195.725 ;
        RECT 138.495 195.265 139.055 195.555 ;
        RECT 137.125 194.905 138.515 195.095 ;
        RECT 138.345 194.815 138.515 194.905 ;
        RECT 133.875 193.345 135.905 193.515 ;
        RECT 136.075 193.175 136.245 194.315 ;
        RECT 136.415 193.345 136.750 194.315 ;
        RECT 136.940 194.485 137.615 194.735 ;
        RECT 137.835 194.485 138.175 194.735 ;
        RECT 138.345 194.485 138.635 194.815 ;
        RECT 136.940 194.125 137.205 194.485 ;
        RECT 138.345 194.235 138.515 194.485 ;
        RECT 137.575 194.065 138.515 194.235 ;
        RECT 137.125 193.175 137.405 193.845 ;
        RECT 137.575 193.515 137.875 194.065 ;
        RECT 138.805 193.895 139.055 195.265 ;
        RECT 139.225 195.000 139.515 195.725 ;
        RECT 139.775 195.175 139.945 195.465 ;
        RECT 140.115 195.345 140.445 195.725 ;
        RECT 139.775 195.005 140.440 195.175 ;
        RECT 138.075 193.175 138.405 193.895 ;
        RECT 138.595 193.345 139.055 193.895 ;
        RECT 139.225 193.175 139.515 194.340 ;
        RECT 139.690 194.185 140.040 194.835 ;
        RECT 140.210 194.015 140.440 195.005 ;
        RECT 139.775 193.845 140.440 194.015 ;
        RECT 139.775 193.345 139.945 193.845 ;
        RECT 140.115 193.175 140.445 193.675 ;
        RECT 140.615 193.345 140.800 195.465 ;
        RECT 141.055 195.265 141.305 195.725 ;
        RECT 141.475 195.275 141.810 195.445 ;
        RECT 142.005 195.275 142.680 195.445 ;
        RECT 141.475 195.135 141.645 195.275 ;
        RECT 140.970 194.145 141.250 195.095 ;
        RECT 141.420 195.005 141.645 195.135 ;
        RECT 141.420 193.900 141.590 195.005 ;
        RECT 141.815 194.855 142.340 195.075 ;
        RECT 141.760 194.090 142.000 194.685 ;
        RECT 142.170 194.155 142.340 194.855 ;
        RECT 142.510 194.495 142.680 195.275 ;
        RECT 143.000 195.225 143.370 195.725 ;
        RECT 143.550 195.275 143.955 195.445 ;
        RECT 144.125 195.275 144.910 195.445 ;
        RECT 143.550 195.045 143.720 195.275 ;
        RECT 142.890 194.745 143.720 195.045 ;
        RECT 144.105 194.775 144.570 195.105 ;
        RECT 142.890 194.715 143.090 194.745 ;
        RECT 143.210 194.495 143.380 194.565 ;
        RECT 142.510 194.325 143.380 194.495 ;
        RECT 142.870 194.235 143.380 194.325 ;
        RECT 141.420 193.770 141.725 193.900 ;
        RECT 142.170 193.790 142.700 194.155 ;
        RECT 141.040 193.175 141.305 193.635 ;
        RECT 141.475 193.345 141.725 193.770 ;
        RECT 142.870 193.620 143.040 194.235 ;
        RECT 141.935 193.450 143.040 193.620 ;
        RECT 143.210 193.175 143.380 193.975 ;
        RECT 143.550 193.675 143.720 194.745 ;
        RECT 143.890 193.845 144.080 194.565 ;
        RECT 144.250 193.815 144.570 194.775 ;
        RECT 144.740 194.815 144.910 195.275 ;
        RECT 145.185 195.195 145.395 195.725 ;
        RECT 145.655 194.985 145.985 195.510 ;
        RECT 146.155 195.115 146.325 195.725 ;
        RECT 146.495 195.070 146.825 195.505 ;
        RECT 146.495 194.985 146.875 195.070 ;
        RECT 145.785 194.815 145.985 194.985 ;
        RECT 146.650 194.945 146.875 194.985 ;
        RECT 144.740 194.485 145.615 194.815 ;
        RECT 145.785 194.485 146.535 194.815 ;
        RECT 143.550 193.345 143.800 193.675 ;
        RECT 144.740 193.645 144.910 194.485 ;
        RECT 145.785 194.280 145.975 194.485 ;
        RECT 146.705 194.365 146.875 194.945 ;
        RECT 147.045 194.955 148.715 195.725 ;
        RECT 148.885 194.975 150.095 195.725 ;
        RECT 147.045 194.435 147.795 194.955 ;
        RECT 146.660 194.315 146.875 194.365 ;
        RECT 145.080 193.905 145.975 194.280 ;
        RECT 146.485 194.235 146.875 194.315 ;
        RECT 147.965 194.265 148.715 194.785 ;
        RECT 144.025 193.475 144.910 193.645 ;
        RECT 145.090 193.175 145.405 193.675 ;
        RECT 145.635 193.345 145.975 193.905 ;
        RECT 146.145 193.175 146.315 194.185 ;
        RECT 146.485 193.390 146.815 194.235 ;
        RECT 147.045 193.175 148.715 194.265 ;
        RECT 148.885 194.265 149.405 194.805 ;
        RECT 149.575 194.435 150.095 194.975 ;
        RECT 148.885 193.175 150.095 194.265 ;
        RECT 36.100 193.005 150.180 193.175 ;
        RECT 36.185 191.915 37.395 193.005 ;
        RECT 37.565 191.915 41.075 193.005 ;
        RECT 42.170 192.205 42.425 193.005 ;
        RECT 42.625 192.155 42.955 192.835 ;
        RECT 36.185 191.205 36.705 191.745 ;
        RECT 36.875 191.375 37.395 191.915 ;
        RECT 37.565 191.225 39.215 191.745 ;
        RECT 39.385 191.395 41.075 191.915 ;
        RECT 42.170 191.665 42.415 192.025 ;
        RECT 42.605 191.875 42.955 192.155 ;
        RECT 42.605 191.495 42.775 191.875 ;
        RECT 43.135 191.695 43.330 192.745 ;
        RECT 43.510 191.865 43.830 193.005 ;
        RECT 44.005 191.915 47.515 193.005 ;
        RECT 47.685 191.915 48.895 193.005 ;
        RECT 42.255 191.325 42.775 191.495 ;
        RECT 42.945 191.365 43.330 191.695 ;
        RECT 43.510 191.645 43.770 191.695 ;
        RECT 43.510 191.475 43.775 191.645 ;
        RECT 43.510 191.365 43.770 191.475 ;
        RECT 36.185 190.455 37.395 191.205 ;
        RECT 37.565 190.455 41.075 191.225 ;
        RECT 42.255 190.760 42.425 191.325 ;
        RECT 44.005 191.225 45.655 191.745 ;
        RECT 45.825 191.395 47.515 191.915 ;
        RECT 42.615 190.985 43.830 191.155 ;
        RECT 42.615 190.680 42.845 190.985 ;
        RECT 43.015 190.455 43.345 190.815 ;
        RECT 43.540 190.635 43.830 190.985 ;
        RECT 44.005 190.455 47.515 191.225 ;
        RECT 47.685 191.205 48.205 191.745 ;
        RECT 48.375 191.375 48.895 191.915 ;
        RECT 49.065 191.840 49.355 193.005 ;
        RECT 49.525 191.915 51.195 193.005 ;
        RECT 49.525 191.225 50.275 191.745 ;
        RECT 50.445 191.395 51.195 191.915 ;
        RECT 51.920 191.810 52.090 193.005 ;
        RECT 52.260 191.865 52.535 192.835 ;
        RECT 52.745 192.205 53.025 193.005 ;
        RECT 53.195 192.495 53.835 192.825 ;
        RECT 54.060 192.575 54.805 192.745 ;
        RECT 55.495 192.575 55.825 193.005 ;
        RECT 54.060 192.325 54.230 192.575 ;
        RECT 55.995 192.405 56.255 192.825 ;
        RECT 53.195 192.155 54.230 192.325 ;
        RECT 54.400 192.235 56.255 192.405 ;
        RECT 53.195 192.035 53.365 192.155 ;
        RECT 52.705 191.865 53.365 192.035 ;
        RECT 54.400 191.955 54.570 192.235 ;
        RECT 47.685 190.455 48.895 191.205 ;
        RECT 49.065 190.455 49.355 191.180 ;
        RECT 49.525 190.455 51.195 191.225 ;
        RECT 51.920 190.455 52.090 191.395 ;
        RECT 52.260 191.130 52.430 191.865 ;
        RECT 52.705 191.695 52.875 191.865 ;
        RECT 53.920 191.785 54.570 191.955 ;
        RECT 54.740 191.895 55.345 192.065 ;
        RECT 52.600 191.365 52.875 191.695 ;
        RECT 53.045 191.365 53.700 191.695 ;
        RECT 53.920 191.365 54.090 191.785 ;
        RECT 54.740 191.615 54.930 191.895 ;
        RECT 54.485 191.445 54.930 191.615 ;
        RECT 52.705 191.195 52.875 191.365 ;
        RECT 54.740 191.195 54.930 191.445 ;
        RECT 55.100 191.365 55.390 191.695 ;
        RECT 55.560 191.365 55.910 192.065 ;
        RECT 56.080 191.195 56.255 192.235 ;
        RECT 52.260 190.785 52.535 191.130 ;
        RECT 52.705 191.025 54.315 191.195 ;
        RECT 54.740 191.025 55.260 191.195 ;
        RECT 52.725 190.455 53.105 190.855 ;
        RECT 53.275 190.675 53.445 191.025 ;
        RECT 53.615 190.455 53.945 190.855 ;
        RECT 54.145 190.675 54.315 191.025 ;
        RECT 54.490 190.455 54.845 190.855 ;
        RECT 55.090 190.820 55.260 191.025 ;
        RECT 55.510 190.455 55.680 191.195 ;
        RECT 55.935 190.820 56.255 191.195 ;
        RECT 56.425 192.535 56.765 192.795 ;
        RECT 56.935 192.545 57.185 193.005 ;
        RECT 56.425 190.930 56.685 192.535 ;
        RECT 57.375 192.365 57.705 192.795 ;
        RECT 56.855 192.195 57.705 192.365 ;
        RECT 57.875 192.335 58.045 192.835 ;
        RECT 58.255 192.545 58.505 193.005 ;
        RECT 58.715 192.335 58.885 192.835 ;
        RECT 59.185 192.545 59.435 193.005 ;
        RECT 59.675 192.335 59.845 192.835 ;
        RECT 56.855 191.275 57.025 192.195 ;
        RECT 57.875 192.165 59.845 192.335 ;
        RECT 57.345 191.445 57.675 192.005 ;
        RECT 57.875 191.985 58.175 191.990 ;
        RECT 57.865 191.815 58.175 191.985 ;
        RECT 57.875 191.695 58.175 191.815 ;
        RECT 57.875 191.365 58.255 191.695 ;
        RECT 56.855 191.180 57.675 191.275 ;
        RECT 56.855 191.105 57.870 191.180 ;
        RECT 56.425 190.670 56.765 190.930 ;
        RECT 56.935 190.455 57.265 190.935 ;
        RECT 57.455 190.670 57.870 191.105 ;
        RECT 58.565 190.970 58.785 191.695 ;
        RECT 59.045 191.365 59.425 191.995 ;
        RECT 59.655 191.365 59.910 191.995 ;
        RECT 60.565 191.930 60.835 192.835 ;
        RECT 61.005 192.245 61.335 193.005 ;
        RECT 61.515 192.075 61.695 192.835 ;
        RECT 58.040 190.785 58.990 190.970 ;
        RECT 59.220 190.765 59.425 191.365 ;
        RECT 59.595 190.455 59.935 191.180 ;
        RECT 60.565 191.130 60.745 191.930 ;
        RECT 61.020 191.905 61.695 192.075 ;
        RECT 61.020 191.760 61.190 191.905 ;
        RECT 60.915 191.430 61.190 191.760 ;
        RECT 61.945 191.865 62.205 192.835 ;
        RECT 62.375 192.580 62.760 193.005 ;
        RECT 62.930 192.410 63.185 192.835 ;
        RECT 62.375 192.215 63.185 192.410 ;
        RECT 61.020 191.175 61.190 191.430 ;
        RECT 61.415 191.355 61.755 191.725 ;
        RECT 61.945 191.195 62.130 191.865 ;
        RECT 62.375 191.695 62.725 192.215 ;
        RECT 63.375 192.045 63.620 192.835 ;
        RECT 63.790 192.580 64.175 193.005 ;
        RECT 64.345 192.410 64.620 192.835 ;
        RECT 62.300 191.365 62.725 191.695 ;
        RECT 62.895 191.865 63.620 192.045 ;
        RECT 63.790 192.215 64.620 192.410 ;
        RECT 62.895 191.365 63.545 191.865 ;
        RECT 63.790 191.695 64.140 192.215 ;
        RECT 64.790 192.045 65.215 192.835 ;
        RECT 65.385 192.580 65.770 193.005 ;
        RECT 65.940 192.410 66.375 192.835 ;
        RECT 66.550 192.580 66.885 193.005 ;
        RECT 63.715 191.365 64.140 191.695 ;
        RECT 64.310 191.865 65.215 192.045 ;
        RECT 65.385 192.240 66.375 192.410 ;
        RECT 67.055 192.400 67.240 192.805 ;
        RECT 64.310 191.365 65.140 191.865 ;
        RECT 65.385 191.695 65.720 192.240 ;
        RECT 66.575 192.225 67.240 192.400 ;
        RECT 67.445 192.225 67.775 193.005 ;
        RECT 65.310 191.365 65.720 191.695 ;
        RECT 65.890 191.365 66.375 192.070 ;
        RECT 62.375 191.195 62.725 191.365 ;
        RECT 63.375 191.195 63.545 191.365 ;
        RECT 63.790 191.195 64.140 191.365 ;
        RECT 64.790 191.195 65.140 191.365 ;
        RECT 65.385 191.195 65.720 191.365 ;
        RECT 66.575 191.195 66.915 192.225 ;
        RECT 67.945 192.035 68.215 192.805 ;
        RECT 68.385 192.570 73.730 193.005 ;
        RECT 67.085 191.865 68.215 192.035 ;
        RECT 67.085 191.365 67.335 191.865 ;
        RECT 60.565 190.625 60.825 191.130 ;
        RECT 61.020 191.005 61.685 191.175 ;
        RECT 61.005 190.455 61.335 190.835 ;
        RECT 61.515 190.625 61.685 191.005 ;
        RECT 61.945 190.625 62.205 191.195 ;
        RECT 62.375 191.025 63.185 191.195 ;
        RECT 62.375 190.455 62.760 190.855 ;
        RECT 62.930 190.625 63.185 191.025 ;
        RECT 63.375 190.625 63.620 191.195 ;
        RECT 63.790 191.025 64.600 191.195 ;
        RECT 63.790 190.455 64.175 190.855 ;
        RECT 64.345 190.625 64.600 191.025 ;
        RECT 64.790 190.625 65.215 191.195 ;
        RECT 65.385 191.025 66.375 191.195 ;
        RECT 66.575 191.025 67.260 191.195 ;
        RECT 67.515 191.115 67.875 191.695 ;
        RECT 65.385 190.455 65.770 190.855 ;
        RECT 65.940 190.625 66.375 191.025 ;
        RECT 66.550 190.455 66.885 190.855 ;
        RECT 67.055 190.625 67.260 191.025 ;
        RECT 68.045 190.955 68.215 191.865 ;
        RECT 69.970 191.000 70.310 191.830 ;
        RECT 71.790 191.320 72.140 192.570 ;
        RECT 74.825 191.840 75.115 193.005 ;
        RECT 67.470 190.455 67.745 190.935 ;
        RECT 67.955 190.625 68.215 190.955 ;
        RECT 68.385 190.455 73.730 191.000 ;
        RECT 74.825 190.455 75.115 191.180 ;
        RECT 75.295 190.635 75.555 192.825 ;
        RECT 75.725 192.275 76.065 193.005 ;
        RECT 76.245 192.095 76.515 192.825 ;
        RECT 75.745 191.875 76.515 192.095 ;
        RECT 76.695 192.115 76.925 192.825 ;
        RECT 77.095 192.295 77.425 193.005 ;
        RECT 77.595 192.115 77.855 192.825 ;
        RECT 78.050 192.205 78.305 193.005 ;
        RECT 78.505 192.155 78.835 192.835 ;
        RECT 76.695 191.875 77.855 192.115 ;
        RECT 75.745 191.205 76.035 191.875 ;
        RECT 76.215 191.385 76.680 191.695 ;
        RECT 76.860 191.385 77.385 191.695 ;
        RECT 75.745 191.005 76.975 191.205 ;
        RECT 75.815 190.455 76.485 190.825 ;
        RECT 76.665 190.635 76.975 191.005 ;
        RECT 77.155 190.745 77.385 191.385 ;
        RECT 77.565 191.365 77.865 191.695 ;
        RECT 78.050 191.665 78.295 192.025 ;
        RECT 78.485 191.875 78.835 192.155 ;
        RECT 78.485 191.495 78.655 191.875 ;
        RECT 79.015 191.695 79.210 192.745 ;
        RECT 79.390 191.865 79.710 193.005 ;
        RECT 79.885 191.930 80.155 192.835 ;
        RECT 80.325 192.245 80.655 193.005 ;
        RECT 80.835 192.075 81.015 192.835 ;
        RECT 81.265 192.570 86.610 193.005 ;
        RECT 78.135 191.325 78.655 191.495 ;
        RECT 78.825 191.365 79.210 191.695 ;
        RECT 79.390 191.365 79.650 191.695 ;
        RECT 77.565 190.455 77.855 191.185 ;
        RECT 78.135 190.760 78.305 191.325 ;
        RECT 78.495 190.985 79.710 191.155 ;
        RECT 78.495 190.680 78.725 190.985 ;
        RECT 78.895 190.455 79.225 190.815 ;
        RECT 79.420 190.635 79.710 190.985 ;
        RECT 79.885 191.130 80.065 191.930 ;
        RECT 80.340 191.905 81.015 192.075 ;
        RECT 80.340 191.760 80.510 191.905 ;
        RECT 80.235 191.430 80.510 191.760 ;
        RECT 80.340 191.175 80.510 191.430 ;
        RECT 80.735 191.355 81.075 191.725 ;
        RECT 79.885 190.625 80.145 191.130 ;
        RECT 80.340 191.005 81.005 191.175 ;
        RECT 80.325 190.455 80.655 190.835 ;
        RECT 80.835 190.625 81.005 191.005 ;
        RECT 82.850 191.000 83.190 191.830 ;
        RECT 84.670 191.320 85.020 192.570 ;
        RECT 87.705 192.245 88.370 192.835 ;
        RECT 87.705 191.275 87.955 192.245 ;
        RECT 88.540 192.165 88.870 193.005 ;
        RECT 89.380 192.415 90.185 192.835 ;
        RECT 89.040 192.245 90.605 192.415 ;
        RECT 89.040 191.995 89.210 192.245 ;
        RECT 88.290 191.825 89.210 191.995 ;
        RECT 88.290 191.655 88.460 191.825 ;
        RECT 89.380 191.655 89.755 192.075 ;
        RECT 88.125 191.445 88.460 191.655 ;
        RECT 88.630 191.445 89.080 191.655 ;
        RECT 89.270 191.645 89.755 191.655 ;
        RECT 89.945 191.695 90.265 192.075 ;
        RECT 90.435 191.995 90.605 192.245 ;
        RECT 90.775 192.165 91.025 193.005 ;
        RECT 91.220 191.995 91.520 192.835 ;
        RECT 90.435 191.825 91.520 191.995 ;
        RECT 89.270 191.475 89.775 191.645 ;
        RECT 89.270 191.445 89.755 191.475 ;
        RECT 89.945 191.445 90.325 191.695 ;
        RECT 90.505 191.445 90.835 191.655 ;
        RECT 81.265 190.455 86.610 191.000 ;
        RECT 87.705 190.635 88.390 191.275 ;
        RECT 88.560 190.455 88.730 191.275 ;
        RECT 88.900 191.105 90.600 191.275 ;
        RECT 88.900 190.640 89.230 191.105 ;
        RECT 90.215 191.015 90.600 191.105 ;
        RECT 91.005 191.195 91.175 191.825 ;
        RECT 91.345 191.365 91.675 191.655 ;
        RECT 91.845 191.400 92.125 192.835 ;
        RECT 92.295 192.230 93.005 193.005 ;
        RECT 93.175 192.060 93.505 192.835 ;
        RECT 92.355 191.845 93.505 192.060 ;
        RECT 91.005 191.015 91.515 191.195 ;
        RECT 89.400 190.455 89.570 190.925 ;
        RECT 89.830 190.675 91.015 190.845 ;
        RECT 91.185 190.625 91.515 191.015 ;
        RECT 91.845 190.625 92.185 191.400 ;
        RECT 92.355 191.275 92.640 191.845 ;
        RECT 92.825 191.445 93.295 191.675 ;
        RECT 93.700 191.645 93.915 192.760 ;
        RECT 94.095 192.285 94.425 193.005 ;
        RECT 94.205 191.645 94.435 191.985 ;
        RECT 93.465 191.465 93.915 191.645 ;
        RECT 93.465 191.445 93.795 191.465 ;
        RECT 94.105 191.445 94.435 191.645 ;
        RECT 95.525 191.930 95.795 192.835 ;
        RECT 95.965 192.245 96.295 193.005 ;
        RECT 96.475 192.075 96.655 192.835 ;
        RECT 92.355 191.085 93.065 191.275 ;
        RECT 92.765 190.945 93.065 191.085 ;
        RECT 93.255 191.085 94.435 191.275 ;
        RECT 93.255 191.005 93.585 191.085 ;
        RECT 92.765 190.935 93.080 190.945 ;
        RECT 92.765 190.925 93.090 190.935 ;
        RECT 92.765 190.920 93.100 190.925 ;
        RECT 92.355 190.455 92.525 190.915 ;
        RECT 92.765 190.910 93.105 190.920 ;
        RECT 92.765 190.905 93.110 190.910 ;
        RECT 92.765 190.895 93.115 190.905 ;
        RECT 92.765 190.890 93.120 190.895 ;
        RECT 92.765 190.625 93.125 190.890 ;
        RECT 93.755 190.455 93.925 190.915 ;
        RECT 94.095 190.625 94.435 191.085 ;
        RECT 95.525 191.130 95.705 191.930 ;
        RECT 95.980 191.905 96.655 192.075 ;
        RECT 95.980 191.760 96.150 191.905 ;
        RECT 95.875 191.430 96.150 191.760 ;
        RECT 96.905 191.865 97.245 192.835 ;
        RECT 97.415 191.865 97.585 193.005 ;
        RECT 97.855 192.205 98.105 193.005 ;
        RECT 98.750 192.035 99.080 192.835 ;
        RECT 99.380 192.205 99.710 193.005 ;
        RECT 99.880 192.035 100.210 192.835 ;
        RECT 97.775 191.865 100.210 192.035 ;
        RECT 95.980 191.175 96.150 191.430 ;
        RECT 96.375 191.355 96.715 191.725 ;
        RECT 96.905 191.255 97.080 191.865 ;
        RECT 97.775 191.615 97.945 191.865 ;
        RECT 97.250 191.445 97.945 191.615 ;
        RECT 98.120 191.445 98.540 191.645 ;
        RECT 98.710 191.445 99.040 191.645 ;
        RECT 99.210 191.445 99.540 191.645 ;
        RECT 95.525 190.625 95.785 191.130 ;
        RECT 95.980 191.005 96.645 191.175 ;
        RECT 95.965 190.455 96.295 190.835 ;
        RECT 96.475 190.625 96.645 191.005 ;
        RECT 96.905 190.625 97.245 191.255 ;
        RECT 97.415 190.455 97.665 191.255 ;
        RECT 97.855 191.105 99.080 191.275 ;
        RECT 97.855 190.625 98.185 191.105 ;
        RECT 98.355 190.455 98.580 190.915 ;
        RECT 98.750 190.625 99.080 191.105 ;
        RECT 99.710 191.235 99.880 191.865 ;
        RECT 100.585 191.840 100.875 193.005 ;
        RECT 101.045 192.245 101.710 192.835 ;
        RECT 100.065 191.445 100.415 191.695 ;
        RECT 101.045 191.275 101.295 192.245 ;
        RECT 101.880 192.165 102.210 193.005 ;
        RECT 102.720 192.415 103.525 192.835 ;
        RECT 102.380 192.245 103.945 192.415 ;
        RECT 102.380 191.995 102.550 192.245 ;
        RECT 101.630 191.825 102.550 191.995 ;
        RECT 101.630 191.655 101.800 191.825 ;
        RECT 102.720 191.655 103.095 192.075 ;
        RECT 101.465 191.445 101.800 191.655 ;
        RECT 101.970 191.445 102.420 191.655 ;
        RECT 102.610 191.645 103.095 191.655 ;
        RECT 103.285 191.695 103.605 192.075 ;
        RECT 103.775 191.995 103.945 192.245 ;
        RECT 104.115 192.165 104.365 193.005 ;
        RECT 104.560 191.995 104.860 192.835 ;
        RECT 103.775 191.825 104.860 191.995 ;
        RECT 105.185 192.165 105.445 192.835 ;
        RECT 105.615 192.605 105.945 193.005 ;
        RECT 106.815 192.605 107.215 193.005 ;
        RECT 107.505 192.425 107.835 192.660 ;
        RECT 105.755 192.255 107.835 192.425 ;
        RECT 102.610 191.475 103.115 191.645 ;
        RECT 102.610 191.445 103.095 191.475 ;
        RECT 103.285 191.445 103.665 191.695 ;
        RECT 103.845 191.445 104.175 191.655 ;
        RECT 99.710 190.625 100.210 191.235 ;
        RECT 100.585 190.455 100.875 191.180 ;
        RECT 101.045 190.635 101.730 191.275 ;
        RECT 101.900 190.455 102.070 191.275 ;
        RECT 102.240 191.105 103.940 191.275 ;
        RECT 102.240 190.640 102.570 191.105 ;
        RECT 103.555 191.015 103.940 191.105 ;
        RECT 104.345 191.195 104.515 191.825 ;
        RECT 104.685 191.365 105.015 191.655 ;
        RECT 105.185 191.195 105.360 192.165 ;
        RECT 105.755 191.985 105.925 192.255 ;
        RECT 105.530 191.815 105.925 191.985 ;
        RECT 106.095 191.865 107.110 192.085 ;
        RECT 105.530 191.365 105.700 191.815 ;
        RECT 106.835 191.725 107.110 191.865 ;
        RECT 107.280 191.865 107.835 192.255 ;
        RECT 105.870 191.445 106.320 191.645 ;
        RECT 106.490 191.275 106.665 191.470 ;
        RECT 104.345 191.015 104.855 191.195 ;
        RECT 102.740 190.455 102.910 190.925 ;
        RECT 103.170 190.675 104.355 190.845 ;
        RECT 104.525 190.625 104.855 191.015 ;
        RECT 105.185 190.625 105.525 191.195 ;
        RECT 105.720 190.455 105.890 191.120 ;
        RECT 106.170 191.105 106.665 191.275 ;
        RECT 106.170 190.965 106.390 191.105 ;
        RECT 106.165 190.795 106.390 190.965 ;
        RECT 106.835 190.935 107.005 191.725 ;
        RECT 107.280 191.615 107.450 191.865 ;
        RECT 108.005 191.695 108.180 192.795 ;
        RECT 108.350 192.185 108.695 193.005 ;
        RECT 107.255 191.445 107.450 191.615 ;
        RECT 107.620 191.445 108.180 191.695 ;
        RECT 108.350 191.445 108.695 192.015 ;
        RECT 108.865 191.865 109.145 193.005 ;
        RECT 109.315 191.855 109.645 192.835 ;
        RECT 109.815 191.865 110.075 193.005 ;
        RECT 110.245 192.410 110.680 192.835 ;
        RECT 110.850 192.580 111.235 193.005 ;
        RECT 110.245 192.240 111.235 192.410 ;
        RECT 107.255 191.060 107.425 191.445 ;
        RECT 108.875 191.425 109.210 191.695 ;
        RECT 106.170 190.750 106.390 190.795 ;
        RECT 106.560 190.765 107.005 190.935 ;
        RECT 107.175 190.690 107.425 191.060 ;
        RECT 107.595 191.095 108.695 191.275 ;
        RECT 109.380 191.255 109.550 191.855 ;
        RECT 109.720 191.445 110.055 191.695 ;
        RECT 110.245 191.365 110.730 192.070 ;
        RECT 110.900 191.695 111.235 192.240 ;
        RECT 111.405 192.045 111.830 192.835 ;
        RECT 112.000 192.410 112.275 192.835 ;
        RECT 112.445 192.580 112.830 193.005 ;
        RECT 112.000 192.215 112.830 192.410 ;
        RECT 111.405 191.865 112.310 192.045 ;
        RECT 110.900 191.365 111.310 191.695 ;
        RECT 111.480 191.365 112.310 191.865 ;
        RECT 112.480 191.695 112.830 192.215 ;
        RECT 113.000 192.045 113.245 192.835 ;
        RECT 113.435 192.410 113.690 192.835 ;
        RECT 113.860 192.580 114.245 193.005 ;
        RECT 113.435 192.215 114.245 192.410 ;
        RECT 113.000 191.865 113.725 192.045 ;
        RECT 112.480 191.365 112.905 191.695 ;
        RECT 113.075 191.365 113.725 191.865 ;
        RECT 113.895 191.695 114.245 192.215 ;
        RECT 114.415 191.865 114.675 192.835 ;
        RECT 113.895 191.365 114.320 191.695 ;
        RECT 107.595 190.690 107.845 191.095 ;
        RECT 108.015 190.455 108.185 190.925 ;
        RECT 108.355 190.690 108.695 191.095 ;
        RECT 108.865 190.455 109.175 191.255 ;
        RECT 109.380 190.625 110.075 191.255 ;
        RECT 110.900 191.195 111.235 191.365 ;
        RECT 111.480 191.195 111.830 191.365 ;
        RECT 112.480 191.195 112.830 191.365 ;
        RECT 113.075 191.195 113.245 191.365 ;
        RECT 113.895 191.195 114.245 191.365 ;
        RECT 114.490 191.195 114.675 191.865 ;
        RECT 110.245 191.025 111.235 191.195 ;
        RECT 110.245 190.625 110.680 191.025 ;
        RECT 110.850 190.455 111.235 190.855 ;
        RECT 111.405 190.625 111.830 191.195 ;
        RECT 112.020 191.025 112.830 191.195 ;
        RECT 112.020 190.625 112.275 191.025 ;
        RECT 112.445 190.455 112.830 190.855 ;
        RECT 113.000 190.625 113.245 191.195 ;
        RECT 113.435 191.025 114.245 191.195 ;
        RECT 113.435 190.625 113.690 191.025 ;
        RECT 113.860 190.455 114.245 190.855 ;
        RECT 114.415 190.625 114.675 191.195 ;
        RECT 114.845 192.205 115.285 192.835 ;
        RECT 114.845 191.195 115.155 192.205 ;
        RECT 115.460 192.155 115.775 193.005 ;
        RECT 115.945 192.665 117.375 192.835 ;
        RECT 115.945 191.985 116.115 192.665 ;
        RECT 115.325 191.815 116.115 191.985 ;
        RECT 115.325 191.365 115.495 191.815 ;
        RECT 116.285 191.695 116.485 192.495 ;
        RECT 115.665 191.365 116.055 191.645 ;
        RECT 116.240 191.365 116.485 191.695 ;
        RECT 116.685 191.365 116.935 192.495 ;
        RECT 117.125 192.035 117.375 192.665 ;
        RECT 117.555 192.205 117.885 193.005 ;
        RECT 119.065 192.075 119.245 192.835 ;
        RECT 119.425 192.245 119.755 193.005 ;
        RECT 117.125 191.865 117.895 192.035 ;
        RECT 119.065 191.905 119.740 192.075 ;
        RECT 119.925 191.930 120.195 192.835 ;
        RECT 117.150 191.365 117.555 191.695 ;
        RECT 117.725 191.195 117.895 191.865 ;
        RECT 119.570 191.760 119.740 191.905 ;
        RECT 119.005 191.355 119.345 191.725 ;
        RECT 119.570 191.430 119.845 191.760 ;
        RECT 114.845 190.635 115.285 191.195 ;
        RECT 115.455 190.455 115.905 191.195 ;
        RECT 116.075 191.025 117.235 191.195 ;
        RECT 116.075 190.625 116.245 191.025 ;
        RECT 116.415 190.455 116.835 190.855 ;
        RECT 117.005 190.625 117.235 191.025 ;
        RECT 117.405 190.625 117.895 191.195 ;
        RECT 119.570 191.175 119.740 191.430 ;
        RECT 119.075 191.005 119.740 191.175 ;
        RECT 120.015 191.130 120.195 191.930 ;
        RECT 120.445 192.075 120.625 192.835 ;
        RECT 120.805 192.245 121.135 193.005 ;
        RECT 120.445 191.905 121.120 192.075 ;
        RECT 121.305 191.930 121.575 192.835 ;
        RECT 120.950 191.760 121.120 191.905 ;
        RECT 120.385 191.355 120.725 191.725 ;
        RECT 120.950 191.430 121.225 191.760 ;
        RECT 120.950 191.175 121.120 191.430 ;
        RECT 119.075 190.625 119.245 191.005 ;
        RECT 119.425 190.455 119.755 190.835 ;
        RECT 119.935 190.625 120.195 191.130 ;
        RECT 120.455 191.005 121.120 191.175 ;
        RECT 121.395 191.130 121.575 191.930 ;
        RECT 121.745 191.915 125.255 193.005 ;
        RECT 120.455 190.625 120.625 191.005 ;
        RECT 120.805 190.455 121.135 190.835 ;
        RECT 121.315 190.625 121.575 191.130 ;
        RECT 121.745 191.225 123.395 191.745 ;
        RECT 123.565 191.395 125.255 191.915 ;
        RECT 126.345 191.840 126.635 193.005 ;
        RECT 127.725 191.930 127.995 192.835 ;
        RECT 128.165 192.245 128.495 193.005 ;
        RECT 128.675 192.075 128.855 192.835 ;
        RECT 121.745 190.455 125.255 191.225 ;
        RECT 126.345 190.455 126.635 191.180 ;
        RECT 127.725 191.130 127.905 191.930 ;
        RECT 128.180 191.905 128.855 192.075 ;
        RECT 129.125 192.115 129.385 192.825 ;
        RECT 129.555 192.295 129.885 193.005 ;
        RECT 130.055 192.115 130.285 192.825 ;
        RECT 128.180 191.760 128.350 191.905 ;
        RECT 129.125 191.875 130.285 192.115 ;
        RECT 130.465 192.095 130.735 192.825 ;
        RECT 130.915 192.275 131.255 193.005 ;
        RECT 130.465 191.875 131.235 192.095 ;
        RECT 128.075 191.430 128.350 191.760 ;
        RECT 128.180 191.175 128.350 191.430 ;
        RECT 128.575 191.355 128.915 191.725 ;
        RECT 129.115 191.365 129.415 191.695 ;
        RECT 129.595 191.385 130.120 191.695 ;
        RECT 130.300 191.385 130.765 191.695 ;
        RECT 127.725 190.625 127.985 191.130 ;
        RECT 128.180 191.005 128.845 191.175 ;
        RECT 128.165 190.455 128.495 190.835 ;
        RECT 128.675 190.625 128.845 191.005 ;
        RECT 129.125 190.455 129.415 191.185 ;
        RECT 129.595 190.745 129.825 191.385 ;
        RECT 130.945 191.205 131.235 191.875 ;
        RECT 130.005 191.005 131.235 191.205 ;
        RECT 130.005 190.635 130.315 191.005 ;
        RECT 130.495 190.455 131.165 190.825 ;
        RECT 131.425 190.635 131.685 192.825 ;
        RECT 131.865 192.135 132.140 192.835 ;
        RECT 132.310 192.460 132.565 193.005 ;
        RECT 132.735 192.495 133.215 192.835 ;
        RECT 133.390 192.450 133.995 193.005 ;
        RECT 133.380 192.350 133.995 192.450 ;
        RECT 133.380 192.325 133.565 192.350 ;
        RECT 131.865 191.105 132.035 192.135 ;
        RECT 132.310 192.005 133.065 192.255 ;
        RECT 133.235 192.080 133.565 192.325 ;
        RECT 132.310 191.970 133.080 192.005 ;
        RECT 132.310 191.960 133.095 191.970 ;
        RECT 132.205 191.945 133.100 191.960 ;
        RECT 132.205 191.930 133.120 191.945 ;
        RECT 132.205 191.920 133.140 191.930 ;
        RECT 132.205 191.910 133.165 191.920 ;
        RECT 132.205 191.880 133.235 191.910 ;
        RECT 132.205 191.850 133.255 191.880 ;
        RECT 132.205 191.820 133.275 191.850 ;
        RECT 132.205 191.795 133.305 191.820 ;
        RECT 132.205 191.760 133.340 191.795 ;
        RECT 132.205 191.755 133.370 191.760 ;
        RECT 132.205 191.360 132.435 191.755 ;
        RECT 132.980 191.750 133.370 191.755 ;
        RECT 133.005 191.740 133.370 191.750 ;
        RECT 133.020 191.735 133.370 191.740 ;
        RECT 133.035 191.730 133.370 191.735 ;
        RECT 133.735 191.730 133.995 192.180 ;
        RECT 134.205 191.865 134.435 193.005 ;
        RECT 134.605 191.855 134.935 192.835 ;
        RECT 135.105 191.865 135.315 193.005 ;
        RECT 135.545 191.915 136.755 193.005 ;
        RECT 133.035 191.725 133.995 191.730 ;
        RECT 133.045 191.715 133.995 191.725 ;
        RECT 133.055 191.710 133.995 191.715 ;
        RECT 133.065 191.700 133.995 191.710 ;
        RECT 133.070 191.690 133.995 191.700 ;
        RECT 133.075 191.685 133.995 191.690 ;
        RECT 133.085 191.670 133.995 191.685 ;
        RECT 133.090 191.655 133.995 191.670 ;
        RECT 133.100 191.630 133.995 191.655 ;
        RECT 132.605 191.160 132.935 191.585 ;
        RECT 131.865 190.625 132.125 191.105 ;
        RECT 132.295 190.455 132.545 190.995 ;
        RECT 132.715 190.675 132.935 191.160 ;
        RECT 133.105 191.560 133.995 191.630 ;
        RECT 133.105 190.835 133.275 191.560 ;
        RECT 134.185 191.445 134.515 191.695 ;
        RECT 133.445 191.005 133.995 191.390 ;
        RECT 133.105 190.665 133.995 190.835 ;
        RECT 134.205 190.455 134.435 191.275 ;
        RECT 134.685 191.255 134.935 191.855 ;
        RECT 134.605 190.625 134.935 191.255 ;
        RECT 135.105 190.455 135.315 191.275 ;
        RECT 135.545 191.205 136.065 191.745 ;
        RECT 136.235 191.375 136.755 191.915 ;
        RECT 137.015 192.075 137.185 192.835 ;
        RECT 137.365 192.245 137.695 193.005 ;
        RECT 137.015 191.905 137.680 192.075 ;
        RECT 137.865 191.930 138.135 192.835 ;
        RECT 137.510 191.760 137.680 191.905 ;
        RECT 136.945 191.355 137.275 191.725 ;
        RECT 137.510 191.430 137.795 191.760 ;
        RECT 135.545 190.455 136.755 191.205 ;
        RECT 137.510 191.175 137.680 191.430 ;
        RECT 137.015 191.005 137.680 191.175 ;
        RECT 137.965 191.130 138.135 191.930 ;
        RECT 137.015 190.625 137.185 191.005 ;
        RECT 137.365 190.455 137.695 190.835 ;
        RECT 137.875 190.625 138.135 191.130 ;
        RECT 138.305 191.865 138.565 192.835 ;
        RECT 138.735 192.580 139.120 193.005 ;
        RECT 139.290 192.410 139.545 192.835 ;
        RECT 138.735 192.215 139.545 192.410 ;
        RECT 138.305 191.195 138.490 191.865 ;
        RECT 138.735 191.695 139.085 192.215 ;
        RECT 139.735 192.045 139.980 192.835 ;
        RECT 140.150 192.580 140.535 193.005 ;
        RECT 140.705 192.410 140.980 192.835 ;
        RECT 138.660 191.365 139.085 191.695 ;
        RECT 139.255 191.865 139.980 192.045 ;
        RECT 140.150 192.215 140.980 192.410 ;
        RECT 139.255 191.365 139.905 191.865 ;
        RECT 140.150 191.695 140.500 192.215 ;
        RECT 141.150 192.045 141.575 192.835 ;
        RECT 141.745 192.580 142.130 193.005 ;
        RECT 142.300 192.410 142.735 192.835 ;
        RECT 140.075 191.365 140.500 191.695 ;
        RECT 140.670 191.865 141.575 192.045 ;
        RECT 141.745 192.240 142.735 192.410 ;
        RECT 140.670 191.365 141.500 191.865 ;
        RECT 141.745 191.695 142.080 192.240 ;
        RECT 141.670 191.365 142.080 191.695 ;
        RECT 142.250 191.365 142.735 192.070 ;
        RECT 142.910 191.865 143.165 193.005 ;
        RECT 143.335 192.035 143.665 192.835 ;
        RECT 143.835 192.205 144.065 193.005 ;
        RECT 144.235 192.035 144.565 192.835 ;
        RECT 143.335 191.865 144.565 192.035 ;
        RECT 144.745 191.915 148.255 193.005 ;
        RECT 138.735 191.195 139.085 191.365 ;
        RECT 139.735 191.195 139.905 191.365 ;
        RECT 140.150 191.195 140.500 191.365 ;
        RECT 141.150 191.195 141.500 191.365 ;
        RECT 141.745 191.195 142.080 191.365 ;
        RECT 138.305 190.625 138.565 191.195 ;
        RECT 138.735 191.025 139.545 191.195 ;
        RECT 138.735 190.455 139.120 190.855 ;
        RECT 139.290 190.625 139.545 191.025 ;
        RECT 139.735 190.625 139.980 191.195 ;
        RECT 140.150 191.025 140.960 191.195 ;
        RECT 140.150 190.455 140.535 190.855 ;
        RECT 140.705 190.625 140.960 191.025 ;
        RECT 141.150 190.625 141.575 191.195 ;
        RECT 141.745 191.025 142.735 191.195 ;
        RECT 142.930 191.115 143.150 191.695 ;
        RECT 141.745 190.455 142.130 190.855 ;
        RECT 142.300 190.625 142.735 191.025 ;
        RECT 143.335 190.965 143.515 191.865 ;
        RECT 143.685 191.135 144.060 191.695 ;
        RECT 144.265 191.365 144.575 191.695 ;
        RECT 144.745 191.225 146.395 191.745 ;
        RECT 146.565 191.395 148.255 191.915 ;
        RECT 148.885 191.915 150.095 193.005 ;
        RECT 148.885 191.375 149.405 191.915 ;
        RECT 144.235 190.965 144.565 191.195 ;
        RECT 142.910 190.455 143.165 190.945 ;
        RECT 143.335 190.625 144.565 190.965 ;
        RECT 144.745 190.455 148.255 191.225 ;
        RECT 149.575 191.205 150.095 191.745 ;
        RECT 148.885 190.455 150.095 191.205 ;
        RECT 36.100 190.285 150.180 190.455 ;
        RECT 36.185 189.535 37.395 190.285 ;
        RECT 36.185 188.995 36.705 189.535 ;
        RECT 37.565 189.515 40.155 190.285 ;
        RECT 40.325 189.610 40.585 190.115 ;
        RECT 40.765 189.905 41.095 190.285 ;
        RECT 41.275 189.735 41.445 190.115 ;
        RECT 36.875 188.825 37.395 189.365 ;
        RECT 37.565 188.995 38.775 189.515 ;
        RECT 38.945 188.825 40.155 189.345 ;
        RECT 36.185 187.735 37.395 188.825 ;
        RECT 37.565 187.735 40.155 188.825 ;
        RECT 40.325 188.810 40.505 189.610 ;
        RECT 40.780 189.565 41.445 189.735 ;
        RECT 41.795 189.735 41.965 190.115 ;
        RECT 42.145 189.905 42.475 190.285 ;
        RECT 41.795 189.565 42.460 189.735 ;
        RECT 42.655 189.610 42.915 190.115 ;
        RECT 43.110 189.895 43.440 190.285 ;
        RECT 43.610 189.725 43.835 190.105 ;
        RECT 40.780 189.310 40.950 189.565 ;
        RECT 40.675 188.980 40.950 189.310 ;
        RECT 41.175 189.015 41.515 189.385 ;
        RECT 41.725 189.015 42.065 189.385 ;
        RECT 42.290 189.310 42.460 189.565 ;
        RECT 40.780 188.835 40.950 188.980 ;
        RECT 42.290 188.980 42.565 189.310 ;
        RECT 42.290 188.835 42.460 188.980 ;
        RECT 40.325 187.905 40.595 188.810 ;
        RECT 40.780 188.665 41.455 188.835 ;
        RECT 40.765 187.735 41.095 188.495 ;
        RECT 41.275 187.905 41.455 188.665 ;
        RECT 41.785 188.665 42.460 188.835 ;
        RECT 42.735 188.810 42.915 189.610 ;
        RECT 43.095 189.045 43.335 189.695 ;
        RECT 43.505 189.545 43.835 189.725 ;
        RECT 43.505 188.875 43.680 189.545 ;
        RECT 44.035 189.375 44.265 189.995 ;
        RECT 44.445 189.555 44.745 190.285 ;
        RECT 44.930 189.810 45.265 190.070 ;
        RECT 45.435 189.885 45.765 190.285 ;
        RECT 45.935 189.885 47.550 190.055 ;
        RECT 43.850 189.045 44.265 189.375 ;
        RECT 44.445 189.045 44.740 189.375 ;
        RECT 41.785 187.905 41.965 188.665 ;
        RECT 42.145 187.735 42.475 188.495 ;
        RECT 42.645 187.905 42.915 188.810 ;
        RECT 43.095 188.685 43.680 188.875 ;
        RECT 43.095 187.915 43.370 188.685 ;
        RECT 43.850 188.515 44.745 188.845 ;
        RECT 43.540 188.345 44.745 188.515 ;
        RECT 43.540 187.915 43.870 188.345 ;
        RECT 44.040 187.735 44.235 188.175 ;
        RECT 44.415 187.915 44.745 188.345 ;
        RECT 44.930 188.455 45.185 189.810 ;
        RECT 45.935 189.715 46.105 189.885 ;
        RECT 45.545 189.545 46.105 189.715 ;
        RECT 45.545 189.375 45.715 189.545 ;
        RECT 45.410 189.045 45.715 189.375 ;
        RECT 45.910 189.265 46.160 189.375 ;
        RECT 46.370 189.265 46.640 189.705 ;
        RECT 46.830 189.605 47.120 189.705 ;
        RECT 46.825 189.435 47.120 189.605 ;
        RECT 45.905 189.095 46.160 189.265 ;
        RECT 46.365 189.095 46.640 189.265 ;
        RECT 45.910 189.045 46.160 189.095 ;
        RECT 46.370 189.045 46.640 189.095 ;
        RECT 46.830 189.045 47.120 189.435 ;
        RECT 47.290 189.045 47.710 189.710 ;
        RECT 48.095 189.565 48.425 190.285 ;
        RECT 48.605 189.635 48.865 190.115 ;
        RECT 49.035 189.745 49.285 190.285 ;
        RECT 48.020 189.045 48.370 189.375 ;
        RECT 45.545 188.875 45.715 189.045 ;
        RECT 48.165 188.925 48.370 189.045 ;
        RECT 45.545 188.705 47.915 188.875 ;
        RECT 48.165 188.755 48.375 188.925 ;
        RECT 44.930 187.945 45.265 188.455 ;
        RECT 45.515 187.735 45.845 188.535 ;
        RECT 46.090 188.325 47.515 188.495 ;
        RECT 46.090 187.905 46.375 188.325 ;
        RECT 46.630 187.735 46.960 188.155 ;
        RECT 47.185 188.075 47.515 188.325 ;
        RECT 47.745 188.245 47.915 188.705 ;
        RECT 48.605 188.605 48.775 189.635 ;
        RECT 49.455 189.580 49.675 190.065 ;
        RECT 48.945 188.985 49.175 189.380 ;
        RECT 49.345 189.155 49.675 189.580 ;
        RECT 49.845 189.905 50.735 190.075 ;
        RECT 49.845 189.180 50.015 189.905 ;
        RECT 50.905 189.740 56.250 190.285 ;
        RECT 50.185 189.350 50.735 189.735 ;
        RECT 49.845 189.110 50.735 189.180 ;
        RECT 49.840 189.085 50.735 189.110 ;
        RECT 49.830 189.070 50.735 189.085 ;
        RECT 49.825 189.055 50.735 189.070 ;
        RECT 49.815 189.050 50.735 189.055 ;
        RECT 49.810 189.040 50.735 189.050 ;
        RECT 49.805 189.030 50.735 189.040 ;
        RECT 49.795 189.025 50.735 189.030 ;
        RECT 49.785 189.015 50.735 189.025 ;
        RECT 49.775 189.010 50.735 189.015 ;
        RECT 49.775 189.005 50.110 189.010 ;
        RECT 49.760 189.000 50.110 189.005 ;
        RECT 49.745 188.990 50.110 189.000 ;
        RECT 49.720 188.985 50.110 188.990 ;
        RECT 48.945 188.980 50.110 188.985 ;
        RECT 48.945 188.945 50.080 188.980 ;
        RECT 48.945 188.920 50.045 188.945 ;
        RECT 48.945 188.890 50.015 188.920 ;
        RECT 48.945 188.860 49.995 188.890 ;
        RECT 48.945 188.830 49.975 188.860 ;
        RECT 48.945 188.820 49.905 188.830 ;
        RECT 48.945 188.810 49.880 188.820 ;
        RECT 48.945 188.795 49.860 188.810 ;
        RECT 48.945 188.780 49.840 188.795 ;
        RECT 49.050 188.770 49.835 188.780 ;
        RECT 49.050 188.735 49.820 188.770 ;
        RECT 48.175 188.075 48.345 188.575 ;
        RECT 47.185 187.905 48.345 188.075 ;
        RECT 48.605 187.905 48.880 188.605 ;
        RECT 49.050 188.485 49.805 188.735 ;
        RECT 49.975 188.415 50.305 188.660 ;
        RECT 50.475 188.560 50.735 189.010 ;
        RECT 52.490 188.910 52.830 189.740 ;
        RECT 56.425 189.485 56.735 190.285 ;
        RECT 56.940 189.485 57.635 190.115 ;
        RECT 57.805 189.515 59.475 190.285 ;
        RECT 60.195 189.735 60.365 190.115 ;
        RECT 60.545 189.905 60.875 190.285 ;
        RECT 60.195 189.565 60.860 189.735 ;
        RECT 61.055 189.610 61.315 190.115 ;
        RECT 50.120 188.390 50.305 188.415 ;
        RECT 50.120 188.290 50.735 188.390 ;
        RECT 49.050 187.735 49.305 188.280 ;
        RECT 49.475 187.905 49.955 188.245 ;
        RECT 50.130 187.735 50.735 188.290 ;
        RECT 54.310 188.170 54.660 189.420 ;
        RECT 56.435 189.045 56.770 189.315 ;
        RECT 56.940 188.885 57.110 189.485 ;
        RECT 57.280 189.045 57.615 189.295 ;
        RECT 57.805 188.995 58.555 189.515 ;
        RECT 50.905 187.735 56.250 188.170 ;
        RECT 56.425 187.735 56.705 188.875 ;
        RECT 56.875 187.905 57.205 188.885 ;
        RECT 57.375 187.735 57.635 188.875 ;
        RECT 58.725 188.825 59.475 189.345 ;
        RECT 60.125 189.015 60.465 189.385 ;
        RECT 60.690 189.310 60.860 189.565 ;
        RECT 60.690 188.980 60.965 189.310 ;
        RECT 60.690 188.835 60.860 188.980 ;
        RECT 57.805 187.735 59.475 188.825 ;
        RECT 60.185 188.665 60.860 188.835 ;
        RECT 61.135 188.810 61.315 189.610 ;
        RECT 61.945 189.560 62.235 190.285 ;
        RECT 62.405 189.535 63.615 190.285 ;
        RECT 63.875 189.805 64.175 190.285 ;
        RECT 64.345 189.635 64.605 190.090 ;
        RECT 64.775 189.805 65.035 190.285 ;
        RECT 65.215 189.635 65.475 190.090 ;
        RECT 65.645 189.805 65.895 190.285 ;
        RECT 66.075 189.635 66.335 190.090 ;
        RECT 66.505 189.805 66.755 190.285 ;
        RECT 66.935 189.635 67.195 190.090 ;
        RECT 67.365 189.805 67.610 190.285 ;
        RECT 67.780 189.635 68.055 190.090 ;
        RECT 68.225 189.805 68.470 190.285 ;
        RECT 68.640 189.635 68.900 190.090 ;
        RECT 69.070 189.805 69.330 190.285 ;
        RECT 69.500 189.635 69.760 190.090 ;
        RECT 69.930 189.805 70.190 190.285 ;
        RECT 70.360 189.635 70.620 190.090 ;
        RECT 70.790 189.725 71.050 190.285 ;
        RECT 62.405 188.995 62.925 189.535 ;
        RECT 63.875 189.465 70.620 189.635 ;
        RECT 60.185 187.905 60.365 188.665 ;
        RECT 60.545 187.735 60.875 188.495 ;
        RECT 61.045 187.905 61.315 188.810 ;
        RECT 61.945 187.735 62.235 188.900 ;
        RECT 63.095 188.825 63.615 189.365 ;
        RECT 62.405 187.735 63.615 188.825 ;
        RECT 63.875 188.875 65.040 189.465 ;
        RECT 71.220 189.295 71.470 190.105 ;
        RECT 71.650 189.760 71.910 190.285 ;
        RECT 72.080 189.295 72.330 190.105 ;
        RECT 72.510 189.775 72.815 190.285 ;
        RECT 65.210 189.045 72.330 189.295 ;
        RECT 72.500 189.045 72.815 189.605 ;
        RECT 72.985 189.535 74.195 190.285 ;
        RECT 74.365 189.635 74.625 190.115 ;
        RECT 74.795 189.745 75.045 190.285 ;
        RECT 63.875 188.650 70.620 188.875 ;
        RECT 63.875 187.735 64.145 188.480 ;
        RECT 64.315 187.910 64.605 188.650 ;
        RECT 65.215 188.635 70.620 188.650 ;
        RECT 64.775 187.740 65.030 188.465 ;
        RECT 65.215 187.910 65.475 188.635 ;
        RECT 65.645 187.740 65.890 188.465 ;
        RECT 66.075 187.910 66.335 188.635 ;
        RECT 66.505 187.740 66.750 188.465 ;
        RECT 66.935 187.910 67.195 188.635 ;
        RECT 67.365 187.740 67.610 188.465 ;
        RECT 67.780 187.910 68.040 188.635 ;
        RECT 68.210 187.740 68.470 188.465 ;
        RECT 68.640 187.910 68.900 188.635 ;
        RECT 69.070 187.740 69.330 188.465 ;
        RECT 69.500 187.910 69.760 188.635 ;
        RECT 69.930 187.740 70.190 188.465 ;
        RECT 70.360 187.910 70.620 188.635 ;
        RECT 70.790 187.740 71.050 188.535 ;
        RECT 71.220 187.910 71.470 189.045 ;
        RECT 64.775 187.735 71.050 187.740 ;
        RECT 71.650 187.735 71.910 188.545 ;
        RECT 72.085 187.905 72.330 189.045 ;
        RECT 72.985 188.995 73.505 189.535 ;
        RECT 73.675 188.825 74.195 189.365 ;
        RECT 72.510 187.735 72.805 188.545 ;
        RECT 72.985 187.735 74.195 188.825 ;
        RECT 74.365 188.605 74.535 189.635 ;
        RECT 75.215 189.580 75.435 190.065 ;
        RECT 74.705 188.985 74.935 189.380 ;
        RECT 75.105 189.155 75.435 189.580 ;
        RECT 75.605 189.905 76.495 190.075 ;
        RECT 75.605 189.180 75.775 189.905 ;
        RECT 76.670 189.755 76.960 190.105 ;
        RECT 77.155 189.925 77.485 190.285 ;
        RECT 77.655 189.755 77.885 190.060 ;
        RECT 75.945 189.350 76.495 189.735 ;
        RECT 76.670 189.585 77.885 189.755 ;
        RECT 78.075 189.415 78.245 189.980 ;
        RECT 76.730 189.265 76.990 189.375 ;
        RECT 75.605 189.110 76.495 189.180 ;
        RECT 75.600 189.085 76.495 189.110 ;
        RECT 76.725 189.095 76.990 189.265 ;
        RECT 75.590 189.070 76.495 189.085 ;
        RECT 75.585 189.055 76.495 189.070 ;
        RECT 75.575 189.050 76.495 189.055 ;
        RECT 75.570 189.040 76.495 189.050 ;
        RECT 76.730 189.045 76.990 189.095 ;
        RECT 77.170 189.045 77.555 189.375 ;
        RECT 77.725 189.245 78.245 189.415 ;
        RECT 78.505 189.610 78.765 190.115 ;
        RECT 78.945 189.905 79.275 190.285 ;
        RECT 79.455 189.735 79.625 190.115 ;
        RECT 75.565 189.030 76.495 189.040 ;
        RECT 75.555 189.025 76.495 189.030 ;
        RECT 75.545 189.015 76.495 189.025 ;
        RECT 75.535 189.010 76.495 189.015 ;
        RECT 75.535 189.005 75.870 189.010 ;
        RECT 75.520 189.000 75.870 189.005 ;
        RECT 75.505 188.990 75.870 189.000 ;
        RECT 75.480 188.985 75.870 188.990 ;
        RECT 74.705 188.980 75.870 188.985 ;
        RECT 74.705 188.945 75.840 188.980 ;
        RECT 74.705 188.920 75.805 188.945 ;
        RECT 74.705 188.890 75.775 188.920 ;
        RECT 74.705 188.860 75.755 188.890 ;
        RECT 74.705 188.830 75.735 188.860 ;
        RECT 74.705 188.820 75.665 188.830 ;
        RECT 74.705 188.810 75.640 188.820 ;
        RECT 74.705 188.795 75.620 188.810 ;
        RECT 74.705 188.780 75.600 188.795 ;
        RECT 74.810 188.770 75.595 188.780 ;
        RECT 74.810 188.735 75.580 188.770 ;
        RECT 74.365 187.905 74.640 188.605 ;
        RECT 74.810 188.485 75.565 188.735 ;
        RECT 75.735 188.415 76.065 188.660 ;
        RECT 76.235 188.560 76.495 189.010 ;
        RECT 75.880 188.390 76.065 188.415 ;
        RECT 75.880 188.290 76.495 188.390 ;
        RECT 74.810 187.735 75.065 188.280 ;
        RECT 75.235 187.905 75.715 188.245 ;
        RECT 75.890 187.735 76.495 188.290 ;
        RECT 76.670 187.735 76.990 188.875 ;
        RECT 77.170 187.995 77.365 189.045 ;
        RECT 77.725 188.865 77.895 189.245 ;
        RECT 77.545 188.585 77.895 188.865 ;
        RECT 78.085 188.715 78.330 189.075 ;
        RECT 78.505 188.810 78.685 189.610 ;
        RECT 78.960 189.565 79.625 189.735 ;
        RECT 78.960 189.310 79.130 189.565 ;
        RECT 79.885 189.515 83.395 190.285 ;
        RECT 84.485 189.675 84.825 190.090 ;
        RECT 84.995 189.845 85.165 190.285 ;
        RECT 85.335 189.895 86.585 190.075 ;
        RECT 85.335 189.675 85.665 189.895 ;
        RECT 86.855 189.825 87.025 190.285 ;
        RECT 78.855 188.980 79.130 189.310 ;
        RECT 79.355 189.015 79.695 189.385 ;
        RECT 79.885 188.995 81.535 189.515 ;
        RECT 84.485 189.505 85.665 189.675 ;
        RECT 85.835 189.655 86.200 189.725 ;
        RECT 85.835 189.475 87.085 189.655 ;
        RECT 78.960 188.835 79.130 188.980 ;
        RECT 77.545 187.905 77.875 188.585 ;
        RECT 78.075 187.735 78.330 188.535 ;
        RECT 78.505 187.905 78.775 188.810 ;
        RECT 78.960 188.665 79.635 188.835 ;
        RECT 81.705 188.825 83.395 189.345 ;
        RECT 84.485 189.095 84.950 189.295 ;
        RECT 85.125 189.045 85.455 189.295 ;
        RECT 85.625 189.265 86.090 189.295 ;
        RECT 85.625 189.095 86.095 189.265 ;
        RECT 85.625 189.045 86.090 189.095 ;
        RECT 86.285 189.045 86.640 189.295 ;
        RECT 85.125 188.925 85.305 189.045 ;
        RECT 78.945 187.735 79.275 188.495 ;
        RECT 79.455 187.905 79.635 188.665 ;
        RECT 79.885 187.735 83.395 188.825 ;
        RECT 84.485 187.735 84.805 188.915 ;
        RECT 84.975 188.755 85.305 188.925 ;
        RECT 86.810 188.875 87.085 189.475 ;
        RECT 84.975 187.965 85.175 188.755 ;
        RECT 85.475 188.665 87.085 188.875 ;
        RECT 85.475 188.565 85.885 188.665 ;
        RECT 85.500 187.905 85.885 188.565 ;
        RECT 86.280 187.735 87.065 188.495 ;
        RECT 87.255 187.905 87.535 190.005 ;
        RECT 87.705 189.560 87.995 190.285 ;
        RECT 88.370 189.505 88.870 190.115 ;
        RECT 88.165 189.045 88.515 189.295 ;
        RECT 87.705 187.735 87.995 188.900 ;
        RECT 88.700 188.875 88.870 189.505 ;
        RECT 89.500 189.635 89.830 190.115 ;
        RECT 90.000 189.825 90.225 190.285 ;
        RECT 90.395 189.635 90.725 190.115 ;
        RECT 89.500 189.465 90.725 189.635 ;
        RECT 90.915 189.485 91.165 190.285 ;
        RECT 91.335 189.485 91.675 190.115 ;
        RECT 91.845 189.740 97.190 190.285 ;
        RECT 89.040 189.095 89.370 189.295 ;
        RECT 89.540 189.095 89.870 189.295 ;
        RECT 90.040 189.095 90.460 189.295 ;
        RECT 90.635 189.125 91.330 189.295 ;
        RECT 90.635 188.875 90.805 189.125 ;
        RECT 91.500 188.875 91.675 189.485 ;
        RECT 93.430 188.910 93.770 189.740 ;
        RECT 97.365 189.535 98.575 190.285 ;
        RECT 98.770 189.895 99.100 190.285 ;
        RECT 99.270 189.725 99.495 190.105 ;
        RECT 88.370 188.705 90.805 188.875 ;
        RECT 88.370 187.905 88.700 188.705 ;
        RECT 88.870 187.735 89.200 188.535 ;
        RECT 89.500 187.905 89.830 188.705 ;
        RECT 90.475 187.735 90.725 188.535 ;
        RECT 90.995 187.735 91.165 188.875 ;
        RECT 91.335 187.905 91.675 188.875 ;
        RECT 95.250 188.170 95.600 189.420 ;
        RECT 97.365 188.995 97.885 189.535 ;
        RECT 98.055 188.825 98.575 189.365 ;
        RECT 98.755 189.045 98.995 189.695 ;
        RECT 99.165 189.545 99.495 189.725 ;
        RECT 99.165 188.875 99.340 189.545 ;
        RECT 99.695 189.375 99.925 189.995 ;
        RECT 100.105 189.555 100.405 190.285 ;
        RECT 100.585 189.485 100.895 190.285 ;
        RECT 101.100 189.485 101.795 190.115 ;
        RECT 101.965 189.515 105.475 190.285 ;
        RECT 106.565 189.610 106.825 190.115 ;
        RECT 107.005 189.905 107.335 190.285 ;
        RECT 107.515 189.735 107.685 190.115 ;
        RECT 107.945 189.740 113.290 190.285 ;
        RECT 101.100 189.435 101.275 189.485 ;
        RECT 99.510 189.045 99.925 189.375 ;
        RECT 100.105 189.045 100.400 189.375 ;
        RECT 100.595 189.045 100.930 189.315 ;
        RECT 101.100 188.885 101.270 189.435 ;
        RECT 101.440 189.045 101.775 189.295 ;
        RECT 101.965 188.995 103.615 189.515 ;
        RECT 91.845 187.735 97.190 188.170 ;
        RECT 97.365 187.735 98.575 188.825 ;
        RECT 98.755 188.685 99.340 188.875 ;
        RECT 98.755 187.915 99.030 188.685 ;
        RECT 99.510 188.515 100.405 188.845 ;
        RECT 99.200 188.345 100.405 188.515 ;
        RECT 99.200 187.915 99.530 188.345 ;
        RECT 99.700 187.735 99.895 188.175 ;
        RECT 100.075 187.915 100.405 188.345 ;
        RECT 100.585 187.735 100.865 188.875 ;
        RECT 101.035 187.905 101.365 188.885 ;
        RECT 101.535 187.735 101.795 188.875 ;
        RECT 103.785 188.825 105.475 189.345 ;
        RECT 101.965 187.735 105.475 188.825 ;
        RECT 106.565 188.810 106.745 189.610 ;
        RECT 107.020 189.565 107.685 189.735 ;
        RECT 107.020 189.310 107.190 189.565 ;
        RECT 106.915 188.980 107.190 189.310 ;
        RECT 107.415 189.015 107.755 189.385 ;
        RECT 107.020 188.835 107.190 188.980 ;
        RECT 109.530 188.910 109.870 189.740 ;
        RECT 113.465 189.560 113.755 190.285 ;
        RECT 113.925 189.515 116.515 190.285 ;
        RECT 116.685 189.810 117.025 190.070 ;
        RECT 106.565 187.905 106.835 188.810 ;
        RECT 107.020 188.665 107.695 188.835 ;
        RECT 107.005 187.735 107.335 188.495 ;
        RECT 107.515 187.905 107.695 188.665 ;
        RECT 111.350 188.170 111.700 189.420 ;
        RECT 113.925 188.995 115.135 189.515 ;
        RECT 107.945 187.735 113.290 188.170 ;
        RECT 113.465 187.735 113.755 188.900 ;
        RECT 115.305 188.825 116.515 189.345 ;
        RECT 113.925 187.735 116.515 188.825 ;
        RECT 116.685 188.205 116.945 189.810 ;
        RECT 117.195 189.805 117.525 190.285 ;
        RECT 117.715 189.635 118.130 190.070 ;
        RECT 118.300 189.770 119.250 189.955 ;
        RECT 117.115 189.560 118.130 189.635 ;
        RECT 117.115 189.465 117.935 189.560 ;
        RECT 117.115 188.545 117.285 189.465 ;
        RECT 117.605 188.735 117.935 189.295 ;
        RECT 118.135 189.045 118.515 189.375 ;
        RECT 118.825 189.265 119.045 189.770 ;
        RECT 119.480 189.375 119.685 189.975 ;
        RECT 119.855 189.560 120.195 190.285 ;
        RECT 120.825 189.775 121.130 190.285 ;
        RECT 118.815 189.095 119.045 189.265 ;
        RECT 118.825 189.045 119.045 189.095 ;
        RECT 118.135 188.925 118.435 189.045 ;
        RECT 118.125 188.755 118.435 188.925 ;
        RECT 118.135 188.750 118.435 188.755 ;
        RECT 119.305 188.745 119.685 189.375 ;
        RECT 119.915 188.745 120.170 189.375 ;
        RECT 120.825 189.045 121.140 189.605 ;
        RECT 121.310 189.295 121.560 190.105 ;
        RECT 121.730 189.760 121.990 190.285 ;
        RECT 122.170 189.295 122.420 190.105 ;
        RECT 122.590 189.725 122.850 190.285 ;
        RECT 123.020 189.635 123.280 190.090 ;
        RECT 123.450 189.805 123.710 190.285 ;
        RECT 123.880 189.635 124.140 190.090 ;
        RECT 124.310 189.805 124.570 190.285 ;
        RECT 124.740 189.635 125.000 190.090 ;
        RECT 125.170 189.805 125.415 190.285 ;
        RECT 125.585 189.635 125.860 190.090 ;
        RECT 126.030 189.805 126.275 190.285 ;
        RECT 126.445 189.635 126.705 190.090 ;
        RECT 126.885 189.805 127.135 190.285 ;
        RECT 127.305 189.635 127.565 190.090 ;
        RECT 127.745 189.805 127.995 190.285 ;
        RECT 128.165 189.635 128.425 190.090 ;
        RECT 128.605 189.805 128.865 190.285 ;
        RECT 129.035 189.635 129.295 190.090 ;
        RECT 129.465 189.805 129.765 190.285 ;
        RECT 130.030 189.885 130.365 190.285 ;
        RECT 130.535 189.715 130.740 190.115 ;
        RECT 130.950 189.805 131.225 190.285 ;
        RECT 131.435 189.785 131.695 190.115 ;
        RECT 123.020 189.465 129.765 189.635 ;
        RECT 121.310 189.045 128.430 189.295 ;
        RECT 117.115 188.375 117.965 188.545 ;
        RECT 116.685 187.945 117.025 188.205 ;
        RECT 117.195 187.735 117.445 188.195 ;
        RECT 117.635 187.945 117.965 188.375 ;
        RECT 118.135 188.405 120.105 188.575 ;
        RECT 118.135 187.905 118.305 188.405 ;
        RECT 118.515 187.735 118.765 188.195 ;
        RECT 118.975 187.905 119.145 188.405 ;
        RECT 119.445 187.735 119.695 188.195 ;
        RECT 119.935 187.905 120.105 188.405 ;
        RECT 120.835 187.735 121.130 188.545 ;
        RECT 121.310 187.905 121.555 189.045 ;
        RECT 121.730 187.735 121.990 188.545 ;
        RECT 122.170 187.910 122.420 189.045 ;
        RECT 128.600 188.875 129.765 189.465 ;
        RECT 123.020 188.650 129.765 188.875 ;
        RECT 130.055 189.545 130.740 189.715 ;
        RECT 123.020 188.635 128.425 188.650 ;
        RECT 122.590 187.740 122.850 188.535 ;
        RECT 123.020 187.910 123.280 188.635 ;
        RECT 123.450 187.740 123.710 188.465 ;
        RECT 123.880 187.910 124.140 188.635 ;
        RECT 124.310 187.740 124.570 188.465 ;
        RECT 124.740 187.910 125.000 188.635 ;
        RECT 125.170 187.740 125.430 188.465 ;
        RECT 125.600 187.910 125.860 188.635 ;
        RECT 126.030 187.740 126.275 188.465 ;
        RECT 126.445 187.910 126.705 188.635 ;
        RECT 126.890 187.740 127.135 188.465 ;
        RECT 127.305 187.910 127.565 188.635 ;
        RECT 127.750 187.740 127.995 188.465 ;
        RECT 128.165 187.910 128.425 188.635 ;
        RECT 128.610 187.740 128.865 188.465 ;
        RECT 129.035 187.910 129.325 188.650 ;
        RECT 130.055 188.515 130.395 189.545 ;
        RECT 130.565 188.875 130.815 189.375 ;
        RECT 130.995 189.045 131.355 189.625 ;
        RECT 131.525 188.875 131.695 189.785 ;
        RECT 131.865 189.515 134.455 190.285 ;
        RECT 134.825 189.655 135.155 190.015 ;
        RECT 135.775 189.825 136.025 190.285 ;
        RECT 136.195 189.825 136.755 190.115 ;
        RECT 131.865 188.995 133.075 189.515 ;
        RECT 134.825 189.465 136.215 189.655 ;
        RECT 136.045 189.375 136.215 189.465 ;
        RECT 130.565 188.705 131.695 188.875 ;
        RECT 133.245 188.825 134.455 189.345 ;
        RECT 122.590 187.735 128.865 187.740 ;
        RECT 129.495 187.735 129.765 188.480 ;
        RECT 130.055 188.340 130.720 188.515 ;
        RECT 130.030 187.735 130.365 188.160 ;
        RECT 130.535 187.935 130.720 188.340 ;
        RECT 130.925 187.735 131.255 188.515 ;
        RECT 131.425 187.935 131.695 188.705 ;
        RECT 131.865 187.735 134.455 188.825 ;
        RECT 134.640 189.045 135.315 189.295 ;
        RECT 135.535 189.045 135.875 189.295 ;
        RECT 136.045 189.045 136.335 189.375 ;
        RECT 134.640 188.685 134.905 189.045 ;
        RECT 136.045 188.795 136.215 189.045 ;
        RECT 135.275 188.625 136.215 188.795 ;
        RECT 134.825 187.735 135.105 188.405 ;
        RECT 135.275 188.075 135.575 188.625 ;
        RECT 136.505 188.455 136.755 189.825 ;
        RECT 136.925 189.515 138.595 190.285 ;
        RECT 139.225 189.560 139.515 190.285 ;
        RECT 136.925 188.995 137.675 189.515 ;
        RECT 139.725 189.465 139.955 190.285 ;
        RECT 140.125 189.485 140.455 190.115 ;
        RECT 137.845 188.825 138.595 189.345 ;
        RECT 139.705 189.045 140.035 189.295 ;
        RECT 135.775 187.735 136.105 188.455 ;
        RECT 136.295 187.905 136.755 188.455 ;
        RECT 136.925 187.735 138.595 188.825 ;
        RECT 139.225 187.735 139.515 188.900 ;
        RECT 140.205 188.885 140.455 189.485 ;
        RECT 140.625 189.465 140.835 190.285 ;
        RECT 141.075 189.560 141.405 190.070 ;
        RECT 141.575 189.885 141.905 190.285 ;
        RECT 142.955 189.715 143.285 190.055 ;
        RECT 143.455 189.885 143.785 190.285 ;
        RECT 144.285 189.825 144.845 190.115 ;
        RECT 145.015 189.825 145.265 190.285 ;
        RECT 139.725 187.735 139.955 188.875 ;
        RECT 140.125 187.905 140.455 188.885 ;
        RECT 140.625 187.735 140.835 188.875 ;
        RECT 141.075 188.795 141.265 189.560 ;
        RECT 141.575 189.545 143.940 189.715 ;
        RECT 141.575 189.375 141.745 189.545 ;
        RECT 141.435 189.045 141.745 189.375 ;
        RECT 141.915 189.045 142.220 189.375 ;
        RECT 141.075 187.945 141.405 188.795 ;
        RECT 141.575 187.735 141.825 188.875 ;
        RECT 142.005 188.715 142.220 189.045 ;
        RECT 142.395 188.715 142.680 189.375 ;
        RECT 142.875 188.715 143.140 189.375 ;
        RECT 143.355 188.715 143.600 189.375 ;
        RECT 143.770 188.545 143.940 189.545 ;
        RECT 142.015 188.375 143.305 188.545 ;
        RECT 142.015 187.955 142.265 188.375 ;
        RECT 142.495 187.735 142.825 188.205 ;
        RECT 143.055 187.955 143.305 188.375 ;
        RECT 143.485 188.375 143.940 188.545 ;
        RECT 144.285 188.455 144.535 189.825 ;
        RECT 145.885 189.655 146.215 190.015 ;
        RECT 144.825 189.465 146.215 189.655 ;
        RECT 146.585 189.515 148.255 190.285 ;
        RECT 148.885 189.535 150.095 190.285 ;
        RECT 144.825 189.375 144.995 189.465 ;
        RECT 144.705 189.045 144.995 189.375 ;
        RECT 145.165 189.045 145.505 189.295 ;
        RECT 145.725 189.045 146.400 189.295 ;
        RECT 144.825 188.795 144.995 189.045 ;
        RECT 144.825 188.625 145.765 188.795 ;
        RECT 146.135 188.685 146.400 189.045 ;
        RECT 146.585 188.995 147.335 189.515 ;
        RECT 147.505 188.825 148.255 189.345 ;
        RECT 143.485 187.945 143.815 188.375 ;
        RECT 144.285 187.905 144.745 188.455 ;
        RECT 144.935 187.735 145.265 188.455 ;
        RECT 145.465 188.075 145.765 188.625 ;
        RECT 145.935 187.735 146.215 188.405 ;
        RECT 146.585 187.735 148.255 188.825 ;
        RECT 148.885 188.825 149.405 189.365 ;
        RECT 149.575 188.995 150.095 189.535 ;
        RECT 148.885 187.735 150.095 188.825 ;
        RECT 36.100 187.565 150.180 187.735 ;
        RECT 36.185 186.475 37.395 187.565 ;
        RECT 37.565 187.130 42.910 187.565 ;
        RECT 36.185 185.765 36.705 186.305 ;
        RECT 36.875 185.935 37.395 186.475 ;
        RECT 36.185 185.015 37.395 185.765 ;
        RECT 39.150 185.560 39.490 186.390 ;
        RECT 40.970 185.880 41.320 187.130 ;
        RECT 43.085 186.475 45.675 187.565 ;
        RECT 43.085 185.785 44.295 186.305 ;
        RECT 44.465 185.955 45.675 186.475 ;
        RECT 45.845 186.765 46.285 187.395 ;
        RECT 37.565 185.015 42.910 185.560 ;
        RECT 43.085 185.015 45.675 185.785 ;
        RECT 45.845 185.755 46.155 186.765 ;
        RECT 46.460 186.715 46.775 187.565 ;
        RECT 46.945 187.225 48.375 187.395 ;
        RECT 46.945 186.545 47.115 187.225 ;
        RECT 46.325 186.375 47.115 186.545 ;
        RECT 46.325 185.925 46.495 186.375 ;
        RECT 47.285 186.255 47.485 187.055 ;
        RECT 46.665 185.925 47.055 186.205 ;
        RECT 47.240 185.925 47.485 186.255 ;
        RECT 47.685 185.925 47.935 187.055 ;
        RECT 48.125 186.595 48.375 187.225 ;
        RECT 48.555 186.765 48.885 187.565 ;
        RECT 48.125 186.425 48.895 186.595 ;
        RECT 48.150 185.925 48.555 186.255 ;
        RECT 48.725 185.755 48.895 186.425 ;
        RECT 49.065 186.400 49.355 187.565 ;
        RECT 49.525 186.425 49.795 187.395 ;
        RECT 50.005 186.765 50.285 187.565 ;
        RECT 50.455 187.055 52.110 187.345 ;
        RECT 52.285 187.130 57.630 187.565 ;
        RECT 50.520 186.715 52.110 186.885 ;
        RECT 50.520 186.595 50.690 186.715 ;
        RECT 49.965 186.425 50.690 186.595 ;
        RECT 45.845 185.195 46.285 185.755 ;
        RECT 46.455 185.015 46.905 185.755 ;
        RECT 47.075 185.585 48.235 185.755 ;
        RECT 47.075 185.185 47.245 185.585 ;
        RECT 47.415 185.015 47.835 185.415 ;
        RECT 48.005 185.185 48.235 185.585 ;
        RECT 48.405 185.185 48.895 185.755 ;
        RECT 49.065 185.015 49.355 185.740 ;
        RECT 49.525 185.690 49.695 186.425 ;
        RECT 49.965 186.255 50.135 186.425 ;
        RECT 49.865 185.925 50.135 186.255 ;
        RECT 50.305 185.925 50.710 186.255 ;
        RECT 50.880 185.925 51.590 186.545 ;
        RECT 51.790 186.425 52.110 186.715 ;
        RECT 49.965 185.755 50.135 185.925 ;
        RECT 49.525 185.345 49.795 185.690 ;
        RECT 49.965 185.585 51.575 185.755 ;
        RECT 51.760 185.685 52.110 186.255 ;
        RECT 49.985 185.015 50.365 185.415 ;
        RECT 50.535 185.235 50.705 185.585 ;
        RECT 50.875 185.015 51.205 185.415 ;
        RECT 51.405 185.235 51.575 185.585 ;
        RECT 53.870 185.560 54.210 186.390 ;
        RECT 55.690 185.880 56.040 187.130 ;
        RECT 58.105 186.925 58.435 187.355 ;
        RECT 57.980 186.755 58.435 186.925 ;
        RECT 58.615 186.925 58.865 187.345 ;
        RECT 59.095 187.095 59.425 187.565 ;
        RECT 59.655 186.925 59.905 187.345 ;
        RECT 58.615 186.755 59.905 186.925 ;
        RECT 57.980 185.755 58.150 186.755 ;
        RECT 58.320 185.925 58.565 186.585 ;
        RECT 58.780 185.925 59.045 186.585 ;
        RECT 59.240 185.925 59.525 186.585 ;
        RECT 59.700 186.255 59.915 186.585 ;
        RECT 60.095 186.425 60.345 187.565 ;
        RECT 60.515 186.505 60.845 187.355 ;
        RECT 61.115 187.015 61.285 187.305 ;
        RECT 61.455 187.185 61.785 187.565 ;
        RECT 62.350 187.055 63.180 187.225 ;
        RECT 61.115 186.885 61.605 187.015 ;
        RECT 61.115 186.845 62.840 186.885 ;
        RECT 61.435 186.715 62.840 186.845 ;
        RECT 59.700 185.925 60.005 186.255 ;
        RECT 60.175 185.925 60.485 186.255 ;
        RECT 60.175 185.755 60.345 185.925 ;
        RECT 57.980 185.585 60.345 185.755 ;
        RECT 60.655 185.740 60.845 186.505 ;
        RECT 61.085 185.905 61.265 186.675 ;
        RECT 51.775 185.015 52.105 185.515 ;
        RECT 52.285 185.015 57.630 185.560 ;
        RECT 58.135 185.015 58.465 185.415 ;
        RECT 58.635 185.245 58.965 185.585 ;
        RECT 60.015 185.015 60.345 185.415 ;
        RECT 60.515 185.230 60.845 185.740 ;
        RECT 61.435 185.735 61.605 186.715 ;
        RECT 61.945 186.375 62.330 186.545 ;
        RECT 62.160 186.215 62.330 186.375 ;
        RECT 62.500 186.505 62.840 186.715 ;
        RECT 61.110 185.565 61.605 185.735 ;
        RECT 61.775 185.695 62.175 186.025 ;
        RECT 62.500 185.965 62.670 186.505 ;
        RECT 63.010 186.335 63.180 187.055 ;
        RECT 63.535 186.985 63.765 187.565 ;
        RECT 64.245 187.055 64.760 187.225 ;
        RECT 63.910 186.715 64.255 186.885 ;
        RECT 64.505 186.740 64.760 187.055 ;
        RECT 64.085 186.590 64.255 186.715 ;
        RECT 64.085 186.420 64.355 186.590 ;
        RECT 61.110 185.275 61.285 185.565 ;
        RECT 61.455 185.015 61.785 185.395 ;
        RECT 61.960 185.325 62.175 185.695 ;
        RECT 62.345 185.635 62.670 185.965 ;
        RECT 62.840 186.165 63.180 186.335 ;
        RECT 64.185 186.320 64.355 186.420 ;
        RECT 62.840 185.465 63.010 186.165 ;
        RECT 63.350 185.945 63.555 186.250 ;
        RECT 63.180 185.645 63.555 185.945 ;
        RECT 63.725 185.645 64.015 186.250 ;
        RECT 64.185 185.990 64.420 186.320 ;
        RECT 62.410 185.295 63.010 185.465 ;
        RECT 63.390 185.015 63.720 185.475 ;
        RECT 64.185 185.395 64.355 185.990 ;
        RECT 64.590 185.605 64.760 186.740 ;
        RECT 63.925 185.225 64.355 185.395 ;
        RECT 64.525 185.275 64.760 185.605 ;
        RECT 64.930 187.055 65.455 187.225 ;
        RECT 64.930 185.275 65.120 187.055 ;
        RECT 65.695 186.935 66.040 187.565 ;
        RECT 66.265 187.085 67.215 187.255 ;
        RECT 65.335 186.665 65.525 186.825 ;
        RECT 66.265 186.665 66.435 187.085 ;
        RECT 67.465 187.055 67.785 187.225 ;
        RECT 65.335 186.495 66.435 186.665 ;
        RECT 65.335 185.515 65.505 186.495 ;
        RECT 65.685 185.645 66.055 186.325 ;
        RECT 65.335 185.185 65.540 185.515 ;
        RECT 65.735 185.015 66.065 185.475 ;
        RECT 66.265 185.395 66.435 186.495 ;
        RECT 66.605 185.965 66.895 186.915 ;
        RECT 67.615 186.595 67.785 187.055 ;
        RECT 67.955 186.765 68.125 187.565 ;
        RECT 68.295 186.765 68.705 187.385 ;
        RECT 67.065 186.175 67.405 186.575 ;
        RECT 67.615 186.425 68.225 186.595 ;
        RECT 68.395 186.425 68.705 186.765 ;
        RECT 68.875 186.425 69.125 187.565 ;
        RECT 69.305 186.475 72.815 187.565 ;
        RECT 68.055 186.255 68.225 186.425 ;
        RECT 67.575 186.005 67.885 186.255 ;
        RECT 66.605 185.635 67.225 185.965 ;
        RECT 67.475 185.925 67.885 186.005 ;
        RECT 68.055 185.925 68.365 186.255 ;
        RECT 66.265 185.225 67.160 185.395 ;
        RECT 67.475 185.305 67.785 185.925 ;
        RECT 67.955 185.015 68.205 185.745 ;
        RECT 68.535 185.655 68.705 186.425 ;
        RECT 68.375 185.195 68.705 185.655 ;
        RECT 68.875 185.015 69.130 185.815 ;
        RECT 69.305 185.785 70.955 186.305 ;
        RECT 71.125 185.955 72.815 186.475 ;
        RECT 72.995 186.955 73.325 187.385 ;
        RECT 73.505 187.125 73.700 187.565 ;
        RECT 73.870 186.955 74.200 187.385 ;
        RECT 72.995 186.785 74.200 186.955 ;
        RECT 72.995 186.455 73.890 186.785 ;
        RECT 74.370 186.615 74.645 187.385 ;
        RECT 74.060 186.425 74.645 186.615 ;
        RECT 73.000 185.925 73.295 186.255 ;
        RECT 73.475 185.925 73.890 186.255 ;
        RECT 69.305 185.015 72.815 185.785 ;
        RECT 72.995 185.015 73.295 185.745 ;
        RECT 73.475 185.305 73.705 185.925 ;
        RECT 74.060 185.755 74.235 186.425 ;
        RECT 74.825 186.400 75.115 187.565 ;
        RECT 75.375 186.895 75.545 187.395 ;
        RECT 75.715 187.065 76.045 187.565 ;
        RECT 75.375 186.725 76.040 186.895 ;
        RECT 73.905 185.575 74.235 185.755 ;
        RECT 74.405 185.605 74.645 186.255 ;
        RECT 75.290 185.905 75.640 186.555 ;
        RECT 73.905 185.195 74.130 185.575 ;
        RECT 74.300 185.015 74.630 185.405 ;
        RECT 74.825 185.015 75.115 185.740 ;
        RECT 75.810 185.735 76.040 186.725 ;
        RECT 75.375 185.565 76.040 185.735 ;
        RECT 75.375 185.275 75.545 185.565 ;
        RECT 75.715 185.015 76.045 185.395 ;
        RECT 76.215 185.275 76.400 187.395 ;
        RECT 76.640 187.105 76.905 187.565 ;
        RECT 77.075 186.970 77.325 187.395 ;
        RECT 77.535 187.120 78.640 187.290 ;
        RECT 77.020 186.840 77.325 186.970 ;
        RECT 76.570 185.645 76.850 186.595 ;
        RECT 77.020 185.735 77.190 186.840 ;
        RECT 77.360 186.055 77.600 186.650 ;
        RECT 77.770 186.585 78.300 186.950 ;
        RECT 77.770 185.885 77.940 186.585 ;
        RECT 78.470 186.505 78.640 187.120 ;
        RECT 78.810 186.765 78.980 187.565 ;
        RECT 79.150 187.065 79.400 187.395 ;
        RECT 79.625 187.095 80.510 187.265 ;
        RECT 78.470 186.415 78.980 186.505 ;
        RECT 77.020 185.605 77.245 185.735 ;
        RECT 77.415 185.665 77.940 185.885 ;
        RECT 78.110 186.245 78.980 186.415 ;
        RECT 76.655 185.015 76.905 185.475 ;
        RECT 77.075 185.465 77.245 185.605 ;
        RECT 78.110 185.465 78.280 186.245 ;
        RECT 78.810 186.175 78.980 186.245 ;
        RECT 78.490 185.995 78.690 186.025 ;
        RECT 79.150 185.995 79.320 187.065 ;
        RECT 79.490 186.175 79.680 186.895 ;
        RECT 78.490 185.695 79.320 185.995 ;
        RECT 79.850 185.965 80.170 186.925 ;
        RECT 77.075 185.295 77.410 185.465 ;
        RECT 77.605 185.295 78.280 185.465 ;
        RECT 78.600 185.015 78.970 185.515 ;
        RECT 79.150 185.465 79.320 185.695 ;
        RECT 79.705 185.635 80.170 185.965 ;
        RECT 80.340 186.255 80.510 187.095 ;
        RECT 80.690 187.065 81.005 187.565 ;
        RECT 81.235 186.835 81.575 187.395 ;
        RECT 80.680 186.460 81.575 186.835 ;
        RECT 81.745 186.555 81.915 187.565 ;
        RECT 81.385 186.255 81.575 186.460 ;
        RECT 82.085 186.505 82.415 187.350 ;
        RECT 82.085 186.425 82.475 186.505 ;
        RECT 82.645 186.475 86.155 187.565 ;
        RECT 86.325 186.475 87.535 187.565 ;
        RECT 82.260 186.375 82.475 186.425 ;
        RECT 80.340 185.925 81.215 186.255 ;
        RECT 81.385 185.925 82.135 186.255 ;
        RECT 80.340 185.465 80.510 185.925 ;
        RECT 81.385 185.755 81.585 185.925 ;
        RECT 82.305 185.795 82.475 186.375 ;
        RECT 82.250 185.755 82.475 185.795 ;
        RECT 79.150 185.295 79.555 185.465 ;
        RECT 79.725 185.295 80.510 185.465 ;
        RECT 80.785 185.015 80.995 185.545 ;
        RECT 81.255 185.230 81.585 185.755 ;
        RECT 82.095 185.670 82.475 185.755 ;
        RECT 82.645 185.785 84.295 186.305 ;
        RECT 84.465 185.955 86.155 186.475 ;
        RECT 81.755 185.015 81.925 185.625 ;
        RECT 82.095 185.235 82.425 185.670 ;
        RECT 82.645 185.015 86.155 185.785 ;
        RECT 86.325 185.765 86.845 186.305 ;
        RECT 87.015 185.935 87.535 186.475 ;
        RECT 87.705 186.490 87.975 187.395 ;
        RECT 88.145 186.805 88.475 187.565 ;
        RECT 88.655 186.635 88.835 187.395 ;
        RECT 89.085 187.130 94.430 187.565 ;
        RECT 86.325 185.015 87.535 185.765 ;
        RECT 87.705 185.690 87.885 186.490 ;
        RECT 88.160 186.465 88.835 186.635 ;
        RECT 88.160 186.320 88.330 186.465 ;
        RECT 88.055 185.990 88.330 186.320 ;
        RECT 88.160 185.735 88.330 185.990 ;
        RECT 88.555 185.915 88.895 186.285 ;
        RECT 87.705 185.185 87.965 185.690 ;
        RECT 88.160 185.565 88.825 185.735 ;
        RECT 88.145 185.015 88.475 185.395 ;
        RECT 88.655 185.185 88.825 185.565 ;
        RECT 90.670 185.560 91.010 186.390 ;
        RECT 92.490 185.880 92.840 187.130 ;
        RECT 94.605 186.970 95.040 187.395 ;
        RECT 95.210 187.140 95.595 187.565 ;
        RECT 94.605 186.800 95.595 186.970 ;
        RECT 94.605 185.925 95.090 186.630 ;
        RECT 95.260 186.255 95.595 186.800 ;
        RECT 95.765 186.605 96.190 187.395 ;
        RECT 96.360 186.970 96.635 187.395 ;
        RECT 96.805 187.140 97.190 187.565 ;
        RECT 96.360 186.775 97.190 186.970 ;
        RECT 95.765 186.425 96.670 186.605 ;
        RECT 95.260 185.925 95.670 186.255 ;
        RECT 95.840 185.925 96.670 186.425 ;
        RECT 96.840 186.255 97.190 186.775 ;
        RECT 97.360 186.605 97.605 187.395 ;
        RECT 97.795 186.970 98.050 187.395 ;
        RECT 98.220 187.140 98.605 187.565 ;
        RECT 97.795 186.775 98.605 186.970 ;
        RECT 97.360 186.425 98.085 186.605 ;
        RECT 96.840 185.925 97.265 186.255 ;
        RECT 97.435 185.925 98.085 186.425 ;
        RECT 98.255 186.255 98.605 186.775 ;
        RECT 98.775 186.425 99.035 187.395 ;
        RECT 99.205 186.475 100.415 187.565 ;
        RECT 98.255 185.925 98.680 186.255 ;
        RECT 95.260 185.755 95.595 185.925 ;
        RECT 95.840 185.755 96.190 185.925 ;
        RECT 96.840 185.755 97.190 185.925 ;
        RECT 97.435 185.755 97.605 185.925 ;
        RECT 98.255 185.755 98.605 185.925 ;
        RECT 98.850 185.755 99.035 186.425 ;
        RECT 94.605 185.585 95.595 185.755 ;
        RECT 89.085 185.015 94.430 185.560 ;
        RECT 94.605 185.185 95.040 185.585 ;
        RECT 95.210 185.015 95.595 185.415 ;
        RECT 95.765 185.185 96.190 185.755 ;
        RECT 96.380 185.585 97.190 185.755 ;
        RECT 96.380 185.185 96.635 185.585 ;
        RECT 96.805 185.015 97.190 185.415 ;
        RECT 97.360 185.185 97.605 185.755 ;
        RECT 97.795 185.585 98.605 185.755 ;
        RECT 97.795 185.185 98.050 185.585 ;
        RECT 98.220 185.015 98.605 185.415 ;
        RECT 98.775 185.185 99.035 185.755 ;
        RECT 99.205 185.765 99.725 186.305 ;
        RECT 99.895 185.935 100.415 186.475 ;
        RECT 100.585 186.400 100.875 187.565 ;
        RECT 101.045 186.970 101.480 187.395 ;
        RECT 101.650 187.140 102.035 187.565 ;
        RECT 101.045 186.800 102.035 186.970 ;
        RECT 101.045 185.925 101.530 186.630 ;
        RECT 101.700 186.255 102.035 186.800 ;
        RECT 102.205 186.605 102.630 187.395 ;
        RECT 102.800 186.970 103.075 187.395 ;
        RECT 103.245 187.140 103.630 187.565 ;
        RECT 102.800 186.775 103.630 186.970 ;
        RECT 102.205 186.425 103.110 186.605 ;
        RECT 101.700 185.925 102.110 186.255 ;
        RECT 102.280 185.925 103.110 186.425 ;
        RECT 103.280 186.255 103.630 186.775 ;
        RECT 103.800 186.605 104.045 187.395 ;
        RECT 104.235 186.970 104.490 187.395 ;
        RECT 104.660 187.140 105.045 187.565 ;
        RECT 104.235 186.775 105.045 186.970 ;
        RECT 103.800 186.425 104.525 186.605 ;
        RECT 103.280 185.925 103.705 186.255 ;
        RECT 103.875 185.925 104.525 186.425 ;
        RECT 104.695 186.255 105.045 186.775 ;
        RECT 105.215 186.425 105.475 187.395 ;
        RECT 104.695 185.925 105.120 186.255 ;
        RECT 99.205 185.015 100.415 185.765 ;
        RECT 101.700 185.755 102.035 185.925 ;
        RECT 102.280 185.755 102.630 185.925 ;
        RECT 103.280 185.755 103.630 185.925 ;
        RECT 103.875 185.755 104.045 185.925 ;
        RECT 104.695 185.755 105.045 185.925 ;
        RECT 105.290 185.755 105.475 186.425 ;
        RECT 100.585 185.015 100.875 185.740 ;
        RECT 101.045 185.585 102.035 185.755 ;
        RECT 101.045 185.185 101.480 185.585 ;
        RECT 101.650 185.015 102.035 185.415 ;
        RECT 102.205 185.185 102.630 185.755 ;
        RECT 102.820 185.585 103.630 185.755 ;
        RECT 102.820 185.185 103.075 185.585 ;
        RECT 103.245 185.015 103.630 185.415 ;
        RECT 103.800 185.185 104.045 185.755 ;
        RECT 104.235 185.585 105.045 185.755 ;
        RECT 104.235 185.185 104.490 185.585 ;
        RECT 104.660 185.015 105.045 185.415 ;
        RECT 105.215 185.185 105.475 185.755 ;
        RECT 105.645 186.425 105.905 187.395 ;
        RECT 106.075 187.140 106.460 187.565 ;
        RECT 106.630 186.970 106.885 187.395 ;
        RECT 106.075 186.775 106.885 186.970 ;
        RECT 105.645 185.755 105.830 186.425 ;
        RECT 106.075 186.255 106.425 186.775 ;
        RECT 107.075 186.605 107.320 187.395 ;
        RECT 107.490 187.140 107.875 187.565 ;
        RECT 108.045 186.970 108.320 187.395 ;
        RECT 106.000 185.925 106.425 186.255 ;
        RECT 106.595 186.425 107.320 186.605 ;
        RECT 107.490 186.775 108.320 186.970 ;
        RECT 106.595 185.925 107.245 186.425 ;
        RECT 107.490 186.255 107.840 186.775 ;
        RECT 108.490 186.605 108.915 187.395 ;
        RECT 109.085 187.140 109.470 187.565 ;
        RECT 109.640 186.970 110.075 187.395 ;
        RECT 107.415 185.925 107.840 186.255 ;
        RECT 108.010 186.425 108.915 186.605 ;
        RECT 109.085 186.800 110.075 186.970 ;
        RECT 110.245 186.970 110.680 187.395 ;
        RECT 110.850 187.140 111.235 187.565 ;
        RECT 110.245 186.800 111.235 186.970 ;
        RECT 108.010 185.925 108.840 186.425 ;
        RECT 109.085 186.255 109.420 186.800 ;
        RECT 109.010 185.925 109.420 186.255 ;
        RECT 109.590 185.925 110.075 186.630 ;
        RECT 110.245 185.925 110.730 186.630 ;
        RECT 110.900 186.255 111.235 186.800 ;
        RECT 111.405 186.605 111.830 187.395 ;
        RECT 112.000 186.970 112.275 187.395 ;
        RECT 112.445 187.140 112.830 187.565 ;
        RECT 112.000 186.775 112.830 186.970 ;
        RECT 111.405 186.425 112.310 186.605 ;
        RECT 110.900 185.925 111.310 186.255 ;
        RECT 111.480 185.925 112.310 186.425 ;
        RECT 112.480 186.255 112.830 186.775 ;
        RECT 113.000 186.605 113.245 187.395 ;
        RECT 113.435 186.970 113.690 187.395 ;
        RECT 113.860 187.140 114.245 187.565 ;
        RECT 113.435 186.775 114.245 186.970 ;
        RECT 113.000 186.425 113.725 186.605 ;
        RECT 112.480 185.925 112.905 186.255 ;
        RECT 113.075 185.925 113.725 186.425 ;
        RECT 113.895 186.255 114.245 186.775 ;
        RECT 114.415 186.425 114.675 187.395 ;
        RECT 114.850 186.425 115.105 187.565 ;
        RECT 115.275 186.595 115.605 187.395 ;
        RECT 115.775 186.765 115.945 187.565 ;
        RECT 116.115 186.595 116.445 187.395 ;
        RECT 116.615 186.765 116.945 187.565 ;
        RECT 117.115 186.595 117.445 187.395 ;
        RECT 117.755 186.765 118.085 187.565 ;
        RECT 118.355 186.595 118.685 187.395 ;
        RECT 113.895 185.925 114.320 186.255 ;
        RECT 106.075 185.755 106.425 185.925 ;
        RECT 107.075 185.755 107.245 185.925 ;
        RECT 107.490 185.755 107.840 185.925 ;
        RECT 108.490 185.755 108.840 185.925 ;
        RECT 109.085 185.755 109.420 185.925 ;
        RECT 110.900 185.755 111.235 185.925 ;
        RECT 111.480 185.755 111.830 185.925 ;
        RECT 112.480 185.755 112.830 185.925 ;
        RECT 113.075 185.755 113.245 185.925 ;
        RECT 113.895 185.755 114.245 185.925 ;
        RECT 114.490 185.755 114.675 186.425 ;
        RECT 115.275 186.375 118.685 186.595 ;
        RECT 118.855 186.375 119.185 187.565 ;
        RECT 120.365 187.135 120.705 187.395 ;
        RECT 114.870 186.005 115.605 186.205 ;
        RECT 115.830 186.005 116.460 186.205 ;
        RECT 116.995 186.005 117.840 186.205 ;
        RECT 118.130 185.985 118.685 186.375 ;
        RECT 118.925 186.005 119.255 186.205 ;
        RECT 105.645 185.185 105.905 185.755 ;
        RECT 106.075 185.585 106.885 185.755 ;
        RECT 106.075 185.015 106.460 185.415 ;
        RECT 106.630 185.185 106.885 185.585 ;
        RECT 107.075 185.185 107.320 185.755 ;
        RECT 107.490 185.585 108.300 185.755 ;
        RECT 107.490 185.015 107.875 185.415 ;
        RECT 108.045 185.185 108.300 185.585 ;
        RECT 108.490 185.185 108.915 185.755 ;
        RECT 109.085 185.585 110.075 185.755 ;
        RECT 109.085 185.015 109.470 185.415 ;
        RECT 109.640 185.185 110.075 185.585 ;
        RECT 110.245 185.585 111.235 185.755 ;
        RECT 110.245 185.185 110.680 185.585 ;
        RECT 110.850 185.015 111.235 185.415 ;
        RECT 111.405 185.185 111.830 185.755 ;
        RECT 112.020 185.585 112.830 185.755 ;
        RECT 112.020 185.185 112.275 185.585 ;
        RECT 112.445 185.015 112.830 185.415 ;
        RECT 113.000 185.185 113.245 185.755 ;
        RECT 113.435 185.585 114.245 185.755 ;
        RECT 113.435 185.185 113.690 185.585 ;
        RECT 113.860 185.015 114.245 185.415 ;
        RECT 114.415 185.185 114.675 185.755 ;
        RECT 114.850 185.665 115.945 185.835 ;
        RECT 114.850 185.185 115.185 185.665 ;
        RECT 115.355 185.015 115.525 185.475 ;
        RECT 115.695 185.395 115.945 185.665 ;
        RECT 116.115 185.565 117.845 185.835 ;
        RECT 118.015 185.395 118.185 185.815 ;
        RECT 118.355 185.565 118.685 185.985 ;
        RECT 118.855 185.395 119.185 185.835 ;
        RECT 115.695 185.185 116.885 185.395 ;
        RECT 117.075 185.185 119.185 185.395 ;
        RECT 120.365 185.735 120.625 187.135 ;
        RECT 120.875 186.765 121.205 187.565 ;
        RECT 121.670 186.595 121.920 187.395 ;
        RECT 122.105 186.845 122.435 187.565 ;
        RECT 122.655 186.595 122.905 187.395 ;
        RECT 123.075 187.185 123.410 187.565 ;
        RECT 120.815 186.425 123.005 186.595 ;
        RECT 120.815 186.255 121.130 186.425 ;
        RECT 120.800 186.005 121.130 186.255 ;
        RECT 120.365 185.225 120.705 185.735 ;
        RECT 120.875 185.015 121.145 185.815 ;
        RECT 121.325 185.285 121.605 186.255 ;
        RECT 121.785 185.285 122.085 186.255 ;
        RECT 122.265 185.290 122.615 186.255 ;
        RECT 122.835 185.515 123.005 186.425 ;
        RECT 123.175 185.695 123.415 187.005 ;
        RECT 123.770 186.595 124.160 186.770 ;
        RECT 124.645 186.765 124.975 187.565 ;
        RECT 125.145 186.775 125.680 187.395 ;
        RECT 123.770 186.425 125.195 186.595 ;
        RECT 123.645 185.695 124.000 186.255 ;
        RECT 124.170 185.525 124.340 186.425 ;
        RECT 124.510 185.695 124.775 186.255 ;
        RECT 125.025 185.925 125.195 186.425 ;
        RECT 125.365 185.755 125.680 186.775 ;
        RECT 126.345 186.400 126.635 187.565 ;
        RECT 126.805 187.010 127.410 187.565 ;
        RECT 127.585 187.055 128.065 187.395 ;
        RECT 128.235 187.020 128.490 187.565 ;
        RECT 126.805 186.910 127.420 187.010 ;
        RECT 127.235 186.885 127.420 186.910 ;
        RECT 126.805 186.290 127.065 186.740 ;
        RECT 127.235 186.640 127.565 186.885 ;
        RECT 127.735 186.565 128.490 186.815 ;
        RECT 128.660 186.695 128.935 187.395 ;
        RECT 127.720 186.530 128.490 186.565 ;
        RECT 127.705 186.520 128.490 186.530 ;
        RECT 127.700 186.505 128.595 186.520 ;
        RECT 127.680 186.490 128.595 186.505 ;
        RECT 127.660 186.480 128.595 186.490 ;
        RECT 127.635 186.470 128.595 186.480 ;
        RECT 127.565 186.440 128.595 186.470 ;
        RECT 127.545 186.410 128.595 186.440 ;
        RECT 127.525 186.380 128.595 186.410 ;
        RECT 127.495 186.355 128.595 186.380 ;
        RECT 127.460 186.320 128.595 186.355 ;
        RECT 127.430 186.315 128.595 186.320 ;
        RECT 127.430 186.310 127.820 186.315 ;
        RECT 127.430 186.300 127.795 186.310 ;
        RECT 127.430 186.295 127.780 186.300 ;
        RECT 127.430 186.290 127.765 186.295 ;
        RECT 126.805 186.285 127.765 186.290 ;
        RECT 126.805 186.275 127.755 186.285 ;
        RECT 126.805 186.270 127.745 186.275 ;
        RECT 126.805 186.260 127.735 186.270 ;
        RECT 126.805 186.250 127.730 186.260 ;
        RECT 126.805 186.245 127.725 186.250 ;
        RECT 126.805 186.230 127.715 186.245 ;
        RECT 126.805 186.215 127.710 186.230 ;
        RECT 126.805 186.190 127.700 186.215 ;
        RECT 126.805 186.120 127.695 186.190 ;
        RECT 122.835 185.185 123.330 185.515 ;
        RECT 123.750 185.015 123.990 185.525 ;
        RECT 124.170 185.195 124.450 185.525 ;
        RECT 124.680 185.015 124.895 185.525 ;
        RECT 125.065 185.185 125.680 185.755 ;
        RECT 126.345 185.015 126.635 185.740 ;
        RECT 126.805 185.565 127.355 185.950 ;
        RECT 127.525 185.395 127.695 186.120 ;
        RECT 126.805 185.225 127.695 185.395 ;
        RECT 127.865 185.720 128.195 186.145 ;
        RECT 128.365 185.920 128.595 186.315 ;
        RECT 127.865 185.235 128.085 185.720 ;
        RECT 128.765 185.665 128.935 186.695 ;
        RECT 128.255 185.015 128.505 185.555 ;
        RECT 128.675 185.185 128.935 185.665 ;
        RECT 129.105 186.845 129.565 187.395 ;
        RECT 129.755 186.845 130.085 187.565 ;
        RECT 129.105 185.475 129.355 186.845 ;
        RECT 130.285 186.675 130.585 187.225 ;
        RECT 130.755 186.895 131.035 187.565 ;
        RECT 131.405 187.010 132.010 187.565 ;
        RECT 132.185 187.055 132.665 187.395 ;
        RECT 132.835 187.020 133.090 187.565 ;
        RECT 131.405 186.910 132.020 187.010 ;
        RECT 131.835 186.885 132.020 186.910 ;
        RECT 129.645 186.505 130.585 186.675 ;
        RECT 129.645 186.255 129.815 186.505 ;
        RECT 130.955 186.255 131.220 186.615 ;
        RECT 129.525 185.925 129.815 186.255 ;
        RECT 129.985 186.005 130.325 186.255 ;
        RECT 130.545 186.005 131.220 186.255 ;
        RECT 131.405 186.290 131.665 186.740 ;
        RECT 131.835 186.640 132.165 186.885 ;
        RECT 132.335 186.565 133.090 186.815 ;
        RECT 133.260 186.695 133.535 187.395 ;
        RECT 132.320 186.530 133.090 186.565 ;
        RECT 132.305 186.520 133.090 186.530 ;
        RECT 132.300 186.505 133.195 186.520 ;
        RECT 132.280 186.490 133.195 186.505 ;
        RECT 132.260 186.480 133.195 186.490 ;
        RECT 132.235 186.470 133.195 186.480 ;
        RECT 132.165 186.440 133.195 186.470 ;
        RECT 132.145 186.410 133.195 186.440 ;
        RECT 132.125 186.380 133.195 186.410 ;
        RECT 132.095 186.355 133.195 186.380 ;
        RECT 132.060 186.320 133.195 186.355 ;
        RECT 132.030 186.315 133.195 186.320 ;
        RECT 132.030 186.310 132.420 186.315 ;
        RECT 132.030 186.300 132.395 186.310 ;
        RECT 132.030 186.295 132.380 186.300 ;
        RECT 132.030 186.290 132.365 186.295 ;
        RECT 131.405 186.285 132.365 186.290 ;
        RECT 131.405 186.275 132.355 186.285 ;
        RECT 131.405 186.270 132.345 186.275 ;
        RECT 131.405 186.260 132.335 186.270 ;
        RECT 131.405 186.250 132.330 186.260 ;
        RECT 131.405 186.245 132.325 186.250 ;
        RECT 131.405 186.230 132.315 186.245 ;
        RECT 131.405 186.215 132.310 186.230 ;
        RECT 131.405 186.190 132.300 186.215 ;
        RECT 131.405 186.120 132.295 186.190 ;
        RECT 129.645 185.835 129.815 185.925 ;
        RECT 129.645 185.645 131.035 185.835 ;
        RECT 129.105 185.185 129.665 185.475 ;
        RECT 129.835 185.015 130.085 185.475 ;
        RECT 130.705 185.285 131.035 185.645 ;
        RECT 131.405 185.565 131.955 185.950 ;
        RECT 132.125 185.395 132.295 186.120 ;
        RECT 131.405 185.225 132.295 185.395 ;
        RECT 132.465 185.720 132.795 186.145 ;
        RECT 132.965 185.920 133.195 186.315 ;
        RECT 132.465 185.235 132.685 185.720 ;
        RECT 133.365 185.665 133.535 186.695 ;
        RECT 133.785 186.635 133.965 187.395 ;
        RECT 134.145 186.805 134.475 187.565 ;
        RECT 133.785 186.465 134.460 186.635 ;
        RECT 134.645 186.490 134.915 187.395 ;
        RECT 134.290 186.320 134.460 186.465 ;
        RECT 133.725 185.915 134.065 186.285 ;
        RECT 134.290 185.990 134.565 186.320 ;
        RECT 134.290 185.735 134.460 185.990 ;
        RECT 132.855 185.015 133.105 185.555 ;
        RECT 133.275 185.185 133.535 185.665 ;
        RECT 133.795 185.565 134.460 185.735 ;
        RECT 134.735 185.690 134.915 186.490 ;
        RECT 135.085 186.475 136.755 187.565 ;
        RECT 133.795 185.185 133.965 185.565 ;
        RECT 134.145 185.015 134.475 185.395 ;
        RECT 134.655 185.185 134.915 185.690 ;
        RECT 135.085 185.785 135.835 186.305 ;
        RECT 136.005 185.955 136.755 186.475 ;
        RECT 136.925 186.385 137.450 187.395 ;
        RECT 137.685 186.845 138.015 187.565 ;
        RECT 138.185 186.675 138.435 187.395 ;
        RECT 137.685 186.385 138.435 186.675 ;
        RECT 136.925 185.815 137.195 186.385 ;
        RECT 137.685 186.215 137.945 186.385 ;
        RECT 137.365 186.005 137.945 186.215 ;
        RECT 138.115 186.005 138.535 186.215 ;
        RECT 138.705 186.005 139.035 187.320 ;
        RECT 139.245 186.005 139.575 187.320 ;
        RECT 139.745 186.005 140.115 187.320 ;
        RECT 140.445 186.445 140.775 187.565 ;
        RECT 141.185 186.445 141.515 187.565 ;
        RECT 140.325 186.005 140.835 186.255 ;
        RECT 141.125 186.005 141.635 186.255 ;
        RECT 141.845 186.005 142.215 187.320 ;
        RECT 142.385 186.005 142.715 187.320 ;
        RECT 142.925 186.005 143.255 187.320 ;
        RECT 143.525 186.675 143.775 187.395 ;
        RECT 143.945 186.845 144.275 187.565 ;
        RECT 143.525 186.385 144.275 186.675 ;
        RECT 144.510 186.385 145.035 187.395 ;
        RECT 144.015 186.215 144.275 186.385 ;
        RECT 143.425 186.005 143.845 186.215 ;
        RECT 144.015 186.005 144.595 186.215 ;
        RECT 137.575 185.835 137.945 186.005 ;
        RECT 144.015 185.835 144.385 186.005 ;
        RECT 135.085 185.015 136.755 185.785 ;
        RECT 136.925 185.185 137.265 185.815 ;
        RECT 137.575 185.645 138.325 185.835 ;
        RECT 137.555 185.015 137.725 185.475 ;
        RECT 137.995 185.200 138.325 185.645 ;
        RECT 138.495 185.665 140.795 185.835 ;
        RECT 138.495 185.345 138.665 185.665 ;
        RECT 138.890 185.015 139.220 185.475 ;
        RECT 139.420 185.185 139.750 185.665 ;
        RECT 139.965 185.015 140.295 185.475 ;
        RECT 140.465 185.185 140.795 185.665 ;
        RECT 141.165 185.665 143.465 185.835 ;
        RECT 141.165 185.185 141.495 185.665 ;
        RECT 141.665 185.015 141.995 185.475 ;
        RECT 142.210 185.185 142.540 185.665 ;
        RECT 142.740 185.015 143.070 185.475 ;
        RECT 143.295 185.345 143.465 185.665 ;
        RECT 143.635 185.645 144.385 185.835 ;
        RECT 144.765 185.815 145.035 186.385 ;
        RECT 143.635 185.200 143.965 185.645 ;
        RECT 144.235 185.015 144.405 185.475 ;
        RECT 144.695 185.185 145.035 185.815 ;
        RECT 145.205 186.695 145.480 187.395 ;
        RECT 145.650 187.020 145.905 187.565 ;
        RECT 146.075 187.055 146.555 187.395 ;
        RECT 146.730 187.010 147.335 187.565 ;
        RECT 146.720 186.910 147.335 187.010 ;
        RECT 146.720 186.885 146.905 186.910 ;
        RECT 145.205 185.665 145.375 186.695 ;
        RECT 145.650 186.565 146.405 186.815 ;
        RECT 146.575 186.640 146.905 186.885 ;
        RECT 145.650 186.530 146.420 186.565 ;
        RECT 145.650 186.520 146.435 186.530 ;
        RECT 145.545 186.505 146.440 186.520 ;
        RECT 145.545 186.490 146.460 186.505 ;
        RECT 145.545 186.480 146.480 186.490 ;
        RECT 145.545 186.470 146.505 186.480 ;
        RECT 145.545 186.440 146.575 186.470 ;
        RECT 145.545 186.410 146.595 186.440 ;
        RECT 145.545 186.380 146.615 186.410 ;
        RECT 145.545 186.355 146.645 186.380 ;
        RECT 145.545 186.320 146.680 186.355 ;
        RECT 145.545 186.315 146.710 186.320 ;
        RECT 145.545 185.920 145.775 186.315 ;
        RECT 146.320 186.310 146.710 186.315 ;
        RECT 146.345 186.300 146.710 186.310 ;
        RECT 146.360 186.295 146.710 186.300 ;
        RECT 146.375 186.290 146.710 186.295 ;
        RECT 147.075 186.290 147.335 186.740 ;
        RECT 147.505 186.475 148.715 187.565 ;
        RECT 146.375 186.285 147.335 186.290 ;
        RECT 146.385 186.275 147.335 186.285 ;
        RECT 146.395 186.270 147.335 186.275 ;
        RECT 146.405 186.260 147.335 186.270 ;
        RECT 146.410 186.250 147.335 186.260 ;
        RECT 146.415 186.245 147.335 186.250 ;
        RECT 146.425 186.230 147.335 186.245 ;
        RECT 146.430 186.215 147.335 186.230 ;
        RECT 146.440 186.190 147.335 186.215 ;
        RECT 145.945 185.720 146.275 186.145 ;
        RECT 145.205 185.185 145.465 185.665 ;
        RECT 145.635 185.015 145.885 185.555 ;
        RECT 146.055 185.235 146.275 185.720 ;
        RECT 146.445 186.120 147.335 186.190 ;
        RECT 146.445 185.395 146.615 186.120 ;
        RECT 146.785 185.565 147.335 185.950 ;
        RECT 147.505 185.765 148.025 186.305 ;
        RECT 148.195 185.935 148.715 186.475 ;
        RECT 148.885 186.475 150.095 187.565 ;
        RECT 148.885 185.935 149.405 186.475 ;
        RECT 149.575 185.765 150.095 186.305 ;
        RECT 146.445 185.225 147.335 185.395 ;
        RECT 147.505 185.015 148.715 185.765 ;
        RECT 148.885 185.015 150.095 185.765 ;
        RECT 36.100 184.845 150.180 185.015 ;
        RECT 36.185 184.095 37.395 184.845 ;
        RECT 37.565 184.300 42.910 184.845 ;
        RECT 43.090 184.355 43.345 184.845 ;
        RECT 43.515 184.335 44.745 184.675 ;
        RECT 45.090 184.335 45.330 184.845 ;
        RECT 45.510 184.335 45.790 184.665 ;
        RECT 46.020 184.335 46.235 184.845 ;
        RECT 36.185 183.555 36.705 184.095 ;
        RECT 36.875 183.385 37.395 183.925 ;
        RECT 39.150 183.470 39.490 184.300 ;
        RECT 36.185 182.295 37.395 183.385 ;
        RECT 40.970 182.730 41.320 183.980 ;
        RECT 43.110 183.605 43.330 184.185 ;
        RECT 43.515 183.435 43.695 184.335 ;
        RECT 43.865 183.605 44.240 184.165 ;
        RECT 44.415 184.105 44.745 184.335 ;
        RECT 44.445 183.605 44.755 183.935 ;
        RECT 44.985 183.605 45.340 184.165 ;
        RECT 45.510 183.435 45.680 184.335 ;
        RECT 45.850 183.605 46.115 184.165 ;
        RECT 46.405 184.105 47.020 184.675 ;
        RECT 46.365 183.435 46.535 183.935 ;
        RECT 37.565 182.295 42.910 182.730 ;
        RECT 43.090 182.295 43.345 183.435 ;
        RECT 43.515 183.265 44.745 183.435 ;
        RECT 43.515 182.465 43.845 183.265 ;
        RECT 44.015 182.295 44.245 183.095 ;
        RECT 44.415 182.465 44.745 183.265 ;
        RECT 45.110 183.265 46.535 183.435 ;
        RECT 45.110 183.090 45.500 183.265 ;
        RECT 45.985 182.295 46.315 183.095 ;
        RECT 46.705 183.085 47.020 184.105 ;
        RECT 46.485 182.465 47.020 183.085 ;
        RECT 47.225 184.170 47.495 184.515 ;
        RECT 47.685 184.445 48.065 184.845 ;
        RECT 48.235 184.275 48.405 184.625 ;
        RECT 48.575 184.445 48.905 184.845 ;
        RECT 49.105 184.275 49.275 184.625 ;
        RECT 49.475 184.345 49.805 184.845 ;
        RECT 47.225 183.435 47.395 184.170 ;
        RECT 47.665 184.105 49.275 184.275 ;
        RECT 50.920 184.275 51.175 184.625 ;
        RECT 51.345 184.445 51.675 184.845 ;
        RECT 51.845 184.275 52.015 184.625 ;
        RECT 52.185 184.445 52.565 184.845 ;
        RECT 47.665 183.935 47.835 184.105 ;
        RECT 47.565 183.605 47.835 183.935 ;
        RECT 48.005 183.605 48.410 183.935 ;
        RECT 47.665 183.435 47.835 183.605 ;
        RECT 47.225 182.465 47.495 183.435 ;
        RECT 47.665 183.265 48.390 183.435 ;
        RECT 48.580 183.315 49.290 183.935 ;
        RECT 49.460 183.605 49.810 184.175 ;
        RECT 50.920 184.105 52.585 184.275 ;
        RECT 52.755 184.170 53.030 184.515 ;
        RECT 52.415 183.935 52.585 184.105 ;
        RECT 50.905 183.605 51.250 183.935 ;
        RECT 51.420 183.605 52.245 183.935 ;
        RECT 52.415 183.605 52.690 183.935 ;
        RECT 48.220 183.145 48.390 183.265 ;
        RECT 49.490 183.145 49.810 183.435 ;
        RECT 47.705 182.295 47.985 183.095 ;
        RECT 48.220 182.975 49.810 183.145 ;
        RECT 50.925 183.145 51.250 183.435 ;
        RECT 51.420 183.315 51.615 183.605 ;
        RECT 52.415 183.435 52.585 183.605 ;
        RECT 52.860 183.435 53.030 184.170 ;
        RECT 53.220 184.275 53.475 184.625 ;
        RECT 53.645 184.445 53.975 184.845 ;
        RECT 54.145 184.275 54.315 184.625 ;
        RECT 54.485 184.445 54.865 184.845 ;
        RECT 53.220 184.105 54.885 184.275 ;
        RECT 55.055 184.170 55.330 184.515 ;
        RECT 54.715 183.935 54.885 184.105 ;
        RECT 53.205 183.605 53.550 183.935 ;
        RECT 53.720 183.605 54.545 183.935 ;
        RECT 54.715 183.605 54.990 183.935 ;
        RECT 51.925 183.265 52.585 183.435 ;
        RECT 51.925 183.145 52.095 183.265 ;
        RECT 50.925 182.975 52.095 183.145 ;
        RECT 48.155 182.515 49.810 182.805 ;
        RECT 50.905 182.515 52.095 182.805 ;
        RECT 52.265 182.295 52.545 183.095 ;
        RECT 52.755 182.465 53.030 183.435 ;
        RECT 53.225 183.145 53.550 183.435 ;
        RECT 53.720 183.315 53.915 183.605 ;
        RECT 54.715 183.435 54.885 183.605 ;
        RECT 55.160 183.435 55.330 184.170 ;
        RECT 55.505 184.075 58.095 184.845 ;
        RECT 58.430 184.335 58.670 184.845 ;
        RECT 58.850 184.335 59.130 184.665 ;
        RECT 59.360 184.335 59.575 184.845 ;
        RECT 55.505 183.555 56.715 184.075 ;
        RECT 54.225 183.265 54.885 183.435 ;
        RECT 54.225 183.145 54.395 183.265 ;
        RECT 53.225 182.975 54.395 183.145 ;
        RECT 53.205 182.515 54.395 182.805 ;
        RECT 54.565 182.295 54.845 183.095 ;
        RECT 55.055 182.465 55.330 183.435 ;
        RECT 56.885 183.385 58.095 183.905 ;
        RECT 58.325 183.605 58.680 184.165 ;
        RECT 58.850 183.435 59.020 184.335 ;
        RECT 59.190 183.605 59.455 184.165 ;
        RECT 59.745 184.105 60.360 184.675 ;
        RECT 59.705 183.435 59.875 183.935 ;
        RECT 55.505 182.295 58.095 183.385 ;
        RECT 58.450 183.265 59.875 183.435 ;
        RECT 58.450 183.090 58.840 183.265 ;
        RECT 59.325 182.295 59.655 183.095 ;
        RECT 60.045 183.085 60.360 184.105 ;
        RECT 60.565 184.095 61.775 184.845 ;
        RECT 61.945 184.120 62.235 184.845 ;
        RECT 63.325 184.170 63.585 184.675 ;
        RECT 63.765 184.465 64.095 184.845 ;
        RECT 64.275 184.295 64.445 184.675 ;
        RECT 64.705 184.300 70.050 184.845 ;
        RECT 70.225 184.300 75.570 184.845 ;
        RECT 60.565 183.555 61.085 184.095 ;
        RECT 61.255 183.385 61.775 183.925 ;
        RECT 59.825 182.465 60.360 183.085 ;
        RECT 60.565 182.295 61.775 183.385 ;
        RECT 61.945 182.295 62.235 183.460 ;
        RECT 63.325 183.370 63.505 184.170 ;
        RECT 63.780 184.125 64.445 184.295 ;
        RECT 63.780 183.870 63.950 184.125 ;
        RECT 63.675 183.540 63.950 183.870 ;
        RECT 64.175 183.575 64.515 183.945 ;
        RECT 63.780 183.395 63.950 183.540 ;
        RECT 66.290 183.470 66.630 184.300 ;
        RECT 63.325 182.465 63.595 183.370 ;
        RECT 63.780 183.225 64.455 183.395 ;
        RECT 63.765 182.295 64.095 183.055 ;
        RECT 64.275 182.465 64.455 183.225 ;
        RECT 68.110 182.730 68.460 183.980 ;
        RECT 71.810 183.470 72.150 184.300 ;
        RECT 75.745 184.075 77.415 184.845 ;
        RECT 77.675 184.295 77.845 184.675 ;
        RECT 78.025 184.465 78.355 184.845 ;
        RECT 77.675 184.125 78.340 184.295 ;
        RECT 78.535 184.170 78.795 184.675 ;
        RECT 73.630 182.730 73.980 183.980 ;
        RECT 75.745 183.555 76.495 184.075 ;
        RECT 76.665 183.385 77.415 183.905 ;
        RECT 77.605 183.575 77.945 183.945 ;
        RECT 78.170 183.870 78.340 184.125 ;
        RECT 78.170 183.540 78.445 183.870 ;
        RECT 78.170 183.395 78.340 183.540 ;
        RECT 64.705 182.295 70.050 182.730 ;
        RECT 70.225 182.295 75.570 182.730 ;
        RECT 75.745 182.295 77.415 183.385 ;
        RECT 77.665 183.225 78.340 183.395 ;
        RECT 78.615 183.370 78.795 184.170 ;
        RECT 77.665 182.465 77.845 183.225 ;
        RECT 78.025 182.295 78.355 183.055 ;
        RECT 78.525 182.465 78.795 183.370 ;
        RECT 78.975 182.475 79.235 184.665 ;
        RECT 79.495 184.475 80.165 184.845 ;
        RECT 80.345 184.295 80.655 184.665 ;
        RECT 79.425 184.095 80.655 184.295 ;
        RECT 79.425 183.425 79.715 184.095 ;
        RECT 80.835 183.915 81.065 184.555 ;
        RECT 81.245 184.115 81.535 184.845 ;
        RECT 81.725 184.385 82.285 184.675 ;
        RECT 82.455 184.385 82.705 184.845 ;
        RECT 79.895 183.605 80.360 183.915 ;
        RECT 80.540 183.605 81.065 183.915 ;
        RECT 81.245 183.605 81.545 183.935 ;
        RECT 79.425 183.205 80.195 183.425 ;
        RECT 79.405 182.295 79.745 183.025 ;
        RECT 79.925 182.475 80.195 183.205 ;
        RECT 80.375 183.185 81.535 183.425 ;
        RECT 80.375 182.475 80.605 183.185 ;
        RECT 80.775 182.295 81.105 183.005 ;
        RECT 81.275 182.475 81.535 183.185 ;
        RECT 81.725 183.015 81.975 184.385 ;
        RECT 83.325 184.215 83.655 184.575 ;
        RECT 82.265 184.025 83.655 184.215 ;
        RECT 84.085 184.025 84.295 184.845 ;
        RECT 84.465 184.045 84.795 184.675 ;
        RECT 82.265 183.935 82.435 184.025 ;
        RECT 82.145 183.605 82.435 183.935 ;
        RECT 82.605 183.605 82.945 183.855 ;
        RECT 83.165 183.605 83.840 183.855 ;
        RECT 82.265 183.355 82.435 183.605 ;
        RECT 82.265 183.185 83.205 183.355 ;
        RECT 83.575 183.245 83.840 183.605 ;
        RECT 84.465 183.445 84.715 184.045 ;
        RECT 84.965 184.025 85.195 184.845 ;
        RECT 85.405 184.075 87.075 184.845 ;
        RECT 87.705 184.120 87.995 184.845 ;
        RECT 84.885 183.605 85.215 183.855 ;
        RECT 85.405 183.555 86.155 184.075 ;
        RECT 88.370 184.065 88.870 184.675 ;
        RECT 81.725 182.465 82.185 183.015 ;
        RECT 82.375 182.295 82.705 183.015 ;
        RECT 82.905 182.635 83.205 183.185 ;
        RECT 83.375 182.295 83.655 182.965 ;
        RECT 84.085 182.295 84.295 183.435 ;
        RECT 84.465 182.465 84.795 183.445 ;
        RECT 84.965 182.295 85.195 183.435 ;
        RECT 86.325 183.385 87.075 183.905 ;
        RECT 88.165 183.605 88.515 183.855 ;
        RECT 85.405 182.295 87.075 183.385 ;
        RECT 87.705 182.295 87.995 183.460 ;
        RECT 88.700 183.435 88.870 184.065 ;
        RECT 89.500 184.195 89.830 184.675 ;
        RECT 90.000 184.385 90.225 184.845 ;
        RECT 90.395 184.195 90.725 184.675 ;
        RECT 89.500 184.025 90.725 184.195 ;
        RECT 90.915 184.045 91.165 184.845 ;
        RECT 91.335 184.045 91.675 184.675 ;
        RECT 89.040 183.655 89.370 183.855 ;
        RECT 89.540 183.655 89.870 183.855 ;
        RECT 90.040 183.655 90.460 183.855 ;
        RECT 90.635 183.685 91.330 183.855 ;
        RECT 90.635 183.435 90.805 183.685 ;
        RECT 91.500 183.435 91.675 184.045 ;
        RECT 88.370 183.265 90.805 183.435 ;
        RECT 88.370 182.465 88.700 183.265 ;
        RECT 88.870 182.295 89.200 183.095 ;
        RECT 89.500 182.465 89.830 183.265 ;
        RECT 90.475 182.295 90.725 183.095 ;
        RECT 90.995 182.295 91.165 183.435 ;
        RECT 91.335 182.465 91.675 183.435 ;
        RECT 91.845 182.465 92.125 184.565 ;
        RECT 92.355 184.385 92.525 184.845 ;
        RECT 92.795 184.455 94.045 184.635 ;
        RECT 93.180 184.215 93.545 184.285 ;
        RECT 92.295 184.035 93.545 184.215 ;
        RECT 93.715 184.235 94.045 184.455 ;
        RECT 94.215 184.405 94.385 184.845 ;
        RECT 94.555 184.235 94.895 184.650 ;
        RECT 93.715 184.065 94.895 184.235 ;
        RECT 95.065 184.170 95.325 184.675 ;
        RECT 95.505 184.465 95.835 184.845 ;
        RECT 96.015 184.295 96.185 184.675 ;
        RECT 92.295 183.435 92.570 184.035 ;
        RECT 92.740 183.605 93.095 183.855 ;
        RECT 93.290 183.825 93.755 183.855 ;
        RECT 93.285 183.655 93.755 183.825 ;
        RECT 93.290 183.605 93.755 183.655 ;
        RECT 93.925 183.605 94.255 183.855 ;
        RECT 94.430 183.655 94.895 183.855 ;
        RECT 94.075 183.485 94.255 183.605 ;
        RECT 92.295 183.225 93.905 183.435 ;
        RECT 94.075 183.315 94.405 183.485 ;
        RECT 93.495 183.125 93.905 183.225 ;
        RECT 92.315 182.295 93.100 183.055 ;
        RECT 93.495 182.465 93.880 183.125 ;
        RECT 94.205 182.525 94.405 183.315 ;
        RECT 94.575 182.295 94.895 183.475 ;
        RECT 95.065 183.370 95.245 184.170 ;
        RECT 95.520 184.125 96.185 184.295 ;
        RECT 96.605 184.285 96.935 184.675 ;
        RECT 97.105 184.455 98.290 184.625 ;
        RECT 98.550 184.375 98.720 184.845 ;
        RECT 95.520 183.870 95.690 184.125 ;
        RECT 96.605 184.105 97.115 184.285 ;
        RECT 95.415 183.540 95.690 183.870 ;
        RECT 95.915 183.575 96.255 183.945 ;
        RECT 96.445 183.645 96.775 183.935 ;
        RECT 95.520 183.395 95.690 183.540 ;
        RECT 96.945 183.475 97.115 184.105 ;
        RECT 97.520 184.195 97.905 184.285 ;
        RECT 98.890 184.195 99.220 184.660 ;
        RECT 97.520 184.025 99.220 184.195 ;
        RECT 99.390 184.025 99.560 184.845 ;
        RECT 99.730 184.025 100.415 184.665 ;
        RECT 97.285 183.645 97.615 183.855 ;
        RECT 97.795 183.605 98.175 183.855 ;
        RECT 95.065 182.465 95.335 183.370 ;
        RECT 95.520 183.225 96.195 183.395 ;
        RECT 95.505 182.295 95.835 183.055 ;
        RECT 96.015 182.465 96.195 183.225 ;
        RECT 96.600 183.305 97.685 183.475 ;
        RECT 96.600 182.465 96.900 183.305 ;
        RECT 97.095 182.295 97.345 183.135 ;
        RECT 97.515 183.055 97.685 183.305 ;
        RECT 97.855 183.225 98.175 183.605 ;
        RECT 98.365 183.645 98.850 183.855 ;
        RECT 99.040 183.645 99.490 183.855 ;
        RECT 99.660 183.645 99.995 183.855 ;
        RECT 98.365 183.485 98.740 183.645 ;
        RECT 98.345 183.315 98.740 183.485 ;
        RECT 99.660 183.475 99.830 183.645 ;
        RECT 98.365 183.225 98.740 183.315 ;
        RECT 98.910 183.305 99.830 183.475 ;
        RECT 98.910 183.055 99.080 183.305 ;
        RECT 97.515 182.885 99.080 183.055 ;
        RECT 97.935 182.465 98.740 182.885 ;
        RECT 99.250 182.295 99.580 183.135 ;
        RECT 100.165 183.055 100.415 184.025 ;
        RECT 99.750 182.465 100.415 183.055 ;
        RECT 100.585 184.025 101.270 184.665 ;
        RECT 101.440 184.025 101.610 184.845 ;
        RECT 101.780 184.195 102.110 184.660 ;
        RECT 102.280 184.375 102.450 184.845 ;
        RECT 102.710 184.455 103.895 184.625 ;
        RECT 104.065 184.285 104.395 184.675 ;
        RECT 103.095 184.195 103.480 184.285 ;
        RECT 101.780 184.025 103.480 184.195 ;
        RECT 103.885 184.105 104.395 184.285 ;
        RECT 104.725 184.170 104.985 184.675 ;
        RECT 105.165 184.465 105.495 184.845 ;
        RECT 105.675 184.295 105.845 184.675 ;
        RECT 100.585 183.055 100.835 184.025 ;
        RECT 101.005 183.645 101.340 183.855 ;
        RECT 101.510 183.645 101.960 183.855 ;
        RECT 102.150 183.645 102.635 183.855 ;
        RECT 101.170 183.475 101.340 183.645 ;
        RECT 101.170 183.305 102.090 183.475 ;
        RECT 100.585 182.465 101.250 183.055 ;
        RECT 101.420 182.295 101.750 183.135 ;
        RECT 101.920 183.055 102.090 183.305 ;
        RECT 102.260 183.225 102.635 183.645 ;
        RECT 102.825 183.605 103.205 183.855 ;
        RECT 103.385 183.645 103.715 183.855 ;
        RECT 102.825 183.225 103.145 183.605 ;
        RECT 103.885 183.475 104.055 184.105 ;
        RECT 104.225 183.645 104.555 183.935 ;
        RECT 103.315 183.305 104.400 183.475 ;
        RECT 103.315 183.055 103.485 183.305 ;
        RECT 101.920 182.885 103.485 183.055 ;
        RECT 102.260 182.465 103.065 182.885 ;
        RECT 103.655 182.295 103.905 183.135 ;
        RECT 104.100 182.465 104.400 183.305 ;
        RECT 104.725 183.370 104.905 184.170 ;
        RECT 105.180 184.125 105.845 184.295 ;
        RECT 105.180 183.870 105.350 184.125 ;
        RECT 107.025 184.045 107.335 184.845 ;
        RECT 107.540 184.045 108.235 184.675 ;
        RECT 108.405 184.275 108.840 184.675 ;
        RECT 109.010 184.445 109.395 184.845 ;
        RECT 108.405 184.105 109.395 184.275 ;
        RECT 109.565 184.105 109.990 184.675 ;
        RECT 110.180 184.275 110.435 184.675 ;
        RECT 110.605 184.445 110.990 184.845 ;
        RECT 110.180 184.105 110.990 184.275 ;
        RECT 111.160 184.105 111.405 184.675 ;
        RECT 111.595 184.275 111.850 184.675 ;
        RECT 112.020 184.445 112.405 184.845 ;
        RECT 111.595 184.105 112.405 184.275 ;
        RECT 112.575 184.105 112.835 184.675 ;
        RECT 113.465 184.120 113.755 184.845 ;
        RECT 113.925 184.345 114.185 184.675 ;
        RECT 114.395 184.365 114.670 184.845 ;
        RECT 105.075 183.540 105.350 183.870 ;
        RECT 105.575 183.575 105.915 183.945 ;
        RECT 107.035 183.605 107.370 183.875 ;
        RECT 105.180 183.395 105.350 183.540 ;
        RECT 107.540 183.445 107.710 184.045 ;
        RECT 109.060 183.935 109.395 184.105 ;
        RECT 109.640 183.935 109.990 184.105 ;
        RECT 110.640 183.935 110.990 184.105 ;
        RECT 111.235 183.935 111.405 184.105 ;
        RECT 112.055 183.935 112.405 184.105 ;
        RECT 107.880 183.605 108.215 183.855 ;
        RECT 104.725 182.465 104.995 183.370 ;
        RECT 105.180 183.225 105.855 183.395 ;
        RECT 105.165 182.295 105.495 183.055 ;
        RECT 105.675 182.465 105.855 183.225 ;
        RECT 107.025 182.295 107.305 183.435 ;
        RECT 107.475 182.465 107.805 183.445 ;
        RECT 107.975 182.295 108.235 183.435 ;
        RECT 108.405 183.230 108.890 183.935 ;
        RECT 109.060 183.605 109.470 183.935 ;
        RECT 109.060 183.060 109.395 183.605 ;
        RECT 109.640 183.435 110.470 183.935 ;
        RECT 108.405 182.890 109.395 183.060 ;
        RECT 109.565 183.255 110.470 183.435 ;
        RECT 110.640 183.605 111.065 183.935 ;
        RECT 108.405 182.465 108.840 182.890 ;
        RECT 109.010 182.295 109.395 182.720 ;
        RECT 109.565 182.465 109.990 183.255 ;
        RECT 110.640 183.085 110.990 183.605 ;
        RECT 111.235 183.435 111.885 183.935 ;
        RECT 110.160 182.890 110.990 183.085 ;
        RECT 111.160 183.255 111.885 183.435 ;
        RECT 112.055 183.605 112.480 183.935 ;
        RECT 110.160 182.465 110.435 182.890 ;
        RECT 110.605 182.295 110.990 182.720 ;
        RECT 111.160 182.465 111.405 183.255 ;
        RECT 112.055 183.085 112.405 183.605 ;
        RECT 112.650 183.435 112.835 184.105 ;
        RECT 111.595 182.890 112.405 183.085 ;
        RECT 111.595 182.465 111.850 182.890 ;
        RECT 112.020 182.295 112.405 182.720 ;
        RECT 112.575 182.465 112.835 183.435 ;
        RECT 113.465 182.295 113.755 183.460 ;
        RECT 113.925 183.435 114.095 184.345 ;
        RECT 114.880 184.275 115.085 184.675 ;
        RECT 115.255 184.445 115.590 184.845 ;
        RECT 114.265 183.605 114.625 184.185 ;
        RECT 114.880 184.105 115.565 184.275 ;
        RECT 114.805 183.435 115.055 183.935 ;
        RECT 113.925 183.265 115.055 183.435 ;
        RECT 113.925 182.495 114.195 183.265 ;
        RECT 115.225 183.075 115.565 184.105 ;
        RECT 115.765 184.095 116.975 184.845 ;
        RECT 117.235 184.295 117.405 184.675 ;
        RECT 117.585 184.465 117.915 184.845 ;
        RECT 117.235 184.125 117.900 184.295 ;
        RECT 118.095 184.170 118.355 184.675 ;
        RECT 115.765 183.555 116.285 184.095 ;
        RECT 116.455 183.385 116.975 183.925 ;
        RECT 117.165 183.575 117.505 183.945 ;
        RECT 117.730 183.870 117.900 184.125 ;
        RECT 117.730 183.540 118.005 183.870 ;
        RECT 117.730 183.395 117.900 183.540 ;
        RECT 114.365 182.295 114.695 183.075 ;
        RECT 114.900 182.900 115.565 183.075 ;
        RECT 114.900 182.495 115.085 182.900 ;
        RECT 115.255 182.295 115.590 182.720 ;
        RECT 115.765 182.295 116.975 183.385 ;
        RECT 117.225 183.225 117.900 183.395 ;
        RECT 118.175 183.370 118.355 184.170 ;
        RECT 118.525 184.025 118.785 184.845 ;
        RECT 118.955 184.025 119.285 184.445 ;
        RECT 119.465 184.275 119.725 184.675 ;
        RECT 119.895 184.445 120.225 184.845 ;
        RECT 120.395 184.275 120.565 184.625 ;
        RECT 120.735 184.445 121.110 184.845 ;
        RECT 119.465 184.105 121.130 184.275 ;
        RECT 121.300 184.170 121.575 184.515 ;
        RECT 121.745 184.465 122.635 184.635 ;
        RECT 119.035 183.935 119.285 184.025 ;
        RECT 120.960 183.935 121.130 184.105 ;
        RECT 118.530 183.605 118.865 183.855 ;
        RECT 119.035 183.605 119.750 183.935 ;
        RECT 119.965 183.605 120.790 183.935 ;
        RECT 120.960 183.605 121.235 183.935 ;
        RECT 117.225 182.465 117.405 183.225 ;
        RECT 117.585 182.295 117.915 183.055 ;
        RECT 118.085 182.465 118.355 183.370 ;
        RECT 118.525 182.295 118.785 183.435 ;
        RECT 119.035 183.045 119.205 183.605 ;
        RECT 119.465 183.145 119.795 183.435 ;
        RECT 119.965 183.315 120.210 183.605 ;
        RECT 120.960 183.435 121.130 183.605 ;
        RECT 121.405 183.435 121.575 184.170 ;
        RECT 121.745 183.910 122.295 184.295 ;
        RECT 122.465 183.740 122.635 184.465 ;
        RECT 120.470 183.265 121.130 183.435 ;
        RECT 120.470 183.145 120.640 183.265 ;
        RECT 119.465 182.975 120.640 183.145 ;
        RECT 119.025 182.475 120.640 182.805 ;
        RECT 120.810 182.295 121.090 183.095 ;
        RECT 121.300 182.465 121.575 183.435 ;
        RECT 121.745 183.670 122.635 183.740 ;
        RECT 122.805 184.140 123.025 184.625 ;
        RECT 123.195 184.305 123.445 184.845 ;
        RECT 123.615 184.195 123.875 184.675 ;
        RECT 122.805 183.715 123.135 184.140 ;
        RECT 121.745 183.645 122.640 183.670 ;
        RECT 121.745 183.630 122.650 183.645 ;
        RECT 121.745 183.615 122.655 183.630 ;
        RECT 121.745 183.610 122.665 183.615 ;
        RECT 121.745 183.600 122.670 183.610 ;
        RECT 121.745 183.590 122.675 183.600 ;
        RECT 121.745 183.585 122.685 183.590 ;
        RECT 121.745 183.575 122.695 183.585 ;
        RECT 121.745 183.570 122.705 183.575 ;
        RECT 121.745 183.120 122.005 183.570 ;
        RECT 122.370 183.565 122.705 183.570 ;
        RECT 122.370 183.560 122.720 183.565 ;
        RECT 122.370 183.550 122.735 183.560 ;
        RECT 122.370 183.545 122.760 183.550 ;
        RECT 123.305 183.545 123.535 183.940 ;
        RECT 122.370 183.540 123.535 183.545 ;
        RECT 122.400 183.505 123.535 183.540 ;
        RECT 122.435 183.480 123.535 183.505 ;
        RECT 122.465 183.450 123.535 183.480 ;
        RECT 122.485 183.420 123.535 183.450 ;
        RECT 122.505 183.390 123.535 183.420 ;
        RECT 122.575 183.380 123.535 183.390 ;
        RECT 122.600 183.370 123.535 183.380 ;
        RECT 122.620 183.355 123.535 183.370 ;
        RECT 122.640 183.340 123.535 183.355 ;
        RECT 122.645 183.330 123.430 183.340 ;
        RECT 122.660 183.295 123.430 183.330 ;
        RECT 122.175 182.975 122.505 183.220 ;
        RECT 122.675 183.045 123.430 183.295 ;
        RECT 123.705 183.165 123.875 184.195 ;
        RECT 125.055 184.295 125.225 184.675 ;
        RECT 125.405 184.465 125.735 184.845 ;
        RECT 125.055 184.125 125.720 184.295 ;
        RECT 125.915 184.170 126.175 184.675 ;
        RECT 124.985 183.575 125.325 183.945 ;
        RECT 125.550 183.870 125.720 184.125 ;
        RECT 125.550 183.540 125.825 183.870 ;
        RECT 125.550 183.395 125.720 183.540 ;
        RECT 122.175 182.950 122.360 182.975 ;
        RECT 121.745 182.850 122.360 182.950 ;
        RECT 121.745 182.295 122.350 182.850 ;
        RECT 122.525 182.465 123.005 182.805 ;
        RECT 123.175 182.295 123.430 182.840 ;
        RECT 123.600 182.465 123.875 183.165 ;
        RECT 125.045 183.225 125.720 183.395 ;
        RECT 125.995 183.370 126.175 184.170 ;
        RECT 125.045 182.465 125.225 183.225 ;
        RECT 125.405 182.295 125.735 183.055 ;
        RECT 125.905 182.465 126.175 183.370 ;
        RECT 126.805 184.345 127.065 184.675 ;
        RECT 127.275 184.365 127.550 184.845 ;
        RECT 126.805 183.435 126.975 184.345 ;
        RECT 127.760 184.275 127.965 184.675 ;
        RECT 128.135 184.445 128.470 184.845 ;
        RECT 127.145 183.605 127.505 184.185 ;
        RECT 127.760 184.105 128.445 184.275 ;
        RECT 127.685 183.435 127.935 183.935 ;
        RECT 126.805 183.265 127.935 183.435 ;
        RECT 126.805 182.495 127.075 183.265 ;
        RECT 128.105 183.075 128.445 184.105 ;
        RECT 127.245 182.295 127.575 183.075 ;
        RECT 127.780 182.900 128.445 183.075 ;
        RECT 128.645 184.170 128.905 184.675 ;
        RECT 129.085 184.465 129.415 184.845 ;
        RECT 129.595 184.295 129.765 184.675 ;
        RECT 128.645 183.370 128.825 184.170 ;
        RECT 129.100 184.125 129.765 184.295 ;
        RECT 129.100 183.870 129.270 184.125 ;
        RECT 130.025 184.095 131.235 184.845 ;
        RECT 128.995 183.540 129.270 183.870 ;
        RECT 129.495 183.575 129.835 183.945 ;
        RECT 130.025 183.555 130.545 184.095 ;
        RECT 131.415 184.035 131.685 184.845 ;
        RECT 131.855 184.035 132.185 184.675 ;
        RECT 132.355 184.035 132.595 184.845 ;
        RECT 129.100 183.395 129.270 183.540 ;
        RECT 127.780 182.495 127.965 182.900 ;
        RECT 128.135 182.295 128.470 182.720 ;
        RECT 128.645 182.465 128.915 183.370 ;
        RECT 129.100 183.225 129.775 183.395 ;
        RECT 130.715 183.385 131.235 183.925 ;
        RECT 131.405 183.605 131.755 183.855 ;
        RECT 131.925 183.435 132.095 184.035 ;
        RECT 132.825 184.025 133.055 184.845 ;
        RECT 133.225 184.045 133.555 184.675 ;
        RECT 132.265 183.605 132.615 183.855 ;
        RECT 132.805 183.605 133.135 183.855 ;
        RECT 133.305 183.445 133.555 184.045 ;
        RECT 133.725 184.025 133.935 184.845 ;
        RECT 134.165 184.170 134.425 184.675 ;
        RECT 134.605 184.465 134.935 184.845 ;
        RECT 135.115 184.295 135.285 184.675 ;
        RECT 129.085 182.295 129.415 183.055 ;
        RECT 129.595 182.465 129.775 183.225 ;
        RECT 130.025 182.295 131.235 183.385 ;
        RECT 131.415 182.295 131.745 183.435 ;
        RECT 131.925 183.265 132.605 183.435 ;
        RECT 132.275 182.480 132.605 183.265 ;
        RECT 132.825 182.295 133.055 183.435 ;
        RECT 133.225 182.465 133.555 183.445 ;
        RECT 133.725 182.295 133.935 183.435 ;
        RECT 134.165 183.370 134.345 184.170 ;
        RECT 134.620 184.125 135.285 184.295 ;
        RECT 134.620 183.870 134.790 184.125 ;
        RECT 135.545 184.075 139.055 184.845 ;
        RECT 139.225 184.120 139.515 184.845 ;
        RECT 139.685 184.105 140.175 184.675 ;
        RECT 140.345 184.275 140.575 184.675 ;
        RECT 140.745 184.445 141.165 184.845 ;
        RECT 141.335 184.275 141.505 184.675 ;
        RECT 140.345 184.105 141.505 184.275 ;
        RECT 141.675 184.105 142.125 184.845 ;
        RECT 142.295 184.105 142.735 184.665 ;
        RECT 134.515 183.540 134.790 183.870 ;
        RECT 135.015 183.575 135.355 183.945 ;
        RECT 135.545 183.555 137.195 184.075 ;
        RECT 134.620 183.395 134.790 183.540 ;
        RECT 134.165 182.465 134.435 183.370 ;
        RECT 134.620 183.225 135.295 183.395 ;
        RECT 137.365 183.385 139.055 183.905 ;
        RECT 134.605 182.295 134.935 183.055 ;
        RECT 135.115 182.465 135.295 183.225 ;
        RECT 135.545 182.295 139.055 183.385 ;
        RECT 139.225 182.295 139.515 183.460 ;
        RECT 139.685 183.435 139.855 184.105 ;
        RECT 140.025 183.605 140.430 183.935 ;
        RECT 139.685 183.265 140.455 183.435 ;
        RECT 139.695 182.295 140.025 183.095 ;
        RECT 140.205 182.635 140.455 183.265 ;
        RECT 140.645 182.805 140.895 183.935 ;
        RECT 141.095 183.605 141.340 183.935 ;
        RECT 141.525 183.655 141.915 183.935 ;
        RECT 141.095 182.805 141.295 183.605 ;
        RECT 142.085 183.485 142.255 183.935 ;
        RECT 141.465 183.315 142.255 183.485 ;
        RECT 141.465 182.635 141.635 183.315 ;
        RECT 140.205 182.465 141.635 182.635 ;
        RECT 141.805 182.295 142.120 183.145 ;
        RECT 142.425 183.095 142.735 184.105 ;
        RECT 142.295 182.465 142.735 183.095 ;
        RECT 142.905 184.170 143.165 184.675 ;
        RECT 143.345 184.465 143.675 184.845 ;
        RECT 143.855 184.295 144.025 184.675 ;
        RECT 142.905 183.370 143.085 184.170 ;
        RECT 143.360 184.125 144.025 184.295 ;
        RECT 143.360 183.870 143.530 184.125 ;
        RECT 144.285 184.075 147.795 184.845 ;
        RECT 148.885 184.095 150.095 184.845 ;
        RECT 143.255 183.540 143.530 183.870 ;
        RECT 143.755 183.575 144.095 183.945 ;
        RECT 144.285 183.555 145.935 184.075 ;
        RECT 143.360 183.395 143.530 183.540 ;
        RECT 142.905 182.465 143.175 183.370 ;
        RECT 143.360 183.225 144.035 183.395 ;
        RECT 146.105 183.385 147.795 183.905 ;
        RECT 143.345 182.295 143.675 183.055 ;
        RECT 143.855 182.465 144.035 183.225 ;
        RECT 144.285 182.295 147.795 183.385 ;
        RECT 148.885 183.385 149.405 183.925 ;
        RECT 149.575 183.555 150.095 184.095 ;
        RECT 148.885 182.295 150.095 183.385 ;
        RECT 36.100 182.125 150.180 182.295 ;
        RECT 36.185 181.035 37.395 182.125 ;
        RECT 37.565 181.690 42.910 182.125 ;
        RECT 36.185 180.325 36.705 180.865 ;
        RECT 36.875 180.495 37.395 181.035 ;
        RECT 36.185 179.575 37.395 180.325 ;
        RECT 39.150 180.120 39.490 180.950 ;
        RECT 40.970 180.440 41.320 181.690 ;
        RECT 43.085 181.035 44.295 182.125 ;
        RECT 43.085 180.325 43.605 180.865 ;
        RECT 43.775 180.495 44.295 181.035 ;
        RECT 44.545 181.195 44.725 181.955 ;
        RECT 44.905 181.365 45.235 182.125 ;
        RECT 44.545 181.025 45.220 181.195 ;
        RECT 45.405 181.050 45.675 181.955 ;
        RECT 45.050 180.880 45.220 181.025 ;
        RECT 44.485 180.475 44.825 180.845 ;
        RECT 45.050 180.550 45.325 180.880 ;
        RECT 37.565 179.575 42.910 180.120 ;
        RECT 43.085 179.575 44.295 180.325 ;
        RECT 45.050 180.295 45.220 180.550 ;
        RECT 44.555 180.125 45.220 180.295 ;
        RECT 45.495 180.250 45.675 181.050 ;
        RECT 45.925 181.195 46.105 181.955 ;
        RECT 46.285 181.365 46.615 182.125 ;
        RECT 45.925 181.025 46.600 181.195 ;
        RECT 46.785 181.050 47.055 181.955 ;
        RECT 46.430 180.880 46.600 181.025 ;
        RECT 45.865 180.475 46.205 180.845 ;
        RECT 46.430 180.550 46.705 180.880 ;
        RECT 46.430 180.295 46.600 180.550 ;
        RECT 44.555 179.745 44.725 180.125 ;
        RECT 44.905 179.575 45.235 179.955 ;
        RECT 45.415 179.745 45.675 180.250 ;
        RECT 45.935 180.125 46.600 180.295 ;
        RECT 46.875 180.250 47.055 181.050 ;
        RECT 47.230 180.985 47.485 182.125 ;
        RECT 47.655 181.155 47.985 181.955 ;
        RECT 48.155 181.325 48.385 182.125 ;
        RECT 48.555 181.155 48.885 181.955 ;
        RECT 47.655 180.985 48.885 181.155 ;
        RECT 45.935 179.745 46.105 180.125 ;
        RECT 46.285 179.575 46.615 179.955 ;
        RECT 46.795 179.745 47.055 180.250 ;
        RECT 47.250 180.235 47.470 180.815 ;
        RECT 47.655 180.085 47.835 180.985 ;
        RECT 49.065 180.960 49.355 182.125 ;
        RECT 49.530 181.615 51.185 181.905 ;
        RECT 49.530 181.275 51.120 181.445 ;
        RECT 51.355 181.325 51.635 182.125 ;
        RECT 49.530 180.985 49.850 181.275 ;
        RECT 50.950 181.155 51.120 181.275 ;
        RECT 48.005 180.255 48.380 180.815 ;
        RECT 48.585 180.485 48.895 180.815 ;
        RECT 48.555 180.085 48.885 180.315 ;
        RECT 47.230 179.575 47.485 180.065 ;
        RECT 47.655 179.745 48.885 180.085 ;
        RECT 49.065 179.575 49.355 180.300 ;
        RECT 49.530 180.245 49.880 180.815 ;
        RECT 50.050 180.485 50.760 181.105 ;
        RECT 50.950 180.985 51.675 181.155 ;
        RECT 51.845 180.985 52.115 181.955 ;
        RECT 52.285 181.035 55.795 182.125 ;
        RECT 51.505 180.815 51.675 180.985 ;
        RECT 50.930 180.485 51.335 180.815 ;
        RECT 51.505 180.485 51.775 180.815 ;
        RECT 51.505 180.315 51.675 180.485 ;
        RECT 50.065 180.145 51.675 180.315 ;
        RECT 51.945 180.250 52.115 180.985 ;
        RECT 49.535 179.575 49.865 180.075 ;
        RECT 50.065 179.795 50.235 180.145 ;
        RECT 50.435 179.575 50.765 179.975 ;
        RECT 50.935 179.795 51.105 180.145 ;
        RECT 51.275 179.575 51.655 179.975 ;
        RECT 51.845 179.905 52.115 180.250 ;
        RECT 52.285 180.345 53.935 180.865 ;
        RECT 54.105 180.515 55.795 181.035 ;
        RECT 56.965 181.195 57.145 181.955 ;
        RECT 57.325 181.365 57.655 182.125 ;
        RECT 56.965 181.025 57.640 181.195 ;
        RECT 57.825 181.050 58.095 181.955 ;
        RECT 57.470 180.880 57.640 181.025 ;
        RECT 56.905 180.475 57.245 180.845 ;
        RECT 57.470 180.550 57.745 180.880 ;
        RECT 52.285 179.575 55.795 180.345 ;
        RECT 57.470 180.295 57.640 180.550 ;
        RECT 56.975 180.125 57.640 180.295 ;
        RECT 57.915 180.250 58.095 181.050 ;
        RECT 58.265 181.035 61.775 182.125 ;
        RECT 62.035 181.575 62.205 181.865 ;
        RECT 62.375 181.745 62.705 182.125 ;
        RECT 63.270 181.615 64.100 181.785 ;
        RECT 62.035 181.445 62.525 181.575 ;
        RECT 62.035 181.405 63.760 181.445 ;
        RECT 62.355 181.275 63.760 181.405 ;
        RECT 56.975 179.745 57.145 180.125 ;
        RECT 57.325 179.575 57.655 179.955 ;
        RECT 57.835 179.745 58.095 180.250 ;
        RECT 58.265 180.345 59.915 180.865 ;
        RECT 60.085 180.515 61.775 181.035 ;
        RECT 62.005 180.465 62.185 181.235 ;
        RECT 58.265 179.575 61.775 180.345 ;
        RECT 62.355 180.295 62.525 181.275 ;
        RECT 62.865 180.935 63.250 181.105 ;
        RECT 63.080 180.775 63.250 180.935 ;
        RECT 63.420 181.065 63.760 181.275 ;
        RECT 62.030 180.125 62.525 180.295 ;
        RECT 62.695 180.255 63.095 180.585 ;
        RECT 63.420 180.525 63.590 181.065 ;
        RECT 63.930 180.895 64.100 181.615 ;
        RECT 64.455 181.545 64.685 182.125 ;
        RECT 65.165 181.615 65.680 181.785 ;
        RECT 64.830 181.275 65.175 181.445 ;
        RECT 65.425 181.300 65.680 181.615 ;
        RECT 65.005 181.150 65.175 181.275 ;
        RECT 65.005 180.980 65.275 181.150 ;
        RECT 62.030 179.835 62.205 180.125 ;
        RECT 62.375 179.575 62.705 179.955 ;
        RECT 62.880 179.885 63.095 180.255 ;
        RECT 63.265 180.195 63.590 180.525 ;
        RECT 63.760 180.725 64.100 180.895 ;
        RECT 65.105 180.880 65.275 180.980 ;
        RECT 63.760 180.025 63.930 180.725 ;
        RECT 64.270 180.505 64.475 180.810 ;
        RECT 64.100 180.205 64.475 180.505 ;
        RECT 64.645 180.205 64.935 180.810 ;
        RECT 65.105 180.550 65.340 180.880 ;
        RECT 63.330 179.855 63.930 180.025 ;
        RECT 64.310 179.575 64.640 180.035 ;
        RECT 65.105 179.955 65.275 180.550 ;
        RECT 65.510 180.165 65.680 181.300 ;
        RECT 64.845 179.785 65.275 179.955 ;
        RECT 65.445 179.835 65.680 180.165 ;
        RECT 65.850 181.615 66.375 181.785 ;
        RECT 65.850 179.835 66.040 181.615 ;
        RECT 66.615 181.495 66.960 182.125 ;
        RECT 67.185 181.645 68.135 181.815 ;
        RECT 66.255 181.225 66.445 181.385 ;
        RECT 67.185 181.225 67.355 181.645 ;
        RECT 68.385 181.615 68.705 181.785 ;
        RECT 66.255 181.055 67.355 181.225 ;
        RECT 66.255 180.075 66.425 181.055 ;
        RECT 66.605 180.205 66.975 180.885 ;
        RECT 66.255 179.745 66.460 180.075 ;
        RECT 66.655 179.575 66.985 180.035 ;
        RECT 67.185 179.955 67.355 181.055 ;
        RECT 67.525 180.525 67.815 181.475 ;
        RECT 68.535 181.155 68.705 181.615 ;
        RECT 68.875 181.325 69.045 182.125 ;
        RECT 69.215 181.325 69.625 181.945 ;
        RECT 67.985 180.735 68.325 181.135 ;
        RECT 68.535 180.985 69.145 181.155 ;
        RECT 69.315 180.985 69.625 181.325 ;
        RECT 69.795 180.985 70.045 182.125 ;
        RECT 70.225 181.035 73.735 182.125 ;
        RECT 68.975 180.815 69.145 180.985 ;
        RECT 68.495 180.565 68.805 180.815 ;
        RECT 67.525 180.195 68.145 180.525 ;
        RECT 68.395 180.485 68.805 180.565 ;
        RECT 68.975 180.485 69.285 180.815 ;
        RECT 67.185 179.785 68.080 179.955 ;
        RECT 68.395 179.865 68.705 180.485 ;
        RECT 68.875 179.575 69.125 180.305 ;
        RECT 69.455 180.215 69.625 180.985 ;
        RECT 69.295 179.755 69.625 180.215 ;
        RECT 69.795 179.575 70.050 180.375 ;
        RECT 70.225 180.345 71.875 180.865 ;
        RECT 72.045 180.515 73.735 181.035 ;
        RECT 74.825 180.960 75.115 182.125 ;
        RECT 75.320 181.625 75.600 181.955 ;
        RECT 75.770 181.625 76.020 182.125 ;
        RECT 76.190 181.785 77.280 181.955 ;
        RECT 76.190 181.625 76.440 181.785 ;
        RECT 77.030 181.625 77.280 181.785 ;
        RECT 75.345 181.615 75.515 181.625 ;
        RECT 76.265 181.615 76.435 181.625 ;
        RECT 77.485 181.615 77.800 181.955 ;
        RECT 77.970 181.625 78.220 182.125 ;
        RECT 76.610 181.445 76.860 181.615 ;
        RECT 77.590 181.445 77.800 181.615 ;
        RECT 78.390 181.445 78.640 181.955 ;
        RECT 78.810 181.625 79.115 182.125 ;
        RECT 79.285 181.785 80.895 181.955 ;
        RECT 79.285 181.445 80.055 181.785 ;
        RECT 75.320 181.275 77.420 181.445 ;
        RECT 77.590 181.275 80.055 181.445 ;
        RECT 75.320 180.395 75.490 181.275 ;
        RECT 77.250 181.105 77.420 181.275 ;
        RECT 80.225 181.115 80.475 181.615 ;
        RECT 80.645 181.285 80.895 181.785 ;
        RECT 81.265 181.690 86.610 182.125 ;
        RECT 75.905 180.935 77.080 181.105 ;
        RECT 77.250 180.935 79.985 181.105 ;
        RECT 75.905 180.765 76.075 180.935 ;
        RECT 76.910 180.765 77.080 180.935 ;
        RECT 75.745 180.565 76.075 180.765 ;
        RECT 76.245 180.565 76.740 180.765 ;
        RECT 76.910 180.565 78.430 180.765 ;
        RECT 78.620 180.565 79.290 180.765 ;
        RECT 79.815 180.735 79.985 180.935 ;
        RECT 80.225 180.905 81.095 181.115 ;
        RECT 79.815 180.565 80.475 180.735 ;
        RECT 79.485 180.395 79.655 180.425 ;
        RECT 80.685 180.395 81.095 180.905 ;
        RECT 70.225 179.575 73.735 180.345 ;
        RECT 74.825 179.575 75.115 180.300 ;
        RECT 75.320 180.215 76.900 180.395 ;
        RECT 75.390 179.575 75.560 180.045 ;
        RECT 75.730 179.745 76.060 180.215 ;
        RECT 76.230 179.575 76.400 180.045 ;
        RECT 76.570 179.745 76.900 180.215 ;
        RECT 77.510 180.215 78.600 180.395 ;
        RECT 77.070 179.575 77.240 180.045 ;
        RECT 77.510 179.745 77.840 180.215 ;
        RECT 78.010 179.575 78.180 180.045 ;
        RECT 78.350 179.965 78.600 180.215 ;
        RECT 78.825 180.215 81.095 180.395 ;
        RECT 78.825 180.135 79.155 180.215 ;
        RECT 80.185 180.135 80.515 180.215 ;
        RECT 82.850 180.120 83.190 180.950 ;
        RECT 84.670 180.440 85.020 181.690 ;
        RECT 86.785 181.035 87.995 182.125 ;
        RECT 86.785 180.325 87.305 180.865 ;
        RECT 87.475 180.495 87.995 181.035 ;
        RECT 78.350 179.745 79.580 179.965 ;
        RECT 79.845 179.575 80.015 180.045 ;
        RECT 80.685 179.575 80.855 180.045 ;
        RECT 81.265 179.575 86.610 180.120 ;
        RECT 86.785 179.575 87.995 180.325 ;
        RECT 88.165 179.855 88.445 181.955 ;
        RECT 88.635 181.365 89.420 182.125 ;
        RECT 89.815 181.295 90.200 181.955 ;
        RECT 89.815 181.195 90.225 181.295 ;
        RECT 88.615 180.985 90.225 181.195 ;
        RECT 90.525 181.105 90.725 181.895 ;
        RECT 88.615 180.385 88.890 180.985 ;
        RECT 90.395 180.935 90.725 181.105 ;
        RECT 90.895 180.945 91.215 182.125 ;
        RECT 91.395 181.405 91.725 182.125 ;
        RECT 90.395 180.815 90.575 180.935 ;
        RECT 89.060 180.565 89.415 180.815 ;
        RECT 89.610 180.765 90.075 180.815 ;
        RECT 89.605 180.595 90.075 180.765 ;
        RECT 89.610 180.565 90.075 180.595 ;
        RECT 90.245 180.565 90.575 180.815 ;
        RECT 91.385 180.765 91.615 181.105 ;
        RECT 91.905 180.765 92.120 181.880 ;
        RECT 92.315 181.180 92.645 181.955 ;
        RECT 92.815 181.350 93.525 182.125 ;
        RECT 92.315 180.965 93.465 181.180 ;
        RECT 90.750 180.565 91.215 180.765 ;
        RECT 91.385 180.565 91.715 180.765 ;
        RECT 91.905 180.585 92.355 180.765 ;
        RECT 92.025 180.565 92.355 180.585 ;
        RECT 92.525 180.565 92.995 180.795 ;
        RECT 93.180 180.395 93.465 180.965 ;
        RECT 93.695 180.520 93.975 181.955 ;
        RECT 88.615 180.205 89.865 180.385 ;
        RECT 89.500 180.135 89.865 180.205 ;
        RECT 90.035 180.185 91.215 180.355 ;
        RECT 88.675 179.575 88.845 180.035 ;
        RECT 90.035 179.965 90.365 180.185 ;
        RECT 89.115 179.785 90.365 179.965 ;
        RECT 90.535 179.575 90.705 180.015 ;
        RECT 90.875 179.770 91.215 180.185 ;
        RECT 91.385 180.205 92.565 180.395 ;
        RECT 91.385 179.745 91.725 180.205 ;
        RECT 92.235 180.125 92.565 180.205 ;
        RECT 92.755 180.205 93.465 180.395 ;
        RECT 92.755 180.065 93.055 180.205 ;
        RECT 92.740 180.055 93.055 180.065 ;
        RECT 92.730 180.045 93.055 180.055 ;
        RECT 92.720 180.040 93.055 180.045 ;
        RECT 91.895 179.575 92.065 180.035 ;
        RECT 92.715 180.030 93.055 180.040 ;
        RECT 92.710 180.025 93.055 180.030 ;
        RECT 92.705 180.015 93.055 180.025 ;
        RECT 92.700 180.010 93.055 180.015 ;
        RECT 92.695 179.745 93.055 180.010 ;
        RECT 93.295 179.575 93.465 180.035 ;
        RECT 93.635 179.745 93.975 180.520 ;
        RECT 94.145 181.050 94.415 181.955 ;
        RECT 94.585 181.365 94.915 182.125 ;
        RECT 95.095 181.195 95.275 181.955 ;
        RECT 94.145 180.250 94.325 181.050 ;
        RECT 94.600 181.025 95.275 181.195 ;
        RECT 95.525 181.035 97.195 182.125 ;
        RECT 94.600 180.880 94.770 181.025 ;
        RECT 94.495 180.550 94.770 180.880 ;
        RECT 94.600 180.295 94.770 180.550 ;
        RECT 94.995 180.475 95.335 180.845 ;
        RECT 95.525 180.345 96.275 180.865 ;
        RECT 96.445 180.515 97.195 181.035 ;
        RECT 97.825 180.520 98.105 181.955 ;
        RECT 98.275 181.350 98.985 182.125 ;
        RECT 99.155 181.180 99.485 181.955 ;
        RECT 98.335 180.965 99.485 181.180 ;
        RECT 94.145 179.745 94.405 180.250 ;
        RECT 94.600 180.125 95.265 180.295 ;
        RECT 94.585 179.575 94.915 179.955 ;
        RECT 95.095 179.745 95.265 180.125 ;
        RECT 95.525 179.575 97.195 180.345 ;
        RECT 97.825 179.745 98.165 180.520 ;
        RECT 98.335 180.395 98.620 180.965 ;
        RECT 98.805 180.565 99.275 180.795 ;
        RECT 99.680 180.765 99.895 181.880 ;
        RECT 100.075 181.405 100.405 182.125 ;
        RECT 100.185 180.765 100.415 181.105 ;
        RECT 100.585 180.960 100.875 182.125 ;
        RECT 101.045 181.035 104.555 182.125 ;
        RECT 99.445 180.585 99.895 180.765 ;
        RECT 99.445 180.565 99.775 180.585 ;
        RECT 100.085 180.565 100.415 180.765 ;
        RECT 98.335 180.205 99.045 180.395 ;
        RECT 98.745 180.065 99.045 180.205 ;
        RECT 99.235 180.205 100.415 180.395 ;
        RECT 101.045 180.345 102.695 180.865 ;
        RECT 102.865 180.515 104.555 181.035 ;
        RECT 104.725 180.985 104.985 181.955 ;
        RECT 105.155 181.700 105.540 182.125 ;
        RECT 105.710 181.530 105.965 181.955 ;
        RECT 105.155 181.335 105.965 181.530 ;
        RECT 99.235 180.125 99.565 180.205 ;
        RECT 98.745 180.055 99.060 180.065 ;
        RECT 98.745 180.045 99.070 180.055 ;
        RECT 98.745 180.040 99.080 180.045 ;
        RECT 98.335 179.575 98.505 180.035 ;
        RECT 98.745 180.030 99.085 180.040 ;
        RECT 98.745 180.025 99.090 180.030 ;
        RECT 98.745 180.015 99.095 180.025 ;
        RECT 98.745 180.010 99.100 180.015 ;
        RECT 98.745 179.745 99.105 180.010 ;
        RECT 99.735 179.575 99.905 180.035 ;
        RECT 100.075 179.745 100.415 180.205 ;
        RECT 100.585 179.575 100.875 180.300 ;
        RECT 101.045 179.575 104.555 180.345 ;
        RECT 104.725 180.315 104.910 180.985 ;
        RECT 105.155 180.815 105.505 181.335 ;
        RECT 106.155 181.165 106.400 181.955 ;
        RECT 106.570 181.700 106.955 182.125 ;
        RECT 107.125 181.530 107.400 181.955 ;
        RECT 105.080 180.485 105.505 180.815 ;
        RECT 105.675 180.985 106.400 181.165 ;
        RECT 106.570 181.335 107.400 181.530 ;
        RECT 105.675 180.485 106.325 180.985 ;
        RECT 106.570 180.815 106.920 181.335 ;
        RECT 107.570 181.165 107.995 181.955 ;
        RECT 108.165 181.700 108.550 182.125 ;
        RECT 108.720 181.530 109.155 181.955 ;
        RECT 106.495 180.485 106.920 180.815 ;
        RECT 107.090 180.985 107.995 181.165 ;
        RECT 108.165 181.360 109.155 181.530 ;
        RECT 109.335 181.405 109.665 182.125 ;
        RECT 107.090 180.485 107.920 180.985 ;
        RECT 108.165 180.815 108.500 181.360 ;
        RECT 108.090 180.485 108.500 180.815 ;
        RECT 108.670 180.485 109.155 181.190 ;
        RECT 109.325 180.765 109.555 181.105 ;
        RECT 109.845 180.765 110.060 181.880 ;
        RECT 110.255 181.180 110.585 181.955 ;
        RECT 110.755 181.350 111.465 182.125 ;
        RECT 110.255 180.965 111.405 181.180 ;
        RECT 109.325 180.565 109.655 180.765 ;
        RECT 109.845 180.585 110.295 180.765 ;
        RECT 109.965 180.565 110.295 180.585 ;
        RECT 110.465 180.565 110.935 180.795 ;
        RECT 105.155 180.315 105.505 180.485 ;
        RECT 106.155 180.315 106.325 180.485 ;
        RECT 106.570 180.315 106.920 180.485 ;
        RECT 107.570 180.315 107.920 180.485 ;
        RECT 108.165 180.315 108.500 180.485 ;
        RECT 111.120 180.395 111.405 180.965 ;
        RECT 111.635 180.520 111.915 181.955 ;
        RECT 112.165 181.195 112.345 181.955 ;
        RECT 112.525 181.365 112.855 182.125 ;
        RECT 112.165 181.025 112.840 181.195 ;
        RECT 113.025 181.050 113.295 181.955 ;
        RECT 112.670 180.880 112.840 181.025 ;
        RECT 104.725 179.745 104.985 180.315 ;
        RECT 105.155 180.145 105.965 180.315 ;
        RECT 105.155 179.575 105.540 179.975 ;
        RECT 105.710 179.745 105.965 180.145 ;
        RECT 106.155 179.745 106.400 180.315 ;
        RECT 106.570 180.145 107.380 180.315 ;
        RECT 106.570 179.575 106.955 179.975 ;
        RECT 107.125 179.745 107.380 180.145 ;
        RECT 107.570 179.745 107.995 180.315 ;
        RECT 108.165 180.145 109.155 180.315 ;
        RECT 108.165 179.575 108.550 179.975 ;
        RECT 108.720 179.745 109.155 180.145 ;
        RECT 109.325 180.205 110.505 180.395 ;
        RECT 109.325 179.745 109.665 180.205 ;
        RECT 110.175 180.125 110.505 180.205 ;
        RECT 110.695 180.205 111.405 180.395 ;
        RECT 110.695 180.065 110.995 180.205 ;
        RECT 110.680 180.055 110.995 180.065 ;
        RECT 110.670 180.045 110.995 180.055 ;
        RECT 110.660 180.040 110.995 180.045 ;
        RECT 109.835 179.575 110.005 180.035 ;
        RECT 110.655 180.030 110.995 180.040 ;
        RECT 110.650 180.025 110.995 180.030 ;
        RECT 110.645 180.015 110.995 180.025 ;
        RECT 110.640 180.010 110.995 180.015 ;
        RECT 110.635 179.745 110.995 180.010 ;
        RECT 111.235 179.575 111.405 180.035 ;
        RECT 111.575 179.745 111.915 180.520 ;
        RECT 112.105 180.475 112.445 180.845 ;
        RECT 112.670 180.550 112.945 180.880 ;
        RECT 112.670 180.295 112.840 180.550 ;
        RECT 112.175 180.125 112.840 180.295 ;
        RECT 113.115 180.250 113.295 181.050 ;
        RECT 112.175 179.745 112.345 180.125 ;
        RECT 112.525 179.575 112.855 179.955 ;
        RECT 113.035 179.745 113.295 180.250 ;
        RECT 113.465 181.050 113.735 181.955 ;
        RECT 113.905 181.365 114.235 182.125 ;
        RECT 114.415 181.195 114.595 181.955 ;
        RECT 113.465 180.250 113.645 181.050 ;
        RECT 113.920 181.025 114.595 181.195 ;
        RECT 114.845 181.050 115.115 181.955 ;
        RECT 115.285 181.365 115.615 182.125 ;
        RECT 115.795 181.195 115.975 181.955 ;
        RECT 113.920 180.880 114.090 181.025 ;
        RECT 113.815 180.550 114.090 180.880 ;
        RECT 113.920 180.295 114.090 180.550 ;
        RECT 114.315 180.475 114.655 180.845 ;
        RECT 113.465 179.745 113.725 180.250 ;
        RECT 113.920 180.125 114.585 180.295 ;
        RECT 113.905 179.575 114.235 179.955 ;
        RECT 114.415 179.745 114.585 180.125 ;
        RECT 114.845 180.250 115.025 181.050 ;
        RECT 115.300 181.025 115.975 181.195 ;
        RECT 116.305 181.195 116.485 181.955 ;
        RECT 116.665 181.365 116.995 182.125 ;
        RECT 116.305 181.025 116.980 181.195 ;
        RECT 117.165 181.050 117.435 181.955 ;
        RECT 117.610 181.615 119.265 181.905 ;
        RECT 115.300 180.880 115.470 181.025 ;
        RECT 115.195 180.550 115.470 180.880 ;
        RECT 116.810 180.880 116.980 181.025 ;
        RECT 115.300 180.295 115.470 180.550 ;
        RECT 115.695 180.475 116.035 180.845 ;
        RECT 116.245 180.475 116.585 180.845 ;
        RECT 116.810 180.550 117.085 180.880 ;
        RECT 116.810 180.295 116.980 180.550 ;
        RECT 114.845 179.745 115.105 180.250 ;
        RECT 115.300 180.125 115.965 180.295 ;
        RECT 115.285 179.575 115.615 179.955 ;
        RECT 115.795 179.745 115.965 180.125 ;
        RECT 116.315 180.125 116.980 180.295 ;
        RECT 117.255 180.250 117.435 181.050 ;
        RECT 117.610 181.275 119.200 181.445 ;
        RECT 119.435 181.325 119.715 182.125 ;
        RECT 117.610 180.985 117.930 181.275 ;
        RECT 119.030 181.155 119.200 181.275 ;
        RECT 116.315 179.745 116.485 180.125 ;
        RECT 116.665 179.575 116.995 179.955 ;
        RECT 117.175 179.745 117.435 180.250 ;
        RECT 117.610 180.245 117.960 180.815 ;
        RECT 118.130 180.485 118.840 181.105 ;
        RECT 119.030 180.985 119.755 181.155 ;
        RECT 119.925 180.985 120.195 181.955 ;
        RECT 120.445 181.195 120.625 181.955 ;
        RECT 120.805 181.365 121.135 182.125 ;
        RECT 120.445 181.025 121.120 181.195 ;
        RECT 121.305 181.050 121.575 181.955 ;
        RECT 119.585 180.815 119.755 180.985 ;
        RECT 119.010 180.485 119.415 180.815 ;
        RECT 119.585 180.485 119.855 180.815 ;
        RECT 119.585 180.315 119.755 180.485 ;
        RECT 118.145 180.145 119.755 180.315 ;
        RECT 120.025 180.250 120.195 180.985 ;
        RECT 120.950 180.880 121.120 181.025 ;
        RECT 120.385 180.475 120.725 180.845 ;
        RECT 120.950 180.550 121.225 180.880 ;
        RECT 120.950 180.295 121.120 180.550 ;
        RECT 117.615 179.575 117.945 180.075 ;
        RECT 118.145 179.795 118.315 180.145 ;
        RECT 118.515 179.575 118.845 179.975 ;
        RECT 119.015 179.795 119.185 180.145 ;
        RECT 119.355 179.575 119.735 179.975 ;
        RECT 119.925 179.905 120.195 180.250 ;
        RECT 120.455 180.125 121.120 180.295 ;
        RECT 121.395 180.250 121.575 181.050 ;
        RECT 121.745 181.035 125.255 182.125 ;
        RECT 120.455 179.745 120.625 180.125 ;
        RECT 120.805 179.575 121.135 179.955 ;
        RECT 121.315 179.745 121.575 180.250 ;
        RECT 121.745 180.345 123.395 180.865 ;
        RECT 123.565 180.515 125.255 181.035 ;
        RECT 126.345 180.960 126.635 182.125 ;
        RECT 126.805 181.405 127.265 181.955 ;
        RECT 127.455 181.405 127.785 182.125 ;
        RECT 121.745 179.575 125.255 180.345 ;
        RECT 126.345 179.575 126.635 180.300 ;
        RECT 126.805 180.035 127.055 181.405 ;
        RECT 127.985 181.235 128.285 181.785 ;
        RECT 128.455 181.455 128.735 182.125 ;
        RECT 127.345 181.065 128.285 181.235 ;
        RECT 127.345 180.815 127.515 181.065 ;
        RECT 128.655 180.815 128.920 181.175 ;
        RECT 129.105 181.035 130.315 182.125 ;
        RECT 127.225 180.485 127.515 180.815 ;
        RECT 127.685 180.565 128.025 180.815 ;
        RECT 128.245 180.565 128.920 180.815 ;
        RECT 127.345 180.395 127.515 180.485 ;
        RECT 127.345 180.205 128.735 180.395 ;
        RECT 126.805 179.745 127.365 180.035 ;
        RECT 127.535 179.575 127.785 180.035 ;
        RECT 128.405 179.845 128.735 180.205 ;
        RECT 129.105 180.325 129.625 180.865 ;
        RECT 129.795 180.495 130.315 181.035 ;
        RECT 130.495 180.985 130.825 182.125 ;
        RECT 131.355 181.155 131.685 181.940 ;
        RECT 131.005 180.985 131.685 181.155 ;
        RECT 132.785 180.985 133.055 181.955 ;
        RECT 133.265 181.325 133.545 182.125 ;
        RECT 133.715 181.615 135.370 181.905 ;
        RECT 133.780 181.275 135.370 181.445 ;
        RECT 133.780 181.155 133.950 181.275 ;
        RECT 133.225 180.985 133.950 181.155 ;
        RECT 130.485 180.565 130.835 180.815 ;
        RECT 131.005 180.385 131.175 180.985 ;
        RECT 131.345 180.565 131.695 180.815 ;
        RECT 129.105 179.575 130.315 180.325 ;
        RECT 130.495 179.575 130.765 180.385 ;
        RECT 130.935 179.745 131.265 180.385 ;
        RECT 131.435 179.575 131.675 180.385 ;
        RECT 132.785 180.250 132.955 180.985 ;
        RECT 133.225 180.815 133.395 180.985 ;
        RECT 134.140 180.935 134.855 181.105 ;
        RECT 135.050 180.985 135.370 181.275 ;
        RECT 135.545 180.985 135.815 181.955 ;
        RECT 136.025 181.325 136.305 182.125 ;
        RECT 136.475 181.615 138.130 181.905 ;
        RECT 139.230 181.615 140.885 181.905 ;
        RECT 136.540 181.275 138.130 181.445 ;
        RECT 136.540 181.155 136.710 181.275 ;
        RECT 135.985 180.985 136.710 181.155 ;
        RECT 133.125 180.485 133.395 180.815 ;
        RECT 133.565 180.485 133.970 180.815 ;
        RECT 134.140 180.485 134.850 180.935 ;
        RECT 133.225 180.315 133.395 180.485 ;
        RECT 132.785 179.905 133.055 180.250 ;
        RECT 133.225 180.145 134.835 180.315 ;
        RECT 135.020 180.245 135.370 180.815 ;
        RECT 135.545 180.250 135.715 180.985 ;
        RECT 135.985 180.815 136.155 180.985 ;
        RECT 136.900 180.935 137.615 181.105 ;
        RECT 137.810 180.985 138.130 181.275 ;
        RECT 139.230 181.275 140.820 181.445 ;
        RECT 141.055 181.325 141.335 182.125 ;
        RECT 139.230 180.985 139.550 181.275 ;
        RECT 140.650 181.155 140.820 181.275 ;
        RECT 139.745 180.935 140.460 181.105 ;
        RECT 140.650 180.985 141.375 181.155 ;
        RECT 141.545 180.985 141.815 181.955 ;
        RECT 141.985 181.530 142.420 181.955 ;
        RECT 142.590 181.700 142.975 182.125 ;
        RECT 141.985 181.360 142.975 181.530 ;
        RECT 135.885 180.485 136.155 180.815 ;
        RECT 136.325 180.485 136.730 180.815 ;
        RECT 136.900 180.485 137.610 180.935 ;
        RECT 135.985 180.315 136.155 180.485 ;
        RECT 133.245 179.575 133.625 179.975 ;
        RECT 133.795 179.795 133.965 180.145 ;
        RECT 134.135 179.575 134.465 179.975 ;
        RECT 134.665 179.795 134.835 180.145 ;
        RECT 135.035 179.575 135.365 180.075 ;
        RECT 135.545 179.905 135.815 180.250 ;
        RECT 135.985 180.145 137.595 180.315 ;
        RECT 137.780 180.245 138.130 180.815 ;
        RECT 139.230 180.245 139.580 180.815 ;
        RECT 139.750 180.485 140.460 180.935 ;
        RECT 141.205 180.815 141.375 180.985 ;
        RECT 140.630 180.485 141.035 180.815 ;
        RECT 141.205 180.485 141.475 180.815 ;
        RECT 141.205 180.315 141.375 180.485 ;
        RECT 136.005 179.575 136.385 179.975 ;
        RECT 136.555 179.795 136.725 180.145 ;
        RECT 136.895 179.575 137.225 179.975 ;
        RECT 137.425 179.795 137.595 180.145 ;
        RECT 139.765 180.145 141.375 180.315 ;
        RECT 141.645 180.250 141.815 180.985 ;
        RECT 141.985 180.485 142.470 181.190 ;
        RECT 142.640 180.815 142.975 181.360 ;
        RECT 143.145 181.165 143.570 181.955 ;
        RECT 143.740 181.530 144.015 181.955 ;
        RECT 144.185 181.700 144.570 182.125 ;
        RECT 143.740 181.335 144.570 181.530 ;
        RECT 143.145 180.985 144.050 181.165 ;
        RECT 142.640 180.485 143.050 180.815 ;
        RECT 143.220 180.485 144.050 180.985 ;
        RECT 144.220 180.815 144.570 181.335 ;
        RECT 144.740 181.165 144.985 181.955 ;
        RECT 145.175 181.530 145.430 181.955 ;
        RECT 145.600 181.700 145.985 182.125 ;
        RECT 145.175 181.335 145.985 181.530 ;
        RECT 144.740 180.985 145.465 181.165 ;
        RECT 144.220 180.485 144.645 180.815 ;
        RECT 144.815 180.485 145.465 180.985 ;
        RECT 145.635 180.815 145.985 181.335 ;
        RECT 146.155 180.985 146.415 181.955 ;
        RECT 146.585 180.985 146.865 182.125 ;
        RECT 145.635 180.485 146.060 180.815 ;
        RECT 142.640 180.315 142.975 180.485 ;
        RECT 143.220 180.315 143.570 180.485 ;
        RECT 144.220 180.315 144.570 180.485 ;
        RECT 144.815 180.315 144.985 180.485 ;
        RECT 145.635 180.315 145.985 180.485 ;
        RECT 146.230 180.315 146.415 180.985 ;
        RECT 147.035 180.975 147.365 181.955 ;
        RECT 147.535 180.985 147.795 182.125 ;
        RECT 148.885 181.035 150.095 182.125 ;
        RECT 146.595 180.545 146.930 180.815 ;
        RECT 147.100 180.375 147.270 180.975 ;
        RECT 147.440 180.565 147.775 180.815 ;
        RECT 148.885 180.495 149.405 181.035 ;
        RECT 137.795 179.575 138.125 180.075 ;
        RECT 139.235 179.575 139.565 180.075 ;
        RECT 139.765 179.795 139.935 180.145 ;
        RECT 140.135 179.575 140.465 179.975 ;
        RECT 140.635 179.795 140.805 180.145 ;
        RECT 140.975 179.575 141.355 179.975 ;
        RECT 141.545 179.905 141.815 180.250 ;
        RECT 141.985 180.145 142.975 180.315 ;
        RECT 141.985 179.745 142.420 180.145 ;
        RECT 142.590 179.575 142.975 179.975 ;
        RECT 143.145 179.745 143.570 180.315 ;
        RECT 143.760 180.145 144.570 180.315 ;
        RECT 143.760 179.745 144.015 180.145 ;
        RECT 144.185 179.575 144.570 179.975 ;
        RECT 144.740 179.745 144.985 180.315 ;
        RECT 145.175 180.145 145.985 180.315 ;
        RECT 145.175 179.745 145.430 180.145 ;
        RECT 145.600 179.575 145.985 179.975 ;
        RECT 146.155 179.745 146.415 180.315 ;
        RECT 146.585 179.575 146.895 180.375 ;
        RECT 147.100 179.745 147.795 180.375 ;
        RECT 149.575 180.325 150.095 180.865 ;
        RECT 148.885 179.575 150.095 180.325 ;
        RECT 36.100 179.405 150.180 179.575 ;
        RECT 36.185 178.655 37.395 179.405 ;
        RECT 37.655 178.855 37.825 179.145 ;
        RECT 37.995 179.025 38.325 179.405 ;
        RECT 37.655 178.685 38.320 178.855 ;
        RECT 36.185 178.115 36.705 178.655 ;
        RECT 36.875 177.945 37.395 178.485 ;
        RECT 36.185 176.855 37.395 177.945 ;
        RECT 37.570 177.865 37.920 178.515 ;
        RECT 38.090 177.695 38.320 178.685 ;
        RECT 37.655 177.525 38.320 177.695 ;
        RECT 37.655 177.025 37.825 177.525 ;
        RECT 37.995 176.855 38.325 177.355 ;
        RECT 38.495 177.025 38.680 179.145 ;
        RECT 38.935 178.945 39.185 179.405 ;
        RECT 39.355 178.955 39.690 179.125 ;
        RECT 39.885 178.955 40.560 179.125 ;
        RECT 39.355 178.815 39.525 178.955 ;
        RECT 38.850 177.825 39.130 178.775 ;
        RECT 39.300 178.685 39.525 178.815 ;
        RECT 39.300 177.580 39.470 178.685 ;
        RECT 39.695 178.535 40.220 178.755 ;
        RECT 39.640 177.770 39.880 178.365 ;
        RECT 40.050 177.835 40.220 178.535 ;
        RECT 40.390 178.175 40.560 178.955 ;
        RECT 40.880 178.905 41.250 179.405 ;
        RECT 41.430 178.955 41.835 179.125 ;
        RECT 42.005 178.955 42.790 179.125 ;
        RECT 41.430 178.725 41.600 178.955 ;
        RECT 40.770 178.425 41.600 178.725 ;
        RECT 41.985 178.455 42.450 178.785 ;
        RECT 40.770 178.395 40.970 178.425 ;
        RECT 41.090 178.175 41.260 178.245 ;
        RECT 40.390 178.005 41.260 178.175 ;
        RECT 40.750 177.915 41.260 178.005 ;
        RECT 39.300 177.450 39.605 177.580 ;
        RECT 40.050 177.470 40.580 177.835 ;
        RECT 38.920 176.855 39.185 177.315 ;
        RECT 39.355 177.025 39.605 177.450 ;
        RECT 40.750 177.300 40.920 177.915 ;
        RECT 39.815 177.130 40.920 177.300 ;
        RECT 41.090 176.855 41.260 177.655 ;
        RECT 41.430 177.355 41.600 178.425 ;
        RECT 41.770 177.525 41.960 178.245 ;
        RECT 42.130 177.495 42.450 178.455 ;
        RECT 42.620 178.495 42.790 178.955 ;
        RECT 43.065 178.875 43.275 179.405 ;
        RECT 43.535 178.665 43.865 179.190 ;
        RECT 44.035 178.795 44.205 179.405 ;
        RECT 44.375 178.750 44.705 179.185 ;
        RECT 44.375 178.665 44.755 178.750 ;
        RECT 43.665 178.495 43.865 178.665 ;
        RECT 44.530 178.625 44.755 178.665 ;
        RECT 42.620 178.165 43.495 178.495 ;
        RECT 43.665 178.165 44.415 178.495 ;
        RECT 41.430 177.025 41.680 177.355 ;
        RECT 42.620 177.325 42.790 178.165 ;
        RECT 43.665 177.960 43.855 178.165 ;
        RECT 44.585 178.045 44.755 178.625 ;
        RECT 44.925 178.635 46.595 179.405 ;
        RECT 47.225 178.905 47.565 179.405 ;
        RECT 44.925 178.115 45.675 178.635 ;
        RECT 44.540 177.995 44.755 178.045 ;
        RECT 42.960 177.585 43.855 177.960 ;
        RECT 44.365 177.915 44.755 177.995 ;
        RECT 45.845 177.945 46.595 178.465 ;
        RECT 47.225 178.165 47.565 178.735 ;
        RECT 47.735 178.495 47.980 179.185 ;
        RECT 48.175 178.905 48.505 179.405 ;
        RECT 48.705 178.835 48.875 179.185 ;
        RECT 49.050 179.005 49.380 179.405 ;
        RECT 49.550 178.835 49.720 179.185 ;
        RECT 49.890 179.005 50.270 179.405 ;
        RECT 48.705 178.665 50.290 178.835 ;
        RECT 50.460 178.730 50.735 179.075 ;
        RECT 50.120 178.495 50.290 178.665 ;
        RECT 47.735 178.165 48.390 178.495 ;
        RECT 41.905 177.155 42.790 177.325 ;
        RECT 42.970 176.855 43.285 177.355 ;
        RECT 43.515 177.025 43.855 177.585 ;
        RECT 44.025 176.855 44.195 177.865 ;
        RECT 44.365 177.070 44.695 177.915 ;
        RECT 44.925 176.855 46.595 177.945 ;
        RECT 47.225 176.855 47.565 177.930 ;
        RECT 47.735 177.570 47.975 178.165 ;
        RECT 48.170 177.705 48.490 177.995 ;
        RECT 48.660 177.875 49.400 178.495 ;
        RECT 49.570 178.165 49.950 178.495 ;
        RECT 50.120 178.165 50.395 178.495 ;
        RECT 50.120 177.995 50.290 178.165 ;
        RECT 50.565 177.995 50.735 178.730 ;
        RECT 50.965 178.585 51.175 179.405 ;
        RECT 51.345 178.605 51.675 179.235 ;
        RECT 51.345 178.005 51.595 178.605 ;
        RECT 51.845 178.585 52.075 179.405 ;
        RECT 52.745 178.730 53.005 179.235 ;
        RECT 53.185 179.025 53.515 179.405 ;
        RECT 53.695 178.855 53.865 179.235 ;
        RECT 51.765 178.165 52.095 178.415 ;
        RECT 49.630 177.825 50.290 177.995 ;
        RECT 49.630 177.705 49.800 177.825 ;
        RECT 48.170 177.535 49.800 177.705 ;
        RECT 47.750 177.075 49.800 177.365 ;
        RECT 49.970 176.855 50.250 177.655 ;
        RECT 50.460 177.025 50.735 177.995 ;
        RECT 50.965 176.855 51.175 177.995 ;
        RECT 51.345 177.025 51.675 178.005 ;
        RECT 51.845 176.855 52.075 177.995 ;
        RECT 52.745 177.930 52.925 178.730 ;
        RECT 53.200 178.685 53.865 178.855 ;
        RECT 53.200 178.430 53.370 178.685 ;
        RECT 54.125 178.635 57.635 179.405 ;
        RECT 58.355 178.855 58.525 179.235 ;
        RECT 58.705 179.025 59.035 179.405 ;
        RECT 58.355 178.685 59.020 178.855 ;
        RECT 59.215 178.730 59.475 179.235 ;
        RECT 53.095 178.100 53.370 178.430 ;
        RECT 53.595 178.135 53.935 178.505 ;
        RECT 54.125 178.115 55.775 178.635 ;
        RECT 53.200 177.955 53.370 178.100 ;
        RECT 52.745 177.025 53.015 177.930 ;
        RECT 53.200 177.785 53.875 177.955 ;
        RECT 55.945 177.945 57.635 178.465 ;
        RECT 58.285 178.135 58.625 178.505 ;
        RECT 58.850 178.430 59.020 178.685 ;
        RECT 58.850 178.100 59.125 178.430 ;
        RECT 58.850 177.955 59.020 178.100 ;
        RECT 53.185 176.855 53.515 177.615 ;
        RECT 53.695 177.025 53.875 177.785 ;
        RECT 54.125 176.855 57.635 177.945 ;
        RECT 58.345 177.785 59.020 177.955 ;
        RECT 59.295 177.930 59.475 178.730 ;
        RECT 59.735 178.855 59.905 179.235 ;
        RECT 60.085 179.025 60.415 179.405 ;
        RECT 59.735 178.685 60.400 178.855 ;
        RECT 60.595 178.730 60.855 179.235 ;
        RECT 59.665 178.135 60.005 178.505 ;
        RECT 60.230 178.430 60.400 178.685 ;
        RECT 60.230 178.100 60.505 178.430 ;
        RECT 60.230 177.955 60.400 178.100 ;
        RECT 58.345 177.025 58.525 177.785 ;
        RECT 58.705 176.855 59.035 177.615 ;
        RECT 59.205 177.025 59.475 177.930 ;
        RECT 59.725 177.785 60.400 177.955 ;
        RECT 60.675 177.930 60.855 178.730 ;
        RECT 61.945 178.680 62.235 179.405 ;
        RECT 62.490 178.855 62.665 179.145 ;
        RECT 62.835 179.025 63.165 179.405 ;
        RECT 62.490 178.685 62.985 178.855 ;
        RECT 63.340 178.725 63.555 179.095 ;
        RECT 63.790 178.955 64.390 179.125 ;
        RECT 59.725 177.025 59.905 177.785 ;
        RECT 60.085 176.855 60.415 177.615 ;
        RECT 60.585 177.025 60.855 177.930 ;
        RECT 61.945 176.855 62.235 178.020 ;
        RECT 62.465 177.745 62.645 178.515 ;
        RECT 62.815 177.705 62.985 178.685 ;
        RECT 63.155 178.395 63.555 178.725 ;
        RECT 63.725 178.455 64.050 178.785 ;
        RECT 63.540 178.045 63.710 178.205 ;
        RECT 63.325 177.875 63.710 178.045 ;
        RECT 63.880 177.915 64.050 178.455 ;
        RECT 64.220 178.255 64.390 178.955 ;
        RECT 64.770 178.945 65.100 179.405 ;
        RECT 65.305 179.025 65.735 179.195 ;
        RECT 64.560 178.475 64.935 178.775 ;
        RECT 64.220 178.085 64.560 178.255 ;
        RECT 64.730 178.170 64.935 178.475 ;
        RECT 65.105 178.170 65.395 178.775 ;
        RECT 65.565 178.430 65.735 179.025 ;
        RECT 65.905 178.815 66.140 179.145 ;
        RECT 63.880 177.705 64.220 177.915 ;
        RECT 62.815 177.575 64.220 177.705 ;
        RECT 62.495 177.535 64.220 177.575 ;
        RECT 62.495 177.405 62.985 177.535 ;
        RECT 62.495 177.115 62.665 177.405 ;
        RECT 64.390 177.365 64.560 178.085 ;
        RECT 65.565 178.100 65.800 178.430 ;
        RECT 65.565 178.000 65.735 178.100 ;
        RECT 65.465 177.830 65.735 178.000 ;
        RECT 65.465 177.705 65.635 177.830 ;
        RECT 65.290 177.535 65.635 177.705 ;
        RECT 65.970 177.680 66.140 178.815 ;
        RECT 62.835 176.855 63.165 177.235 ;
        RECT 63.730 177.195 64.560 177.365 ;
        RECT 64.915 176.855 65.145 177.435 ;
        RECT 65.885 177.365 66.140 177.680 ;
        RECT 65.625 177.195 66.140 177.365 ;
        RECT 66.310 177.365 66.500 179.145 ;
        RECT 66.715 178.905 66.920 179.235 ;
        RECT 67.115 178.945 67.445 179.405 ;
        RECT 67.645 179.025 68.540 179.195 ;
        RECT 66.715 177.925 66.885 178.905 ;
        RECT 67.065 178.095 67.435 178.775 ;
        RECT 67.645 177.925 67.815 179.025 ;
        RECT 66.715 177.755 67.815 177.925 ;
        RECT 66.715 177.595 66.905 177.755 ;
        RECT 66.310 177.195 66.835 177.365 ;
        RECT 67.075 176.855 67.420 177.485 ;
        RECT 67.645 177.335 67.815 177.755 ;
        RECT 67.985 178.455 68.605 178.785 ;
        RECT 68.855 178.495 69.165 179.115 ;
        RECT 69.335 178.675 69.585 179.405 ;
        RECT 69.755 178.765 70.085 179.225 ;
        RECT 67.985 177.505 68.275 178.455 ;
        RECT 68.855 178.415 69.265 178.495 ;
        RECT 68.445 177.845 68.785 178.245 ;
        RECT 68.955 178.165 69.265 178.415 ;
        RECT 69.435 178.165 69.745 178.495 ;
        RECT 69.435 177.995 69.605 178.165 ;
        RECT 69.915 177.995 70.085 178.765 ;
        RECT 70.255 178.605 70.510 179.405 ;
        RECT 70.685 178.860 76.030 179.405 ;
        RECT 77.125 179.015 78.435 179.185 ;
        RECT 72.270 178.030 72.610 178.860 ;
        RECT 68.995 177.825 69.605 177.995 ;
        RECT 68.995 177.365 69.165 177.825 ;
        RECT 69.775 177.655 70.085 177.995 ;
        RECT 67.645 177.165 68.595 177.335 ;
        RECT 68.845 177.195 69.165 177.365 ;
        RECT 69.335 176.855 69.505 177.655 ;
        RECT 69.675 177.035 70.085 177.655 ;
        RECT 70.255 176.855 70.505 177.995 ;
        RECT 74.090 177.290 74.440 178.540 ;
        RECT 77.125 178.075 77.515 179.015 ;
        RECT 78.705 178.935 78.875 179.405 ;
        RECT 77.685 178.765 78.015 178.845 ;
        RECT 79.045 178.765 79.410 179.235 ;
        RECT 79.580 178.935 79.750 179.405 ;
        RECT 79.920 178.765 80.250 179.235 ;
        RECT 77.685 178.585 80.250 178.765 ;
        RECT 80.420 178.585 80.590 179.405 ;
        RECT 80.900 178.765 81.230 179.235 ;
        RECT 81.400 178.935 81.570 179.405 ;
        RECT 81.740 179.015 82.915 179.235 ;
        RECT 81.740 178.765 81.990 179.015 ;
        RECT 80.900 178.585 81.990 178.765 ;
        RECT 82.160 178.595 82.935 178.845 ;
        RECT 77.725 178.245 78.385 178.415 ;
        RECT 77.125 177.865 77.975 178.075 ;
        RECT 78.215 178.035 78.385 178.245 ;
        RECT 79.065 178.385 80.090 178.415 ;
        RECT 79.065 178.215 80.115 178.385 ;
        RECT 80.315 178.215 81.765 178.415 ;
        RECT 79.065 178.205 80.090 178.215 ;
        RECT 79.920 178.045 80.090 178.205 ;
        RECT 82.060 178.205 82.535 178.415 ;
        RECT 82.060 178.045 82.230 178.205 ;
        RECT 78.215 177.865 79.710 178.035 ;
        RECT 79.920 177.875 82.230 178.045 ;
        RECT 77.725 177.695 77.975 177.865 ;
        RECT 79.540 177.705 79.710 177.865 ;
        RECT 82.705 177.705 82.935 178.595 ;
        RECT 83.105 178.635 86.615 179.405 ;
        RECT 87.705 178.680 87.995 179.405 ;
        RECT 83.105 178.115 84.755 178.635 ;
        RECT 89.085 178.585 89.770 179.225 ;
        RECT 89.940 178.585 90.110 179.405 ;
        RECT 90.280 178.755 90.610 179.220 ;
        RECT 90.780 178.935 90.950 179.405 ;
        RECT 91.210 179.015 92.395 179.185 ;
        RECT 92.565 178.845 92.895 179.235 ;
        RECT 93.315 178.925 93.615 179.405 ;
        RECT 91.595 178.755 91.980 178.845 ;
        RECT 90.280 178.585 91.980 178.755 ;
        RECT 92.385 178.665 92.895 178.845 ;
        RECT 93.785 178.755 94.045 179.210 ;
        RECT 94.215 178.925 94.475 179.405 ;
        RECT 94.655 178.755 94.915 179.210 ;
        RECT 95.085 178.925 95.335 179.405 ;
        RECT 95.515 178.755 95.775 179.210 ;
        RECT 95.945 178.925 96.195 179.405 ;
        RECT 96.375 178.755 96.635 179.210 ;
        RECT 96.805 178.925 97.050 179.405 ;
        RECT 97.220 178.755 97.495 179.210 ;
        RECT 97.665 178.925 97.910 179.405 ;
        RECT 98.080 178.755 98.340 179.210 ;
        RECT 98.510 178.925 98.770 179.405 ;
        RECT 98.940 178.755 99.200 179.210 ;
        RECT 99.370 178.925 99.630 179.405 ;
        RECT 99.800 178.755 100.060 179.210 ;
        RECT 100.230 178.845 100.490 179.405 ;
        RECT 84.925 177.945 86.615 178.465 ;
        RECT 70.685 176.855 76.030 177.290 ;
        RECT 77.125 176.855 77.555 177.695 ;
        RECT 77.725 177.525 79.295 177.695 ;
        RECT 79.540 177.535 82.935 177.705 ;
        RECT 77.725 177.365 77.975 177.525 ;
        RECT 79.085 177.365 79.295 177.525 ;
        RECT 80.940 177.525 82.935 177.535 ;
        RECT 78.145 176.855 78.395 177.355 ;
        RECT 78.665 177.195 78.915 177.355 ;
        RECT 79.465 177.195 79.790 177.365 ;
        RECT 78.665 177.025 79.790 177.195 ;
        RECT 79.960 176.855 80.210 177.355 ;
        RECT 80.380 177.025 80.630 177.365 ;
        RECT 80.940 177.025 81.190 177.525 ;
        RECT 81.360 176.855 81.610 177.355 ;
        RECT 81.780 177.025 82.030 177.525 ;
        RECT 82.200 176.855 82.450 177.355 ;
        RECT 82.620 177.025 82.935 177.525 ;
        RECT 83.105 176.855 86.615 177.945 ;
        RECT 87.705 176.855 87.995 178.020 ;
        RECT 89.085 177.615 89.335 178.585 ;
        RECT 89.505 178.205 89.840 178.415 ;
        RECT 90.010 178.205 90.460 178.415 ;
        RECT 90.650 178.205 91.135 178.415 ;
        RECT 89.670 178.035 89.840 178.205 ;
        RECT 90.760 178.045 91.135 178.205 ;
        RECT 91.325 178.165 91.705 178.415 ;
        RECT 91.885 178.205 92.215 178.415 ;
        RECT 89.670 177.865 90.590 178.035 ;
        RECT 89.085 177.025 89.750 177.615 ;
        RECT 89.920 176.855 90.250 177.695 ;
        RECT 90.420 177.615 90.590 177.865 ;
        RECT 90.760 177.875 91.155 178.045 ;
        RECT 90.760 177.785 91.135 177.875 ;
        RECT 91.325 177.785 91.645 178.165 ;
        RECT 92.385 178.035 92.555 178.665 ;
        RECT 93.315 178.585 100.060 178.755 ;
        RECT 92.725 178.205 93.055 178.495 ;
        RECT 91.815 177.865 92.900 178.035 ;
        RECT 91.815 177.615 91.985 177.865 ;
        RECT 90.420 177.445 91.985 177.615 ;
        RECT 90.760 177.025 91.565 177.445 ;
        RECT 92.155 176.855 92.405 177.695 ;
        RECT 92.600 177.025 92.900 177.865 ;
        RECT 93.315 177.995 94.480 178.585 ;
        RECT 100.660 178.415 100.910 179.225 ;
        RECT 101.090 178.880 101.350 179.405 ;
        RECT 101.520 178.415 101.770 179.225 ;
        RECT 101.950 178.895 102.255 179.405 ;
        RECT 102.585 178.845 102.915 179.235 ;
        RECT 103.085 179.015 104.270 179.185 ;
        RECT 104.530 178.935 104.700 179.405 ;
        RECT 94.650 178.165 101.770 178.415 ;
        RECT 101.940 178.165 102.255 178.725 ;
        RECT 102.585 178.665 103.095 178.845 ;
        RECT 102.425 178.205 102.755 178.495 ;
        RECT 93.315 177.770 100.060 177.995 ;
        RECT 93.315 176.855 93.585 177.600 ;
        RECT 93.755 177.030 94.045 177.770 ;
        RECT 94.655 177.755 100.060 177.770 ;
        RECT 94.215 176.860 94.470 177.585 ;
        RECT 94.655 177.030 94.915 177.755 ;
        RECT 95.085 176.860 95.330 177.585 ;
        RECT 95.515 177.030 95.775 177.755 ;
        RECT 95.945 176.860 96.190 177.585 ;
        RECT 96.375 177.030 96.635 177.755 ;
        RECT 96.805 176.860 97.050 177.585 ;
        RECT 97.220 177.030 97.480 177.755 ;
        RECT 97.650 176.860 97.910 177.585 ;
        RECT 98.080 177.030 98.340 177.755 ;
        RECT 98.510 176.860 98.770 177.585 ;
        RECT 98.940 177.030 99.200 177.755 ;
        RECT 99.370 176.860 99.630 177.585 ;
        RECT 99.800 177.030 100.060 177.755 ;
        RECT 100.230 176.860 100.490 177.655 ;
        RECT 100.660 177.030 100.910 178.165 ;
        RECT 94.215 176.855 100.490 176.860 ;
        RECT 101.090 176.855 101.350 177.665 ;
        RECT 101.525 177.025 101.770 178.165 ;
        RECT 102.925 178.035 103.095 178.665 ;
        RECT 103.500 178.755 103.885 178.845 ;
        RECT 104.870 178.755 105.200 179.220 ;
        RECT 103.500 178.585 105.200 178.755 ;
        RECT 105.370 178.585 105.540 179.405 ;
        RECT 105.710 178.585 106.395 179.225 ;
        RECT 106.730 178.895 106.970 179.405 ;
        RECT 107.150 178.895 107.430 179.225 ;
        RECT 107.660 178.895 107.875 179.405 ;
        RECT 103.265 178.205 103.595 178.415 ;
        RECT 103.775 178.165 104.155 178.415 ;
        RECT 104.345 178.385 104.830 178.415 ;
        RECT 104.325 178.215 104.830 178.385 ;
        RECT 102.580 177.865 103.665 178.035 ;
        RECT 101.950 176.855 102.245 177.665 ;
        RECT 102.580 177.025 102.880 177.865 ;
        RECT 103.075 176.855 103.325 177.695 ;
        RECT 103.495 177.615 103.665 177.865 ;
        RECT 103.835 177.785 104.155 178.165 ;
        RECT 104.345 178.205 104.830 178.215 ;
        RECT 105.020 178.205 105.470 178.415 ;
        RECT 105.640 178.205 105.975 178.415 ;
        RECT 104.345 177.785 104.720 178.205 ;
        RECT 105.640 178.035 105.810 178.205 ;
        RECT 104.890 177.865 105.810 178.035 ;
        RECT 104.890 177.615 105.060 177.865 ;
        RECT 103.495 177.445 105.060 177.615 ;
        RECT 103.915 177.025 104.720 177.445 ;
        RECT 105.230 176.855 105.560 177.695 ;
        RECT 106.145 177.615 106.395 178.585 ;
        RECT 106.625 178.165 106.980 178.725 ;
        RECT 107.150 177.995 107.320 178.895 ;
        RECT 107.490 178.165 107.755 178.725 ;
        RECT 108.045 178.665 108.660 179.235 ;
        RECT 108.005 177.995 108.175 178.495 ;
        RECT 106.750 177.825 108.175 177.995 ;
        RECT 106.750 177.650 107.140 177.825 ;
        RECT 105.730 177.025 106.395 177.615 ;
        RECT 107.625 176.855 107.955 177.655 ;
        RECT 108.345 177.645 108.660 178.665 ;
        RECT 108.125 177.025 108.660 177.645 ;
        RECT 108.865 178.730 109.125 179.235 ;
        RECT 109.305 179.025 109.635 179.405 ;
        RECT 109.815 178.855 109.985 179.235 ;
        RECT 108.865 177.930 109.045 178.730 ;
        RECT 109.320 178.685 109.985 178.855 ;
        RECT 110.335 178.855 110.505 179.235 ;
        RECT 110.685 179.025 111.015 179.405 ;
        RECT 110.335 178.685 111.000 178.855 ;
        RECT 111.195 178.730 111.455 179.235 ;
        RECT 109.320 178.430 109.490 178.685 ;
        RECT 109.215 178.100 109.490 178.430 ;
        RECT 109.715 178.135 110.055 178.505 ;
        RECT 110.265 178.135 110.605 178.505 ;
        RECT 110.830 178.430 111.000 178.685 ;
        RECT 109.320 177.955 109.490 178.100 ;
        RECT 110.830 178.100 111.105 178.430 ;
        RECT 110.830 177.955 111.000 178.100 ;
        RECT 108.865 177.025 109.135 177.930 ;
        RECT 109.320 177.785 109.995 177.955 ;
        RECT 109.305 176.855 109.635 177.615 ;
        RECT 109.815 177.025 109.995 177.785 ;
        RECT 110.325 177.785 111.000 177.955 ;
        RECT 111.275 177.930 111.455 178.730 ;
        RECT 111.625 178.635 113.295 179.405 ;
        RECT 113.465 178.680 113.755 179.405 ;
        RECT 113.925 178.635 116.515 179.405 ;
        RECT 117.015 179.005 117.345 179.405 ;
        RECT 117.515 178.835 117.845 179.175 ;
        RECT 118.895 179.005 119.225 179.405 ;
        RECT 116.860 178.665 119.225 178.835 ;
        RECT 119.395 178.680 119.725 179.190 ;
        RECT 119.905 178.895 120.210 179.405 ;
        RECT 111.625 178.115 112.375 178.635 ;
        RECT 112.545 177.945 113.295 178.465 ;
        RECT 113.925 178.115 115.135 178.635 ;
        RECT 110.325 177.025 110.505 177.785 ;
        RECT 110.685 176.855 111.015 177.615 ;
        RECT 111.185 177.025 111.455 177.930 ;
        RECT 111.625 176.855 113.295 177.945 ;
        RECT 113.465 176.855 113.755 178.020 ;
        RECT 115.305 177.945 116.515 178.465 ;
        RECT 113.925 176.855 116.515 177.945 ;
        RECT 116.860 177.665 117.030 178.665 ;
        RECT 119.055 178.495 119.225 178.665 ;
        RECT 117.200 177.835 117.445 178.495 ;
        RECT 117.660 177.835 117.925 178.495 ;
        RECT 118.120 177.835 118.405 178.495 ;
        RECT 118.580 178.165 118.885 178.495 ;
        RECT 119.055 178.165 119.365 178.495 ;
        RECT 118.580 177.835 118.795 178.165 ;
        RECT 116.860 177.495 117.315 177.665 ;
        RECT 116.985 177.065 117.315 177.495 ;
        RECT 117.495 177.495 118.785 177.665 ;
        RECT 117.495 177.075 117.745 177.495 ;
        RECT 117.975 176.855 118.305 177.325 ;
        RECT 118.535 177.075 118.785 177.495 ;
        RECT 118.975 176.855 119.225 177.995 ;
        RECT 119.535 177.915 119.725 178.680 ;
        RECT 119.905 178.165 120.220 178.725 ;
        RECT 120.390 178.415 120.640 179.225 ;
        RECT 120.810 178.880 121.070 179.405 ;
        RECT 121.250 178.415 121.500 179.225 ;
        RECT 121.670 178.845 121.930 179.405 ;
        RECT 122.100 178.755 122.360 179.210 ;
        RECT 122.530 178.925 122.790 179.405 ;
        RECT 122.960 178.755 123.220 179.210 ;
        RECT 123.390 178.925 123.650 179.405 ;
        RECT 123.820 178.755 124.080 179.210 ;
        RECT 124.250 178.925 124.495 179.405 ;
        RECT 124.665 178.755 124.940 179.210 ;
        RECT 125.110 178.925 125.355 179.405 ;
        RECT 125.525 178.755 125.785 179.210 ;
        RECT 125.965 178.925 126.215 179.405 ;
        RECT 126.385 178.755 126.645 179.210 ;
        RECT 126.825 178.925 127.075 179.405 ;
        RECT 127.245 178.755 127.505 179.210 ;
        RECT 127.685 178.925 127.945 179.405 ;
        RECT 128.115 178.755 128.375 179.210 ;
        RECT 128.545 178.925 128.845 179.405 ;
        RECT 122.100 178.585 128.845 178.755 ;
        RECT 120.390 178.165 127.510 178.415 ;
        RECT 119.395 177.065 119.725 177.915 ;
        RECT 119.915 176.855 120.210 177.665 ;
        RECT 120.390 177.025 120.635 178.165 ;
        RECT 120.810 176.855 121.070 177.665 ;
        RECT 121.250 177.030 121.500 178.165 ;
        RECT 127.680 177.995 128.845 178.585 ;
        RECT 122.100 177.770 128.845 177.995 ;
        RECT 122.100 177.755 127.505 177.770 ;
        RECT 121.670 176.860 121.930 177.655 ;
        RECT 122.100 177.030 122.360 177.755 ;
        RECT 122.530 176.860 122.790 177.585 ;
        RECT 122.960 177.030 123.220 177.755 ;
        RECT 123.390 176.860 123.650 177.585 ;
        RECT 123.820 177.030 124.080 177.755 ;
        RECT 124.250 176.860 124.510 177.585 ;
        RECT 124.680 177.030 124.940 177.755 ;
        RECT 125.110 176.860 125.355 177.585 ;
        RECT 125.525 177.030 125.785 177.755 ;
        RECT 125.970 176.860 126.215 177.585 ;
        RECT 126.385 177.030 126.645 177.755 ;
        RECT 126.830 176.860 127.075 177.585 ;
        RECT 127.245 177.030 127.505 177.755 ;
        RECT 127.690 176.860 127.945 177.585 ;
        RECT 128.115 177.030 128.405 177.770 ;
        RECT 121.670 176.855 127.945 176.860 ;
        RECT 128.575 176.855 128.845 177.600 ;
        RECT 130.025 177.025 130.775 179.235 ;
        RECT 131.865 178.905 132.205 179.405 ;
        RECT 131.865 178.165 132.205 178.735 ;
        RECT 132.375 178.495 132.620 179.185 ;
        RECT 132.815 178.905 133.145 179.405 ;
        RECT 133.345 178.835 133.515 179.185 ;
        RECT 133.690 179.005 134.020 179.405 ;
        RECT 134.190 178.835 134.360 179.185 ;
        RECT 134.530 179.005 134.910 179.405 ;
        RECT 133.345 178.665 134.930 178.835 ;
        RECT 135.100 178.730 135.375 179.075 ;
        RECT 134.760 178.495 134.930 178.665 ;
        RECT 132.375 178.165 133.030 178.495 ;
        RECT 131.865 176.855 132.205 177.930 ;
        RECT 132.375 177.570 132.615 178.165 ;
        RECT 132.810 177.705 133.130 177.995 ;
        RECT 133.300 177.875 134.040 178.495 ;
        RECT 134.210 178.165 134.590 178.495 ;
        RECT 134.760 178.165 135.035 178.495 ;
        RECT 134.760 177.995 134.930 178.165 ;
        RECT 135.205 177.995 135.375 178.730 ;
        RECT 135.630 178.835 135.805 179.235 ;
        RECT 135.975 179.025 136.305 179.405 ;
        RECT 136.550 178.905 136.780 179.235 ;
        RECT 135.630 178.665 136.260 178.835 ;
        RECT 136.090 178.495 136.260 178.665 ;
        RECT 134.270 177.825 134.930 177.995 ;
        RECT 134.270 177.705 134.440 177.825 ;
        RECT 132.810 177.535 134.440 177.705 ;
        RECT 132.390 177.075 134.440 177.365 ;
        RECT 134.610 176.855 134.890 177.655 ;
        RECT 135.100 177.025 135.375 177.995 ;
        RECT 135.545 177.815 135.910 178.495 ;
        RECT 136.090 178.165 136.440 178.495 ;
        RECT 136.090 177.645 136.260 178.165 ;
        RECT 135.630 177.475 136.260 177.645 ;
        RECT 136.610 177.615 136.780 178.905 ;
        RECT 136.980 177.795 137.260 179.070 ;
        RECT 137.485 179.065 137.755 179.070 ;
        RECT 137.445 178.895 137.755 179.065 ;
        RECT 138.215 179.025 138.545 179.405 ;
        RECT 138.715 179.150 139.050 179.195 ;
        RECT 137.485 177.795 137.755 178.895 ;
        RECT 137.945 177.795 138.285 178.825 ;
        RECT 138.715 178.685 139.055 179.150 ;
        RECT 138.455 178.165 138.715 178.495 ;
        RECT 138.455 177.615 138.625 178.165 ;
        RECT 138.885 177.995 139.055 178.685 ;
        RECT 139.225 178.680 139.515 179.405 ;
        RECT 140.235 178.855 140.405 179.145 ;
        RECT 140.575 179.025 140.905 179.405 ;
        RECT 140.235 178.685 140.900 178.855 ;
        RECT 135.630 177.025 135.805 177.475 ;
        RECT 136.610 177.445 138.625 177.615 ;
        RECT 135.975 176.855 136.305 177.295 ;
        RECT 136.610 177.025 136.780 177.445 ;
        RECT 137.015 176.855 137.685 177.265 ;
        RECT 137.900 177.025 138.070 177.445 ;
        RECT 138.270 176.855 138.600 177.265 ;
        RECT 138.795 177.025 139.055 177.995 ;
        RECT 139.225 176.855 139.515 178.020 ;
        RECT 140.150 177.865 140.500 178.515 ;
        RECT 140.670 177.695 140.900 178.685 ;
        RECT 140.235 177.525 140.900 177.695 ;
        RECT 140.235 177.025 140.405 177.525 ;
        RECT 140.575 176.855 140.905 177.355 ;
        RECT 141.075 177.025 141.260 179.145 ;
        RECT 141.515 178.945 141.765 179.405 ;
        RECT 141.935 178.955 142.270 179.125 ;
        RECT 142.465 178.955 143.140 179.125 ;
        RECT 141.935 178.815 142.105 178.955 ;
        RECT 141.430 177.825 141.710 178.775 ;
        RECT 141.880 178.685 142.105 178.815 ;
        RECT 141.880 177.580 142.050 178.685 ;
        RECT 142.275 178.535 142.800 178.755 ;
        RECT 142.220 177.770 142.460 178.365 ;
        RECT 142.630 177.835 142.800 178.535 ;
        RECT 142.970 178.175 143.140 178.955 ;
        RECT 143.460 178.905 143.830 179.405 ;
        RECT 144.010 178.955 144.415 179.125 ;
        RECT 144.585 178.955 145.370 179.125 ;
        RECT 144.010 178.725 144.180 178.955 ;
        RECT 143.350 178.425 144.180 178.725 ;
        RECT 144.565 178.455 145.030 178.785 ;
        RECT 143.350 178.395 143.550 178.425 ;
        RECT 143.670 178.175 143.840 178.245 ;
        RECT 142.970 178.005 143.840 178.175 ;
        RECT 143.330 177.915 143.840 178.005 ;
        RECT 141.880 177.450 142.185 177.580 ;
        RECT 142.630 177.470 143.160 177.835 ;
        RECT 141.500 176.855 141.765 177.315 ;
        RECT 141.935 177.025 142.185 177.450 ;
        RECT 143.330 177.300 143.500 177.915 ;
        RECT 142.395 177.130 143.500 177.300 ;
        RECT 143.670 176.855 143.840 177.655 ;
        RECT 144.010 177.355 144.180 178.425 ;
        RECT 144.350 177.525 144.540 178.245 ;
        RECT 144.710 177.495 145.030 178.455 ;
        RECT 145.200 178.495 145.370 178.955 ;
        RECT 145.645 178.875 145.855 179.405 ;
        RECT 146.115 178.665 146.445 179.190 ;
        RECT 146.615 178.795 146.785 179.405 ;
        RECT 146.955 178.750 147.285 179.185 ;
        RECT 146.955 178.665 147.335 178.750 ;
        RECT 146.245 178.495 146.445 178.665 ;
        RECT 147.110 178.625 147.335 178.665 ;
        RECT 145.200 178.165 146.075 178.495 ;
        RECT 146.245 178.165 146.995 178.495 ;
        RECT 144.010 177.025 144.260 177.355 ;
        RECT 145.200 177.325 145.370 178.165 ;
        RECT 146.245 177.960 146.435 178.165 ;
        RECT 147.165 178.045 147.335 178.625 ;
        RECT 147.505 178.655 148.715 179.405 ;
        RECT 148.885 178.655 150.095 179.405 ;
        RECT 147.505 178.115 148.025 178.655 ;
        RECT 147.120 177.995 147.335 178.045 ;
        RECT 145.540 177.585 146.435 177.960 ;
        RECT 146.945 177.915 147.335 177.995 ;
        RECT 148.195 177.945 148.715 178.485 ;
        RECT 144.485 177.155 145.370 177.325 ;
        RECT 145.550 176.855 145.865 177.355 ;
        RECT 146.095 177.025 146.435 177.585 ;
        RECT 146.605 176.855 146.775 177.865 ;
        RECT 146.945 177.070 147.275 177.915 ;
        RECT 147.505 176.855 148.715 177.945 ;
        RECT 148.885 177.945 149.405 178.485 ;
        RECT 149.575 178.115 150.095 178.655 ;
        RECT 148.885 176.855 150.095 177.945 ;
        RECT 36.100 176.685 150.180 176.855 ;
        RECT 36.185 175.595 37.395 176.685 ;
        RECT 37.565 175.595 40.155 176.685 ;
        RECT 36.185 174.885 36.705 175.425 ;
        RECT 36.875 175.055 37.395 175.595 ;
        RECT 37.565 174.905 38.775 175.425 ;
        RECT 38.945 175.075 40.155 175.595 ;
        RECT 40.335 175.715 40.665 176.500 ;
        RECT 40.335 175.545 41.015 175.715 ;
        RECT 41.195 175.545 41.525 176.685 ;
        RECT 41.705 175.595 44.295 176.685 ;
        RECT 40.325 175.125 40.675 175.375 ;
        RECT 40.845 174.945 41.015 175.545 ;
        RECT 41.185 175.125 41.535 175.375 ;
        RECT 36.185 174.135 37.395 174.885 ;
        RECT 37.565 174.135 40.155 174.905 ;
        RECT 40.345 174.135 40.585 174.945 ;
        RECT 40.755 174.305 41.085 174.945 ;
        RECT 41.255 174.135 41.525 174.945 ;
        RECT 41.705 174.905 42.915 175.425 ;
        RECT 43.085 175.075 44.295 175.595 ;
        RECT 44.465 175.545 44.725 176.515 ;
        RECT 44.895 176.260 45.280 176.685 ;
        RECT 45.450 176.090 45.705 176.515 ;
        RECT 44.895 175.895 45.705 176.090 ;
        RECT 41.705 174.135 44.295 174.905 ;
        RECT 44.465 174.875 44.650 175.545 ;
        RECT 44.895 175.375 45.245 175.895 ;
        RECT 45.895 175.725 46.140 176.515 ;
        RECT 46.310 176.260 46.695 176.685 ;
        RECT 46.865 176.090 47.140 176.515 ;
        RECT 44.820 175.045 45.245 175.375 ;
        RECT 45.415 175.545 46.140 175.725 ;
        RECT 46.310 175.895 47.140 176.090 ;
        RECT 45.415 175.045 46.065 175.545 ;
        RECT 46.310 175.375 46.660 175.895 ;
        RECT 47.310 175.725 47.735 176.515 ;
        RECT 47.905 176.260 48.290 176.685 ;
        RECT 48.460 176.090 48.895 176.515 ;
        RECT 46.235 175.045 46.660 175.375 ;
        RECT 46.830 175.545 47.735 175.725 ;
        RECT 47.905 175.920 48.895 176.090 ;
        RECT 46.830 175.045 47.660 175.545 ;
        RECT 47.905 175.375 48.240 175.920 ;
        RECT 47.830 175.045 48.240 175.375 ;
        RECT 48.410 175.045 48.895 175.750 ;
        RECT 49.065 175.520 49.355 176.685 ;
        RECT 49.525 175.545 49.795 176.515 ;
        RECT 50.005 175.885 50.285 176.685 ;
        RECT 50.455 176.175 52.110 176.465 ;
        RECT 50.520 175.835 52.110 176.005 ;
        RECT 50.520 175.715 50.690 175.835 ;
        RECT 49.965 175.545 50.690 175.715 ;
        RECT 44.895 174.875 45.245 175.045 ;
        RECT 45.895 174.875 46.065 175.045 ;
        RECT 46.310 174.875 46.660 175.045 ;
        RECT 47.310 174.875 47.660 175.045 ;
        RECT 47.905 174.875 48.240 175.045 ;
        RECT 44.465 174.305 44.725 174.875 ;
        RECT 44.895 174.705 45.705 174.875 ;
        RECT 44.895 174.135 45.280 174.535 ;
        RECT 45.450 174.305 45.705 174.705 ;
        RECT 45.895 174.305 46.140 174.875 ;
        RECT 46.310 174.705 47.120 174.875 ;
        RECT 46.310 174.135 46.695 174.535 ;
        RECT 46.865 174.305 47.120 174.705 ;
        RECT 47.310 174.305 47.735 174.875 ;
        RECT 47.905 174.705 48.895 174.875 ;
        RECT 47.905 174.135 48.290 174.535 ;
        RECT 48.460 174.305 48.895 174.705 ;
        RECT 49.065 174.135 49.355 174.860 ;
        RECT 49.525 174.810 49.695 175.545 ;
        RECT 49.965 175.375 50.135 175.545 ;
        RECT 49.865 175.045 50.135 175.375 ;
        RECT 50.305 175.045 50.710 175.375 ;
        RECT 50.880 175.045 51.590 175.665 ;
        RECT 51.790 175.545 52.110 175.835 ;
        RECT 52.365 175.755 52.545 176.515 ;
        RECT 52.725 175.925 53.055 176.685 ;
        RECT 52.365 175.585 53.040 175.755 ;
        RECT 53.225 175.610 53.495 176.515 ;
        RECT 52.870 175.440 53.040 175.585 ;
        RECT 49.965 174.875 50.135 175.045 ;
        RECT 49.525 174.465 49.795 174.810 ;
        RECT 49.965 174.705 51.575 174.875 ;
        RECT 51.760 174.805 52.110 175.375 ;
        RECT 52.305 175.035 52.645 175.405 ;
        RECT 52.870 175.110 53.145 175.440 ;
        RECT 52.870 174.855 53.040 175.110 ;
        RECT 49.985 174.135 50.365 174.535 ;
        RECT 50.535 174.355 50.705 174.705 ;
        RECT 50.875 174.135 51.205 174.535 ;
        RECT 51.405 174.355 51.575 174.705 ;
        RECT 52.375 174.685 53.040 174.855 ;
        RECT 53.315 174.810 53.495 175.610 ;
        RECT 53.675 175.545 53.925 176.685 ;
        RECT 54.095 175.885 54.505 176.505 ;
        RECT 54.675 175.885 54.845 176.685 ;
        RECT 55.015 176.175 55.335 176.345 ;
        RECT 55.585 176.205 56.535 176.375 ;
        RECT 54.095 175.545 54.405 175.885 ;
        RECT 55.015 175.715 55.185 176.175 ;
        RECT 54.575 175.545 55.185 175.715 ;
        RECT 51.775 174.135 52.105 174.635 ;
        RECT 52.375 174.305 52.545 174.685 ;
        RECT 52.725 174.135 53.055 174.515 ;
        RECT 53.235 174.305 53.495 174.810 ;
        RECT 53.670 174.135 53.925 174.935 ;
        RECT 54.095 174.775 54.265 175.545 ;
        RECT 54.575 175.375 54.745 175.545 ;
        RECT 54.435 175.045 54.745 175.375 ;
        RECT 54.915 175.125 55.225 175.375 ;
        RECT 55.395 175.295 55.735 175.695 ;
        RECT 54.915 175.045 55.325 175.125 ;
        RECT 55.905 175.085 56.195 176.035 ;
        RECT 54.095 174.315 54.425 174.775 ;
        RECT 54.595 174.135 54.845 174.865 ;
        RECT 55.015 174.425 55.325 175.045 ;
        RECT 55.575 174.755 56.195 175.085 ;
        RECT 56.365 175.785 56.535 176.205 ;
        RECT 56.760 176.055 57.105 176.685 ;
        RECT 57.345 176.175 57.870 176.345 ;
        RECT 57.275 175.785 57.465 175.945 ;
        RECT 56.365 175.615 57.465 175.785 ;
        RECT 56.365 174.515 56.535 175.615 ;
        RECT 56.745 174.765 57.115 175.445 ;
        RECT 57.295 174.635 57.465 175.615 ;
        RECT 55.640 174.345 56.535 174.515 ;
        RECT 56.735 174.135 57.065 174.595 ;
        RECT 57.260 174.305 57.465 174.635 ;
        RECT 57.680 174.395 57.870 176.175 ;
        RECT 58.040 176.175 58.555 176.345 ;
        RECT 58.040 175.860 58.295 176.175 ;
        RECT 59.035 176.105 59.265 176.685 ;
        RECT 59.620 176.175 60.450 176.345 ;
        RECT 61.015 176.305 61.345 176.685 ;
        RECT 58.040 174.725 58.210 175.860 ;
        RECT 58.545 175.835 58.890 176.005 ;
        RECT 58.545 175.710 58.715 175.835 ;
        RECT 58.445 175.540 58.715 175.710 ;
        RECT 58.445 175.440 58.615 175.540 ;
        RECT 58.380 175.110 58.615 175.440 ;
        RECT 59.620 175.455 59.790 176.175 ;
        RECT 61.515 176.135 61.685 176.425 ;
        RECT 61.195 176.005 61.685 176.135 ;
        RECT 59.960 175.965 61.685 176.005 ;
        RECT 59.960 175.835 61.365 175.965 ;
        RECT 62.035 175.940 62.305 176.685 ;
        RECT 62.935 176.680 69.210 176.685 ;
        RECT 59.960 175.625 60.300 175.835 ;
        RECT 58.040 174.395 58.275 174.725 ;
        RECT 58.445 174.515 58.615 175.110 ;
        RECT 58.785 174.765 59.075 175.370 ;
        RECT 59.245 175.065 59.450 175.370 ;
        RECT 59.620 175.285 59.960 175.455 ;
        RECT 59.245 174.765 59.620 175.065 ;
        RECT 58.445 174.345 58.875 174.515 ;
        RECT 59.080 174.135 59.410 174.595 ;
        RECT 59.790 174.585 59.960 175.285 ;
        RECT 60.130 175.085 60.300 175.625 ;
        RECT 60.470 175.495 60.855 175.665 ;
        RECT 60.470 175.335 60.640 175.495 ;
        RECT 60.130 174.755 60.455 175.085 ;
        RECT 60.625 174.815 61.025 175.145 ;
        RECT 61.195 174.855 61.365 175.835 ;
        RECT 61.535 175.025 61.715 175.795 ;
        RECT 62.475 175.770 62.765 176.510 ;
        RECT 62.935 175.955 63.190 176.680 ;
        RECT 63.375 175.785 63.635 176.510 ;
        RECT 63.805 175.955 64.050 176.680 ;
        RECT 64.235 175.785 64.495 176.510 ;
        RECT 64.665 175.955 64.910 176.680 ;
        RECT 65.095 175.785 65.355 176.510 ;
        RECT 65.525 175.955 65.770 176.680 ;
        RECT 65.940 175.785 66.200 176.510 ;
        RECT 66.370 175.955 66.630 176.680 ;
        RECT 66.800 175.785 67.060 176.510 ;
        RECT 67.230 175.955 67.490 176.680 ;
        RECT 67.660 175.785 67.920 176.510 ;
        RECT 68.090 175.955 68.350 176.680 ;
        RECT 68.520 175.785 68.780 176.510 ;
        RECT 68.950 175.885 69.210 176.680 ;
        RECT 63.375 175.770 68.780 175.785 ;
        RECT 62.035 175.545 68.780 175.770 ;
        RECT 62.035 174.955 63.200 175.545 ;
        RECT 69.380 175.375 69.630 176.510 ;
        RECT 69.810 175.875 70.070 176.685 ;
        RECT 70.245 175.375 70.490 176.515 ;
        RECT 70.670 175.875 70.965 176.685 ;
        RECT 71.145 175.595 74.655 176.685 ;
        RECT 63.370 175.125 70.490 175.375 ;
        RECT 59.790 174.415 60.390 174.585 ;
        RECT 60.625 174.445 60.840 174.815 ;
        RECT 61.195 174.685 61.690 174.855 ;
        RECT 62.035 174.785 68.780 174.955 ;
        RECT 61.015 174.135 61.345 174.515 ;
        RECT 61.515 174.395 61.690 174.685 ;
        RECT 62.035 174.135 62.335 174.615 ;
        RECT 62.505 174.330 62.765 174.785 ;
        RECT 62.935 174.135 63.195 174.615 ;
        RECT 63.375 174.330 63.635 174.785 ;
        RECT 63.805 174.135 64.055 174.615 ;
        RECT 64.235 174.330 64.495 174.785 ;
        RECT 64.665 174.135 64.915 174.615 ;
        RECT 65.095 174.330 65.355 174.785 ;
        RECT 65.525 174.135 65.770 174.615 ;
        RECT 65.940 174.330 66.215 174.785 ;
        RECT 66.385 174.135 66.630 174.615 ;
        RECT 66.800 174.330 67.060 174.785 ;
        RECT 67.230 174.135 67.490 174.615 ;
        RECT 67.660 174.330 67.920 174.785 ;
        RECT 68.090 174.135 68.350 174.615 ;
        RECT 68.520 174.330 68.780 174.785 ;
        RECT 68.950 174.135 69.210 174.695 ;
        RECT 69.380 174.315 69.630 175.125 ;
        RECT 69.810 174.135 70.070 174.660 ;
        RECT 70.240 174.315 70.490 175.125 ;
        RECT 70.660 174.815 70.975 175.375 ;
        RECT 71.145 174.905 72.795 175.425 ;
        RECT 72.965 175.075 74.655 175.595 ;
        RECT 74.825 175.520 75.115 176.685 ;
        RECT 75.285 176.250 80.630 176.685 ;
        RECT 70.670 174.135 70.975 174.645 ;
        RECT 71.145 174.135 74.655 174.905 ;
        RECT 74.825 174.135 75.115 174.860 ;
        RECT 76.870 174.680 77.210 175.510 ;
        RECT 78.690 175.000 79.040 176.250 ;
        RECT 80.805 175.595 82.475 176.685 ;
        RECT 80.805 174.905 81.555 175.425 ;
        RECT 81.725 175.075 82.475 175.595 ;
        RECT 83.290 175.715 83.680 175.890 ;
        RECT 84.165 175.885 84.495 176.685 ;
        RECT 84.665 175.895 85.200 176.515 ;
        RECT 83.290 175.545 84.715 175.715 ;
        RECT 75.285 174.135 80.630 174.680 ;
        RECT 80.805 174.135 82.475 174.905 ;
        RECT 83.165 174.815 83.520 175.375 ;
        RECT 83.690 174.645 83.860 175.545 ;
        RECT 84.030 174.815 84.295 175.375 ;
        RECT 84.545 175.045 84.715 175.545 ;
        RECT 84.885 174.875 85.200 175.895 ;
        RECT 85.590 175.715 85.980 175.890 ;
        RECT 86.465 175.885 86.795 176.685 ;
        RECT 86.965 175.895 87.500 176.515 ;
        RECT 85.590 175.545 87.015 175.715 ;
        RECT 83.270 174.135 83.510 174.645 ;
        RECT 83.690 174.315 83.970 174.645 ;
        RECT 84.200 174.135 84.415 174.645 ;
        RECT 84.585 174.305 85.200 174.875 ;
        RECT 85.465 174.815 85.820 175.375 ;
        RECT 85.990 174.645 86.160 175.545 ;
        RECT 86.330 174.815 86.595 175.375 ;
        RECT 86.845 175.045 87.015 175.545 ;
        RECT 87.185 174.875 87.500 175.895 ;
        RECT 87.910 175.715 88.240 176.515 ;
        RECT 88.410 175.885 88.740 176.685 ;
        RECT 89.040 175.715 89.370 176.515 ;
        RECT 90.015 175.885 90.265 176.685 ;
        RECT 87.910 175.545 90.345 175.715 ;
        RECT 90.535 175.545 90.705 176.685 ;
        RECT 90.875 175.545 91.215 176.515 ;
        RECT 91.685 176.045 92.015 176.475 ;
        RECT 87.705 175.125 88.055 175.375 ;
        RECT 88.240 174.915 88.410 175.545 ;
        RECT 88.580 175.125 88.910 175.325 ;
        RECT 89.080 175.125 89.410 175.325 ;
        RECT 89.580 175.125 90.000 175.325 ;
        RECT 90.175 175.295 90.345 175.545 ;
        RECT 90.175 175.125 90.870 175.295 ;
        RECT 85.570 174.135 85.810 174.645 ;
        RECT 85.990 174.315 86.270 174.645 ;
        RECT 86.500 174.135 86.715 174.645 ;
        RECT 86.885 174.305 87.500 174.875 ;
        RECT 87.910 174.305 88.410 174.915 ;
        RECT 89.040 174.785 90.265 174.955 ;
        RECT 91.040 174.935 91.215 175.545 ;
        RECT 89.040 174.305 89.370 174.785 ;
        RECT 89.540 174.135 89.765 174.595 ;
        RECT 89.935 174.305 90.265 174.785 ;
        RECT 90.455 174.135 90.705 174.935 ;
        RECT 90.875 174.305 91.215 174.935 ;
        RECT 91.560 175.875 92.015 176.045 ;
        RECT 92.195 176.045 92.445 176.465 ;
        RECT 92.675 176.215 93.005 176.685 ;
        RECT 93.235 176.045 93.485 176.465 ;
        RECT 92.195 175.875 93.485 176.045 ;
        RECT 91.560 174.875 91.730 175.875 ;
        RECT 91.900 175.045 92.145 175.705 ;
        RECT 92.360 175.045 92.625 175.705 ;
        RECT 92.820 175.045 93.105 175.705 ;
        RECT 93.280 175.375 93.495 175.705 ;
        RECT 93.675 175.545 93.925 176.685 ;
        RECT 94.095 175.625 94.425 176.475 ;
        RECT 93.280 175.045 93.585 175.375 ;
        RECT 93.755 175.045 94.065 175.375 ;
        RECT 93.755 174.875 93.925 175.045 ;
        RECT 91.560 174.705 93.925 174.875 ;
        RECT 94.235 174.860 94.425 175.625 ;
        RECT 94.605 175.595 95.815 176.685 ;
        RECT 91.715 174.135 92.045 174.535 ;
        RECT 92.215 174.365 92.545 174.705 ;
        RECT 93.595 174.135 93.925 174.535 ;
        RECT 94.095 174.350 94.425 174.860 ;
        RECT 94.605 174.885 95.125 175.425 ;
        RECT 95.295 175.055 95.815 175.595 ;
        RECT 95.985 175.545 96.245 176.515 ;
        RECT 96.415 176.260 96.800 176.685 ;
        RECT 96.970 176.090 97.225 176.515 ;
        RECT 96.415 175.895 97.225 176.090 ;
        RECT 94.605 174.135 95.815 174.885 ;
        RECT 95.985 174.875 96.170 175.545 ;
        RECT 96.415 175.375 96.765 175.895 ;
        RECT 97.415 175.725 97.660 176.515 ;
        RECT 97.830 176.260 98.215 176.685 ;
        RECT 98.385 176.090 98.660 176.515 ;
        RECT 96.340 175.045 96.765 175.375 ;
        RECT 96.935 175.545 97.660 175.725 ;
        RECT 97.830 175.895 98.660 176.090 ;
        RECT 96.935 175.045 97.585 175.545 ;
        RECT 97.830 175.375 98.180 175.895 ;
        RECT 98.830 175.725 99.255 176.515 ;
        RECT 99.425 176.260 99.810 176.685 ;
        RECT 99.980 176.090 100.415 176.515 ;
        RECT 97.755 175.045 98.180 175.375 ;
        RECT 98.350 175.545 99.255 175.725 ;
        RECT 99.425 175.920 100.415 176.090 ;
        RECT 98.350 175.045 99.180 175.545 ;
        RECT 99.425 175.375 99.760 175.920 ;
        RECT 99.350 175.045 99.760 175.375 ;
        RECT 99.930 175.045 100.415 175.750 ;
        RECT 100.585 175.520 100.875 176.685 ;
        RECT 101.200 175.675 101.500 176.515 ;
        RECT 101.695 175.845 101.945 176.685 ;
        RECT 102.535 176.095 103.340 176.515 ;
        RECT 102.115 175.925 103.680 176.095 ;
        RECT 102.115 175.675 102.285 175.925 ;
        RECT 101.200 175.505 102.285 175.675 ;
        RECT 101.045 175.045 101.375 175.335 ;
        RECT 96.415 174.875 96.765 175.045 ;
        RECT 97.415 174.875 97.585 175.045 ;
        RECT 97.830 174.875 98.180 175.045 ;
        RECT 98.830 174.875 99.180 175.045 ;
        RECT 99.425 174.875 99.760 175.045 ;
        RECT 101.545 174.875 101.715 175.505 ;
        RECT 102.455 175.375 102.775 175.755 ;
        RECT 102.965 175.665 103.340 175.755 ;
        RECT 102.945 175.495 103.340 175.665 ;
        RECT 103.510 175.675 103.680 175.925 ;
        RECT 103.850 175.845 104.180 176.685 ;
        RECT 104.350 175.925 105.015 176.515 ;
        RECT 105.485 176.045 105.815 176.475 ;
        RECT 103.510 175.505 104.430 175.675 ;
        RECT 101.885 175.125 102.215 175.335 ;
        RECT 102.395 175.125 102.775 175.375 ;
        RECT 102.965 175.335 103.340 175.495 ;
        RECT 104.260 175.335 104.430 175.505 ;
        RECT 102.965 175.125 103.450 175.335 ;
        RECT 103.640 175.125 104.090 175.335 ;
        RECT 104.260 175.125 104.595 175.335 ;
        RECT 104.765 174.955 105.015 175.925 ;
        RECT 95.985 174.305 96.245 174.875 ;
        RECT 96.415 174.705 97.225 174.875 ;
        RECT 96.415 174.135 96.800 174.535 ;
        RECT 96.970 174.305 97.225 174.705 ;
        RECT 97.415 174.305 97.660 174.875 ;
        RECT 97.830 174.705 98.640 174.875 ;
        RECT 97.830 174.135 98.215 174.535 ;
        RECT 98.385 174.305 98.640 174.705 ;
        RECT 98.830 174.305 99.255 174.875 ;
        RECT 99.425 174.705 100.415 174.875 ;
        RECT 99.425 174.135 99.810 174.535 ;
        RECT 99.980 174.305 100.415 174.705 ;
        RECT 100.585 174.135 100.875 174.860 ;
        RECT 101.205 174.695 101.715 174.875 ;
        RECT 102.120 174.785 103.820 174.955 ;
        RECT 102.120 174.695 102.505 174.785 ;
        RECT 101.205 174.305 101.535 174.695 ;
        RECT 101.705 174.355 102.890 174.525 ;
        RECT 103.150 174.135 103.320 174.605 ;
        RECT 103.490 174.320 103.820 174.785 ;
        RECT 103.990 174.135 104.160 174.955 ;
        RECT 104.330 174.315 105.015 174.955 ;
        RECT 105.360 175.875 105.815 176.045 ;
        RECT 105.995 176.045 106.245 176.465 ;
        RECT 106.475 176.215 106.805 176.685 ;
        RECT 107.035 176.045 107.285 176.465 ;
        RECT 105.995 175.875 107.285 176.045 ;
        RECT 105.360 174.875 105.530 175.875 ;
        RECT 105.700 175.045 105.945 175.705 ;
        RECT 106.160 175.045 106.425 175.705 ;
        RECT 106.620 175.045 106.905 175.705 ;
        RECT 107.080 175.375 107.295 175.705 ;
        RECT 107.475 175.545 107.725 176.685 ;
        RECT 107.895 175.625 108.225 176.475 ;
        RECT 107.080 175.045 107.385 175.375 ;
        RECT 107.555 175.045 107.865 175.375 ;
        RECT 107.555 174.875 107.725 175.045 ;
        RECT 105.360 174.705 107.725 174.875 ;
        RECT 108.035 174.860 108.225 175.625 ;
        RECT 105.515 174.135 105.845 174.535 ;
        RECT 106.015 174.365 106.345 174.705 ;
        RECT 107.395 174.135 107.725 174.535 ;
        RECT 107.895 174.350 108.225 174.860 ;
        RECT 108.405 174.415 108.685 176.515 ;
        RECT 108.875 175.925 109.660 176.685 ;
        RECT 110.055 175.855 110.440 176.515 ;
        RECT 110.055 175.755 110.465 175.855 ;
        RECT 108.855 175.545 110.465 175.755 ;
        RECT 110.765 175.665 110.965 176.455 ;
        RECT 108.855 174.945 109.130 175.545 ;
        RECT 110.635 175.495 110.965 175.665 ;
        RECT 111.135 175.505 111.455 176.685 ;
        RECT 111.625 175.595 114.215 176.685 ;
        RECT 114.385 176.090 114.820 176.515 ;
        RECT 114.990 176.260 115.375 176.685 ;
        RECT 114.385 175.920 115.375 176.090 ;
        RECT 110.635 175.375 110.815 175.495 ;
        RECT 109.300 175.125 109.655 175.375 ;
        RECT 109.850 175.325 110.315 175.375 ;
        RECT 109.845 175.155 110.315 175.325 ;
        RECT 109.850 175.125 110.315 175.155 ;
        RECT 110.485 175.125 110.815 175.375 ;
        RECT 110.990 175.125 111.455 175.325 ;
        RECT 108.855 174.765 110.105 174.945 ;
        RECT 109.740 174.695 110.105 174.765 ;
        RECT 110.275 174.745 111.455 174.915 ;
        RECT 108.915 174.135 109.085 174.595 ;
        RECT 110.275 174.525 110.605 174.745 ;
        RECT 109.355 174.345 110.605 174.525 ;
        RECT 110.775 174.135 110.945 174.575 ;
        RECT 111.115 174.330 111.455 174.745 ;
        RECT 111.625 174.905 112.835 175.425 ;
        RECT 113.005 175.075 114.215 175.595 ;
        RECT 114.385 175.045 114.870 175.750 ;
        RECT 115.040 175.375 115.375 175.920 ;
        RECT 115.545 175.725 115.970 176.515 ;
        RECT 116.140 176.090 116.415 176.515 ;
        RECT 116.585 176.260 116.970 176.685 ;
        RECT 116.140 175.895 116.970 176.090 ;
        RECT 115.545 175.545 116.450 175.725 ;
        RECT 115.040 175.045 115.450 175.375 ;
        RECT 115.620 175.045 116.450 175.545 ;
        RECT 116.620 175.375 116.970 175.895 ;
        RECT 117.140 175.725 117.385 176.515 ;
        RECT 117.575 176.090 117.830 176.515 ;
        RECT 118.000 176.260 118.385 176.685 ;
        RECT 117.575 175.895 118.385 176.090 ;
        RECT 117.140 175.545 117.865 175.725 ;
        RECT 116.620 175.045 117.045 175.375 ;
        RECT 117.215 175.045 117.865 175.545 ;
        RECT 118.035 175.375 118.385 175.895 ;
        RECT 118.555 175.545 118.815 176.515 ;
        RECT 118.995 176.075 119.325 176.505 ;
        RECT 119.505 176.245 119.700 176.685 ;
        RECT 119.870 176.075 120.200 176.505 ;
        RECT 118.995 175.905 120.200 176.075 ;
        RECT 118.995 175.575 119.890 175.905 ;
        RECT 120.370 175.735 120.645 176.505 ;
        RECT 118.035 175.045 118.460 175.375 ;
        RECT 111.625 174.135 114.215 174.905 ;
        RECT 115.040 174.875 115.375 175.045 ;
        RECT 115.620 174.875 115.970 175.045 ;
        RECT 116.620 174.875 116.970 175.045 ;
        RECT 117.215 174.875 117.385 175.045 ;
        RECT 118.035 174.875 118.385 175.045 ;
        RECT 118.630 174.875 118.815 175.545 ;
        RECT 120.060 175.545 120.645 175.735 ;
        RECT 120.830 175.545 121.150 176.685 ;
        RECT 119.000 175.045 119.295 175.375 ;
        RECT 119.475 175.045 119.890 175.375 ;
        RECT 114.385 174.705 115.375 174.875 ;
        RECT 114.385 174.305 114.820 174.705 ;
        RECT 114.990 174.135 115.375 174.535 ;
        RECT 115.545 174.305 115.970 174.875 ;
        RECT 116.160 174.705 116.970 174.875 ;
        RECT 116.160 174.305 116.415 174.705 ;
        RECT 116.585 174.135 116.970 174.535 ;
        RECT 117.140 174.305 117.385 174.875 ;
        RECT 117.575 174.705 118.385 174.875 ;
        RECT 117.575 174.305 117.830 174.705 ;
        RECT 118.000 174.135 118.385 174.535 ;
        RECT 118.555 174.305 118.815 174.875 ;
        RECT 118.995 174.135 119.295 174.865 ;
        RECT 119.475 174.425 119.705 175.045 ;
        RECT 120.060 174.875 120.235 175.545 ;
        RECT 121.330 175.375 121.525 176.425 ;
        RECT 121.705 175.835 122.035 176.515 ;
        RECT 122.235 175.885 122.490 176.685 ;
        RECT 123.130 176.295 123.465 176.515 ;
        RECT 124.470 176.305 124.825 176.685 ;
        RECT 121.705 175.555 122.055 175.835 ;
        RECT 119.905 174.695 120.235 174.875 ;
        RECT 120.405 174.725 120.645 175.375 ;
        RECT 120.890 175.325 121.150 175.375 ;
        RECT 120.885 175.155 121.150 175.325 ;
        RECT 120.890 175.045 121.150 175.155 ;
        RECT 121.330 175.045 121.715 175.375 ;
        RECT 121.885 175.175 122.055 175.555 ;
        RECT 122.245 175.345 122.490 175.705 ;
        RECT 123.130 175.675 123.385 176.295 ;
        RECT 123.635 176.135 123.865 176.175 ;
        RECT 124.995 176.135 125.245 176.515 ;
        RECT 123.635 175.935 125.245 176.135 ;
        RECT 123.635 175.845 123.820 175.935 ;
        RECT 124.410 175.925 125.245 175.935 ;
        RECT 125.495 175.905 125.745 176.685 ;
        RECT 125.915 175.835 126.175 176.515 ;
        RECT 123.975 175.735 124.305 175.765 ;
        RECT 123.975 175.675 125.775 175.735 ;
        RECT 123.130 175.565 125.835 175.675 ;
        RECT 123.130 175.505 124.305 175.565 ;
        RECT 125.635 175.530 125.835 175.565 ;
        RECT 121.885 175.005 122.405 175.175 ;
        RECT 123.125 175.125 123.615 175.325 ;
        RECT 123.805 175.125 124.280 175.335 ;
        RECT 122.235 174.985 122.405 175.005 ;
        RECT 119.905 174.315 120.130 174.695 ;
        RECT 120.830 174.665 122.045 174.835 ;
        RECT 120.300 174.135 120.630 174.525 ;
        RECT 120.830 174.315 121.120 174.665 ;
        RECT 121.315 174.135 121.645 174.495 ;
        RECT 121.815 174.360 122.045 174.665 ;
        RECT 122.235 174.815 122.435 174.985 ;
        RECT 122.235 174.440 122.405 174.815 ;
        RECT 123.130 174.135 123.585 174.900 ;
        RECT 124.060 174.725 124.280 175.125 ;
        RECT 124.525 175.125 124.855 175.335 ;
        RECT 124.525 174.725 124.735 175.125 ;
        RECT 125.025 175.090 125.435 175.395 ;
        RECT 125.665 174.955 125.835 175.530 ;
        RECT 125.565 174.835 125.835 174.955 ;
        RECT 124.990 174.790 125.835 174.835 ;
        RECT 124.990 174.665 125.745 174.790 ;
        RECT 124.990 174.515 125.160 174.665 ;
        RECT 126.005 174.645 126.175 175.835 ;
        RECT 126.345 175.520 126.635 176.685 ;
        RECT 126.815 175.545 127.145 176.685 ;
        RECT 127.675 175.715 128.005 176.500 ;
        RECT 128.275 176.015 128.445 176.515 ;
        RECT 128.615 176.185 128.945 176.685 ;
        RECT 128.275 175.845 128.940 176.015 ;
        RECT 127.325 175.545 128.005 175.715 ;
        RECT 126.805 175.125 127.155 175.375 ;
        RECT 127.325 174.945 127.495 175.545 ;
        RECT 127.665 175.125 128.015 175.375 ;
        RECT 128.190 175.025 128.540 175.675 ;
        RECT 125.945 174.635 126.175 174.645 ;
        RECT 123.860 174.305 125.160 174.515 ;
        RECT 125.415 174.135 125.745 174.495 ;
        RECT 125.915 174.305 126.175 174.635 ;
        RECT 126.345 174.135 126.635 174.860 ;
        RECT 126.815 174.135 127.085 174.945 ;
        RECT 127.255 174.305 127.585 174.945 ;
        RECT 127.755 174.135 127.995 174.945 ;
        RECT 128.710 174.855 128.940 175.845 ;
        RECT 128.275 174.685 128.940 174.855 ;
        RECT 128.275 174.395 128.445 174.685 ;
        RECT 128.615 174.135 128.945 174.515 ;
        RECT 129.115 174.395 129.300 176.515 ;
        RECT 129.540 176.225 129.805 176.685 ;
        RECT 129.975 176.090 130.225 176.515 ;
        RECT 130.435 176.240 131.540 176.410 ;
        RECT 129.920 175.960 130.225 176.090 ;
        RECT 129.470 174.765 129.750 175.715 ;
        RECT 129.920 174.855 130.090 175.960 ;
        RECT 130.260 175.175 130.500 175.770 ;
        RECT 130.670 175.705 131.200 176.070 ;
        RECT 130.670 175.005 130.840 175.705 ;
        RECT 131.370 175.625 131.540 176.240 ;
        RECT 131.710 175.885 131.880 176.685 ;
        RECT 132.050 176.185 132.300 176.515 ;
        RECT 132.525 176.215 133.410 176.385 ;
        RECT 131.370 175.535 131.880 175.625 ;
        RECT 129.920 174.725 130.145 174.855 ;
        RECT 130.315 174.785 130.840 175.005 ;
        RECT 131.010 175.365 131.880 175.535 ;
        RECT 129.555 174.135 129.805 174.595 ;
        RECT 129.975 174.585 130.145 174.725 ;
        RECT 131.010 174.585 131.180 175.365 ;
        RECT 131.710 175.295 131.880 175.365 ;
        RECT 131.390 175.115 131.590 175.145 ;
        RECT 132.050 175.115 132.220 176.185 ;
        RECT 132.390 175.295 132.580 176.015 ;
        RECT 131.390 174.815 132.220 175.115 ;
        RECT 132.750 175.085 133.070 176.045 ;
        RECT 129.975 174.415 130.310 174.585 ;
        RECT 130.505 174.415 131.180 174.585 ;
        RECT 131.500 174.135 131.870 174.635 ;
        RECT 132.050 174.585 132.220 174.815 ;
        RECT 132.605 174.755 133.070 175.085 ;
        RECT 133.240 175.375 133.410 176.215 ;
        RECT 133.590 176.185 133.905 176.685 ;
        RECT 134.135 175.955 134.475 176.515 ;
        RECT 133.580 175.580 134.475 175.955 ;
        RECT 134.645 175.675 134.815 176.685 ;
        RECT 134.285 175.375 134.475 175.580 ;
        RECT 134.985 175.625 135.315 176.470 ;
        RECT 135.485 175.770 135.655 176.685 ;
        RECT 136.555 175.755 136.725 176.515 ;
        RECT 136.905 175.925 137.235 176.685 ;
        RECT 134.985 175.545 135.375 175.625 ;
        RECT 136.555 175.585 137.220 175.755 ;
        RECT 137.405 175.610 137.675 176.515 ;
        RECT 135.160 175.495 135.375 175.545 ;
        RECT 133.240 175.045 134.115 175.375 ;
        RECT 134.285 175.045 135.035 175.375 ;
        RECT 133.240 174.585 133.410 175.045 ;
        RECT 134.285 174.875 134.485 175.045 ;
        RECT 135.205 174.915 135.375 175.495 ;
        RECT 137.050 175.440 137.220 175.585 ;
        RECT 136.485 175.035 136.815 175.405 ;
        RECT 137.050 175.110 137.335 175.440 ;
        RECT 135.150 174.875 135.375 174.915 ;
        RECT 132.050 174.415 132.455 174.585 ;
        RECT 132.625 174.415 133.410 174.585 ;
        RECT 133.685 174.135 133.895 174.665 ;
        RECT 134.155 174.350 134.485 174.875 ;
        RECT 134.995 174.790 135.375 174.875 ;
        RECT 137.050 174.855 137.220 175.110 ;
        RECT 134.655 174.135 134.825 174.745 ;
        RECT 134.995 174.355 135.325 174.790 ;
        RECT 136.555 174.685 137.220 174.855 ;
        RECT 137.505 174.810 137.675 175.610 ;
        RECT 137.905 175.545 138.115 176.685 ;
        RECT 138.285 175.535 138.615 176.515 ;
        RECT 138.785 175.545 139.015 176.685 ;
        RECT 139.225 176.250 144.570 176.685 ;
        RECT 135.495 174.135 135.665 174.650 ;
        RECT 136.555 174.305 136.725 174.685 ;
        RECT 136.905 174.135 137.235 174.515 ;
        RECT 137.415 174.305 137.675 174.810 ;
        RECT 137.905 174.135 138.115 174.955 ;
        RECT 138.285 174.935 138.535 175.535 ;
        RECT 138.705 175.125 139.035 175.375 ;
        RECT 138.285 174.305 138.615 174.935 ;
        RECT 138.785 174.135 139.015 174.955 ;
        RECT 140.810 174.680 141.150 175.510 ;
        RECT 142.630 175.000 142.980 176.250 ;
        RECT 144.745 175.595 148.255 176.685 ;
        RECT 144.745 174.905 146.395 175.425 ;
        RECT 146.565 175.075 148.255 175.595 ;
        RECT 148.885 175.595 150.095 176.685 ;
        RECT 148.885 175.055 149.405 175.595 ;
        RECT 139.225 174.135 144.570 174.680 ;
        RECT 144.745 174.135 148.255 174.905 ;
        RECT 149.575 174.885 150.095 175.425 ;
        RECT 148.885 174.135 150.095 174.885 ;
        RECT 36.100 173.965 150.180 174.135 ;
        RECT 36.185 173.215 37.395 173.965 ;
        RECT 36.185 172.675 36.705 173.215 ;
        RECT 37.565 173.195 41.075 173.965 ;
        RECT 42.255 173.625 42.425 173.660 ;
        RECT 42.225 173.455 42.425 173.625 ;
        RECT 36.875 172.505 37.395 173.045 ;
        RECT 37.565 172.675 39.215 173.195 ;
        RECT 42.255 173.095 42.425 173.455 ;
        RECT 42.615 173.435 42.845 173.740 ;
        RECT 43.015 173.605 43.345 173.965 ;
        RECT 43.540 173.435 43.830 173.785 ;
        RECT 42.615 173.265 43.830 173.435 ;
        RECT 44.005 173.215 45.215 173.965 ;
        RECT 45.385 173.315 45.645 173.795 ;
        RECT 45.815 173.425 46.065 173.965 ;
        RECT 39.385 172.505 41.075 173.025 ;
        RECT 42.255 172.925 42.775 173.095 ;
        RECT 36.185 171.415 37.395 172.505 ;
        RECT 37.565 171.415 41.075 172.505 ;
        RECT 42.170 172.395 42.415 172.755 ;
        RECT 42.605 172.545 42.775 172.925 ;
        RECT 42.945 172.725 43.330 173.055 ;
        RECT 43.510 172.945 43.770 173.055 ;
        RECT 43.510 172.775 43.775 172.945 ;
        RECT 43.510 172.725 43.770 172.775 ;
        RECT 42.605 172.265 42.955 172.545 ;
        RECT 42.170 171.415 42.425 172.215 ;
        RECT 42.625 171.585 42.955 172.265 ;
        RECT 43.135 171.675 43.330 172.725 ;
        RECT 44.005 172.675 44.525 173.215 ;
        RECT 43.510 171.415 43.830 172.555 ;
        RECT 44.695 172.505 45.215 173.045 ;
        RECT 44.005 171.415 45.215 172.505 ;
        RECT 45.385 172.285 45.555 173.315 ;
        RECT 46.235 173.260 46.455 173.745 ;
        RECT 45.725 172.665 45.955 173.060 ;
        RECT 46.125 172.835 46.455 173.260 ;
        RECT 46.625 173.585 47.515 173.755 ;
        RECT 46.625 172.860 46.795 173.585 ;
        RECT 47.775 173.415 47.945 173.795 ;
        RECT 48.125 173.585 48.455 173.965 ;
        RECT 46.965 173.030 47.515 173.415 ;
        RECT 47.775 173.245 48.440 173.415 ;
        RECT 48.635 173.290 48.895 173.795 ;
        RECT 46.625 172.790 47.515 172.860 ;
        RECT 46.620 172.765 47.515 172.790 ;
        RECT 46.610 172.750 47.515 172.765 ;
        RECT 46.605 172.735 47.515 172.750 ;
        RECT 46.595 172.730 47.515 172.735 ;
        RECT 46.590 172.720 47.515 172.730 ;
        RECT 46.585 172.710 47.515 172.720 ;
        RECT 46.575 172.705 47.515 172.710 ;
        RECT 46.565 172.695 47.515 172.705 ;
        RECT 47.705 172.695 48.045 173.065 ;
        RECT 48.270 172.990 48.440 173.245 ;
        RECT 46.555 172.690 47.515 172.695 ;
        RECT 46.555 172.685 46.890 172.690 ;
        RECT 46.540 172.680 46.890 172.685 ;
        RECT 46.525 172.670 46.890 172.680 ;
        RECT 46.500 172.665 46.890 172.670 ;
        RECT 45.725 172.660 46.890 172.665 ;
        RECT 45.725 172.625 46.860 172.660 ;
        RECT 45.725 172.600 46.825 172.625 ;
        RECT 45.725 172.570 46.795 172.600 ;
        RECT 45.725 172.540 46.775 172.570 ;
        RECT 45.725 172.510 46.755 172.540 ;
        RECT 45.725 172.500 46.685 172.510 ;
        RECT 45.725 172.490 46.660 172.500 ;
        RECT 45.725 172.475 46.640 172.490 ;
        RECT 45.725 172.460 46.620 172.475 ;
        RECT 45.830 172.450 46.615 172.460 ;
        RECT 45.830 172.415 46.600 172.450 ;
        RECT 45.385 171.585 45.660 172.285 ;
        RECT 45.830 172.165 46.585 172.415 ;
        RECT 46.755 172.095 47.085 172.340 ;
        RECT 47.255 172.240 47.515 172.690 ;
        RECT 48.270 172.660 48.545 172.990 ;
        RECT 48.270 172.515 48.440 172.660 ;
        RECT 47.765 172.345 48.440 172.515 ;
        RECT 48.715 172.490 48.895 173.290 ;
        RECT 49.065 173.165 49.375 173.965 ;
        RECT 49.580 173.165 50.275 173.795 ;
        RECT 50.535 173.415 50.705 173.795 ;
        RECT 50.885 173.585 51.215 173.965 ;
        RECT 50.535 173.245 51.200 173.415 ;
        RECT 51.395 173.290 51.655 173.795 ;
        RECT 49.075 172.725 49.410 172.995 ;
        RECT 49.580 172.565 49.750 173.165 ;
        RECT 49.920 172.725 50.255 172.975 ;
        RECT 50.465 172.695 50.805 173.065 ;
        RECT 51.030 172.990 51.200 173.245 ;
        RECT 51.030 172.660 51.305 172.990 ;
        RECT 46.900 172.070 47.085 172.095 ;
        RECT 46.900 171.970 47.515 172.070 ;
        RECT 45.830 171.415 46.085 171.960 ;
        RECT 46.255 171.585 46.735 171.925 ;
        RECT 46.910 171.415 47.515 171.970 ;
        RECT 47.765 171.585 47.945 172.345 ;
        RECT 48.125 171.415 48.455 172.175 ;
        RECT 48.625 171.585 48.895 172.490 ;
        RECT 49.065 171.415 49.345 172.555 ;
        RECT 49.515 171.585 49.845 172.565 ;
        RECT 50.015 171.415 50.275 172.555 ;
        RECT 51.030 172.515 51.200 172.660 ;
        RECT 50.525 172.345 51.200 172.515 ;
        RECT 51.475 172.490 51.655 173.290 ;
        RECT 50.525 171.585 50.705 172.345 ;
        RECT 50.885 171.415 51.215 172.175 ;
        RECT 51.385 171.585 51.655 172.490 ;
        RECT 52.285 173.290 52.545 173.795 ;
        RECT 52.725 173.585 53.055 173.965 ;
        RECT 53.235 173.415 53.405 173.795 ;
        RECT 52.285 172.490 52.465 173.290 ;
        RECT 52.740 173.245 53.405 173.415 ;
        RECT 54.215 173.415 54.385 173.795 ;
        RECT 54.565 173.585 54.895 173.965 ;
        RECT 54.215 173.245 54.880 173.415 ;
        RECT 55.075 173.290 55.335 173.795 ;
        RECT 52.740 172.990 52.910 173.245 ;
        RECT 52.635 172.660 52.910 172.990 ;
        RECT 53.135 172.695 53.475 173.065 ;
        RECT 54.145 172.695 54.485 173.065 ;
        RECT 54.710 172.990 54.880 173.245 ;
        RECT 52.740 172.515 52.910 172.660 ;
        RECT 54.710 172.660 54.985 172.990 ;
        RECT 54.710 172.515 54.880 172.660 ;
        RECT 52.285 171.585 52.555 172.490 ;
        RECT 52.740 172.345 53.415 172.515 ;
        RECT 52.725 171.415 53.055 172.175 ;
        RECT 53.235 171.585 53.415 172.345 ;
        RECT 54.205 172.345 54.880 172.515 ;
        RECT 55.155 172.490 55.335 173.290 ;
        RECT 54.205 171.585 54.385 172.345 ;
        RECT 54.565 171.415 54.895 172.175 ;
        RECT 55.065 171.585 55.335 172.490 ;
        RECT 55.505 173.290 55.765 173.795 ;
        RECT 55.945 173.585 56.275 173.965 ;
        RECT 56.455 173.415 56.625 173.795 ;
        RECT 55.505 172.490 55.685 173.290 ;
        RECT 55.960 173.245 56.625 173.415 ;
        RECT 55.960 172.990 56.130 173.245 ;
        RECT 56.885 173.195 60.395 173.965 ;
        RECT 60.565 173.215 61.775 173.965 ;
        RECT 61.945 173.240 62.235 173.965 ;
        RECT 62.405 173.215 63.615 173.965 ;
        RECT 63.870 173.415 64.045 173.705 ;
        RECT 64.215 173.585 64.545 173.965 ;
        RECT 63.870 173.245 64.365 173.415 ;
        RECT 64.720 173.285 64.935 173.655 ;
        RECT 65.170 173.515 65.770 173.685 ;
        RECT 55.855 172.660 56.130 172.990 ;
        RECT 56.355 172.695 56.695 173.065 ;
        RECT 56.885 172.675 58.535 173.195 ;
        RECT 55.960 172.515 56.130 172.660 ;
        RECT 55.505 171.585 55.775 172.490 ;
        RECT 55.960 172.345 56.635 172.515 ;
        RECT 58.705 172.505 60.395 173.025 ;
        RECT 60.565 172.675 61.085 173.215 ;
        RECT 61.255 172.505 61.775 173.045 ;
        RECT 62.405 172.675 62.925 173.215 ;
        RECT 55.945 171.415 56.275 172.175 ;
        RECT 56.455 171.585 56.635 172.345 ;
        RECT 56.885 171.415 60.395 172.505 ;
        RECT 60.565 171.415 61.775 172.505 ;
        RECT 61.945 171.415 62.235 172.580 ;
        RECT 63.095 172.505 63.615 173.045 ;
        RECT 62.405 171.415 63.615 172.505 ;
        RECT 63.845 172.305 64.025 173.075 ;
        RECT 64.195 172.265 64.365 173.245 ;
        RECT 64.535 172.955 64.935 173.285 ;
        RECT 65.105 173.015 65.430 173.345 ;
        RECT 64.920 172.605 65.090 172.765 ;
        RECT 64.705 172.435 65.090 172.605 ;
        RECT 65.260 172.475 65.430 173.015 ;
        RECT 65.600 172.815 65.770 173.515 ;
        RECT 66.150 173.505 66.480 173.965 ;
        RECT 66.685 173.585 67.115 173.755 ;
        RECT 65.940 173.035 66.315 173.335 ;
        RECT 65.600 172.645 65.940 172.815 ;
        RECT 66.110 172.730 66.315 173.035 ;
        RECT 66.485 172.730 66.775 173.335 ;
        RECT 66.945 172.990 67.115 173.585 ;
        RECT 67.285 173.375 67.520 173.705 ;
        RECT 65.260 172.265 65.600 172.475 ;
        RECT 64.195 172.135 65.600 172.265 ;
        RECT 63.875 172.095 65.600 172.135 ;
        RECT 63.875 171.965 64.365 172.095 ;
        RECT 63.875 171.675 64.045 171.965 ;
        RECT 65.770 171.925 65.940 172.645 ;
        RECT 66.945 172.660 67.180 172.990 ;
        RECT 66.945 172.560 67.115 172.660 ;
        RECT 66.845 172.390 67.115 172.560 ;
        RECT 66.845 172.265 67.015 172.390 ;
        RECT 66.670 172.095 67.015 172.265 ;
        RECT 67.350 172.240 67.520 173.375 ;
        RECT 64.215 171.415 64.545 171.795 ;
        RECT 65.110 171.755 65.940 171.925 ;
        RECT 66.295 171.415 66.525 171.995 ;
        RECT 67.265 171.925 67.520 172.240 ;
        RECT 67.005 171.755 67.520 171.925 ;
        RECT 67.690 171.925 67.880 173.705 ;
        RECT 68.095 173.465 68.300 173.795 ;
        RECT 68.495 173.505 68.825 173.965 ;
        RECT 69.025 173.585 69.920 173.755 ;
        RECT 68.095 172.485 68.265 173.465 ;
        RECT 68.445 172.655 68.815 173.335 ;
        RECT 69.025 172.485 69.195 173.585 ;
        RECT 68.095 172.315 69.195 172.485 ;
        RECT 68.095 172.155 68.285 172.315 ;
        RECT 67.690 171.755 68.215 171.925 ;
        RECT 68.455 171.415 68.800 172.045 ;
        RECT 69.025 171.895 69.195 172.315 ;
        RECT 69.365 173.015 69.985 173.345 ;
        RECT 70.235 173.055 70.545 173.675 ;
        RECT 70.715 173.235 70.965 173.965 ;
        RECT 71.135 173.325 71.465 173.785 ;
        RECT 69.365 172.065 69.655 173.015 ;
        RECT 70.235 172.975 70.645 173.055 ;
        RECT 69.825 172.405 70.165 172.805 ;
        RECT 70.335 172.725 70.645 172.975 ;
        RECT 70.815 172.725 71.125 173.055 ;
        RECT 70.815 172.555 70.985 172.725 ;
        RECT 71.295 172.555 71.465 173.325 ;
        RECT 71.635 173.165 71.890 173.965 ;
        RECT 72.615 173.415 72.785 173.795 ;
        RECT 72.965 173.585 73.295 173.965 ;
        RECT 72.615 173.245 73.280 173.415 ;
        RECT 73.475 173.290 73.735 173.795 ;
        RECT 72.545 172.695 72.885 173.065 ;
        RECT 73.110 172.990 73.280 173.245 ;
        RECT 73.110 172.660 73.385 172.990 ;
        RECT 70.375 172.385 70.985 172.555 ;
        RECT 70.375 171.925 70.545 172.385 ;
        RECT 71.155 172.215 71.465 172.555 ;
        RECT 69.025 171.725 69.975 171.895 ;
        RECT 70.225 171.755 70.545 171.925 ;
        RECT 70.715 171.415 70.885 172.215 ;
        RECT 71.055 171.595 71.465 172.215 ;
        RECT 71.635 171.415 71.885 172.555 ;
        RECT 73.110 172.515 73.280 172.660 ;
        RECT 72.605 172.345 73.280 172.515 ;
        RECT 73.555 172.490 73.735 173.290 ;
        RECT 73.995 173.415 74.165 173.705 ;
        RECT 74.335 173.585 74.665 173.965 ;
        RECT 73.995 173.245 74.660 173.415 ;
        RECT 72.605 171.585 72.785 172.345 ;
        RECT 72.965 171.415 73.295 172.175 ;
        RECT 73.465 171.585 73.735 172.490 ;
        RECT 73.910 172.425 74.260 173.075 ;
        RECT 74.430 172.255 74.660 173.245 ;
        RECT 73.995 172.085 74.660 172.255 ;
        RECT 73.995 171.585 74.165 172.085 ;
        RECT 74.335 171.415 74.665 171.915 ;
        RECT 74.835 171.585 75.020 173.705 ;
        RECT 75.275 173.505 75.525 173.965 ;
        RECT 75.695 173.515 76.030 173.685 ;
        RECT 76.225 173.515 76.900 173.685 ;
        RECT 75.695 173.375 75.865 173.515 ;
        RECT 75.190 172.385 75.470 173.335 ;
        RECT 75.640 173.245 75.865 173.375 ;
        RECT 75.640 172.140 75.810 173.245 ;
        RECT 76.035 173.095 76.560 173.315 ;
        RECT 75.980 172.330 76.220 172.925 ;
        RECT 76.390 172.395 76.560 173.095 ;
        RECT 76.730 172.735 76.900 173.515 ;
        RECT 77.220 173.465 77.590 173.965 ;
        RECT 77.770 173.515 78.175 173.685 ;
        RECT 78.345 173.515 79.130 173.685 ;
        RECT 77.770 173.285 77.940 173.515 ;
        RECT 77.110 172.985 77.940 173.285 ;
        RECT 78.325 173.015 78.790 173.345 ;
        RECT 77.110 172.955 77.310 172.985 ;
        RECT 77.430 172.735 77.600 172.805 ;
        RECT 76.730 172.565 77.600 172.735 ;
        RECT 77.090 172.475 77.600 172.565 ;
        RECT 75.640 172.010 75.945 172.140 ;
        RECT 76.390 172.030 76.920 172.395 ;
        RECT 75.260 171.415 75.525 171.875 ;
        RECT 75.695 171.585 75.945 172.010 ;
        RECT 77.090 171.860 77.260 172.475 ;
        RECT 76.155 171.690 77.260 171.860 ;
        RECT 77.430 171.415 77.600 172.215 ;
        RECT 77.770 171.915 77.940 172.985 ;
        RECT 78.110 172.085 78.300 172.805 ;
        RECT 78.470 172.055 78.790 173.015 ;
        RECT 78.960 173.055 79.130 173.515 ;
        RECT 79.405 173.435 79.615 173.965 ;
        RECT 79.875 173.225 80.205 173.750 ;
        RECT 80.375 173.355 80.545 173.965 ;
        RECT 80.715 173.310 81.045 173.745 ;
        RECT 80.715 173.225 81.095 173.310 ;
        RECT 80.005 173.055 80.205 173.225 ;
        RECT 80.870 173.185 81.095 173.225 ;
        RECT 78.960 172.725 79.835 173.055 ;
        RECT 80.005 172.725 80.755 173.055 ;
        RECT 77.770 171.585 78.020 171.915 ;
        RECT 78.960 171.885 79.130 172.725 ;
        RECT 80.005 172.520 80.195 172.725 ;
        RECT 80.925 172.605 81.095 173.185 ;
        RECT 81.265 173.195 84.775 173.965 ;
        RECT 84.945 173.215 86.155 173.965 ;
        RECT 81.265 172.675 82.915 173.195 ;
        RECT 80.880 172.555 81.095 172.605 ;
        RECT 79.300 172.145 80.195 172.520 ;
        RECT 80.705 172.475 81.095 172.555 ;
        RECT 83.085 172.505 84.775 173.025 ;
        RECT 84.945 172.675 85.465 173.215 ;
        RECT 86.325 173.165 86.635 173.965 ;
        RECT 86.840 173.165 87.535 173.795 ;
        RECT 87.705 173.240 87.995 173.965 ;
        RECT 88.325 173.405 88.655 173.795 ;
        RECT 88.825 173.575 90.010 173.745 ;
        RECT 90.270 173.495 90.440 173.965 ;
        RECT 88.325 173.225 88.835 173.405 ;
        RECT 85.635 172.505 86.155 173.045 ;
        RECT 86.335 172.725 86.670 172.995 ;
        RECT 86.840 172.565 87.010 173.165 ;
        RECT 87.180 172.725 87.515 172.975 ;
        RECT 88.165 172.765 88.495 173.055 ;
        RECT 88.665 172.595 88.835 173.225 ;
        RECT 89.240 173.315 89.625 173.405 ;
        RECT 90.610 173.315 90.940 173.780 ;
        RECT 89.240 173.145 90.940 173.315 ;
        RECT 91.110 173.145 91.280 173.965 ;
        RECT 91.450 173.145 92.135 173.785 ;
        RECT 89.005 172.765 89.335 172.975 ;
        RECT 89.515 172.725 89.895 172.975 ;
        RECT 90.085 172.945 90.570 172.975 ;
        RECT 90.065 172.775 90.570 172.945 ;
        RECT 78.245 171.715 79.130 171.885 ;
        RECT 79.310 171.415 79.625 171.915 ;
        RECT 79.855 171.585 80.195 172.145 ;
        RECT 80.365 171.415 80.535 172.425 ;
        RECT 80.705 171.630 81.035 172.475 ;
        RECT 81.265 171.415 84.775 172.505 ;
        RECT 84.945 171.415 86.155 172.505 ;
        RECT 86.325 171.415 86.605 172.555 ;
        RECT 86.775 171.585 87.105 172.565 ;
        RECT 87.275 171.415 87.535 172.555 ;
        RECT 87.705 171.415 87.995 172.580 ;
        RECT 88.320 172.425 89.405 172.595 ;
        RECT 88.320 171.585 88.620 172.425 ;
        RECT 88.815 171.415 89.065 172.255 ;
        RECT 89.235 172.175 89.405 172.425 ;
        RECT 89.575 172.345 89.895 172.725 ;
        RECT 90.085 172.765 90.570 172.775 ;
        RECT 90.760 172.765 91.210 172.975 ;
        RECT 91.380 172.765 91.715 172.975 ;
        RECT 90.085 172.345 90.460 172.765 ;
        RECT 91.380 172.595 91.550 172.765 ;
        RECT 90.630 172.425 91.550 172.595 ;
        RECT 90.630 172.175 90.800 172.425 ;
        RECT 89.235 172.005 90.800 172.175 ;
        RECT 89.655 171.585 90.460 172.005 ;
        RECT 90.970 171.415 91.300 172.255 ;
        RECT 91.885 172.175 92.135 173.145 ;
        RECT 91.470 171.585 92.135 172.175 ;
        RECT 92.315 173.240 92.645 173.750 ;
        RECT 92.815 173.565 93.145 173.965 ;
        RECT 94.195 173.395 94.525 173.735 ;
        RECT 94.695 173.565 95.025 173.965 ;
        RECT 92.315 172.475 92.505 173.240 ;
        RECT 92.815 173.225 95.180 173.395 ;
        RECT 92.815 173.055 92.985 173.225 ;
        RECT 92.675 172.725 92.985 173.055 ;
        RECT 93.155 172.725 93.460 173.055 ;
        RECT 92.315 171.625 92.645 172.475 ;
        RECT 92.815 171.415 93.065 172.555 ;
        RECT 93.245 172.395 93.460 172.725 ;
        RECT 93.635 172.395 93.920 173.055 ;
        RECT 94.115 172.395 94.380 173.055 ;
        RECT 94.595 172.395 94.840 173.055 ;
        RECT 95.010 172.225 95.180 173.225 ;
        RECT 95.525 173.195 99.035 173.965 ;
        RECT 99.825 173.405 100.155 173.795 ;
        RECT 100.325 173.575 101.510 173.745 ;
        RECT 101.770 173.495 101.940 173.965 ;
        RECT 99.825 173.225 100.335 173.405 ;
        RECT 95.525 172.675 97.175 173.195 ;
        RECT 97.345 172.505 99.035 173.025 ;
        RECT 99.665 172.765 99.995 173.055 ;
        RECT 100.165 172.595 100.335 173.225 ;
        RECT 100.740 173.315 101.125 173.405 ;
        RECT 102.110 173.315 102.440 173.780 ;
        RECT 100.740 173.145 102.440 173.315 ;
        RECT 102.610 173.145 102.780 173.965 ;
        RECT 102.950 173.145 103.635 173.785 ;
        RECT 103.805 173.165 104.115 173.965 ;
        RECT 104.320 173.165 105.015 173.795 ;
        RECT 106.105 173.335 106.445 173.795 ;
        RECT 106.615 173.505 106.785 173.965 ;
        RECT 107.415 173.530 107.775 173.795 ;
        RECT 107.420 173.525 107.775 173.530 ;
        RECT 107.425 173.515 107.775 173.525 ;
        RECT 107.430 173.510 107.775 173.515 ;
        RECT 107.435 173.500 107.775 173.510 ;
        RECT 108.015 173.505 108.185 173.965 ;
        RECT 107.440 173.495 107.775 173.500 ;
        RECT 107.450 173.485 107.775 173.495 ;
        RECT 107.460 173.475 107.775 173.485 ;
        RECT 106.955 173.335 107.285 173.415 ;
        RECT 100.505 172.765 100.835 172.975 ;
        RECT 101.015 172.725 101.395 172.975 ;
        RECT 93.255 172.055 94.545 172.225 ;
        RECT 93.255 171.635 93.505 172.055 ;
        RECT 93.735 171.415 94.065 171.885 ;
        RECT 94.295 171.635 94.545 172.055 ;
        RECT 94.725 172.055 95.180 172.225 ;
        RECT 94.725 171.625 95.055 172.055 ;
        RECT 95.525 171.415 99.035 172.505 ;
        RECT 99.820 172.425 100.905 172.595 ;
        RECT 99.820 171.585 100.120 172.425 ;
        RECT 100.315 171.415 100.565 172.255 ;
        RECT 100.735 172.175 100.905 172.425 ;
        RECT 101.075 172.345 101.395 172.725 ;
        RECT 101.585 172.765 102.070 172.975 ;
        RECT 102.260 172.765 102.710 172.975 ;
        RECT 102.880 172.765 103.215 172.975 ;
        RECT 101.585 172.605 101.960 172.765 ;
        RECT 101.565 172.435 101.960 172.605 ;
        RECT 102.880 172.595 103.050 172.765 ;
        RECT 101.585 172.345 101.960 172.435 ;
        RECT 102.130 172.425 103.050 172.595 ;
        RECT 102.130 172.175 102.300 172.425 ;
        RECT 100.735 172.005 102.300 172.175 ;
        RECT 101.155 171.585 101.960 172.005 ;
        RECT 102.470 171.415 102.800 172.255 ;
        RECT 103.385 172.175 103.635 173.145 ;
        RECT 103.815 172.725 104.150 172.995 ;
        RECT 104.320 172.565 104.490 173.165 ;
        RECT 106.105 173.145 107.285 173.335 ;
        RECT 107.475 173.335 107.775 173.475 ;
        RECT 107.475 173.145 108.185 173.335 ;
        RECT 104.660 172.725 104.995 172.975 ;
        RECT 106.105 172.775 106.435 172.975 ;
        RECT 106.745 172.955 107.075 172.975 ;
        RECT 106.625 172.775 107.075 172.955 ;
        RECT 102.970 171.585 103.635 172.175 ;
        RECT 103.805 171.415 104.085 172.555 ;
        RECT 104.255 171.585 104.585 172.565 ;
        RECT 104.755 171.415 105.015 172.555 ;
        RECT 106.105 172.435 106.335 172.775 ;
        RECT 106.115 171.415 106.445 172.135 ;
        RECT 106.625 171.660 106.840 172.775 ;
        RECT 107.245 172.745 107.715 172.975 ;
        RECT 107.900 172.575 108.185 173.145 ;
        RECT 108.355 173.020 108.695 173.795 ;
        RECT 107.035 172.360 108.185 172.575 ;
        RECT 107.035 171.585 107.365 172.360 ;
        RECT 107.535 171.415 108.245 172.190 ;
        RECT 108.415 171.585 108.695 173.020 ;
        RECT 108.865 173.195 112.375 173.965 ;
        RECT 113.465 173.240 113.755 173.965 ;
        RECT 113.925 173.195 115.595 173.965 ;
        RECT 116.315 173.415 116.485 173.795 ;
        RECT 116.665 173.585 116.995 173.965 ;
        RECT 116.315 173.245 116.980 173.415 ;
        RECT 117.175 173.290 117.435 173.795 ;
        RECT 108.865 172.675 110.515 173.195 ;
        RECT 110.685 172.505 112.375 173.025 ;
        RECT 113.925 172.675 114.675 173.195 ;
        RECT 108.865 171.415 112.375 172.505 ;
        RECT 113.465 171.415 113.755 172.580 ;
        RECT 114.845 172.505 115.595 173.025 ;
        RECT 116.245 172.695 116.585 173.065 ;
        RECT 116.810 172.990 116.980 173.245 ;
        RECT 116.810 172.660 117.085 172.990 ;
        RECT 116.810 172.515 116.980 172.660 ;
        RECT 113.925 171.415 115.595 172.505 ;
        RECT 116.305 172.345 116.980 172.515 ;
        RECT 117.255 172.490 117.435 173.290 ;
        RECT 117.605 173.195 119.275 173.965 ;
        RECT 119.930 173.575 120.260 173.965 ;
        RECT 120.430 173.405 120.655 173.785 ;
        RECT 117.605 172.675 118.355 173.195 ;
        RECT 118.525 172.505 119.275 173.025 ;
        RECT 119.915 172.725 120.155 173.375 ;
        RECT 120.325 173.225 120.655 173.405 ;
        RECT 120.325 172.555 120.500 173.225 ;
        RECT 120.855 173.055 121.085 173.675 ;
        RECT 121.265 173.235 121.565 173.965 ;
        RECT 121.745 173.420 127.090 173.965 ;
        RECT 127.265 173.420 132.610 173.965 ;
        RECT 120.670 172.725 121.085 173.055 ;
        RECT 121.265 172.725 121.560 173.055 ;
        RECT 123.330 172.590 123.670 173.420 ;
        RECT 116.305 171.585 116.485 172.345 ;
        RECT 116.665 171.415 116.995 172.175 ;
        RECT 117.165 171.585 117.435 172.490 ;
        RECT 117.605 171.415 119.275 172.505 ;
        RECT 119.915 172.365 120.500 172.555 ;
        RECT 119.915 171.595 120.190 172.365 ;
        RECT 120.670 172.195 121.565 172.525 ;
        RECT 120.360 172.025 121.565 172.195 ;
        RECT 120.360 171.595 120.690 172.025 ;
        RECT 120.860 171.415 121.055 171.855 ;
        RECT 121.235 171.595 121.565 172.025 ;
        RECT 125.150 171.850 125.500 173.100 ;
        RECT 128.850 172.590 129.190 173.420 ;
        RECT 132.785 173.195 136.295 173.965 ;
        RECT 136.465 173.215 137.675 173.965 ;
        RECT 137.845 173.290 138.105 173.795 ;
        RECT 138.285 173.585 138.615 173.965 ;
        RECT 138.795 173.415 138.965 173.795 ;
        RECT 130.670 171.850 131.020 173.100 ;
        RECT 132.785 172.675 134.435 173.195 ;
        RECT 134.605 172.505 136.295 173.025 ;
        RECT 136.465 172.675 136.985 173.215 ;
        RECT 137.155 172.505 137.675 173.045 ;
        RECT 121.745 171.415 127.090 171.850 ;
        RECT 127.265 171.415 132.610 171.850 ;
        RECT 132.785 171.415 136.295 172.505 ;
        RECT 136.465 171.415 137.675 172.505 ;
        RECT 137.845 172.490 138.025 173.290 ;
        RECT 138.300 173.245 138.965 173.415 ;
        RECT 138.300 172.990 138.470 173.245 ;
        RECT 139.225 173.240 139.515 173.965 ;
        RECT 139.685 173.165 140.025 173.795 ;
        RECT 140.315 173.505 140.485 173.965 ;
        RECT 140.755 173.335 141.085 173.780 ;
        RECT 138.195 172.660 138.470 172.990 ;
        RECT 138.695 172.695 139.035 173.065 ;
        RECT 138.300 172.515 138.470 172.660 ;
        RECT 139.685 172.595 139.955 173.165 ;
        RECT 140.335 173.145 141.085 173.335 ;
        RECT 141.255 173.315 141.425 173.635 ;
        RECT 141.650 173.505 141.980 173.965 ;
        RECT 142.180 173.315 142.510 173.795 ;
        RECT 142.725 173.505 143.055 173.965 ;
        RECT 143.225 173.315 143.555 173.795 ;
        RECT 141.255 173.145 143.555 173.315 ;
        RECT 143.825 173.195 147.335 173.965 ;
        RECT 147.505 173.215 148.715 173.965 ;
        RECT 148.885 173.215 150.095 173.965 ;
        RECT 140.335 172.975 140.705 173.145 ;
        RECT 140.125 172.765 140.705 172.975 ;
        RECT 140.875 172.765 141.295 172.975 ;
        RECT 140.445 172.595 140.705 172.765 ;
        RECT 137.845 171.585 138.115 172.490 ;
        RECT 138.300 172.345 138.975 172.515 ;
        RECT 138.285 171.415 138.615 172.175 ;
        RECT 138.795 171.585 138.975 172.345 ;
        RECT 139.225 171.415 139.515 172.580 ;
        RECT 139.685 171.585 140.210 172.595 ;
        RECT 140.445 172.305 141.195 172.595 ;
        RECT 140.445 171.415 140.775 172.135 ;
        RECT 140.945 171.585 141.195 172.305 ;
        RECT 141.465 171.660 141.795 172.975 ;
        RECT 142.005 171.660 142.335 172.975 ;
        RECT 142.505 171.660 142.875 172.975 ;
        RECT 143.085 172.725 143.595 172.975 ;
        RECT 143.825 172.675 145.475 173.195 ;
        RECT 143.205 171.415 143.535 172.535 ;
        RECT 145.645 172.505 147.335 173.025 ;
        RECT 147.505 172.675 148.025 173.215 ;
        RECT 148.195 172.505 148.715 173.045 ;
        RECT 143.825 171.415 147.335 172.505 ;
        RECT 147.505 171.415 148.715 172.505 ;
        RECT 148.885 172.505 149.405 173.045 ;
        RECT 149.575 172.675 150.095 173.215 ;
        RECT 148.885 171.415 150.095 172.505 ;
        RECT 36.100 171.245 150.180 171.415 ;
        RECT 36.185 170.155 37.395 171.245 ;
        RECT 37.565 170.155 40.155 171.245 ;
        RECT 36.185 169.445 36.705 169.985 ;
        RECT 36.875 169.615 37.395 170.155 ;
        RECT 37.565 169.465 38.775 169.985 ;
        RECT 38.945 169.635 40.155 170.155 ;
        RECT 40.790 170.105 41.110 171.245 ;
        RECT 41.290 169.935 41.485 170.985 ;
        RECT 41.665 170.395 41.995 171.075 ;
        RECT 42.195 170.445 42.450 171.245 ;
        RECT 42.825 170.575 43.105 171.245 ;
        RECT 41.665 170.115 42.015 170.395 ;
        RECT 43.275 170.355 43.575 170.905 ;
        RECT 43.775 170.525 44.105 171.245 ;
        RECT 44.295 170.525 44.755 171.075 ;
        RECT 40.850 169.885 41.110 169.935 ;
        RECT 40.845 169.715 41.110 169.885 ;
        RECT 40.850 169.605 41.110 169.715 ;
        RECT 41.290 169.605 41.675 169.935 ;
        RECT 41.845 169.735 42.015 170.115 ;
        RECT 42.205 169.905 42.450 170.265 ;
        RECT 42.640 169.935 42.905 170.295 ;
        RECT 43.275 170.185 44.215 170.355 ;
        RECT 44.045 169.935 44.215 170.185 ;
        RECT 41.845 169.565 42.365 169.735 ;
        RECT 42.640 169.685 43.315 169.935 ;
        RECT 43.535 169.685 43.875 169.935 ;
        RECT 42.195 169.545 42.365 169.565 ;
        RECT 44.045 169.605 44.335 169.935 ;
        RECT 36.185 168.695 37.395 169.445 ;
        RECT 37.565 168.695 40.155 169.465 ;
        RECT 40.790 169.225 42.005 169.395 ;
        RECT 40.790 168.875 41.080 169.225 ;
        RECT 41.275 168.695 41.605 169.055 ;
        RECT 41.775 168.920 42.005 169.225 ;
        RECT 42.195 169.375 42.395 169.545 ;
        RECT 44.045 169.515 44.215 169.605 ;
        RECT 42.195 169.000 42.365 169.375 ;
        RECT 42.825 169.325 44.215 169.515 ;
        RECT 42.825 168.965 43.155 169.325 ;
        RECT 44.505 169.155 44.755 170.525 ;
        RECT 44.935 170.105 45.265 171.245 ;
        RECT 45.795 170.275 46.125 171.060 ;
        RECT 45.445 170.105 46.125 170.275 ;
        RECT 46.305 170.375 46.580 171.075 ;
        RECT 46.750 170.700 47.005 171.245 ;
        RECT 47.175 170.735 47.655 171.075 ;
        RECT 47.830 170.690 48.435 171.245 ;
        RECT 47.820 170.590 48.435 170.690 ;
        RECT 47.820 170.565 48.005 170.590 ;
        RECT 44.925 169.685 45.275 169.935 ;
        RECT 45.445 169.505 45.615 170.105 ;
        RECT 45.785 169.685 46.135 169.935 ;
        RECT 43.775 168.695 44.025 169.155 ;
        RECT 44.195 168.865 44.755 169.155 ;
        RECT 44.935 168.695 45.205 169.505 ;
        RECT 45.375 168.865 45.705 169.505 ;
        RECT 45.875 168.695 46.115 169.505 ;
        RECT 46.305 169.345 46.475 170.375 ;
        RECT 46.750 170.245 47.505 170.495 ;
        RECT 47.675 170.320 48.005 170.565 ;
        RECT 46.750 170.210 47.520 170.245 ;
        RECT 46.750 170.200 47.535 170.210 ;
        RECT 46.645 170.185 47.540 170.200 ;
        RECT 46.645 170.170 47.560 170.185 ;
        RECT 46.645 170.160 47.580 170.170 ;
        RECT 46.645 170.150 47.605 170.160 ;
        RECT 46.645 170.120 47.675 170.150 ;
        RECT 46.645 170.090 47.695 170.120 ;
        RECT 46.645 170.060 47.715 170.090 ;
        RECT 46.645 170.035 47.745 170.060 ;
        RECT 46.645 170.000 47.780 170.035 ;
        RECT 46.645 169.995 47.810 170.000 ;
        RECT 46.645 169.600 46.875 169.995 ;
        RECT 47.420 169.990 47.810 169.995 ;
        RECT 47.445 169.980 47.810 169.990 ;
        RECT 47.460 169.975 47.810 169.980 ;
        RECT 47.475 169.970 47.810 169.975 ;
        RECT 48.175 169.970 48.435 170.420 ;
        RECT 49.065 170.080 49.355 171.245 ;
        RECT 49.525 170.810 54.870 171.245 ;
        RECT 55.045 170.810 60.390 171.245 ;
        RECT 47.475 169.965 48.435 169.970 ;
        RECT 47.485 169.955 48.435 169.965 ;
        RECT 47.495 169.950 48.435 169.955 ;
        RECT 47.505 169.940 48.435 169.950 ;
        RECT 47.510 169.930 48.435 169.940 ;
        RECT 47.515 169.925 48.435 169.930 ;
        RECT 47.525 169.910 48.435 169.925 ;
        RECT 47.530 169.895 48.435 169.910 ;
        RECT 47.540 169.870 48.435 169.895 ;
        RECT 47.045 169.400 47.375 169.825 ;
        RECT 46.305 168.865 46.565 169.345 ;
        RECT 46.735 168.695 46.985 169.235 ;
        RECT 47.155 168.915 47.375 169.400 ;
        RECT 47.545 169.800 48.435 169.870 ;
        RECT 47.545 169.075 47.715 169.800 ;
        RECT 47.885 169.245 48.435 169.630 ;
        RECT 47.545 168.905 48.435 169.075 ;
        RECT 49.065 168.695 49.355 169.420 ;
        RECT 51.110 169.240 51.450 170.070 ;
        RECT 52.930 169.560 53.280 170.810 ;
        RECT 56.630 169.240 56.970 170.070 ;
        RECT 58.450 169.560 58.800 170.810 ;
        RECT 61.105 170.315 61.285 171.075 ;
        RECT 61.465 170.485 61.795 171.245 ;
        RECT 61.105 170.145 61.780 170.315 ;
        RECT 61.965 170.170 62.235 171.075 ;
        RECT 62.495 170.695 62.665 170.985 ;
        RECT 62.835 170.865 63.165 171.245 ;
        RECT 63.730 170.735 64.560 170.905 ;
        RECT 62.495 170.565 62.985 170.695 ;
        RECT 62.495 170.525 64.220 170.565 ;
        RECT 62.815 170.395 64.220 170.525 ;
        RECT 61.610 170.000 61.780 170.145 ;
        RECT 61.045 169.595 61.385 169.965 ;
        RECT 61.610 169.670 61.885 170.000 ;
        RECT 61.610 169.415 61.780 169.670 ;
        RECT 61.115 169.245 61.780 169.415 ;
        RECT 62.055 169.370 62.235 170.170 ;
        RECT 62.465 169.585 62.645 170.355 ;
        RECT 62.815 169.415 62.985 170.395 ;
        RECT 63.325 170.055 63.710 170.225 ;
        RECT 63.540 169.895 63.710 170.055 ;
        RECT 63.880 170.185 64.220 170.395 ;
        RECT 49.525 168.695 54.870 169.240 ;
        RECT 55.045 168.695 60.390 169.240 ;
        RECT 61.115 168.865 61.285 169.245 ;
        RECT 61.465 168.695 61.795 169.075 ;
        RECT 61.975 168.865 62.235 169.370 ;
        RECT 62.490 169.245 62.985 169.415 ;
        RECT 63.155 169.375 63.555 169.705 ;
        RECT 63.880 169.645 64.050 170.185 ;
        RECT 64.390 170.015 64.560 170.735 ;
        RECT 64.915 170.665 65.145 171.245 ;
        RECT 65.625 170.735 66.140 170.905 ;
        RECT 65.290 170.395 65.635 170.565 ;
        RECT 65.885 170.420 66.140 170.735 ;
        RECT 65.465 170.270 65.635 170.395 ;
        RECT 65.465 170.100 65.735 170.270 ;
        RECT 62.490 168.955 62.665 169.245 ;
        RECT 62.835 168.695 63.165 169.075 ;
        RECT 63.340 169.005 63.555 169.375 ;
        RECT 63.725 169.315 64.050 169.645 ;
        RECT 64.220 169.845 64.560 170.015 ;
        RECT 65.565 170.000 65.735 170.100 ;
        RECT 64.220 169.145 64.390 169.845 ;
        RECT 64.730 169.625 64.935 169.930 ;
        RECT 64.560 169.325 64.935 169.625 ;
        RECT 65.105 169.325 65.395 169.930 ;
        RECT 65.565 169.670 65.800 170.000 ;
        RECT 63.790 168.975 64.390 169.145 ;
        RECT 64.770 168.695 65.100 169.155 ;
        RECT 65.565 169.075 65.735 169.670 ;
        RECT 65.970 169.285 66.140 170.420 ;
        RECT 65.305 168.905 65.735 169.075 ;
        RECT 65.905 168.955 66.140 169.285 ;
        RECT 66.310 170.735 66.835 170.905 ;
        RECT 66.310 168.955 66.500 170.735 ;
        RECT 67.075 170.615 67.420 171.245 ;
        RECT 67.645 170.765 68.595 170.935 ;
        RECT 66.715 170.345 66.905 170.505 ;
        RECT 67.645 170.345 67.815 170.765 ;
        RECT 68.845 170.735 69.165 170.905 ;
        RECT 66.715 170.175 67.815 170.345 ;
        RECT 66.715 169.195 66.885 170.175 ;
        RECT 67.065 169.325 67.435 170.005 ;
        RECT 66.715 168.865 66.920 169.195 ;
        RECT 67.115 168.695 67.445 169.155 ;
        RECT 67.645 169.075 67.815 170.175 ;
        RECT 67.985 169.645 68.275 170.595 ;
        RECT 68.995 170.275 69.165 170.735 ;
        RECT 69.335 170.445 69.505 171.245 ;
        RECT 69.675 170.445 70.085 171.065 ;
        RECT 68.445 169.855 68.785 170.255 ;
        RECT 68.995 170.105 69.605 170.275 ;
        RECT 69.775 170.105 70.085 170.445 ;
        RECT 70.255 170.105 70.505 171.245 ;
        RECT 70.685 170.155 74.195 171.245 ;
        RECT 69.435 169.935 69.605 170.105 ;
        RECT 68.955 169.685 69.265 169.935 ;
        RECT 67.985 169.315 68.605 169.645 ;
        RECT 68.855 169.605 69.265 169.685 ;
        RECT 69.435 169.605 69.745 169.935 ;
        RECT 67.645 168.905 68.540 169.075 ;
        RECT 68.855 168.985 69.165 169.605 ;
        RECT 69.335 168.695 69.585 169.425 ;
        RECT 69.915 169.335 70.085 170.105 ;
        RECT 69.755 168.875 70.085 169.335 ;
        RECT 70.255 168.695 70.510 169.495 ;
        RECT 70.685 169.465 72.335 169.985 ;
        RECT 72.505 169.635 74.195 170.155 ;
        RECT 74.825 170.080 75.115 171.245 ;
        RECT 75.285 170.375 75.560 171.075 ;
        RECT 75.770 170.700 75.985 171.245 ;
        RECT 76.155 170.735 76.630 171.075 ;
        RECT 76.800 170.740 77.415 171.245 ;
        RECT 76.800 170.565 76.995 170.740 ;
        RECT 70.685 168.695 74.195 169.465 ;
        RECT 74.825 168.695 75.115 169.420 ;
        RECT 75.285 169.345 75.455 170.375 ;
        RECT 75.730 170.205 76.445 170.500 ;
        RECT 76.665 170.375 76.995 170.565 ;
        RECT 77.165 170.205 77.415 170.570 ;
        RECT 75.625 170.035 77.415 170.205 ;
        RECT 75.625 169.605 75.855 170.035 ;
        RECT 75.285 168.865 75.545 169.345 ;
        RECT 76.025 169.335 76.435 169.855 ;
        RECT 75.715 168.695 76.045 169.155 ;
        RECT 76.235 168.915 76.435 169.335 ;
        RECT 76.605 169.180 76.860 170.035 ;
        RECT 77.655 169.855 77.825 171.075 ;
        RECT 78.075 170.735 78.335 171.245 ;
        RECT 78.505 170.810 83.850 171.245 ;
        RECT 77.030 169.605 77.825 169.855 ;
        RECT 77.995 169.685 78.335 170.565 ;
        RECT 77.575 169.515 77.825 169.605 ;
        RECT 76.605 168.915 77.395 169.180 ;
        RECT 77.575 169.095 77.905 169.515 ;
        RECT 78.075 168.695 78.335 169.515 ;
        RECT 80.090 169.240 80.430 170.070 ;
        RECT 81.910 169.560 82.260 170.810 ;
        RECT 84.025 170.155 87.535 171.245 ;
        RECT 84.025 169.465 85.675 169.985 ;
        RECT 85.845 169.635 87.535 170.155 ;
        RECT 87.715 170.185 88.045 171.035 ;
        RECT 78.505 168.695 83.850 169.240 ;
        RECT 84.025 168.695 87.535 169.465 ;
        RECT 87.715 169.420 87.905 170.185 ;
        RECT 88.215 170.105 88.465 171.245 ;
        RECT 88.655 170.605 88.905 171.025 ;
        RECT 89.135 170.775 89.465 171.245 ;
        RECT 89.695 170.605 89.945 171.025 ;
        RECT 88.655 170.435 89.945 170.605 ;
        RECT 90.125 170.605 90.455 171.035 ;
        RECT 91.225 170.605 91.555 171.035 ;
        RECT 90.125 170.435 90.580 170.605 ;
        RECT 88.645 169.935 88.860 170.265 ;
        RECT 88.075 169.605 88.385 169.935 ;
        RECT 88.555 169.605 88.860 169.935 ;
        RECT 89.035 169.605 89.320 170.265 ;
        RECT 89.515 169.605 89.780 170.265 ;
        RECT 89.995 169.605 90.240 170.265 ;
        RECT 88.215 169.435 88.385 169.605 ;
        RECT 90.410 169.435 90.580 170.435 ;
        RECT 87.715 168.910 88.045 169.420 ;
        RECT 88.215 169.265 90.580 169.435 ;
        RECT 91.100 170.435 91.555 170.605 ;
        RECT 91.735 170.605 91.985 171.025 ;
        RECT 92.215 170.775 92.545 171.245 ;
        RECT 92.775 170.605 93.025 171.025 ;
        RECT 91.735 170.435 93.025 170.605 ;
        RECT 91.100 169.435 91.270 170.435 ;
        RECT 91.440 169.605 91.685 170.265 ;
        RECT 91.900 169.605 92.165 170.265 ;
        RECT 92.360 169.605 92.645 170.265 ;
        RECT 92.820 169.935 93.035 170.265 ;
        RECT 93.215 170.105 93.465 171.245 ;
        RECT 93.635 170.185 93.965 171.035 ;
        RECT 92.820 169.605 93.125 169.935 ;
        RECT 93.295 169.605 93.605 169.935 ;
        RECT 93.295 169.435 93.465 169.605 ;
        RECT 91.100 169.265 93.465 169.435 ;
        RECT 93.775 169.420 93.965 170.185 ;
        RECT 94.330 170.275 94.720 170.450 ;
        RECT 95.205 170.445 95.535 171.245 ;
        RECT 95.705 170.455 96.240 171.075 ;
        RECT 94.330 170.105 95.755 170.275 ;
        RECT 88.215 168.695 88.545 169.095 ;
        RECT 89.595 168.925 89.925 169.265 ;
        RECT 90.095 168.695 90.425 169.095 ;
        RECT 91.255 168.695 91.585 169.095 ;
        RECT 91.755 168.925 92.085 169.265 ;
        RECT 93.135 168.695 93.465 169.095 ;
        RECT 93.635 168.910 93.965 169.420 ;
        RECT 94.205 169.375 94.560 169.935 ;
        RECT 94.730 169.205 94.900 170.105 ;
        RECT 95.070 169.375 95.335 169.935 ;
        RECT 95.585 169.605 95.755 170.105 ;
        RECT 95.925 169.435 96.240 170.455 ;
        RECT 96.445 170.155 99.955 171.245 ;
        RECT 94.310 168.695 94.550 169.205 ;
        RECT 94.730 168.875 95.010 169.205 ;
        RECT 95.240 168.695 95.455 169.205 ;
        RECT 95.625 168.865 96.240 169.435 ;
        RECT 96.445 169.465 98.095 169.985 ;
        RECT 98.265 169.635 99.955 170.155 ;
        RECT 100.585 170.080 100.875 171.245 ;
        RECT 101.045 169.640 101.325 171.075 ;
        RECT 101.495 170.470 102.205 171.245 ;
        RECT 102.375 170.300 102.705 171.075 ;
        RECT 101.555 170.085 102.705 170.300 ;
        RECT 96.445 168.695 99.955 169.465 ;
        RECT 100.585 168.695 100.875 169.420 ;
        RECT 101.045 168.865 101.385 169.640 ;
        RECT 101.555 169.515 101.840 170.085 ;
        RECT 102.025 169.685 102.495 169.915 ;
        RECT 102.900 169.885 103.115 171.000 ;
        RECT 103.295 170.525 103.625 171.245 ;
        RECT 103.405 169.885 103.635 170.225 ;
        RECT 103.805 170.155 107.315 171.245 ;
        RECT 102.665 169.705 103.115 169.885 ;
        RECT 102.665 169.685 102.995 169.705 ;
        RECT 103.305 169.685 103.635 169.885 ;
        RECT 101.555 169.325 102.265 169.515 ;
        RECT 101.965 169.185 102.265 169.325 ;
        RECT 102.455 169.325 103.635 169.515 ;
        RECT 102.455 169.245 102.785 169.325 ;
        RECT 101.965 169.175 102.280 169.185 ;
        RECT 101.965 169.165 102.290 169.175 ;
        RECT 101.965 169.160 102.300 169.165 ;
        RECT 101.555 168.695 101.725 169.155 ;
        RECT 101.965 169.150 102.305 169.160 ;
        RECT 101.965 169.145 102.310 169.150 ;
        RECT 101.965 169.135 102.315 169.145 ;
        RECT 101.965 169.130 102.320 169.135 ;
        RECT 101.965 168.865 102.325 169.130 ;
        RECT 102.955 168.695 103.125 169.155 ;
        RECT 103.295 168.865 103.635 169.325 ;
        RECT 103.805 169.465 105.455 169.985 ;
        RECT 105.625 169.635 107.315 170.155 ;
        RECT 107.485 170.105 107.765 171.245 ;
        RECT 107.935 170.095 108.265 171.075 ;
        RECT 108.435 170.105 108.695 171.245 ;
        RECT 109.165 170.605 109.495 171.035 ;
        RECT 109.040 170.435 109.495 170.605 ;
        RECT 109.675 170.605 109.925 171.025 ;
        RECT 110.155 170.775 110.485 171.245 ;
        RECT 110.715 170.605 110.965 171.025 ;
        RECT 109.675 170.435 110.965 170.605 ;
        RECT 107.495 169.665 107.830 169.935 ;
        RECT 108.000 169.545 108.170 170.095 ;
        RECT 108.340 169.685 108.675 169.935 ;
        RECT 108.000 169.495 108.175 169.545 ;
        RECT 103.805 168.695 107.315 169.465 ;
        RECT 107.485 168.695 107.795 169.495 ;
        RECT 108.000 168.865 108.695 169.495 ;
        RECT 109.040 169.435 109.210 170.435 ;
        RECT 109.380 169.605 109.625 170.265 ;
        RECT 109.840 169.605 110.105 170.265 ;
        RECT 110.300 169.605 110.585 170.265 ;
        RECT 110.760 169.935 110.975 170.265 ;
        RECT 111.155 170.105 111.405 171.245 ;
        RECT 111.575 170.185 111.905 171.035 ;
        RECT 110.760 169.605 111.065 169.935 ;
        RECT 111.235 169.605 111.545 169.935 ;
        RECT 111.235 169.435 111.405 169.605 ;
        RECT 109.040 169.265 111.405 169.435 ;
        RECT 111.715 169.420 111.905 170.185 ;
        RECT 112.270 170.275 112.660 170.450 ;
        RECT 113.145 170.445 113.475 171.245 ;
        RECT 113.645 170.455 114.180 171.075 ;
        RECT 112.270 170.105 113.695 170.275 ;
        RECT 109.195 168.695 109.525 169.095 ;
        RECT 109.695 168.925 110.025 169.265 ;
        RECT 111.075 168.695 111.405 169.095 ;
        RECT 111.575 168.910 111.905 169.420 ;
        RECT 112.145 169.375 112.500 169.935 ;
        RECT 112.670 169.205 112.840 170.105 ;
        RECT 113.010 169.375 113.275 169.935 ;
        RECT 113.525 169.605 113.695 170.105 ;
        RECT 113.865 169.435 114.180 170.455 ;
        RECT 112.250 168.695 112.490 169.205 ;
        RECT 112.670 168.875 112.950 169.205 ;
        RECT 113.180 168.695 113.395 169.205 ;
        RECT 113.565 168.865 114.180 169.435 ;
        RECT 114.385 170.170 114.655 171.075 ;
        RECT 114.825 170.485 115.155 171.245 ;
        RECT 115.335 170.315 115.515 171.075 ;
        RECT 115.765 170.810 121.110 171.245 ;
        RECT 114.385 169.370 114.565 170.170 ;
        RECT 114.840 170.145 115.515 170.315 ;
        RECT 114.840 170.000 115.010 170.145 ;
        RECT 114.735 169.670 115.010 170.000 ;
        RECT 114.840 169.415 115.010 169.670 ;
        RECT 115.235 169.595 115.575 169.965 ;
        RECT 114.385 168.865 114.645 169.370 ;
        RECT 114.840 169.245 115.505 169.415 ;
        RECT 114.825 168.695 115.155 169.075 ;
        RECT 115.335 168.865 115.505 169.245 ;
        RECT 117.350 169.240 117.690 170.070 ;
        RECT 119.170 169.560 119.520 170.810 ;
        RECT 121.285 170.155 122.955 171.245 ;
        RECT 121.285 169.465 122.035 169.985 ;
        RECT 122.205 169.635 122.955 170.155 ;
        RECT 123.135 170.105 123.465 171.245 ;
        RECT 123.995 170.275 124.325 171.060 ;
        RECT 123.645 170.105 124.325 170.275 ;
        RECT 124.505 170.155 126.175 171.245 ;
        RECT 123.125 169.685 123.475 169.935 ;
        RECT 123.645 169.505 123.815 170.105 ;
        RECT 123.985 169.685 124.335 169.935 ;
        RECT 115.765 168.695 121.110 169.240 ;
        RECT 121.285 168.695 122.955 169.465 ;
        RECT 123.135 168.695 123.405 169.505 ;
        RECT 123.575 168.865 123.905 169.505 ;
        RECT 124.075 168.695 124.315 169.505 ;
        RECT 124.505 169.465 125.255 169.985 ;
        RECT 125.425 169.635 126.175 170.155 ;
        RECT 126.345 170.080 126.635 171.245 ;
        RECT 126.810 170.855 127.145 171.075 ;
        RECT 128.150 170.865 128.505 171.245 ;
        RECT 126.810 170.235 127.065 170.855 ;
        RECT 127.315 170.695 127.545 170.735 ;
        RECT 128.675 170.695 128.925 171.075 ;
        RECT 127.315 170.495 128.925 170.695 ;
        RECT 127.315 170.405 127.500 170.495 ;
        RECT 128.090 170.485 128.925 170.495 ;
        RECT 129.175 170.465 129.425 171.245 ;
        RECT 129.595 170.395 129.855 171.075 ;
        RECT 130.025 170.810 135.370 171.245 ;
        RECT 127.655 170.295 127.985 170.325 ;
        RECT 127.655 170.235 129.455 170.295 ;
        RECT 126.810 170.125 129.515 170.235 ;
        RECT 126.810 170.065 127.985 170.125 ;
        RECT 129.315 170.090 129.515 170.125 ;
        RECT 126.805 169.685 127.295 169.885 ;
        RECT 127.485 169.685 127.960 169.895 ;
        RECT 124.505 168.695 126.175 169.465 ;
        RECT 126.345 168.695 126.635 169.420 ;
        RECT 126.810 168.695 127.265 169.460 ;
        RECT 127.740 169.285 127.960 169.685 ;
        RECT 128.205 169.685 128.535 169.895 ;
        RECT 128.205 169.285 128.415 169.685 ;
        RECT 128.705 169.650 129.115 169.955 ;
        RECT 129.345 169.515 129.515 170.090 ;
        RECT 129.245 169.395 129.515 169.515 ;
        RECT 128.670 169.350 129.515 169.395 ;
        RECT 128.670 169.225 129.425 169.350 ;
        RECT 128.670 169.075 128.840 169.225 ;
        RECT 129.685 169.205 129.855 170.395 ;
        RECT 131.610 169.240 131.950 170.070 ;
        RECT 133.430 169.560 133.780 170.810 ;
        RECT 135.545 170.155 137.215 171.245 ;
        RECT 137.850 170.735 139.505 171.025 ;
        RECT 135.545 169.465 136.295 169.985 ;
        RECT 136.465 169.635 137.215 170.155 ;
        RECT 137.850 170.395 139.440 170.565 ;
        RECT 139.675 170.445 139.955 171.245 ;
        RECT 137.850 170.105 138.170 170.395 ;
        RECT 139.270 170.275 139.440 170.395 ;
        RECT 138.365 170.055 139.080 170.225 ;
        RECT 139.270 170.105 139.995 170.275 ;
        RECT 140.165 170.105 140.435 171.075 ;
        RECT 140.695 170.575 140.865 171.075 ;
        RECT 141.035 170.745 141.365 171.245 ;
        RECT 140.695 170.405 141.360 170.575 ;
        RECT 129.625 169.195 129.855 169.205 ;
        RECT 127.540 168.865 128.840 169.075 ;
        RECT 129.095 168.695 129.425 169.055 ;
        RECT 129.595 168.865 129.855 169.195 ;
        RECT 130.025 168.695 135.370 169.240 ;
        RECT 135.545 168.695 137.215 169.465 ;
        RECT 137.850 169.365 138.200 169.935 ;
        RECT 138.370 169.605 139.080 170.055 ;
        RECT 139.825 169.935 139.995 170.105 ;
        RECT 139.250 169.605 139.655 169.935 ;
        RECT 139.825 169.605 140.095 169.935 ;
        RECT 139.825 169.435 139.995 169.605 ;
        RECT 138.385 169.265 139.995 169.435 ;
        RECT 140.265 169.370 140.435 170.105 ;
        RECT 140.610 169.585 140.960 170.235 ;
        RECT 141.130 169.415 141.360 170.405 ;
        RECT 137.855 168.695 138.185 169.195 ;
        RECT 138.385 168.915 138.555 169.265 ;
        RECT 138.755 168.695 139.085 169.095 ;
        RECT 139.255 168.915 139.425 169.265 ;
        RECT 139.595 168.695 139.975 169.095 ;
        RECT 140.165 169.025 140.435 169.370 ;
        RECT 140.695 169.245 141.360 169.415 ;
        RECT 140.695 168.955 140.865 169.245 ;
        RECT 141.035 168.695 141.365 169.075 ;
        RECT 141.535 168.955 141.720 171.075 ;
        RECT 141.960 170.785 142.225 171.245 ;
        RECT 142.395 170.650 142.645 171.075 ;
        RECT 142.855 170.800 143.960 170.970 ;
        RECT 142.340 170.520 142.645 170.650 ;
        RECT 141.890 169.325 142.170 170.275 ;
        RECT 142.340 169.415 142.510 170.520 ;
        RECT 142.680 169.735 142.920 170.330 ;
        RECT 143.090 170.265 143.620 170.630 ;
        RECT 143.090 169.565 143.260 170.265 ;
        RECT 143.790 170.185 143.960 170.800 ;
        RECT 144.130 170.445 144.300 171.245 ;
        RECT 144.470 170.745 144.720 171.075 ;
        RECT 144.945 170.775 145.830 170.945 ;
        RECT 143.790 170.095 144.300 170.185 ;
        RECT 142.340 169.285 142.565 169.415 ;
        RECT 142.735 169.345 143.260 169.565 ;
        RECT 143.430 169.925 144.300 170.095 ;
        RECT 141.975 168.695 142.225 169.155 ;
        RECT 142.395 169.145 142.565 169.285 ;
        RECT 143.430 169.145 143.600 169.925 ;
        RECT 144.130 169.855 144.300 169.925 ;
        RECT 143.810 169.675 144.010 169.705 ;
        RECT 144.470 169.675 144.640 170.745 ;
        RECT 144.810 169.855 145.000 170.575 ;
        RECT 143.810 169.375 144.640 169.675 ;
        RECT 145.170 169.645 145.490 170.605 ;
        RECT 142.395 168.975 142.730 169.145 ;
        RECT 142.925 168.975 143.600 169.145 ;
        RECT 143.920 168.695 144.290 169.195 ;
        RECT 144.470 169.145 144.640 169.375 ;
        RECT 145.025 169.315 145.490 169.645 ;
        RECT 145.660 169.935 145.830 170.775 ;
        RECT 146.010 170.745 146.325 171.245 ;
        RECT 146.555 170.515 146.895 171.075 ;
        RECT 146.000 170.140 146.895 170.515 ;
        RECT 147.065 170.235 147.235 171.245 ;
        RECT 146.705 169.935 146.895 170.140 ;
        RECT 147.405 170.185 147.735 171.030 ;
        RECT 147.405 170.105 147.795 170.185 ;
        RECT 147.580 170.055 147.795 170.105 ;
        RECT 145.660 169.605 146.535 169.935 ;
        RECT 146.705 169.605 147.455 169.935 ;
        RECT 145.660 169.145 145.830 169.605 ;
        RECT 146.705 169.435 146.905 169.605 ;
        RECT 147.625 169.475 147.795 170.055 ;
        RECT 148.885 170.155 150.095 171.245 ;
        RECT 148.885 169.615 149.405 170.155 ;
        RECT 147.570 169.435 147.795 169.475 ;
        RECT 149.575 169.445 150.095 169.985 ;
        RECT 144.470 168.975 144.875 169.145 ;
        RECT 145.045 168.975 145.830 169.145 ;
        RECT 146.105 168.695 146.315 169.225 ;
        RECT 146.575 168.910 146.905 169.435 ;
        RECT 147.415 169.350 147.795 169.435 ;
        RECT 147.075 168.695 147.245 169.305 ;
        RECT 147.415 168.915 147.745 169.350 ;
        RECT 148.885 168.695 150.095 169.445 ;
        RECT 36.100 168.525 150.180 168.695 ;
        RECT 36.185 167.775 37.395 168.525 ;
        RECT 36.185 167.235 36.705 167.775 ;
        RECT 37.565 167.755 41.075 168.525 ;
        RECT 36.875 167.065 37.395 167.605 ;
        RECT 37.565 167.235 39.215 167.755 ;
        RECT 41.705 167.705 41.965 168.525 ;
        RECT 42.135 167.705 42.465 168.125 ;
        RECT 42.645 168.040 43.435 168.305 ;
        RECT 42.215 167.615 42.465 167.705 ;
        RECT 39.385 167.065 41.075 167.585 ;
        RECT 36.185 165.975 37.395 167.065 ;
        RECT 37.565 165.975 41.075 167.065 ;
        RECT 41.705 166.655 42.045 167.535 ;
        RECT 42.215 167.365 43.010 167.615 ;
        RECT 41.705 165.975 41.965 166.485 ;
        RECT 42.215 166.145 42.385 167.365 ;
        RECT 43.180 167.185 43.435 168.040 ;
        RECT 43.605 167.885 43.805 168.305 ;
        RECT 43.995 168.065 44.325 168.525 ;
        RECT 43.605 167.365 44.015 167.885 ;
        RECT 44.495 167.875 44.755 168.355 ;
        RECT 44.185 167.185 44.415 167.615 ;
        RECT 42.625 167.015 44.415 167.185 ;
        RECT 42.625 166.650 42.875 167.015 ;
        RECT 43.045 166.655 43.375 166.845 ;
        RECT 43.595 166.720 44.310 167.015 ;
        RECT 44.585 166.845 44.755 167.875 ;
        RECT 45.015 167.975 45.185 168.265 ;
        RECT 45.355 168.145 45.685 168.525 ;
        RECT 45.015 167.805 45.680 167.975 ;
        RECT 44.930 166.985 45.280 167.635 ;
        RECT 43.045 166.480 43.240 166.655 ;
        RECT 42.625 165.975 43.240 166.480 ;
        RECT 43.410 166.145 43.885 166.485 ;
        RECT 44.055 165.975 44.270 166.520 ;
        RECT 44.480 166.145 44.755 166.845 ;
        RECT 45.450 166.815 45.680 167.805 ;
        RECT 45.015 166.645 45.680 166.815 ;
        RECT 45.015 166.145 45.185 166.645 ;
        RECT 45.355 165.975 45.685 166.475 ;
        RECT 45.855 166.145 46.040 168.265 ;
        RECT 46.295 168.065 46.545 168.525 ;
        RECT 46.715 168.075 47.050 168.245 ;
        RECT 47.245 168.075 47.920 168.245 ;
        RECT 46.715 167.935 46.885 168.075 ;
        RECT 46.210 166.945 46.490 167.895 ;
        RECT 46.660 167.805 46.885 167.935 ;
        RECT 46.660 166.700 46.830 167.805 ;
        RECT 47.055 167.655 47.580 167.875 ;
        RECT 47.000 166.890 47.240 167.485 ;
        RECT 47.410 166.955 47.580 167.655 ;
        RECT 47.750 167.295 47.920 168.075 ;
        RECT 48.240 168.025 48.610 168.525 ;
        RECT 48.790 168.075 49.195 168.245 ;
        RECT 49.365 168.075 50.150 168.245 ;
        RECT 48.790 167.845 48.960 168.075 ;
        RECT 48.130 167.545 48.960 167.845 ;
        RECT 49.345 167.575 49.810 167.905 ;
        RECT 48.130 167.515 48.330 167.545 ;
        RECT 48.450 167.295 48.620 167.365 ;
        RECT 47.750 167.125 48.620 167.295 ;
        RECT 48.110 167.035 48.620 167.125 ;
        RECT 46.660 166.570 46.965 166.700 ;
        RECT 47.410 166.590 47.940 166.955 ;
        RECT 46.280 165.975 46.545 166.435 ;
        RECT 46.715 166.145 46.965 166.570 ;
        RECT 48.110 166.420 48.280 167.035 ;
        RECT 47.175 166.250 48.280 166.420 ;
        RECT 48.450 165.975 48.620 166.775 ;
        RECT 48.790 166.475 48.960 167.545 ;
        RECT 49.130 166.645 49.320 167.365 ;
        RECT 49.490 166.615 49.810 167.575 ;
        RECT 49.980 167.615 50.150 168.075 ;
        RECT 50.425 167.995 50.635 168.525 ;
        RECT 50.895 167.785 51.225 168.310 ;
        RECT 51.395 167.915 51.565 168.525 ;
        RECT 51.735 167.870 52.065 168.305 ;
        RECT 52.285 167.980 57.630 168.525 ;
        RECT 51.735 167.785 52.115 167.870 ;
        RECT 51.025 167.615 51.225 167.785 ;
        RECT 51.890 167.745 52.115 167.785 ;
        RECT 49.980 167.285 50.855 167.615 ;
        RECT 51.025 167.285 51.775 167.615 ;
        RECT 48.790 166.145 49.040 166.475 ;
        RECT 49.980 166.445 50.150 167.285 ;
        RECT 51.025 167.080 51.215 167.285 ;
        RECT 51.945 167.165 52.115 167.745 ;
        RECT 51.900 167.115 52.115 167.165 ;
        RECT 53.870 167.150 54.210 167.980 ;
        RECT 57.815 167.800 58.145 168.310 ;
        RECT 58.315 168.125 58.645 168.525 ;
        RECT 59.695 167.955 60.025 168.295 ;
        RECT 60.195 168.125 60.525 168.525 ;
        RECT 50.320 166.705 51.215 167.080 ;
        RECT 51.725 167.035 52.115 167.115 ;
        RECT 49.265 166.275 50.150 166.445 ;
        RECT 50.330 165.975 50.645 166.475 ;
        RECT 50.875 166.145 51.215 166.705 ;
        RECT 51.385 165.975 51.555 166.985 ;
        RECT 51.725 166.190 52.055 167.035 ;
        RECT 55.690 166.410 56.040 167.660 ;
        RECT 57.815 167.035 58.005 167.800 ;
        RECT 58.315 167.785 60.680 167.955 ;
        RECT 61.945 167.800 62.235 168.525 ;
        RECT 62.495 167.975 62.665 168.265 ;
        RECT 62.835 168.145 63.165 168.525 ;
        RECT 62.495 167.805 63.160 167.975 ;
        RECT 58.315 167.615 58.485 167.785 ;
        RECT 58.175 167.285 58.485 167.615 ;
        RECT 58.655 167.285 58.960 167.615 ;
        RECT 52.285 165.975 57.630 166.410 ;
        RECT 57.815 166.185 58.145 167.035 ;
        RECT 58.315 165.975 58.565 167.115 ;
        RECT 58.745 166.955 58.960 167.285 ;
        RECT 59.135 166.955 59.420 167.615 ;
        RECT 59.615 166.955 59.880 167.615 ;
        RECT 60.095 166.955 60.340 167.615 ;
        RECT 60.510 166.785 60.680 167.785 ;
        RECT 58.755 166.615 60.045 166.785 ;
        RECT 58.755 166.195 59.005 166.615 ;
        RECT 59.235 165.975 59.565 166.445 ;
        RECT 59.795 166.195 60.045 166.615 ;
        RECT 60.225 166.615 60.680 166.785 ;
        RECT 60.225 166.185 60.555 166.615 ;
        RECT 61.945 165.975 62.235 167.140 ;
        RECT 62.410 166.985 62.760 167.635 ;
        RECT 62.930 166.815 63.160 167.805 ;
        RECT 62.495 166.645 63.160 166.815 ;
        RECT 62.495 166.145 62.665 166.645 ;
        RECT 62.835 165.975 63.165 166.475 ;
        RECT 63.335 166.145 63.520 168.265 ;
        RECT 63.775 168.065 64.025 168.525 ;
        RECT 64.195 168.075 64.530 168.245 ;
        RECT 64.725 168.075 65.400 168.245 ;
        RECT 64.195 167.935 64.365 168.075 ;
        RECT 63.690 166.945 63.970 167.895 ;
        RECT 64.140 167.805 64.365 167.935 ;
        RECT 64.140 166.700 64.310 167.805 ;
        RECT 64.535 167.655 65.060 167.875 ;
        RECT 64.480 166.890 64.720 167.485 ;
        RECT 64.890 166.955 65.060 167.655 ;
        RECT 65.230 167.295 65.400 168.075 ;
        RECT 65.720 168.025 66.090 168.525 ;
        RECT 66.270 168.075 66.675 168.245 ;
        RECT 66.845 168.075 67.630 168.245 ;
        RECT 66.270 167.845 66.440 168.075 ;
        RECT 65.610 167.545 66.440 167.845 ;
        RECT 66.825 167.575 67.290 167.905 ;
        RECT 65.610 167.515 65.810 167.545 ;
        RECT 65.930 167.295 66.100 167.365 ;
        RECT 65.230 167.125 66.100 167.295 ;
        RECT 65.590 167.035 66.100 167.125 ;
        RECT 64.140 166.570 64.445 166.700 ;
        RECT 64.890 166.590 65.420 166.955 ;
        RECT 63.760 165.975 64.025 166.435 ;
        RECT 64.195 166.145 64.445 166.570 ;
        RECT 65.590 166.420 65.760 167.035 ;
        RECT 64.655 166.250 65.760 166.420 ;
        RECT 65.930 165.975 66.100 166.775 ;
        RECT 66.270 166.475 66.440 167.545 ;
        RECT 66.610 166.645 66.800 167.365 ;
        RECT 66.970 166.615 67.290 167.575 ;
        RECT 67.460 167.615 67.630 168.075 ;
        RECT 67.905 167.995 68.115 168.525 ;
        RECT 68.375 167.785 68.705 168.310 ;
        RECT 68.875 167.915 69.045 168.525 ;
        RECT 69.215 167.870 69.545 168.305 ;
        RECT 69.215 167.785 69.595 167.870 ;
        RECT 68.505 167.615 68.705 167.785 ;
        RECT 69.370 167.745 69.595 167.785 ;
        RECT 67.460 167.285 68.335 167.615 ;
        RECT 68.505 167.285 69.255 167.615 ;
        RECT 66.270 166.145 66.520 166.475 ;
        RECT 67.460 166.445 67.630 167.285 ;
        RECT 68.505 167.080 68.695 167.285 ;
        RECT 69.425 167.165 69.595 167.745 ;
        RECT 69.765 167.775 70.975 168.525 ;
        RECT 71.235 167.975 71.405 168.355 ;
        RECT 71.585 168.145 71.915 168.525 ;
        RECT 71.235 167.805 71.900 167.975 ;
        RECT 72.095 167.850 72.355 168.355 ;
        RECT 72.610 168.025 73.105 168.355 ;
        RECT 69.765 167.235 70.285 167.775 ;
        RECT 69.380 167.115 69.595 167.165 ;
        RECT 67.800 166.705 68.695 167.080 ;
        RECT 69.205 167.035 69.595 167.115 ;
        RECT 70.455 167.065 70.975 167.605 ;
        RECT 71.165 167.255 71.505 167.625 ;
        RECT 71.730 167.550 71.900 167.805 ;
        RECT 71.730 167.220 72.005 167.550 ;
        RECT 71.730 167.075 71.900 167.220 ;
        RECT 66.745 166.275 67.630 166.445 ;
        RECT 67.810 165.975 68.125 166.475 ;
        RECT 68.355 166.145 68.695 166.705 ;
        RECT 68.865 165.975 69.035 166.985 ;
        RECT 69.205 166.190 69.535 167.035 ;
        RECT 69.765 165.975 70.975 167.065 ;
        RECT 71.225 166.905 71.900 167.075 ;
        RECT 72.175 167.050 72.355 167.850 ;
        RECT 71.225 166.145 71.405 166.905 ;
        RECT 71.585 165.975 71.915 166.735 ;
        RECT 72.085 166.145 72.355 167.050 ;
        RECT 72.525 166.535 72.765 167.845 ;
        RECT 72.935 167.115 73.105 168.025 ;
        RECT 73.325 167.285 73.675 168.250 ;
        RECT 73.855 167.285 74.155 168.255 ;
        RECT 74.335 167.285 74.615 168.255 ;
        RECT 74.795 167.725 75.065 168.525 ;
        RECT 75.235 167.805 75.575 168.315 ;
        RECT 74.810 167.285 75.140 167.535 ;
        RECT 74.810 167.115 75.125 167.285 ;
        RECT 72.935 166.945 75.125 167.115 ;
        RECT 72.530 165.975 72.865 166.355 ;
        RECT 73.035 166.145 73.285 166.945 ;
        RECT 73.505 165.975 73.835 166.695 ;
        RECT 74.020 166.145 74.270 166.945 ;
        RECT 74.735 165.975 75.065 166.775 ;
        RECT 75.315 166.405 75.575 167.805 ;
        RECT 75.235 166.145 75.575 166.405 ;
        RECT 75.755 167.800 76.085 168.310 ;
        RECT 76.255 168.125 76.585 168.525 ;
        RECT 77.635 167.955 77.965 168.295 ;
        RECT 78.135 168.125 78.465 168.525 ;
        RECT 75.755 167.035 75.945 167.800 ;
        RECT 76.255 167.785 78.620 167.955 ;
        RECT 76.255 167.615 76.425 167.785 ;
        RECT 76.115 167.285 76.425 167.615 ;
        RECT 76.595 167.285 76.900 167.615 ;
        RECT 75.755 166.185 76.085 167.035 ;
        RECT 76.255 165.975 76.505 167.115 ;
        RECT 76.685 166.955 76.900 167.285 ;
        RECT 77.075 166.955 77.360 167.615 ;
        RECT 77.555 166.955 77.820 167.615 ;
        RECT 78.035 166.955 78.280 167.615 ;
        RECT 78.450 166.785 78.620 167.785 ;
        RECT 79.005 167.705 79.235 168.525 ;
        RECT 79.405 167.725 79.735 168.355 ;
        RECT 78.985 167.285 79.315 167.535 ;
        RECT 79.485 167.125 79.735 167.725 ;
        RECT 79.905 167.705 80.115 168.525 ;
        RECT 80.345 167.980 85.690 168.525 ;
        RECT 81.930 167.150 82.270 167.980 ;
        RECT 86.325 167.850 86.585 168.355 ;
        RECT 86.765 168.145 87.095 168.525 ;
        RECT 87.275 167.975 87.445 168.355 ;
        RECT 76.695 166.615 77.985 166.785 ;
        RECT 76.695 166.195 76.945 166.615 ;
        RECT 77.175 165.975 77.505 166.445 ;
        RECT 77.735 166.195 77.985 166.615 ;
        RECT 78.165 166.615 78.620 166.785 ;
        RECT 78.165 166.185 78.495 166.615 ;
        RECT 79.005 165.975 79.235 167.115 ;
        RECT 79.405 166.145 79.735 167.125 ;
        RECT 79.905 165.975 80.115 167.115 ;
        RECT 83.750 166.410 84.100 167.660 ;
        RECT 86.325 167.050 86.505 167.850 ;
        RECT 86.780 167.805 87.445 167.975 ;
        RECT 86.780 167.550 86.950 167.805 ;
        RECT 87.705 167.800 87.995 168.525 ;
        RECT 88.370 167.745 88.870 168.355 ;
        RECT 86.675 167.220 86.950 167.550 ;
        RECT 87.175 167.255 87.515 167.625 ;
        RECT 88.165 167.285 88.515 167.535 ;
        RECT 86.780 167.075 86.950 167.220 ;
        RECT 80.345 165.975 85.690 166.410 ;
        RECT 86.325 166.145 86.595 167.050 ;
        RECT 86.780 166.905 87.455 167.075 ;
        RECT 86.765 165.975 87.095 166.735 ;
        RECT 87.275 166.145 87.455 166.905 ;
        RECT 87.705 165.975 87.995 167.140 ;
        RECT 88.700 167.115 88.870 167.745 ;
        RECT 89.500 167.875 89.830 168.355 ;
        RECT 90.000 168.065 90.225 168.525 ;
        RECT 90.395 167.875 90.725 168.355 ;
        RECT 89.500 167.705 90.725 167.875 ;
        RECT 90.915 167.725 91.165 168.525 ;
        RECT 91.335 167.725 91.675 168.355 ;
        RECT 89.040 167.335 89.370 167.535 ;
        RECT 89.540 167.335 89.870 167.535 ;
        RECT 90.040 167.335 90.460 167.535 ;
        RECT 90.635 167.365 91.330 167.535 ;
        RECT 90.635 167.115 90.805 167.365 ;
        RECT 91.500 167.115 91.675 167.725 ;
        RECT 91.845 167.755 93.515 168.525 ;
        RECT 94.015 168.125 94.345 168.525 ;
        RECT 94.515 167.955 94.845 168.295 ;
        RECT 95.895 168.125 96.225 168.525 ;
        RECT 93.860 167.785 96.225 167.955 ;
        RECT 96.395 167.800 96.725 168.310 ;
        RECT 91.845 167.235 92.595 167.755 ;
        RECT 88.370 166.945 90.805 167.115 ;
        RECT 88.370 166.145 88.700 166.945 ;
        RECT 88.870 165.975 89.200 166.775 ;
        RECT 89.500 166.145 89.830 166.945 ;
        RECT 90.475 165.975 90.725 166.775 ;
        RECT 90.995 165.975 91.165 167.115 ;
        RECT 91.335 166.145 91.675 167.115 ;
        RECT 92.765 167.065 93.515 167.585 ;
        RECT 91.845 165.975 93.515 167.065 ;
        RECT 93.860 166.785 94.030 167.785 ;
        RECT 96.055 167.615 96.225 167.785 ;
        RECT 94.200 166.955 94.445 167.615 ;
        RECT 94.660 166.955 94.925 167.615 ;
        RECT 95.120 166.955 95.405 167.615 ;
        RECT 95.580 167.285 95.885 167.615 ;
        RECT 96.055 167.285 96.365 167.615 ;
        RECT 95.580 166.955 95.795 167.285 ;
        RECT 93.860 166.615 94.315 166.785 ;
        RECT 93.985 166.185 94.315 166.615 ;
        RECT 94.495 166.615 95.785 166.785 ;
        RECT 94.495 166.195 94.745 166.615 ;
        RECT 94.975 165.975 95.305 166.445 ;
        RECT 95.535 166.195 95.785 166.615 ;
        RECT 95.975 165.975 96.225 167.115 ;
        RECT 96.535 167.035 96.725 167.800 ;
        RECT 97.065 167.965 97.395 168.355 ;
        RECT 97.565 168.135 98.750 168.305 ;
        RECT 99.010 168.055 99.180 168.525 ;
        RECT 97.065 167.785 97.575 167.965 ;
        RECT 96.905 167.325 97.235 167.615 ;
        RECT 97.405 167.155 97.575 167.785 ;
        RECT 97.980 167.875 98.365 167.965 ;
        RECT 99.350 167.875 99.680 168.340 ;
        RECT 97.980 167.705 99.680 167.875 ;
        RECT 99.850 167.705 100.020 168.525 ;
        RECT 100.190 167.705 100.875 168.345 ;
        RECT 97.745 167.325 98.075 167.535 ;
        RECT 98.255 167.285 98.635 167.535 ;
        RECT 96.395 166.185 96.725 167.035 ;
        RECT 97.060 166.985 98.145 167.155 ;
        RECT 97.060 166.145 97.360 166.985 ;
        RECT 97.555 165.975 97.805 166.815 ;
        RECT 97.975 166.735 98.145 166.985 ;
        RECT 98.315 166.905 98.635 167.285 ;
        RECT 98.825 167.325 99.310 167.535 ;
        RECT 99.500 167.325 99.950 167.535 ;
        RECT 100.120 167.325 100.455 167.535 ;
        RECT 98.825 167.165 99.200 167.325 ;
        RECT 98.805 166.995 99.200 167.165 ;
        RECT 100.120 167.155 100.290 167.325 ;
        RECT 98.825 166.905 99.200 166.995 ;
        RECT 99.370 166.985 100.290 167.155 ;
        RECT 99.370 166.735 99.540 166.985 ;
        RECT 97.975 166.565 99.540 166.735 ;
        RECT 98.395 166.145 99.200 166.565 ;
        RECT 99.710 165.975 100.040 166.815 ;
        RECT 100.625 166.735 100.875 167.705 ;
        RECT 100.210 166.145 100.875 166.735 ;
        RECT 101.045 167.580 101.385 168.355 ;
        RECT 101.555 168.065 101.725 168.525 ;
        RECT 101.965 168.090 102.325 168.355 ;
        RECT 101.965 168.085 102.320 168.090 ;
        RECT 101.965 168.075 102.315 168.085 ;
        RECT 101.965 168.070 102.310 168.075 ;
        RECT 101.965 168.060 102.305 168.070 ;
        RECT 102.955 168.065 103.125 168.525 ;
        RECT 101.965 168.055 102.300 168.060 ;
        RECT 101.965 168.045 102.290 168.055 ;
        RECT 101.965 168.035 102.280 168.045 ;
        RECT 101.965 167.895 102.265 168.035 ;
        RECT 101.555 167.705 102.265 167.895 ;
        RECT 102.455 167.895 102.785 167.975 ;
        RECT 103.295 167.895 103.635 168.355 ;
        RECT 103.805 167.980 109.150 168.525 ;
        RECT 102.455 167.705 103.635 167.895 ;
        RECT 101.045 166.145 101.325 167.580 ;
        RECT 101.555 167.135 101.840 167.705 ;
        RECT 102.025 167.305 102.495 167.535 ;
        RECT 102.665 167.515 102.995 167.535 ;
        RECT 102.665 167.335 103.115 167.515 ;
        RECT 103.305 167.335 103.635 167.535 ;
        RECT 101.555 166.920 102.705 167.135 ;
        RECT 101.495 165.975 102.205 166.750 ;
        RECT 102.375 166.145 102.705 166.920 ;
        RECT 102.900 166.220 103.115 167.335 ;
        RECT 103.405 166.995 103.635 167.335 ;
        RECT 105.390 167.150 105.730 167.980 ;
        RECT 109.325 167.850 109.585 168.355 ;
        RECT 109.765 168.145 110.095 168.525 ;
        RECT 110.275 167.975 110.445 168.355 ;
        RECT 103.295 165.975 103.625 166.695 ;
        RECT 107.210 166.410 107.560 167.660 ;
        RECT 109.325 167.050 109.505 167.850 ;
        RECT 109.780 167.805 110.445 167.975 ;
        RECT 110.705 167.850 110.965 168.355 ;
        RECT 111.145 168.145 111.475 168.525 ;
        RECT 111.655 167.975 111.825 168.355 ;
        RECT 109.780 167.550 109.950 167.805 ;
        RECT 109.675 167.220 109.950 167.550 ;
        RECT 110.175 167.255 110.515 167.625 ;
        RECT 109.780 167.075 109.950 167.220 ;
        RECT 103.805 165.975 109.150 166.410 ;
        RECT 109.325 166.145 109.595 167.050 ;
        RECT 109.780 166.905 110.455 167.075 ;
        RECT 109.765 165.975 110.095 166.735 ;
        RECT 110.275 166.145 110.455 166.905 ;
        RECT 110.705 167.050 110.885 167.850 ;
        RECT 111.160 167.805 111.825 167.975 ;
        RECT 111.160 167.550 111.330 167.805 ;
        RECT 112.085 167.775 113.295 168.525 ;
        RECT 113.465 167.800 113.755 168.525 ;
        RECT 111.055 167.220 111.330 167.550 ;
        RECT 111.555 167.255 111.895 167.625 ;
        RECT 112.085 167.235 112.605 167.775 ;
        RECT 113.925 167.755 117.435 168.525 ;
        RECT 117.605 167.850 117.865 168.355 ;
        RECT 118.045 168.145 118.375 168.525 ;
        RECT 118.555 167.975 118.725 168.355 ;
        RECT 111.160 167.075 111.330 167.220 ;
        RECT 110.705 166.145 110.975 167.050 ;
        RECT 111.160 166.905 111.835 167.075 ;
        RECT 112.775 167.065 113.295 167.605 ;
        RECT 113.925 167.235 115.575 167.755 ;
        RECT 111.145 165.975 111.475 166.735 ;
        RECT 111.655 166.145 111.835 166.905 ;
        RECT 112.085 165.975 113.295 167.065 ;
        RECT 113.465 165.975 113.755 167.140 ;
        RECT 115.745 167.065 117.435 167.585 ;
        RECT 113.925 165.975 117.435 167.065 ;
        RECT 117.605 167.050 117.785 167.850 ;
        RECT 118.060 167.805 118.725 167.975 ;
        RECT 119.075 167.975 119.245 168.355 ;
        RECT 119.425 168.145 119.755 168.525 ;
        RECT 119.075 167.805 119.740 167.975 ;
        RECT 119.935 167.850 120.195 168.355 ;
        RECT 118.060 167.550 118.230 167.805 ;
        RECT 117.955 167.220 118.230 167.550 ;
        RECT 118.455 167.255 118.795 167.625 ;
        RECT 119.005 167.255 119.345 167.625 ;
        RECT 119.570 167.550 119.740 167.805 ;
        RECT 118.060 167.075 118.230 167.220 ;
        RECT 119.570 167.220 119.845 167.550 ;
        RECT 119.570 167.075 119.740 167.220 ;
        RECT 117.605 166.145 117.875 167.050 ;
        RECT 118.060 166.905 118.735 167.075 ;
        RECT 118.045 165.975 118.375 166.735 ;
        RECT 118.555 166.145 118.735 166.905 ;
        RECT 119.065 166.905 119.740 167.075 ;
        RECT 120.015 167.050 120.195 167.850 ;
        RECT 121.295 167.715 121.565 168.525 ;
        RECT 121.735 167.715 122.065 168.355 ;
        RECT 122.235 167.715 122.475 168.525 ;
        RECT 122.665 168.065 123.225 168.355 ;
        RECT 123.395 168.065 123.645 168.525 ;
        RECT 121.285 167.285 121.635 167.535 ;
        RECT 121.805 167.115 121.975 167.715 ;
        RECT 122.145 167.285 122.495 167.535 ;
        RECT 119.065 166.145 119.245 166.905 ;
        RECT 119.425 165.975 119.755 166.735 ;
        RECT 119.925 166.145 120.195 167.050 ;
        RECT 121.295 165.975 121.625 167.115 ;
        RECT 121.805 166.945 122.485 167.115 ;
        RECT 122.155 166.160 122.485 166.945 ;
        RECT 122.665 166.695 122.915 168.065 ;
        RECT 124.265 167.895 124.595 168.255 ;
        RECT 123.205 167.705 124.595 167.895 ;
        RECT 124.970 167.760 125.425 168.525 ;
        RECT 125.700 168.145 127.000 168.355 ;
        RECT 127.255 168.165 127.585 168.525 ;
        RECT 126.830 167.995 127.000 168.145 ;
        RECT 127.755 168.025 128.015 168.355 ;
        RECT 127.785 168.015 128.015 168.025 ;
        RECT 123.205 167.615 123.375 167.705 ;
        RECT 123.085 167.285 123.375 167.615 ;
        RECT 125.900 167.535 126.120 167.935 ;
        RECT 123.545 167.285 123.885 167.535 ;
        RECT 124.105 167.285 124.780 167.535 ;
        RECT 124.965 167.335 125.455 167.535 ;
        RECT 125.645 167.325 126.120 167.535 ;
        RECT 126.365 167.535 126.575 167.935 ;
        RECT 126.830 167.870 127.585 167.995 ;
        RECT 126.830 167.825 127.675 167.870 ;
        RECT 127.405 167.705 127.675 167.825 ;
        RECT 126.365 167.325 126.695 167.535 ;
        RECT 123.205 167.035 123.375 167.285 ;
        RECT 123.205 166.865 124.145 167.035 ;
        RECT 124.515 166.925 124.780 167.285 ;
        RECT 126.865 167.265 127.275 167.570 ;
        RECT 124.970 167.095 126.145 167.155 ;
        RECT 127.505 167.130 127.675 167.705 ;
        RECT 127.475 167.095 127.675 167.130 ;
        RECT 124.970 166.985 127.675 167.095 ;
        RECT 122.665 166.145 123.125 166.695 ;
        RECT 123.315 165.975 123.645 166.695 ;
        RECT 123.845 166.315 124.145 166.865 ;
        RECT 124.315 165.975 124.595 166.645 ;
        RECT 124.970 166.365 125.225 166.985 ;
        RECT 125.815 166.925 127.615 166.985 ;
        RECT 125.815 166.895 126.145 166.925 ;
        RECT 127.845 166.825 128.015 168.015 ;
        RECT 128.205 167.715 128.445 168.525 ;
        RECT 128.615 167.715 128.945 168.355 ;
        RECT 129.115 167.715 129.385 168.525 ;
        RECT 129.565 167.755 131.235 168.525 ;
        RECT 131.955 167.975 132.125 168.265 ;
        RECT 132.295 168.145 132.625 168.525 ;
        RECT 131.955 167.805 132.620 167.975 ;
        RECT 128.185 167.285 128.535 167.535 ;
        RECT 128.705 167.115 128.875 167.715 ;
        RECT 129.045 167.285 129.395 167.535 ;
        RECT 129.565 167.235 130.315 167.755 ;
        RECT 125.475 166.725 125.660 166.815 ;
        RECT 126.250 166.725 127.085 166.735 ;
        RECT 125.475 166.525 127.085 166.725 ;
        RECT 125.475 166.485 125.705 166.525 ;
        RECT 124.970 166.145 125.305 166.365 ;
        RECT 126.310 165.975 126.665 166.355 ;
        RECT 126.835 166.145 127.085 166.525 ;
        RECT 127.335 165.975 127.585 166.755 ;
        RECT 127.755 166.145 128.015 166.825 ;
        RECT 128.195 166.945 128.875 167.115 ;
        RECT 128.195 166.160 128.525 166.945 ;
        RECT 129.055 165.975 129.385 167.115 ;
        RECT 130.485 167.065 131.235 167.585 ;
        RECT 129.565 165.975 131.235 167.065 ;
        RECT 131.870 166.985 132.220 167.635 ;
        RECT 132.390 166.815 132.620 167.805 ;
        RECT 131.955 166.645 132.620 166.815 ;
        RECT 131.955 166.145 132.125 166.645 ;
        RECT 132.295 165.975 132.625 166.475 ;
        RECT 132.795 166.145 132.980 168.265 ;
        RECT 133.235 168.065 133.485 168.525 ;
        RECT 133.655 168.075 133.990 168.245 ;
        RECT 134.185 168.075 134.860 168.245 ;
        RECT 133.655 167.935 133.825 168.075 ;
        RECT 133.150 166.945 133.430 167.895 ;
        RECT 133.600 167.805 133.825 167.935 ;
        RECT 133.600 166.700 133.770 167.805 ;
        RECT 133.995 167.655 134.520 167.875 ;
        RECT 133.940 166.890 134.180 167.485 ;
        RECT 134.350 166.955 134.520 167.655 ;
        RECT 134.690 167.295 134.860 168.075 ;
        RECT 135.180 168.025 135.550 168.525 ;
        RECT 135.730 168.075 136.135 168.245 ;
        RECT 136.305 168.075 137.090 168.245 ;
        RECT 135.730 167.845 135.900 168.075 ;
        RECT 135.070 167.545 135.900 167.845 ;
        RECT 136.285 167.575 136.750 167.905 ;
        RECT 135.070 167.515 135.270 167.545 ;
        RECT 135.390 167.295 135.560 167.365 ;
        RECT 134.690 167.125 135.560 167.295 ;
        RECT 135.050 167.035 135.560 167.125 ;
        RECT 133.600 166.570 133.905 166.700 ;
        RECT 134.350 166.590 134.880 166.955 ;
        RECT 133.220 165.975 133.485 166.435 ;
        RECT 133.655 166.145 133.905 166.570 ;
        RECT 135.050 166.420 135.220 167.035 ;
        RECT 134.115 166.250 135.220 166.420 ;
        RECT 135.390 165.975 135.560 166.775 ;
        RECT 135.730 166.475 135.900 167.545 ;
        RECT 136.070 166.645 136.260 167.365 ;
        RECT 136.430 166.615 136.750 167.575 ;
        RECT 136.920 167.615 137.090 168.075 ;
        RECT 137.365 167.995 137.575 168.525 ;
        RECT 137.835 167.785 138.165 168.310 ;
        RECT 138.335 167.915 138.505 168.525 ;
        RECT 138.675 167.870 139.005 168.305 ;
        RECT 138.675 167.785 139.055 167.870 ;
        RECT 139.225 167.800 139.515 168.525 ;
        RECT 137.965 167.615 138.165 167.785 ;
        RECT 138.830 167.745 139.055 167.785 ;
        RECT 136.920 167.285 137.795 167.615 ;
        RECT 137.965 167.285 138.715 167.615 ;
        RECT 135.730 166.145 135.980 166.475 ;
        RECT 136.920 166.445 137.090 167.285 ;
        RECT 137.965 167.080 138.155 167.285 ;
        RECT 138.885 167.165 139.055 167.745 ;
        RECT 138.840 167.115 139.055 167.165 ;
        RECT 140.145 167.785 140.460 168.160 ;
        RECT 140.715 167.785 140.885 168.525 ;
        RECT 141.135 167.955 141.305 168.160 ;
        RECT 141.530 168.125 141.905 168.525 ;
        RECT 142.075 167.955 142.245 168.305 ;
        RECT 142.430 168.125 142.760 168.525 ;
        RECT 142.930 167.955 143.100 168.305 ;
        RECT 143.270 168.125 143.650 168.525 ;
        RECT 141.135 167.785 141.635 167.955 ;
        RECT 142.075 167.785 143.670 167.955 ;
        RECT 143.840 167.850 144.115 168.195 ;
        RECT 137.260 166.705 138.155 167.080 ;
        RECT 138.665 167.035 139.055 167.115 ;
        RECT 136.205 166.275 137.090 166.445 ;
        RECT 137.270 165.975 137.585 166.475 ;
        RECT 137.815 166.145 138.155 166.705 ;
        RECT 138.325 165.975 138.495 166.985 ;
        RECT 138.665 166.190 138.995 167.035 ;
        RECT 139.225 165.975 139.515 167.140 ;
        RECT 140.145 166.745 140.315 167.785 ;
        RECT 140.485 166.915 140.835 167.615 ;
        RECT 141.005 167.285 141.295 167.615 ;
        RECT 141.465 167.535 141.635 167.785 ;
        RECT 143.500 167.615 143.670 167.785 ;
        RECT 141.465 167.365 141.890 167.535 ;
        RECT 141.465 167.085 141.635 167.365 ;
        RECT 142.285 167.195 142.455 167.615 ;
        RECT 142.675 167.285 143.330 167.615 ;
        RECT 143.500 167.285 143.775 167.615 ;
        RECT 141.050 166.915 141.635 167.085 ;
        RECT 141.805 167.025 142.455 167.195 ;
        RECT 143.500 167.115 143.670 167.285 ;
        RECT 143.945 167.115 144.115 167.850 ;
        RECT 144.375 167.975 144.545 168.355 ;
        RECT 144.760 168.145 145.090 168.525 ;
        RECT 144.375 167.805 145.090 167.975 ;
        RECT 144.285 167.255 144.640 167.625 ;
        RECT 144.920 167.615 145.090 167.805 ;
        RECT 145.260 167.780 145.515 168.355 ;
        RECT 144.920 167.285 145.175 167.615 ;
        RECT 141.805 166.745 141.975 167.025 ;
        RECT 143.010 166.945 143.670 167.115 ;
        RECT 143.010 166.825 143.180 166.945 ;
        RECT 140.145 166.575 141.975 166.745 ;
        RECT 142.145 166.655 143.180 166.825 ;
        RECT 140.145 166.155 140.405 166.575 ;
        RECT 142.145 166.405 142.315 166.655 ;
        RECT 140.575 165.975 140.905 166.405 ;
        RECT 141.570 166.235 142.315 166.405 ;
        RECT 142.540 166.155 143.180 166.485 ;
        RECT 143.350 165.975 143.630 166.775 ;
        RECT 143.840 166.145 144.115 167.115 ;
        RECT 144.920 167.075 145.090 167.285 ;
        RECT 144.375 166.905 145.090 167.075 ;
        RECT 145.345 167.050 145.515 167.780 ;
        RECT 145.690 167.685 145.950 168.525 ;
        RECT 146.125 167.755 148.715 168.525 ;
        RECT 148.885 167.775 150.095 168.525 ;
        RECT 146.125 167.235 147.335 167.755 ;
        RECT 144.375 166.145 144.545 166.905 ;
        RECT 144.760 165.975 145.090 166.735 ;
        RECT 145.260 166.145 145.515 167.050 ;
        RECT 145.690 165.975 145.950 167.125 ;
        RECT 147.505 167.065 148.715 167.585 ;
        RECT 146.125 165.975 148.715 167.065 ;
        RECT 148.885 167.065 149.405 167.605 ;
        RECT 149.575 167.235 150.095 167.775 ;
        RECT 148.885 165.975 150.095 167.065 ;
        RECT 36.100 165.805 150.180 165.975 ;
        RECT 36.185 164.715 37.395 165.805 ;
        RECT 37.565 165.370 42.910 165.805 ;
        RECT 36.185 164.005 36.705 164.545 ;
        RECT 36.875 164.175 37.395 164.715 ;
        RECT 36.185 163.255 37.395 164.005 ;
        RECT 39.150 163.800 39.490 164.630 ;
        RECT 40.970 164.120 41.320 165.370 ;
        RECT 43.090 165.005 43.345 165.805 ;
        RECT 43.545 164.955 43.875 165.635 ;
        RECT 43.090 164.465 43.335 164.825 ;
        RECT 43.525 164.675 43.875 164.955 ;
        RECT 43.525 164.295 43.695 164.675 ;
        RECT 44.055 164.495 44.250 165.545 ;
        RECT 44.430 164.665 44.750 165.805 ;
        RECT 44.925 164.730 45.195 165.635 ;
        RECT 45.365 165.045 45.695 165.805 ;
        RECT 45.875 164.875 46.045 165.635 ;
        RECT 43.175 164.125 43.695 164.295 ;
        RECT 43.865 164.165 44.250 164.495 ;
        RECT 44.430 164.445 44.690 164.495 ;
        RECT 44.430 164.275 44.695 164.445 ;
        RECT 44.430 164.165 44.690 164.275 ;
        RECT 37.565 163.255 42.910 163.800 ;
        RECT 43.175 163.765 43.345 164.125 ;
        RECT 43.145 163.595 43.345 163.765 ;
        RECT 43.175 163.560 43.345 163.595 ;
        RECT 43.535 163.785 44.750 163.955 ;
        RECT 43.535 163.480 43.765 163.785 ;
        RECT 43.935 163.255 44.265 163.615 ;
        RECT 44.460 163.435 44.750 163.785 ;
        RECT 44.925 163.930 45.095 164.730 ;
        RECT 45.380 164.705 46.045 164.875 ;
        RECT 46.305 164.715 48.895 165.805 ;
        RECT 45.380 164.560 45.550 164.705 ;
        RECT 45.265 164.230 45.550 164.560 ;
        RECT 45.380 163.975 45.550 164.230 ;
        RECT 45.785 164.155 46.115 164.525 ;
        RECT 46.305 164.025 47.515 164.545 ;
        RECT 47.685 164.195 48.895 164.715 ;
        RECT 49.065 164.640 49.355 165.805 ;
        RECT 49.525 164.715 53.035 165.805 ;
        RECT 49.525 164.025 51.175 164.545 ;
        RECT 51.345 164.195 53.035 164.715 ;
        RECT 53.205 164.665 53.465 165.635 ;
        RECT 53.635 165.380 54.020 165.805 ;
        RECT 54.190 165.210 54.445 165.635 ;
        RECT 53.635 165.015 54.445 165.210 ;
        RECT 44.925 163.425 45.185 163.930 ;
        RECT 45.380 163.805 46.045 163.975 ;
        RECT 45.365 163.255 45.695 163.635 ;
        RECT 45.875 163.425 46.045 163.805 ;
        RECT 46.305 163.255 48.895 164.025 ;
        RECT 49.065 163.255 49.355 163.980 ;
        RECT 49.525 163.255 53.035 164.025 ;
        RECT 53.205 163.995 53.390 164.665 ;
        RECT 53.635 164.495 53.985 165.015 ;
        RECT 54.635 164.845 54.880 165.635 ;
        RECT 55.050 165.380 55.435 165.805 ;
        RECT 55.605 165.210 55.880 165.635 ;
        RECT 53.560 164.165 53.985 164.495 ;
        RECT 54.155 164.665 54.880 164.845 ;
        RECT 55.050 165.015 55.880 165.210 ;
        RECT 54.155 164.165 54.805 164.665 ;
        RECT 55.050 164.495 55.400 165.015 ;
        RECT 56.050 164.845 56.475 165.635 ;
        RECT 56.645 165.380 57.030 165.805 ;
        RECT 57.200 165.210 57.635 165.635 ;
        RECT 54.975 164.165 55.400 164.495 ;
        RECT 55.570 164.665 56.475 164.845 ;
        RECT 56.645 165.040 57.635 165.210 ;
        RECT 55.570 164.165 56.400 164.665 ;
        RECT 56.645 164.495 56.980 165.040 ;
        RECT 56.570 164.165 56.980 164.495 ;
        RECT 57.150 164.165 57.635 164.870 ;
        RECT 57.805 164.715 59.015 165.805 ;
        RECT 53.635 163.995 53.985 164.165 ;
        RECT 54.635 163.995 54.805 164.165 ;
        RECT 55.050 163.995 55.400 164.165 ;
        RECT 56.050 163.995 56.400 164.165 ;
        RECT 56.645 163.995 56.980 164.165 ;
        RECT 57.805 164.005 58.325 164.545 ;
        RECT 58.495 164.175 59.015 164.715 ;
        RECT 59.275 164.875 59.445 165.635 ;
        RECT 59.625 165.045 59.955 165.805 ;
        RECT 59.275 164.705 59.940 164.875 ;
        RECT 60.125 164.730 60.395 165.635 ;
        RECT 60.565 165.210 61.000 165.635 ;
        RECT 61.170 165.380 61.555 165.805 ;
        RECT 60.565 165.040 61.555 165.210 ;
        RECT 59.770 164.560 59.940 164.705 ;
        RECT 59.205 164.155 59.535 164.525 ;
        RECT 59.770 164.230 60.055 164.560 ;
        RECT 53.205 163.425 53.465 163.995 ;
        RECT 53.635 163.825 54.445 163.995 ;
        RECT 53.635 163.255 54.020 163.655 ;
        RECT 54.190 163.425 54.445 163.825 ;
        RECT 54.635 163.425 54.880 163.995 ;
        RECT 55.050 163.825 55.860 163.995 ;
        RECT 55.050 163.255 55.435 163.655 ;
        RECT 55.605 163.425 55.860 163.825 ;
        RECT 56.050 163.425 56.475 163.995 ;
        RECT 56.645 163.825 57.635 163.995 ;
        RECT 56.645 163.255 57.030 163.655 ;
        RECT 57.200 163.425 57.635 163.825 ;
        RECT 57.805 163.255 59.015 164.005 ;
        RECT 59.770 163.975 59.940 164.230 ;
        RECT 59.275 163.805 59.940 163.975 ;
        RECT 60.225 163.930 60.395 164.730 ;
        RECT 60.565 164.165 61.050 164.870 ;
        RECT 61.220 164.495 61.555 165.040 ;
        RECT 61.725 164.845 62.150 165.635 ;
        RECT 62.320 165.210 62.595 165.635 ;
        RECT 62.765 165.380 63.150 165.805 ;
        RECT 62.320 165.015 63.150 165.210 ;
        RECT 61.725 164.665 62.630 164.845 ;
        RECT 61.220 164.165 61.630 164.495 ;
        RECT 61.800 164.165 62.630 164.665 ;
        RECT 62.800 164.495 63.150 165.015 ;
        RECT 63.320 164.845 63.565 165.635 ;
        RECT 63.755 165.210 64.010 165.635 ;
        RECT 64.180 165.380 64.565 165.805 ;
        RECT 63.755 165.015 64.565 165.210 ;
        RECT 63.320 164.665 64.045 164.845 ;
        RECT 62.800 164.165 63.225 164.495 ;
        RECT 63.395 164.165 64.045 164.665 ;
        RECT 64.215 164.495 64.565 165.015 ;
        RECT 64.735 164.665 64.995 165.635 ;
        RECT 65.165 165.210 65.600 165.635 ;
        RECT 65.770 165.380 66.155 165.805 ;
        RECT 65.165 165.040 66.155 165.210 ;
        RECT 64.215 164.165 64.640 164.495 ;
        RECT 61.220 163.995 61.555 164.165 ;
        RECT 61.800 163.995 62.150 164.165 ;
        RECT 62.800 163.995 63.150 164.165 ;
        RECT 63.395 163.995 63.565 164.165 ;
        RECT 64.215 163.995 64.565 164.165 ;
        RECT 64.810 163.995 64.995 164.665 ;
        RECT 65.165 164.165 65.650 164.870 ;
        RECT 65.820 164.495 66.155 165.040 ;
        RECT 66.325 164.845 66.750 165.635 ;
        RECT 66.920 165.210 67.195 165.635 ;
        RECT 67.365 165.380 67.750 165.805 ;
        RECT 66.920 165.015 67.750 165.210 ;
        RECT 66.325 164.665 67.230 164.845 ;
        RECT 65.820 164.165 66.230 164.495 ;
        RECT 66.400 164.165 67.230 164.665 ;
        RECT 67.400 164.495 67.750 165.015 ;
        RECT 67.920 164.845 68.165 165.635 ;
        RECT 68.355 165.210 68.610 165.635 ;
        RECT 68.780 165.380 69.165 165.805 ;
        RECT 68.355 165.015 69.165 165.210 ;
        RECT 67.920 164.665 68.645 164.845 ;
        RECT 67.400 164.165 67.825 164.495 ;
        RECT 67.995 164.165 68.645 164.665 ;
        RECT 68.815 164.495 69.165 165.015 ;
        RECT 69.335 164.665 69.595 165.635 ;
        RECT 70.225 165.295 70.525 165.805 ;
        RECT 70.695 165.125 71.025 165.635 ;
        RECT 71.195 165.295 71.825 165.805 ;
        RECT 72.405 165.295 72.785 165.465 ;
        RECT 72.955 165.295 73.255 165.805 ;
        RECT 72.615 165.125 72.785 165.295 ;
        RECT 68.815 164.165 69.240 164.495 ;
        RECT 65.820 163.995 66.155 164.165 ;
        RECT 66.400 163.995 66.750 164.165 ;
        RECT 67.400 163.995 67.750 164.165 ;
        RECT 67.995 163.995 68.165 164.165 ;
        RECT 68.815 163.995 69.165 164.165 ;
        RECT 69.410 163.995 69.595 164.665 ;
        RECT 59.275 163.425 59.445 163.805 ;
        RECT 59.625 163.255 59.955 163.635 ;
        RECT 60.135 163.425 60.395 163.930 ;
        RECT 60.565 163.825 61.555 163.995 ;
        RECT 60.565 163.425 61.000 163.825 ;
        RECT 61.170 163.255 61.555 163.655 ;
        RECT 61.725 163.425 62.150 163.995 ;
        RECT 62.340 163.825 63.150 163.995 ;
        RECT 62.340 163.425 62.595 163.825 ;
        RECT 62.765 163.255 63.150 163.655 ;
        RECT 63.320 163.425 63.565 163.995 ;
        RECT 63.755 163.825 64.565 163.995 ;
        RECT 63.755 163.425 64.010 163.825 ;
        RECT 64.180 163.255 64.565 163.655 ;
        RECT 64.735 163.425 64.995 163.995 ;
        RECT 65.165 163.825 66.155 163.995 ;
        RECT 65.165 163.425 65.600 163.825 ;
        RECT 65.770 163.255 66.155 163.655 ;
        RECT 66.325 163.425 66.750 163.995 ;
        RECT 66.940 163.825 67.750 163.995 ;
        RECT 66.940 163.425 67.195 163.825 ;
        RECT 67.365 163.255 67.750 163.655 ;
        RECT 67.920 163.425 68.165 163.995 ;
        RECT 68.355 163.825 69.165 163.995 ;
        RECT 68.355 163.425 68.610 163.825 ;
        RECT 68.780 163.255 69.165 163.655 ;
        RECT 69.335 163.425 69.595 163.995 ;
        RECT 70.225 164.955 72.445 165.125 ;
        RECT 70.225 163.995 70.395 164.955 ;
        RECT 70.565 164.615 72.105 164.785 ;
        RECT 70.565 164.165 70.810 164.615 ;
        RECT 71.070 164.245 71.765 164.445 ;
        RECT 71.935 164.415 72.105 164.615 ;
        RECT 72.275 164.755 72.445 164.955 ;
        RECT 72.615 164.925 73.275 165.125 ;
        RECT 72.275 164.585 72.935 164.755 ;
        RECT 71.935 164.245 72.535 164.415 ;
        RECT 72.765 164.165 72.935 164.585 ;
        RECT 70.225 163.450 70.690 163.995 ;
        RECT 71.195 163.255 71.365 164.075 ;
        RECT 71.535 163.995 72.445 164.075 ;
        RECT 73.105 163.995 73.275 164.925 ;
        RECT 73.445 164.715 74.655 165.805 ;
        RECT 71.535 163.905 72.785 163.995 ;
        RECT 71.535 163.425 71.865 163.905 ;
        RECT 72.275 163.825 72.785 163.905 ;
        RECT 72.035 163.255 72.385 163.645 ;
        RECT 72.555 163.425 72.785 163.825 ;
        RECT 72.955 163.515 73.275 163.995 ;
        RECT 73.445 164.005 73.965 164.545 ;
        RECT 74.135 164.175 74.655 164.715 ;
        RECT 74.825 164.640 75.115 165.805 ;
        RECT 75.305 164.915 75.565 165.625 ;
        RECT 75.735 165.095 76.065 165.805 ;
        RECT 76.235 164.915 76.465 165.625 ;
        RECT 75.305 164.675 76.465 164.915 ;
        RECT 76.645 164.895 76.915 165.625 ;
        RECT 77.095 165.075 77.435 165.805 ;
        RECT 76.645 164.675 77.415 164.895 ;
        RECT 75.295 164.165 75.595 164.495 ;
        RECT 75.775 164.185 76.300 164.495 ;
        RECT 76.480 164.185 76.945 164.495 ;
        RECT 73.445 163.255 74.655 164.005 ;
        RECT 74.825 163.255 75.115 163.980 ;
        RECT 75.305 163.255 75.595 163.985 ;
        RECT 75.775 163.545 76.005 164.185 ;
        RECT 77.125 164.005 77.415 164.675 ;
        RECT 76.185 163.805 77.415 164.005 ;
        RECT 76.185 163.435 76.495 163.805 ;
        RECT 76.675 163.255 77.345 163.625 ;
        RECT 77.605 163.435 77.865 165.625 ;
        RECT 78.045 165.370 83.390 165.805 ;
        RECT 79.630 163.800 79.970 164.630 ;
        RECT 81.450 164.120 81.800 165.370 ;
        RECT 83.565 164.715 84.775 165.805 ;
        RECT 83.565 164.005 84.085 164.545 ;
        RECT 84.255 164.175 84.775 164.715 ;
        RECT 85.130 164.835 85.520 165.010 ;
        RECT 86.005 165.005 86.335 165.805 ;
        RECT 86.505 165.015 87.040 165.635 ;
        RECT 85.130 164.665 86.555 164.835 ;
        RECT 78.045 163.255 83.390 163.800 ;
        RECT 83.565 163.255 84.775 164.005 ;
        RECT 85.005 163.935 85.360 164.495 ;
        RECT 85.530 163.765 85.700 164.665 ;
        RECT 85.870 163.935 86.135 164.495 ;
        RECT 86.385 164.165 86.555 164.665 ;
        RECT 86.725 163.995 87.040 165.015 ;
        RECT 87.400 164.795 87.700 165.635 ;
        RECT 87.895 164.965 88.145 165.805 ;
        RECT 88.735 165.215 89.540 165.635 ;
        RECT 88.315 165.045 89.880 165.215 ;
        RECT 88.315 164.795 88.485 165.045 ;
        RECT 87.400 164.625 88.485 164.795 ;
        RECT 87.245 164.165 87.575 164.455 ;
        RECT 87.745 163.995 87.915 164.625 ;
        RECT 88.655 164.495 88.975 164.875 ;
        RECT 88.085 164.245 88.415 164.455 ;
        RECT 88.595 164.245 88.975 164.495 ;
        RECT 89.165 164.455 89.540 164.875 ;
        RECT 89.710 164.795 89.880 165.045 ;
        RECT 90.050 164.965 90.380 165.805 ;
        RECT 90.550 165.045 91.215 165.635 ;
        RECT 91.685 165.165 92.015 165.595 ;
        RECT 89.710 164.625 90.630 164.795 ;
        RECT 90.460 164.455 90.630 164.625 ;
        RECT 89.165 164.445 89.650 164.455 ;
        RECT 89.145 164.275 89.650 164.445 ;
        RECT 89.165 164.245 89.650 164.275 ;
        RECT 89.840 164.245 90.290 164.455 ;
        RECT 90.460 164.245 90.795 164.455 ;
        RECT 90.965 164.075 91.215 165.045 ;
        RECT 85.110 163.255 85.350 163.765 ;
        RECT 85.530 163.435 85.810 163.765 ;
        RECT 86.040 163.255 86.255 163.765 ;
        RECT 86.425 163.425 87.040 163.995 ;
        RECT 87.405 163.815 87.915 163.995 ;
        RECT 88.320 163.905 90.020 164.075 ;
        RECT 88.320 163.815 88.705 163.905 ;
        RECT 87.405 163.425 87.735 163.815 ;
        RECT 87.905 163.475 89.090 163.645 ;
        RECT 89.350 163.255 89.520 163.725 ;
        RECT 89.690 163.440 90.020 163.905 ;
        RECT 90.190 163.255 90.360 164.075 ;
        RECT 90.530 163.435 91.215 164.075 ;
        RECT 91.560 164.995 92.015 165.165 ;
        RECT 92.195 165.165 92.445 165.585 ;
        RECT 92.675 165.335 93.005 165.805 ;
        RECT 93.235 165.165 93.485 165.585 ;
        RECT 92.195 164.995 93.485 165.165 ;
        RECT 91.560 163.995 91.730 164.995 ;
        RECT 91.900 164.165 92.145 164.825 ;
        RECT 92.360 164.165 92.625 164.825 ;
        RECT 92.820 164.165 93.105 164.825 ;
        RECT 93.280 164.495 93.495 164.825 ;
        RECT 93.675 164.665 93.925 165.805 ;
        RECT 94.095 164.745 94.425 165.595 ;
        RECT 93.280 164.165 93.585 164.495 ;
        RECT 93.755 164.165 94.065 164.495 ;
        RECT 93.755 163.995 93.925 164.165 ;
        RECT 91.560 163.825 93.925 163.995 ;
        RECT 94.235 163.980 94.425 164.745 ;
        RECT 91.715 163.255 92.045 163.655 ;
        RECT 92.215 163.485 92.545 163.825 ;
        RECT 93.595 163.255 93.925 163.655 ;
        RECT 94.095 163.470 94.425 163.980 ;
        RECT 95.065 164.665 95.405 165.635 ;
        RECT 95.575 164.665 95.745 165.805 ;
        RECT 96.015 165.005 96.265 165.805 ;
        RECT 96.910 164.835 97.240 165.635 ;
        RECT 97.540 165.005 97.870 165.805 ;
        RECT 98.040 164.835 98.370 165.635 ;
        RECT 95.935 164.665 98.370 164.835 ;
        RECT 98.745 164.715 100.415 165.805 ;
        RECT 95.065 164.055 95.240 164.665 ;
        RECT 95.935 164.415 96.105 164.665 ;
        RECT 95.410 164.245 96.105 164.415 ;
        RECT 96.280 164.245 96.700 164.445 ;
        RECT 96.870 164.245 97.200 164.445 ;
        RECT 97.370 164.245 97.700 164.445 ;
        RECT 95.065 163.425 95.405 164.055 ;
        RECT 95.575 163.255 95.825 164.055 ;
        RECT 96.015 163.905 97.240 164.075 ;
        RECT 96.015 163.425 96.345 163.905 ;
        RECT 96.515 163.255 96.740 163.715 ;
        RECT 96.910 163.425 97.240 163.905 ;
        RECT 97.870 164.035 98.040 164.665 ;
        RECT 98.225 164.245 98.575 164.495 ;
        RECT 97.870 163.425 98.370 164.035 ;
        RECT 98.745 164.025 99.495 164.545 ;
        RECT 99.665 164.195 100.415 164.715 ;
        RECT 100.585 164.640 100.875 165.805 ;
        RECT 101.045 165.210 101.480 165.635 ;
        RECT 101.650 165.380 102.035 165.805 ;
        RECT 101.045 165.040 102.035 165.210 ;
        RECT 101.045 164.165 101.530 164.870 ;
        RECT 101.700 164.495 102.035 165.040 ;
        RECT 102.205 164.845 102.630 165.635 ;
        RECT 102.800 165.210 103.075 165.635 ;
        RECT 103.245 165.380 103.630 165.805 ;
        RECT 102.800 165.015 103.630 165.210 ;
        RECT 102.205 164.665 103.110 164.845 ;
        RECT 101.700 164.165 102.110 164.495 ;
        RECT 102.280 164.165 103.110 164.665 ;
        RECT 103.280 164.495 103.630 165.015 ;
        RECT 103.800 164.845 104.045 165.635 ;
        RECT 104.235 165.210 104.490 165.635 ;
        RECT 104.660 165.380 105.045 165.805 ;
        RECT 104.235 165.015 105.045 165.210 ;
        RECT 103.800 164.665 104.525 164.845 ;
        RECT 103.280 164.165 103.705 164.495 ;
        RECT 103.875 164.165 104.525 164.665 ;
        RECT 104.695 164.495 105.045 165.015 ;
        RECT 105.215 164.665 105.475 165.635 ;
        RECT 105.645 164.715 106.855 165.805 ;
        RECT 104.695 164.165 105.120 164.495 ;
        RECT 98.745 163.255 100.415 164.025 ;
        RECT 101.700 163.995 102.035 164.165 ;
        RECT 102.280 163.995 102.630 164.165 ;
        RECT 103.280 163.995 103.630 164.165 ;
        RECT 103.875 163.995 104.045 164.165 ;
        RECT 104.695 163.995 105.045 164.165 ;
        RECT 105.290 163.995 105.475 164.665 ;
        RECT 100.585 163.255 100.875 163.980 ;
        RECT 101.045 163.825 102.035 163.995 ;
        RECT 101.045 163.425 101.480 163.825 ;
        RECT 101.650 163.255 102.035 163.655 ;
        RECT 102.205 163.425 102.630 163.995 ;
        RECT 102.820 163.825 103.630 163.995 ;
        RECT 102.820 163.425 103.075 163.825 ;
        RECT 103.245 163.255 103.630 163.655 ;
        RECT 103.800 163.425 104.045 163.995 ;
        RECT 104.235 163.825 105.045 163.995 ;
        RECT 104.235 163.425 104.490 163.825 ;
        RECT 104.660 163.255 105.045 163.655 ;
        RECT 105.215 163.425 105.475 163.995 ;
        RECT 105.645 164.005 106.165 164.545 ;
        RECT 106.335 164.175 106.855 164.715 ;
        RECT 107.025 164.730 107.295 165.635 ;
        RECT 107.465 165.045 107.795 165.805 ;
        RECT 107.975 164.875 108.155 165.635 ;
        RECT 105.645 163.255 106.855 164.005 ;
        RECT 107.025 163.930 107.205 164.730 ;
        RECT 107.480 164.705 108.155 164.875 ;
        RECT 107.480 164.560 107.650 164.705 ;
        RECT 107.375 164.230 107.650 164.560 ;
        RECT 107.480 163.975 107.650 164.230 ;
        RECT 107.875 164.155 108.215 164.525 ;
        RECT 107.025 163.425 107.285 163.930 ;
        RECT 107.480 163.805 108.145 163.975 ;
        RECT 107.465 163.255 107.795 163.635 ;
        RECT 107.975 163.425 108.145 163.805 ;
        RECT 108.405 163.535 108.685 165.635 ;
        RECT 108.875 165.045 109.660 165.805 ;
        RECT 110.055 164.975 110.440 165.635 ;
        RECT 110.055 164.875 110.465 164.975 ;
        RECT 108.855 164.665 110.465 164.875 ;
        RECT 110.765 164.785 110.965 165.575 ;
        RECT 108.855 164.065 109.130 164.665 ;
        RECT 110.635 164.615 110.965 164.785 ;
        RECT 111.135 164.625 111.455 165.805 ;
        RECT 110.635 164.495 110.815 164.615 ;
        RECT 109.300 164.245 109.655 164.495 ;
        RECT 109.850 164.445 110.315 164.495 ;
        RECT 109.845 164.275 110.315 164.445 ;
        RECT 109.850 164.245 110.315 164.275 ;
        RECT 110.485 164.245 110.815 164.495 ;
        RECT 110.990 164.245 111.455 164.445 ;
        RECT 108.855 163.885 110.105 164.065 ;
        RECT 109.740 163.815 110.105 163.885 ;
        RECT 110.275 163.865 111.455 164.035 ;
        RECT 108.915 163.255 109.085 163.715 ;
        RECT 110.275 163.645 110.605 163.865 ;
        RECT 109.355 163.465 110.605 163.645 ;
        RECT 110.775 163.255 110.945 163.695 ;
        RECT 111.115 163.450 111.455 163.865 ;
        RECT 111.640 163.435 111.920 165.625 ;
        RECT 112.110 164.665 112.395 165.805 ;
        RECT 112.660 165.155 112.830 165.625 ;
        RECT 113.005 165.325 113.335 165.805 ;
        RECT 113.505 165.155 113.685 165.625 ;
        RECT 112.660 164.955 113.685 165.155 ;
        RECT 112.120 163.985 112.380 164.495 ;
        RECT 112.590 164.165 112.850 164.785 ;
        RECT 113.045 164.165 113.470 164.785 ;
        RECT 113.855 164.515 114.185 165.625 ;
        RECT 114.355 165.395 114.705 165.805 ;
        RECT 114.875 165.215 115.115 165.605 ;
        RECT 115.305 165.370 120.650 165.805 ;
        RECT 113.640 164.215 114.185 164.515 ;
        RECT 114.365 165.015 115.115 165.215 ;
        RECT 114.365 164.335 114.705 165.015 ;
        RECT 113.640 163.985 113.860 164.215 ;
        RECT 112.120 163.795 113.860 163.985 ;
        RECT 112.120 163.255 112.850 163.625 ;
        RECT 113.430 163.435 113.860 163.795 ;
        RECT 114.030 163.255 114.275 164.035 ;
        RECT 114.475 163.435 114.705 164.335 ;
        RECT 114.885 163.495 115.115 164.835 ;
        RECT 116.890 163.800 117.230 164.630 ;
        RECT 118.710 164.120 119.060 165.370 ;
        RECT 121.825 164.875 122.005 165.635 ;
        RECT 122.185 165.045 122.515 165.805 ;
        RECT 121.825 164.705 122.500 164.875 ;
        RECT 122.685 164.730 122.955 165.635 ;
        RECT 124.245 165.135 124.525 165.805 ;
        RECT 124.695 164.915 124.995 165.465 ;
        RECT 125.195 165.085 125.525 165.805 ;
        RECT 125.715 165.085 126.175 165.635 ;
        RECT 122.330 164.560 122.500 164.705 ;
        RECT 121.765 164.155 122.105 164.525 ;
        RECT 122.330 164.230 122.605 164.560 ;
        RECT 122.330 163.975 122.500 164.230 ;
        RECT 121.835 163.805 122.500 163.975 ;
        RECT 122.775 163.930 122.955 164.730 ;
        RECT 124.060 164.495 124.325 164.855 ;
        RECT 124.695 164.745 125.635 164.915 ;
        RECT 125.465 164.495 125.635 164.745 ;
        RECT 124.060 164.245 124.735 164.495 ;
        RECT 124.955 164.245 125.295 164.495 ;
        RECT 125.465 164.165 125.755 164.495 ;
        RECT 125.465 164.075 125.635 164.165 ;
        RECT 115.305 163.255 120.650 163.800 ;
        RECT 121.835 163.425 122.005 163.805 ;
        RECT 122.185 163.255 122.515 163.635 ;
        RECT 122.695 163.425 122.955 163.930 ;
        RECT 124.245 163.885 125.635 164.075 ;
        RECT 124.245 163.525 124.575 163.885 ;
        RECT 125.925 163.715 126.175 165.085 ;
        RECT 126.345 164.640 126.635 165.805 ;
        RECT 126.815 164.665 127.145 165.805 ;
        RECT 127.675 164.835 128.005 165.620 ;
        RECT 128.185 165.370 133.530 165.805 ;
        RECT 127.325 164.665 128.005 164.835 ;
        RECT 126.805 164.245 127.155 164.495 ;
        RECT 127.325 164.065 127.495 164.665 ;
        RECT 127.665 164.245 128.015 164.495 ;
        RECT 125.195 163.255 125.445 163.715 ;
        RECT 125.615 163.425 126.175 163.715 ;
        RECT 126.345 163.255 126.635 163.980 ;
        RECT 126.815 163.255 127.085 164.065 ;
        RECT 127.255 163.425 127.585 164.065 ;
        RECT 127.755 163.255 127.995 164.065 ;
        RECT 129.770 163.800 130.110 164.630 ;
        RECT 131.590 164.120 131.940 165.370 ;
        RECT 133.705 164.715 137.215 165.805 ;
        RECT 137.385 164.715 138.595 165.805 ;
        RECT 133.705 164.025 135.355 164.545 ;
        RECT 135.525 164.195 137.215 164.715 ;
        RECT 128.185 163.255 133.530 163.800 ;
        RECT 133.705 163.255 137.215 164.025 ;
        RECT 137.385 164.005 137.905 164.545 ;
        RECT 138.075 164.175 138.595 164.715 ;
        RECT 138.770 164.665 139.045 165.635 ;
        RECT 139.255 165.005 139.535 165.805 ;
        RECT 139.705 165.295 140.895 165.585 ;
        RECT 141.070 165.380 141.405 165.805 ;
        RECT 141.575 165.200 141.760 165.605 ;
        RECT 139.705 164.955 140.875 165.125 ;
        RECT 139.705 164.835 139.875 164.955 ;
        RECT 139.215 164.665 139.875 164.835 ;
        RECT 137.385 163.255 138.595 164.005 ;
        RECT 138.770 163.930 138.940 164.665 ;
        RECT 139.215 164.495 139.385 164.665 ;
        RECT 140.185 164.495 140.380 164.785 ;
        RECT 140.550 164.665 140.875 164.955 ;
        RECT 141.095 165.025 141.760 165.200 ;
        RECT 141.965 165.025 142.295 165.805 ;
        RECT 139.110 164.165 139.385 164.495 ;
        RECT 139.555 164.165 140.380 164.495 ;
        RECT 140.550 164.165 140.895 164.495 ;
        RECT 139.215 163.995 139.385 164.165 ;
        RECT 141.095 163.995 141.435 165.025 ;
        RECT 142.465 164.835 142.735 165.605 ;
        RECT 141.605 164.665 142.735 164.835 ;
        RECT 142.905 164.665 143.165 165.805 ;
        RECT 141.605 164.165 141.855 164.665 ;
        RECT 138.770 163.585 139.045 163.930 ;
        RECT 139.215 163.825 140.880 163.995 ;
        RECT 141.095 163.825 141.780 163.995 ;
        RECT 142.035 163.915 142.395 164.495 ;
        RECT 139.235 163.255 139.615 163.655 ;
        RECT 139.785 163.475 139.955 163.825 ;
        RECT 140.125 163.255 140.455 163.655 ;
        RECT 140.625 163.475 140.880 163.825 ;
        RECT 141.070 163.255 141.405 163.655 ;
        RECT 141.575 163.425 141.780 163.825 ;
        RECT 142.565 163.755 142.735 164.665 ;
        RECT 143.335 164.655 143.665 165.635 ;
        RECT 143.835 164.665 144.115 165.805 ;
        RECT 144.285 164.715 147.795 165.805 ;
        RECT 142.925 164.245 143.260 164.495 ;
        RECT 143.430 164.055 143.600 164.655 ;
        RECT 143.770 164.225 144.105 164.495 ;
        RECT 141.990 163.255 142.265 163.735 ;
        RECT 142.475 163.425 142.735 163.755 ;
        RECT 142.905 163.425 143.600 164.055 ;
        RECT 143.805 163.255 144.115 164.055 ;
        RECT 144.285 164.025 145.935 164.545 ;
        RECT 146.105 164.195 147.795 164.715 ;
        RECT 148.885 164.715 150.095 165.805 ;
        RECT 148.885 164.175 149.405 164.715 ;
        RECT 144.285 163.255 147.795 164.025 ;
        RECT 149.575 164.005 150.095 164.545 ;
        RECT 148.885 163.255 150.095 164.005 ;
        RECT 36.100 163.085 150.180 163.255 ;
        RECT 36.185 162.335 37.395 163.085 ;
        RECT 36.185 161.795 36.705 162.335 ;
        RECT 37.565 162.315 39.235 163.085 ;
        RECT 39.955 162.535 40.125 162.825 ;
        RECT 40.295 162.705 40.625 163.085 ;
        RECT 39.955 162.365 40.620 162.535 ;
        RECT 36.875 161.625 37.395 162.165 ;
        RECT 37.565 161.795 38.315 162.315 ;
        RECT 38.485 161.625 39.235 162.145 ;
        RECT 36.185 160.535 37.395 161.625 ;
        RECT 37.565 160.535 39.235 161.625 ;
        RECT 39.870 161.545 40.220 162.195 ;
        RECT 40.390 161.375 40.620 162.365 ;
        RECT 39.955 161.205 40.620 161.375 ;
        RECT 39.955 160.705 40.125 161.205 ;
        RECT 40.295 160.535 40.625 161.035 ;
        RECT 40.795 160.705 40.980 162.825 ;
        RECT 41.235 162.625 41.485 163.085 ;
        RECT 41.655 162.635 41.990 162.805 ;
        RECT 42.185 162.635 42.860 162.805 ;
        RECT 41.655 162.495 41.825 162.635 ;
        RECT 41.150 161.505 41.430 162.455 ;
        RECT 41.600 162.365 41.825 162.495 ;
        RECT 41.600 161.260 41.770 162.365 ;
        RECT 41.995 162.215 42.520 162.435 ;
        RECT 41.940 161.450 42.180 162.045 ;
        RECT 42.350 161.515 42.520 162.215 ;
        RECT 42.690 161.855 42.860 162.635 ;
        RECT 43.180 162.585 43.550 163.085 ;
        RECT 43.730 162.635 44.135 162.805 ;
        RECT 44.305 162.635 45.090 162.805 ;
        RECT 43.730 162.405 43.900 162.635 ;
        RECT 43.070 162.105 43.900 162.405 ;
        RECT 44.285 162.135 44.750 162.465 ;
        RECT 43.070 162.075 43.270 162.105 ;
        RECT 43.390 161.855 43.560 161.925 ;
        RECT 42.690 161.685 43.560 161.855 ;
        RECT 43.050 161.595 43.560 161.685 ;
        RECT 41.600 161.130 41.905 161.260 ;
        RECT 42.350 161.150 42.880 161.515 ;
        RECT 41.220 160.535 41.485 160.995 ;
        RECT 41.655 160.705 41.905 161.130 ;
        RECT 43.050 160.980 43.220 161.595 ;
        RECT 42.115 160.810 43.220 160.980 ;
        RECT 43.390 160.535 43.560 161.335 ;
        RECT 43.730 161.035 43.900 162.105 ;
        RECT 44.070 161.205 44.260 161.925 ;
        RECT 44.430 161.175 44.750 162.135 ;
        RECT 44.920 162.175 45.090 162.635 ;
        RECT 45.365 162.555 45.575 163.085 ;
        RECT 45.835 162.345 46.165 162.870 ;
        RECT 46.335 162.475 46.505 163.085 ;
        RECT 46.675 162.430 47.005 162.865 ;
        RECT 46.675 162.345 47.055 162.430 ;
        RECT 45.965 162.175 46.165 162.345 ;
        RECT 46.830 162.305 47.055 162.345 ;
        RECT 44.920 161.845 45.795 162.175 ;
        RECT 45.965 161.845 46.715 162.175 ;
        RECT 43.730 160.705 43.980 161.035 ;
        RECT 44.920 161.005 45.090 161.845 ;
        RECT 45.965 161.640 46.155 161.845 ;
        RECT 46.885 161.725 47.055 162.305 ;
        RECT 47.225 162.315 49.815 163.085 ;
        RECT 50.445 162.410 50.705 162.915 ;
        RECT 50.885 162.705 51.215 163.085 ;
        RECT 51.395 162.535 51.565 162.915 ;
        RECT 47.225 161.795 48.435 162.315 ;
        RECT 46.840 161.675 47.055 161.725 ;
        RECT 45.260 161.265 46.155 161.640 ;
        RECT 46.665 161.595 47.055 161.675 ;
        RECT 48.605 161.625 49.815 162.145 ;
        RECT 44.205 160.835 45.090 161.005 ;
        RECT 45.270 160.535 45.585 161.035 ;
        RECT 45.815 160.705 46.155 161.265 ;
        RECT 46.325 160.535 46.495 161.545 ;
        RECT 46.665 160.750 46.995 161.595 ;
        RECT 47.225 160.535 49.815 161.625 ;
        RECT 50.445 161.610 50.625 162.410 ;
        RECT 50.900 162.365 51.565 162.535 ;
        RECT 51.825 162.515 52.260 162.915 ;
        RECT 52.430 162.685 52.815 163.085 ;
        RECT 50.900 162.110 51.070 162.365 ;
        RECT 51.825 162.345 52.815 162.515 ;
        RECT 52.985 162.345 53.410 162.915 ;
        RECT 53.600 162.515 53.855 162.915 ;
        RECT 54.025 162.685 54.410 163.085 ;
        RECT 53.600 162.345 54.410 162.515 ;
        RECT 54.580 162.345 54.825 162.915 ;
        RECT 55.015 162.515 55.270 162.915 ;
        RECT 55.440 162.685 55.825 163.085 ;
        RECT 55.015 162.345 55.825 162.515 ;
        RECT 55.995 162.345 56.255 162.915 ;
        RECT 50.795 161.780 51.070 162.110 ;
        RECT 51.295 161.815 51.635 162.185 ;
        RECT 52.480 162.175 52.815 162.345 ;
        RECT 53.060 162.175 53.410 162.345 ;
        RECT 54.060 162.175 54.410 162.345 ;
        RECT 54.655 162.175 54.825 162.345 ;
        RECT 55.475 162.175 55.825 162.345 ;
        RECT 50.900 161.635 51.070 161.780 ;
        RECT 50.445 160.705 50.715 161.610 ;
        RECT 50.900 161.465 51.575 161.635 ;
        RECT 51.825 161.470 52.310 162.175 ;
        RECT 52.480 161.845 52.890 162.175 ;
        RECT 50.885 160.535 51.215 161.295 ;
        RECT 51.395 160.705 51.575 161.465 ;
        RECT 52.480 161.300 52.815 161.845 ;
        RECT 53.060 161.675 53.890 162.175 ;
        RECT 51.825 161.130 52.815 161.300 ;
        RECT 52.985 161.495 53.890 161.675 ;
        RECT 54.060 161.845 54.485 162.175 ;
        RECT 51.825 160.705 52.260 161.130 ;
        RECT 52.430 160.535 52.815 160.960 ;
        RECT 52.985 160.705 53.410 161.495 ;
        RECT 54.060 161.325 54.410 161.845 ;
        RECT 54.655 161.675 55.305 162.175 ;
        RECT 53.580 161.130 54.410 161.325 ;
        RECT 54.580 161.495 55.305 161.675 ;
        RECT 55.475 161.845 55.900 162.175 ;
        RECT 53.580 160.705 53.855 161.130 ;
        RECT 54.025 160.535 54.410 160.960 ;
        RECT 54.580 160.705 54.825 161.495 ;
        RECT 55.475 161.325 55.825 161.845 ;
        RECT 56.070 161.675 56.255 162.345 ;
        RECT 56.625 162.455 56.955 162.815 ;
        RECT 57.575 162.625 57.825 163.085 ;
        RECT 57.995 162.625 58.555 162.915 ;
        RECT 56.625 162.265 58.015 162.455 ;
        RECT 57.845 162.175 58.015 162.265 ;
        RECT 55.015 161.130 55.825 161.325 ;
        RECT 55.015 160.705 55.270 161.130 ;
        RECT 55.440 160.535 55.825 160.960 ;
        RECT 55.995 160.705 56.255 161.675 ;
        RECT 56.440 161.845 57.115 162.095 ;
        RECT 57.335 161.845 57.675 162.095 ;
        RECT 57.845 161.845 58.135 162.175 ;
        RECT 56.440 161.485 56.705 161.845 ;
        RECT 57.845 161.595 58.015 161.845 ;
        RECT 57.075 161.425 58.015 161.595 ;
        RECT 56.625 160.535 56.905 161.205 ;
        RECT 57.075 160.875 57.375 161.425 ;
        RECT 58.305 161.255 58.555 162.625 ;
        RECT 58.725 162.335 59.935 163.085 ;
        RECT 60.195 162.535 60.365 162.915 ;
        RECT 60.545 162.705 60.875 163.085 ;
        RECT 60.195 162.365 60.860 162.535 ;
        RECT 61.055 162.410 61.315 162.915 ;
        RECT 58.725 161.795 59.245 162.335 ;
        RECT 59.415 161.625 59.935 162.165 ;
        RECT 60.125 161.815 60.465 162.185 ;
        RECT 60.690 162.110 60.860 162.365 ;
        RECT 60.690 161.780 60.965 162.110 ;
        RECT 60.690 161.635 60.860 161.780 ;
        RECT 57.575 160.535 57.905 161.255 ;
        RECT 58.095 160.705 58.555 161.255 ;
        RECT 58.725 160.535 59.935 161.625 ;
        RECT 60.185 161.465 60.860 161.635 ;
        RECT 61.135 161.610 61.315 162.410 ;
        RECT 61.945 162.360 62.235 163.085 ;
        RECT 62.445 162.265 62.675 163.085 ;
        RECT 62.845 162.285 63.175 162.915 ;
        RECT 62.425 161.845 62.755 162.095 ;
        RECT 60.185 160.705 60.365 161.465 ;
        RECT 60.545 160.535 60.875 161.295 ;
        RECT 61.045 160.705 61.315 161.610 ;
        RECT 61.945 160.535 62.235 161.700 ;
        RECT 62.925 161.685 63.175 162.285 ;
        RECT 63.345 162.265 63.555 163.085 ;
        RECT 63.785 162.315 66.375 163.085 ;
        RECT 67.055 162.695 67.385 163.085 ;
        RECT 67.555 162.515 67.725 162.835 ;
        RECT 67.895 162.695 68.225 163.085 ;
        RECT 68.640 162.685 69.595 162.855 ;
        RECT 67.005 162.345 69.255 162.515 ;
        RECT 63.785 161.795 64.995 162.315 ;
        RECT 62.445 160.535 62.675 161.675 ;
        RECT 62.845 160.705 63.175 161.685 ;
        RECT 63.345 160.535 63.555 161.675 ;
        RECT 65.165 161.625 66.375 162.145 ;
        RECT 63.785 160.535 66.375 161.625 ;
        RECT 67.005 161.385 67.175 162.345 ;
        RECT 67.345 161.725 67.590 162.175 ;
        RECT 67.760 161.895 68.310 162.095 ;
        RECT 68.480 161.925 68.855 162.095 ;
        RECT 68.480 161.725 68.650 161.925 ;
        RECT 69.025 161.845 69.255 162.345 ;
        RECT 67.345 161.555 68.650 161.725 ;
        RECT 69.425 161.805 69.595 162.685 ;
        RECT 69.765 162.250 70.055 163.085 ;
        RECT 70.425 162.455 70.755 162.815 ;
        RECT 71.375 162.625 71.625 163.085 ;
        RECT 71.795 162.625 72.355 162.915 ;
        RECT 70.425 162.265 71.815 162.455 ;
        RECT 71.645 162.175 71.815 162.265 ;
        RECT 70.240 161.845 70.915 162.095 ;
        RECT 71.135 161.845 71.475 162.095 ;
        RECT 71.645 161.845 71.935 162.175 ;
        RECT 69.425 161.635 70.055 161.805 ;
        RECT 67.005 160.705 67.385 161.385 ;
        RECT 67.975 160.535 68.145 161.385 ;
        RECT 68.315 161.215 69.555 161.385 ;
        RECT 68.315 160.705 68.645 161.215 ;
        RECT 68.815 160.535 68.985 161.045 ;
        RECT 69.155 160.705 69.555 161.215 ;
        RECT 69.735 160.705 70.055 161.635 ;
        RECT 70.240 161.485 70.505 161.845 ;
        RECT 71.645 161.595 71.815 161.845 ;
        RECT 70.875 161.425 71.815 161.595 ;
        RECT 70.425 160.535 70.705 161.205 ;
        RECT 70.875 160.875 71.175 161.425 ;
        RECT 72.105 161.255 72.355 162.625 ;
        RECT 72.525 162.540 77.870 163.085 ;
        RECT 78.045 162.540 83.390 163.085 ;
        RECT 74.110 161.710 74.450 162.540 ;
        RECT 71.375 160.535 71.705 161.255 ;
        RECT 71.895 160.705 72.355 161.255 ;
        RECT 75.930 160.970 76.280 162.220 ;
        RECT 79.630 161.710 79.970 162.540 ;
        RECT 83.565 162.315 86.155 163.085 ;
        RECT 86.415 162.535 86.585 162.915 ;
        RECT 86.765 162.705 87.095 163.085 ;
        RECT 86.415 162.365 87.080 162.535 ;
        RECT 87.275 162.410 87.535 162.915 ;
        RECT 81.450 160.970 81.800 162.220 ;
        RECT 83.565 161.795 84.775 162.315 ;
        RECT 84.945 161.625 86.155 162.145 ;
        RECT 86.345 161.815 86.685 162.185 ;
        RECT 86.910 162.110 87.080 162.365 ;
        RECT 86.910 161.780 87.185 162.110 ;
        RECT 86.910 161.635 87.080 161.780 ;
        RECT 72.525 160.535 77.870 160.970 ;
        RECT 78.045 160.535 83.390 160.970 ;
        RECT 83.565 160.535 86.155 161.625 ;
        RECT 86.405 161.465 87.080 161.635 ;
        RECT 87.355 161.610 87.535 162.410 ;
        RECT 87.705 162.360 87.995 163.085 ;
        RECT 88.165 162.315 91.675 163.085 ;
        RECT 88.165 161.795 89.815 162.315 ;
        RECT 91.845 162.285 92.155 163.085 ;
        RECT 92.360 162.285 93.055 162.915 ;
        RECT 93.225 162.315 96.735 163.085 ;
        RECT 97.365 162.455 97.705 162.915 ;
        RECT 97.875 162.625 98.045 163.085 ;
        RECT 98.675 162.650 99.035 162.915 ;
        RECT 98.680 162.645 99.035 162.650 ;
        RECT 98.685 162.635 99.035 162.645 ;
        RECT 98.690 162.630 99.035 162.635 ;
        RECT 98.695 162.620 99.035 162.630 ;
        RECT 99.275 162.625 99.445 163.085 ;
        RECT 98.700 162.615 99.035 162.620 ;
        RECT 98.710 162.605 99.035 162.615 ;
        RECT 98.720 162.595 99.035 162.605 ;
        RECT 98.215 162.455 98.545 162.535 ;
        RECT 86.405 160.705 86.585 161.465 ;
        RECT 86.765 160.535 87.095 161.295 ;
        RECT 87.265 160.705 87.535 161.610 ;
        RECT 87.705 160.535 87.995 161.700 ;
        RECT 89.985 161.625 91.675 162.145 ;
        RECT 91.855 161.845 92.190 162.115 ;
        RECT 92.360 161.685 92.530 162.285 ;
        RECT 92.700 161.845 93.035 162.095 ;
        RECT 93.225 161.795 94.875 162.315 ;
        RECT 97.365 162.265 98.545 162.455 ;
        RECT 98.735 162.455 99.035 162.595 ;
        RECT 98.735 162.265 99.445 162.455 ;
        RECT 88.165 160.535 91.675 161.625 ;
        RECT 91.845 160.535 92.125 161.675 ;
        RECT 92.295 160.705 92.625 161.685 ;
        RECT 92.795 160.535 93.055 161.675 ;
        RECT 95.045 161.625 96.735 162.145 ;
        RECT 93.225 160.535 96.735 161.625 ;
        RECT 97.365 161.895 97.695 162.095 ;
        RECT 98.005 162.075 98.335 162.095 ;
        RECT 97.885 161.895 98.335 162.075 ;
        RECT 97.365 161.555 97.595 161.895 ;
        RECT 97.375 160.535 97.705 161.255 ;
        RECT 97.885 160.780 98.100 161.895 ;
        RECT 98.505 161.865 98.975 162.095 ;
        RECT 99.160 161.695 99.445 162.265 ;
        RECT 99.615 162.140 99.955 162.915 ;
        RECT 98.295 161.480 99.445 161.695 ;
        RECT 98.295 160.705 98.625 161.480 ;
        RECT 98.795 160.535 99.505 161.310 ;
        RECT 99.675 160.705 99.955 162.140 ;
        RECT 101.045 160.705 101.325 162.805 ;
        RECT 101.555 162.625 101.725 163.085 ;
        RECT 101.995 162.695 103.245 162.875 ;
        RECT 102.380 162.455 102.745 162.525 ;
        RECT 101.495 162.275 102.745 162.455 ;
        RECT 102.915 162.475 103.245 162.695 ;
        RECT 103.415 162.645 103.585 163.085 ;
        RECT 103.755 162.475 104.095 162.890 ;
        RECT 102.915 162.305 104.095 162.475 ;
        RECT 104.265 162.410 104.525 162.915 ;
        RECT 104.705 162.705 105.035 163.085 ;
        RECT 105.215 162.535 105.385 162.915 ;
        RECT 101.495 161.675 101.770 162.275 ;
        RECT 101.940 161.845 102.295 162.095 ;
        RECT 102.490 162.065 102.955 162.095 ;
        RECT 102.485 161.895 102.955 162.065 ;
        RECT 102.490 161.845 102.955 161.895 ;
        RECT 103.125 161.845 103.455 162.095 ;
        RECT 103.630 161.895 104.095 162.095 ;
        RECT 103.275 161.725 103.455 161.845 ;
        RECT 101.495 161.465 103.105 161.675 ;
        RECT 103.275 161.555 103.605 161.725 ;
        RECT 102.695 161.365 103.105 161.465 ;
        RECT 101.515 160.535 102.300 161.295 ;
        RECT 102.695 160.705 103.080 161.365 ;
        RECT 103.405 160.765 103.605 161.555 ;
        RECT 103.775 160.535 104.095 161.715 ;
        RECT 104.265 161.610 104.445 162.410 ;
        RECT 104.720 162.365 105.385 162.535 ;
        RECT 104.720 162.110 104.890 162.365 ;
        RECT 105.645 162.315 109.155 163.085 ;
        RECT 109.485 162.525 109.815 162.915 ;
        RECT 109.985 162.695 111.170 162.865 ;
        RECT 111.430 162.615 111.600 163.085 ;
        RECT 109.485 162.345 109.995 162.525 ;
        RECT 104.615 161.780 104.890 162.110 ;
        RECT 105.115 161.815 105.455 162.185 ;
        RECT 105.645 161.795 107.295 162.315 ;
        RECT 104.720 161.635 104.890 161.780 ;
        RECT 104.265 160.705 104.535 161.610 ;
        RECT 104.720 161.465 105.395 161.635 ;
        RECT 107.465 161.625 109.155 162.145 ;
        RECT 109.325 161.885 109.655 162.175 ;
        RECT 109.825 161.715 109.995 162.345 ;
        RECT 110.400 162.435 110.785 162.525 ;
        RECT 111.770 162.435 112.100 162.900 ;
        RECT 110.400 162.265 112.100 162.435 ;
        RECT 112.270 162.265 112.440 163.085 ;
        RECT 112.610 162.265 113.295 162.905 ;
        RECT 113.465 162.360 113.755 163.085 ;
        RECT 114.085 162.525 114.415 162.915 ;
        RECT 114.585 162.695 115.770 162.865 ;
        RECT 116.030 162.615 116.200 163.085 ;
        RECT 114.085 162.345 114.595 162.525 ;
        RECT 110.165 161.885 110.495 162.095 ;
        RECT 110.675 161.845 111.055 162.095 ;
        RECT 111.245 162.065 111.730 162.095 ;
        RECT 111.225 161.895 111.730 162.065 ;
        RECT 104.705 160.535 105.035 161.295 ;
        RECT 105.215 160.705 105.395 161.465 ;
        RECT 105.645 160.535 109.155 161.625 ;
        RECT 109.480 161.545 110.565 161.715 ;
        RECT 109.480 160.705 109.780 161.545 ;
        RECT 109.975 160.535 110.225 161.375 ;
        RECT 110.395 161.295 110.565 161.545 ;
        RECT 110.735 161.465 111.055 161.845 ;
        RECT 111.245 161.885 111.730 161.895 ;
        RECT 111.920 161.885 112.370 162.095 ;
        RECT 112.540 161.885 112.875 162.095 ;
        RECT 111.245 161.465 111.620 161.885 ;
        RECT 112.540 161.715 112.710 161.885 ;
        RECT 111.790 161.545 112.710 161.715 ;
        RECT 111.790 161.295 111.960 161.545 ;
        RECT 110.395 161.125 111.960 161.295 ;
        RECT 110.815 160.705 111.620 161.125 ;
        RECT 112.130 160.535 112.460 161.375 ;
        RECT 113.045 161.295 113.295 162.265 ;
        RECT 113.925 161.885 114.255 162.175 ;
        RECT 114.425 161.715 114.595 162.345 ;
        RECT 115.000 162.435 115.385 162.525 ;
        RECT 116.370 162.435 116.700 162.900 ;
        RECT 115.000 162.265 116.700 162.435 ;
        RECT 116.870 162.265 117.040 163.085 ;
        RECT 117.210 162.265 117.895 162.905 ;
        RECT 118.065 162.540 123.410 163.085 ;
        RECT 123.595 162.585 123.925 163.085 ;
        RECT 114.765 161.885 115.095 162.095 ;
        RECT 115.275 161.845 115.655 162.095 ;
        RECT 115.845 162.065 116.330 162.095 ;
        RECT 115.825 161.895 116.330 162.065 ;
        RECT 112.630 160.705 113.295 161.295 ;
        RECT 113.465 160.535 113.755 161.700 ;
        RECT 114.080 161.545 115.165 161.715 ;
        RECT 114.080 160.705 114.380 161.545 ;
        RECT 114.575 160.535 114.825 161.375 ;
        RECT 114.995 161.295 115.165 161.545 ;
        RECT 115.335 161.465 115.655 161.845 ;
        RECT 115.845 161.885 116.330 161.895 ;
        RECT 116.520 161.885 116.970 162.095 ;
        RECT 117.140 161.885 117.475 162.095 ;
        RECT 115.845 161.465 116.220 161.885 ;
        RECT 117.140 161.715 117.310 161.885 ;
        RECT 116.390 161.545 117.310 161.715 ;
        RECT 116.390 161.295 116.560 161.545 ;
        RECT 114.995 161.125 116.560 161.295 ;
        RECT 115.415 160.705 116.220 161.125 ;
        RECT 116.730 160.535 117.060 161.375 ;
        RECT 117.645 161.295 117.895 162.265 ;
        RECT 119.650 161.710 119.990 162.540 ;
        RECT 124.125 162.515 124.295 162.865 ;
        RECT 124.495 162.685 124.825 163.085 ;
        RECT 124.995 162.515 125.165 162.865 ;
        RECT 125.335 162.685 125.715 163.085 ;
        RECT 117.230 160.705 117.895 161.295 ;
        RECT 121.470 160.970 121.820 162.220 ;
        RECT 123.590 161.845 123.940 162.415 ;
        RECT 124.125 162.345 125.735 162.515 ;
        RECT 125.905 162.410 126.175 162.755 ;
        RECT 125.565 162.175 125.735 162.345 ;
        RECT 123.590 161.385 123.910 161.675 ;
        RECT 124.110 161.555 124.820 162.175 ;
        RECT 124.990 161.845 125.395 162.175 ;
        RECT 125.565 161.845 125.835 162.175 ;
        RECT 125.565 161.675 125.735 161.845 ;
        RECT 126.005 161.675 126.175 162.410 ;
        RECT 126.345 162.335 127.555 163.085 ;
        RECT 127.725 162.410 127.985 162.915 ;
        RECT 128.165 162.705 128.495 163.085 ;
        RECT 128.675 162.535 128.845 162.915 ;
        RECT 126.345 161.795 126.865 162.335 ;
        RECT 125.010 161.505 125.735 161.675 ;
        RECT 125.010 161.385 125.180 161.505 ;
        RECT 123.590 161.215 125.180 161.385 ;
        RECT 118.065 160.535 123.410 160.970 ;
        RECT 123.590 160.755 125.245 161.045 ;
        RECT 125.415 160.535 125.695 161.335 ;
        RECT 125.905 160.705 126.175 161.675 ;
        RECT 127.035 161.625 127.555 162.165 ;
        RECT 126.345 160.535 127.555 161.625 ;
        RECT 127.725 161.610 127.905 162.410 ;
        RECT 128.180 162.365 128.845 162.535 ;
        RECT 128.180 162.110 128.350 162.365 ;
        RECT 129.105 162.315 130.775 163.085 ;
        RECT 130.950 162.555 131.240 162.905 ;
        RECT 131.435 162.725 131.765 163.085 ;
        RECT 131.935 162.555 132.165 162.860 ;
        RECT 130.950 162.385 132.165 162.555 ;
        RECT 128.075 161.780 128.350 162.110 ;
        RECT 128.575 161.815 128.915 162.185 ;
        RECT 129.105 161.795 129.855 162.315 ;
        RECT 132.355 162.215 132.525 162.780 ;
        RECT 128.180 161.635 128.350 161.780 ;
        RECT 127.725 160.705 127.995 161.610 ;
        RECT 128.180 161.465 128.855 161.635 ;
        RECT 130.025 161.625 130.775 162.145 ;
        RECT 131.010 162.065 131.270 162.175 ;
        RECT 131.005 161.895 131.270 162.065 ;
        RECT 131.010 161.845 131.270 161.895 ;
        RECT 131.450 161.845 131.835 162.175 ;
        RECT 132.005 162.045 132.525 162.215 ;
        RECT 132.785 162.315 134.455 163.085 ;
        RECT 128.165 160.535 128.495 161.295 ;
        RECT 128.675 160.705 128.855 161.465 ;
        RECT 129.105 160.535 130.775 161.625 ;
        RECT 130.950 160.535 131.270 161.675 ;
        RECT 131.450 160.795 131.645 161.845 ;
        RECT 132.005 161.665 132.175 162.045 ;
        RECT 131.825 161.385 132.175 161.665 ;
        RECT 132.365 161.515 132.610 161.875 ;
        RECT 132.785 161.795 133.535 162.315 ;
        RECT 133.705 161.625 134.455 162.145 ;
        RECT 131.825 160.705 132.155 161.385 ;
        RECT 132.355 160.535 132.610 161.335 ;
        RECT 132.785 160.535 134.455 161.625 ;
        RECT 134.625 160.705 135.375 162.915 ;
        RECT 136.475 162.585 136.805 163.085 ;
        RECT 137.005 162.515 137.175 162.865 ;
        RECT 137.375 162.685 137.705 163.085 ;
        RECT 137.875 162.515 138.045 162.865 ;
        RECT 138.215 162.685 138.595 163.085 ;
        RECT 136.470 161.845 136.820 162.415 ;
        RECT 137.005 162.345 138.615 162.515 ;
        RECT 138.785 162.410 139.055 162.755 ;
        RECT 138.445 162.175 138.615 162.345 ;
        RECT 136.470 161.385 136.790 161.675 ;
        RECT 136.990 161.555 137.700 162.175 ;
        RECT 137.870 161.845 138.275 162.175 ;
        RECT 138.445 161.845 138.715 162.175 ;
        RECT 138.445 161.675 138.615 161.845 ;
        RECT 138.885 161.675 139.055 162.410 ;
        RECT 139.225 162.360 139.515 163.085 ;
        RECT 139.775 162.535 139.945 162.825 ;
        RECT 140.115 162.705 140.445 163.085 ;
        RECT 139.775 162.365 140.440 162.535 ;
        RECT 137.890 161.505 138.615 161.675 ;
        RECT 137.890 161.385 138.060 161.505 ;
        RECT 136.470 161.215 138.060 161.385 ;
        RECT 136.470 160.755 138.125 161.045 ;
        RECT 138.295 160.535 138.575 161.335 ;
        RECT 138.785 160.705 139.055 161.675 ;
        RECT 139.225 160.535 139.515 161.700 ;
        RECT 139.690 161.545 140.040 162.195 ;
        RECT 140.210 161.375 140.440 162.365 ;
        RECT 139.775 161.205 140.440 161.375 ;
        RECT 139.775 160.705 139.945 161.205 ;
        RECT 140.115 160.535 140.445 161.035 ;
        RECT 140.615 160.705 140.800 162.825 ;
        RECT 141.055 162.625 141.305 163.085 ;
        RECT 141.475 162.635 141.810 162.805 ;
        RECT 142.005 162.635 142.680 162.805 ;
        RECT 141.475 162.495 141.645 162.635 ;
        RECT 140.970 161.505 141.250 162.455 ;
        RECT 141.420 162.365 141.645 162.495 ;
        RECT 141.420 161.260 141.590 162.365 ;
        RECT 141.815 162.215 142.340 162.435 ;
        RECT 141.760 161.450 142.000 162.045 ;
        RECT 142.170 161.515 142.340 162.215 ;
        RECT 142.510 161.855 142.680 162.635 ;
        RECT 143.000 162.585 143.370 163.085 ;
        RECT 143.550 162.635 143.955 162.805 ;
        RECT 144.125 162.635 144.910 162.805 ;
        RECT 143.550 162.405 143.720 162.635 ;
        RECT 142.890 162.105 143.720 162.405 ;
        RECT 144.105 162.135 144.570 162.465 ;
        RECT 142.890 162.075 143.090 162.105 ;
        RECT 143.210 161.855 143.380 161.925 ;
        RECT 142.510 161.685 143.380 161.855 ;
        RECT 142.870 161.595 143.380 161.685 ;
        RECT 141.420 161.130 141.725 161.260 ;
        RECT 142.170 161.150 142.700 161.515 ;
        RECT 141.040 160.535 141.305 160.995 ;
        RECT 141.475 160.705 141.725 161.130 ;
        RECT 142.870 160.980 143.040 161.595 ;
        RECT 141.935 160.810 143.040 160.980 ;
        RECT 143.210 160.535 143.380 161.335 ;
        RECT 143.550 161.035 143.720 162.105 ;
        RECT 143.890 161.205 144.080 161.925 ;
        RECT 144.250 161.175 144.570 162.135 ;
        RECT 144.740 162.175 144.910 162.635 ;
        RECT 145.185 162.555 145.395 163.085 ;
        RECT 145.655 162.345 145.985 162.870 ;
        RECT 146.155 162.475 146.325 163.085 ;
        RECT 146.495 162.430 146.825 162.865 ;
        RECT 146.495 162.345 146.875 162.430 ;
        RECT 145.785 162.175 145.985 162.345 ;
        RECT 146.650 162.305 146.875 162.345 ;
        RECT 144.740 161.845 145.615 162.175 ;
        RECT 145.785 161.845 146.535 162.175 ;
        RECT 143.550 160.705 143.800 161.035 ;
        RECT 144.740 161.005 144.910 161.845 ;
        RECT 145.785 161.640 145.975 161.845 ;
        RECT 146.705 161.725 146.875 162.305 ;
        RECT 147.045 162.315 148.715 163.085 ;
        RECT 148.885 162.335 150.095 163.085 ;
        RECT 147.045 161.795 147.795 162.315 ;
        RECT 146.660 161.675 146.875 161.725 ;
        RECT 145.080 161.265 145.975 161.640 ;
        RECT 146.485 161.595 146.875 161.675 ;
        RECT 147.965 161.625 148.715 162.145 ;
        RECT 144.025 160.835 144.910 161.005 ;
        RECT 145.090 160.535 145.405 161.035 ;
        RECT 145.635 160.705 145.975 161.265 ;
        RECT 146.145 160.535 146.315 161.545 ;
        RECT 146.485 160.750 146.815 161.595 ;
        RECT 147.045 160.535 148.715 161.625 ;
        RECT 148.885 161.625 149.405 162.165 ;
        RECT 149.575 161.795 150.095 162.335 ;
        RECT 148.885 160.535 150.095 161.625 ;
        RECT 36.100 160.365 150.180 160.535 ;
        RECT 36.185 159.275 37.395 160.365 ;
        RECT 37.565 159.275 41.075 160.365 ;
        RECT 36.185 158.565 36.705 159.105 ;
        RECT 36.875 158.735 37.395 159.275 ;
        RECT 37.565 158.585 39.215 159.105 ;
        RECT 39.385 158.755 41.075 159.275 ;
        RECT 42.175 159.415 42.450 160.185 ;
        RECT 42.620 159.755 42.950 160.185 ;
        RECT 43.120 159.925 43.315 160.365 ;
        RECT 43.495 159.755 43.825 160.185 ;
        RECT 42.620 159.585 43.825 159.755 ;
        RECT 45.125 159.695 45.405 160.365 ;
        RECT 42.175 159.225 42.760 159.415 ;
        RECT 42.930 159.255 43.825 159.585 ;
        RECT 45.575 159.475 45.875 160.025 ;
        RECT 46.075 159.645 46.405 160.365 ;
        RECT 46.595 159.645 47.055 160.195 ;
        RECT 36.185 157.815 37.395 158.565 ;
        RECT 37.565 157.815 41.075 158.585 ;
        RECT 42.175 158.405 42.415 159.055 ;
        RECT 42.585 158.555 42.760 159.225 ;
        RECT 44.940 159.055 45.205 159.415 ;
        RECT 45.575 159.305 46.515 159.475 ;
        RECT 46.345 159.055 46.515 159.305 ;
        RECT 42.930 158.725 43.345 159.055 ;
        RECT 43.525 158.725 43.820 159.055 ;
        RECT 44.940 158.805 45.615 159.055 ;
        RECT 45.835 158.805 46.175 159.055 ;
        RECT 46.345 158.725 46.635 159.055 ;
        RECT 42.585 158.375 42.915 158.555 ;
        RECT 42.190 157.815 42.520 158.205 ;
        RECT 42.690 157.995 42.915 158.375 ;
        RECT 43.115 158.105 43.345 158.725 ;
        RECT 46.345 158.635 46.515 158.725 ;
        RECT 43.525 157.815 43.825 158.545 ;
        RECT 45.125 158.445 46.515 158.635 ;
        RECT 45.125 158.085 45.455 158.445 ;
        RECT 46.805 158.275 47.055 159.645 ;
        RECT 47.225 159.275 48.895 160.365 ;
        RECT 46.075 157.815 46.325 158.275 ;
        RECT 46.495 157.985 47.055 158.275 ;
        RECT 47.225 158.585 47.975 159.105 ;
        RECT 48.145 158.755 48.895 159.275 ;
        RECT 49.065 159.200 49.355 160.365 ;
        RECT 49.525 159.275 53.035 160.365 ;
        RECT 49.525 158.585 51.175 159.105 ;
        RECT 51.345 158.755 53.035 159.275 ;
        RECT 53.665 159.515 54.045 160.195 ;
        RECT 54.635 159.515 54.805 160.365 ;
        RECT 54.975 159.685 55.305 160.195 ;
        RECT 55.475 159.855 55.645 160.365 ;
        RECT 55.815 159.685 56.215 160.195 ;
        RECT 54.975 159.515 56.215 159.685 ;
        RECT 47.225 157.815 48.895 158.585 ;
        RECT 49.065 157.815 49.355 158.540 ;
        RECT 49.525 157.815 53.035 158.585 ;
        RECT 53.665 158.555 53.835 159.515 ;
        RECT 54.005 159.175 55.310 159.345 ;
        RECT 56.395 159.265 56.715 160.195 ;
        RECT 56.885 159.275 58.095 160.365 ;
        RECT 54.005 158.725 54.250 159.175 ;
        RECT 54.420 158.805 54.970 159.005 ;
        RECT 55.140 158.975 55.310 159.175 ;
        RECT 56.085 159.095 56.715 159.265 ;
        RECT 55.140 158.805 55.515 158.975 ;
        RECT 55.685 158.555 55.915 159.055 ;
        RECT 53.665 158.385 55.915 158.555 ;
        RECT 53.715 157.815 54.045 158.205 ;
        RECT 54.215 158.065 54.385 158.385 ;
        RECT 56.085 158.215 56.255 159.095 ;
        RECT 54.555 157.815 54.885 158.205 ;
        RECT 55.300 158.045 56.255 158.215 ;
        RECT 56.425 157.815 56.715 158.650 ;
        RECT 56.885 158.565 57.405 159.105 ;
        RECT 57.575 158.735 58.095 159.275 ;
        RECT 58.285 159.475 58.545 160.185 ;
        RECT 58.715 159.655 59.045 160.365 ;
        RECT 59.215 159.475 59.445 160.185 ;
        RECT 58.285 159.235 59.445 159.475 ;
        RECT 59.625 159.455 59.895 160.185 ;
        RECT 60.075 159.635 60.415 160.365 ;
        RECT 59.625 159.235 60.395 159.455 ;
        RECT 58.275 158.725 58.575 159.055 ;
        RECT 58.755 158.745 59.280 159.055 ;
        RECT 59.460 158.745 59.925 159.055 ;
        RECT 56.885 157.815 58.095 158.565 ;
        RECT 58.285 157.815 58.575 158.545 ;
        RECT 58.755 158.105 58.985 158.745 ;
        RECT 60.105 158.565 60.395 159.235 ;
        RECT 59.165 158.365 60.395 158.565 ;
        RECT 59.165 157.995 59.475 158.365 ;
        RECT 59.655 157.815 60.325 158.185 ;
        RECT 60.585 157.995 60.845 160.185 ;
        RECT 61.025 159.930 66.370 160.365 ;
        RECT 62.610 158.360 62.950 159.190 ;
        RECT 64.430 158.680 64.780 159.930 ;
        RECT 66.545 159.275 70.055 160.365 ;
        RECT 70.225 159.275 71.435 160.365 ;
        RECT 71.805 159.695 72.085 160.365 ;
        RECT 72.255 159.475 72.555 160.025 ;
        RECT 72.755 159.645 73.085 160.365 ;
        RECT 73.275 159.645 73.735 160.195 ;
        RECT 66.545 158.585 68.195 159.105 ;
        RECT 68.365 158.755 70.055 159.275 ;
        RECT 61.025 157.815 66.370 158.360 ;
        RECT 66.545 157.815 70.055 158.585 ;
        RECT 70.225 158.565 70.745 159.105 ;
        RECT 70.915 158.735 71.435 159.275 ;
        RECT 71.620 159.055 71.885 159.415 ;
        RECT 72.255 159.305 73.195 159.475 ;
        RECT 73.025 159.055 73.195 159.305 ;
        RECT 71.620 158.805 72.295 159.055 ;
        RECT 72.515 158.805 72.855 159.055 ;
        RECT 73.025 158.725 73.315 159.055 ;
        RECT 73.025 158.635 73.195 158.725 ;
        RECT 70.225 157.815 71.435 158.565 ;
        RECT 71.805 158.445 73.195 158.635 ;
        RECT 71.805 158.085 72.135 158.445 ;
        RECT 73.485 158.275 73.735 159.645 ;
        RECT 74.825 159.200 75.115 160.365 ;
        RECT 75.295 159.395 75.625 160.180 ;
        RECT 75.295 159.225 75.975 159.395 ;
        RECT 76.155 159.225 76.485 160.365 ;
        RECT 76.665 159.275 78.335 160.365 ;
        RECT 78.540 159.865 78.820 160.195 ;
        RECT 78.990 159.865 79.240 160.365 ;
        RECT 79.410 160.025 80.500 160.195 ;
        RECT 79.410 159.865 79.660 160.025 ;
        RECT 80.250 159.865 80.500 160.025 ;
        RECT 78.565 159.855 78.735 159.865 ;
        RECT 79.485 159.855 79.655 159.865 ;
        RECT 80.705 159.855 81.020 160.195 ;
        RECT 81.190 159.865 81.440 160.365 ;
        RECT 79.830 159.685 80.080 159.855 ;
        RECT 80.810 159.685 81.020 159.855 ;
        RECT 81.610 159.685 81.860 160.195 ;
        RECT 82.030 159.865 82.335 160.365 ;
        RECT 82.505 160.025 84.115 160.195 ;
        RECT 82.505 159.685 83.275 160.025 ;
        RECT 75.285 158.805 75.635 159.055 ;
        RECT 75.805 158.625 75.975 159.225 ;
        RECT 76.145 158.805 76.495 159.055 ;
        RECT 72.755 157.815 73.005 158.275 ;
        RECT 73.175 157.985 73.735 158.275 ;
        RECT 74.825 157.815 75.115 158.540 ;
        RECT 75.305 157.815 75.545 158.625 ;
        RECT 75.715 157.985 76.045 158.625 ;
        RECT 76.215 157.815 76.485 158.625 ;
        RECT 76.665 158.585 77.415 159.105 ;
        RECT 77.585 158.755 78.335 159.275 ;
        RECT 78.540 159.515 80.640 159.685 ;
        RECT 80.810 159.515 83.275 159.685 ;
        RECT 78.540 158.635 78.710 159.515 ;
        RECT 80.470 159.345 80.640 159.515 ;
        RECT 83.445 159.355 83.695 159.855 ;
        RECT 83.865 159.525 84.115 160.025 ;
        RECT 84.485 159.930 89.830 160.365 ;
        RECT 90.005 159.930 95.350 160.365 ;
        RECT 79.125 159.175 80.300 159.345 ;
        RECT 80.470 159.175 83.205 159.345 ;
        RECT 79.125 159.005 79.295 159.175 ;
        RECT 80.130 159.005 80.300 159.175 ;
        RECT 78.965 158.805 79.295 159.005 ;
        RECT 79.465 158.805 79.960 159.005 ;
        RECT 80.130 158.805 81.650 159.005 ;
        RECT 81.840 158.805 82.510 159.005 ;
        RECT 83.035 158.975 83.205 159.175 ;
        RECT 83.445 159.145 84.315 159.355 ;
        RECT 83.035 158.805 83.695 158.975 ;
        RECT 83.905 158.635 84.315 159.145 ;
        RECT 76.665 157.815 78.335 158.585 ;
        RECT 78.540 158.455 80.120 158.635 ;
        RECT 78.610 157.815 78.780 158.285 ;
        RECT 78.950 157.985 79.280 158.455 ;
        RECT 79.450 157.815 79.620 158.285 ;
        RECT 79.790 157.985 80.120 158.455 ;
        RECT 80.730 158.455 81.820 158.635 ;
        RECT 80.290 157.815 80.460 158.285 ;
        RECT 80.730 157.985 81.060 158.455 ;
        RECT 81.230 157.815 81.400 158.285 ;
        RECT 81.570 158.205 81.820 158.455 ;
        RECT 82.045 158.455 84.315 158.635 ;
        RECT 82.045 158.375 82.375 158.455 ;
        RECT 83.405 158.375 83.735 158.455 ;
        RECT 86.070 158.360 86.410 159.190 ;
        RECT 87.890 158.680 88.240 159.930 ;
        RECT 91.590 158.360 91.930 159.190 ;
        RECT 93.410 158.680 93.760 159.930 ;
        RECT 95.525 159.275 96.735 160.365 ;
        RECT 95.525 158.565 96.045 159.105 ;
        RECT 96.215 158.735 96.735 159.275 ;
        RECT 97.110 159.395 97.440 160.195 ;
        RECT 97.610 159.565 97.940 160.365 ;
        RECT 98.240 159.395 98.570 160.195 ;
        RECT 99.215 159.565 99.465 160.365 ;
        RECT 97.110 159.225 99.545 159.395 ;
        RECT 99.735 159.225 99.905 160.365 ;
        RECT 100.075 159.225 100.415 160.195 ;
        RECT 96.905 158.805 97.255 159.055 ;
        RECT 97.440 158.595 97.610 159.225 ;
        RECT 97.780 158.805 98.110 159.005 ;
        RECT 98.280 158.805 98.610 159.005 ;
        RECT 98.780 158.805 99.200 159.005 ;
        RECT 99.375 158.975 99.545 159.225 ;
        RECT 100.185 159.175 100.415 159.225 ;
        RECT 100.585 159.200 100.875 160.365 ;
        RECT 101.200 159.355 101.500 160.195 ;
        RECT 101.695 159.525 101.945 160.365 ;
        RECT 102.535 159.775 103.340 160.195 ;
        RECT 102.115 159.605 103.680 159.775 ;
        RECT 102.115 159.355 102.285 159.605 ;
        RECT 101.200 159.185 102.285 159.355 ;
        RECT 99.375 158.805 100.070 158.975 ;
        RECT 81.570 157.985 82.800 158.205 ;
        RECT 83.065 157.815 83.235 158.285 ;
        RECT 83.905 157.815 84.075 158.285 ;
        RECT 84.485 157.815 89.830 158.360 ;
        RECT 90.005 157.815 95.350 158.360 ;
        RECT 95.525 157.815 96.735 158.565 ;
        RECT 97.110 157.985 97.610 158.595 ;
        RECT 98.240 158.465 99.465 158.635 ;
        RECT 100.240 158.615 100.415 159.175 ;
        RECT 101.045 158.725 101.375 159.015 ;
        RECT 98.240 157.985 98.570 158.465 ;
        RECT 98.740 157.815 98.965 158.275 ;
        RECT 99.135 157.985 99.465 158.465 ;
        RECT 99.655 157.815 99.905 158.615 ;
        RECT 100.075 157.985 100.415 158.615 ;
        RECT 101.545 158.555 101.715 159.185 ;
        RECT 102.455 159.055 102.775 159.435 ;
        RECT 102.965 159.345 103.340 159.435 ;
        RECT 102.945 159.175 103.340 159.345 ;
        RECT 103.510 159.355 103.680 159.605 ;
        RECT 103.850 159.525 104.180 160.365 ;
        RECT 104.350 159.605 105.015 160.195 ;
        RECT 105.195 159.645 105.525 160.365 ;
        RECT 103.510 159.185 104.430 159.355 ;
        RECT 101.885 158.805 102.215 159.015 ;
        RECT 102.395 158.805 102.775 159.055 ;
        RECT 102.965 159.015 103.340 159.175 ;
        RECT 104.260 159.015 104.430 159.185 ;
        RECT 102.965 158.805 103.450 159.015 ;
        RECT 103.640 158.805 104.090 159.015 ;
        RECT 104.260 158.805 104.595 159.015 ;
        RECT 104.765 158.635 105.015 159.605 ;
        RECT 105.185 159.005 105.415 159.345 ;
        RECT 105.705 159.005 105.920 160.120 ;
        RECT 106.115 159.420 106.445 160.195 ;
        RECT 106.615 159.590 107.325 160.365 ;
        RECT 106.115 159.205 107.265 159.420 ;
        RECT 105.185 158.805 105.515 159.005 ;
        RECT 105.705 158.825 106.155 159.005 ;
        RECT 105.825 158.805 106.155 158.825 ;
        RECT 106.325 158.805 106.795 159.035 ;
        RECT 106.980 158.635 107.265 159.205 ;
        RECT 107.495 158.760 107.775 160.195 ;
        RECT 107.945 159.275 109.155 160.365 ;
        RECT 100.585 157.815 100.875 158.540 ;
        RECT 101.205 158.375 101.715 158.555 ;
        RECT 102.120 158.465 103.820 158.635 ;
        RECT 102.120 158.375 102.505 158.465 ;
        RECT 101.205 157.985 101.535 158.375 ;
        RECT 101.705 158.035 102.890 158.205 ;
        RECT 103.150 157.815 103.320 158.285 ;
        RECT 103.490 158.000 103.820 158.465 ;
        RECT 103.990 157.815 104.160 158.635 ;
        RECT 104.330 157.995 105.015 158.635 ;
        RECT 105.185 158.445 106.365 158.635 ;
        RECT 105.185 157.985 105.525 158.445 ;
        RECT 106.035 158.365 106.365 158.445 ;
        RECT 106.555 158.445 107.265 158.635 ;
        RECT 106.555 158.305 106.855 158.445 ;
        RECT 106.540 158.295 106.855 158.305 ;
        RECT 106.530 158.285 106.855 158.295 ;
        RECT 106.520 158.280 106.855 158.285 ;
        RECT 105.695 157.815 105.865 158.275 ;
        RECT 106.515 158.270 106.855 158.280 ;
        RECT 106.510 158.265 106.855 158.270 ;
        RECT 106.505 158.255 106.855 158.265 ;
        RECT 106.500 158.250 106.855 158.255 ;
        RECT 106.495 157.985 106.855 158.250 ;
        RECT 107.095 157.815 107.265 158.275 ;
        RECT 107.435 157.985 107.775 158.760 ;
        RECT 107.945 158.565 108.465 159.105 ;
        RECT 108.635 158.735 109.155 159.275 ;
        RECT 109.325 159.605 109.990 160.195 ;
        RECT 109.325 158.635 109.575 159.605 ;
        RECT 110.160 159.525 110.490 160.365 ;
        RECT 111.000 159.775 111.805 160.195 ;
        RECT 110.660 159.605 112.225 159.775 ;
        RECT 110.660 159.355 110.830 159.605 ;
        RECT 109.910 159.185 110.830 159.355 ;
        RECT 109.910 159.015 110.080 159.185 ;
        RECT 111.000 159.015 111.375 159.435 ;
        RECT 109.745 158.805 110.080 159.015 ;
        RECT 110.250 158.805 110.700 159.015 ;
        RECT 110.890 159.005 111.375 159.015 ;
        RECT 111.565 159.055 111.885 159.435 ;
        RECT 112.055 159.355 112.225 159.605 ;
        RECT 112.395 159.525 112.645 160.365 ;
        RECT 112.840 159.355 113.140 160.195 ;
        RECT 113.475 159.645 113.805 160.365 ;
        RECT 112.055 159.185 113.140 159.355 ;
        RECT 110.890 158.835 111.395 159.005 ;
        RECT 110.890 158.805 111.375 158.835 ;
        RECT 111.565 158.805 111.945 159.055 ;
        RECT 112.125 158.805 112.455 159.015 ;
        RECT 107.945 157.815 109.155 158.565 ;
        RECT 109.325 157.995 110.010 158.635 ;
        RECT 110.180 157.815 110.350 158.635 ;
        RECT 110.520 158.465 112.220 158.635 ;
        RECT 110.520 158.000 110.850 158.465 ;
        RECT 111.835 158.375 112.220 158.465 ;
        RECT 112.625 158.555 112.795 159.185 ;
        RECT 112.965 158.725 113.295 159.015 ;
        RECT 113.465 159.005 113.695 159.345 ;
        RECT 113.985 159.005 114.200 160.120 ;
        RECT 114.395 159.420 114.725 160.195 ;
        RECT 114.895 159.590 115.605 160.365 ;
        RECT 114.395 159.205 115.545 159.420 ;
        RECT 113.465 158.805 113.795 159.005 ;
        RECT 113.985 158.825 114.435 159.005 ;
        RECT 114.105 158.805 114.435 158.825 ;
        RECT 114.605 158.805 115.075 159.035 ;
        RECT 115.260 158.635 115.545 159.205 ;
        RECT 115.775 158.760 116.055 160.195 ;
        RECT 116.225 159.930 121.570 160.365 ;
        RECT 112.625 158.375 113.135 158.555 ;
        RECT 111.020 157.815 111.190 158.285 ;
        RECT 111.450 158.035 112.635 158.205 ;
        RECT 112.805 157.985 113.135 158.375 ;
        RECT 113.465 158.445 114.645 158.635 ;
        RECT 113.465 157.985 113.805 158.445 ;
        RECT 114.315 158.365 114.645 158.445 ;
        RECT 114.835 158.445 115.545 158.635 ;
        RECT 114.835 158.305 115.135 158.445 ;
        RECT 114.820 158.295 115.135 158.305 ;
        RECT 114.810 158.285 115.135 158.295 ;
        RECT 114.800 158.280 115.135 158.285 ;
        RECT 113.975 157.815 114.145 158.275 ;
        RECT 114.795 158.270 115.135 158.280 ;
        RECT 114.790 158.265 115.135 158.270 ;
        RECT 114.785 158.255 115.135 158.265 ;
        RECT 114.780 158.250 115.135 158.255 ;
        RECT 114.775 157.985 115.135 158.250 ;
        RECT 115.375 157.815 115.545 158.275 ;
        RECT 115.715 157.985 116.055 158.760 ;
        RECT 117.810 158.360 118.150 159.190 ;
        RECT 119.630 158.680 119.980 159.930 ;
        RECT 121.745 159.275 124.335 160.365 ;
        RECT 121.745 158.585 122.955 159.105 ;
        RECT 123.125 158.755 124.335 159.275 ;
        RECT 124.965 159.290 125.235 160.195 ;
        RECT 125.405 159.605 125.735 160.365 ;
        RECT 125.915 159.435 126.095 160.195 ;
        RECT 116.225 157.815 121.570 158.360 ;
        RECT 121.745 157.815 124.335 158.585 ;
        RECT 124.965 158.490 125.145 159.290 ;
        RECT 125.420 159.265 126.095 159.435 ;
        RECT 125.420 159.120 125.590 159.265 ;
        RECT 126.345 159.200 126.635 160.365 ;
        RECT 126.805 159.770 127.240 160.195 ;
        RECT 127.410 159.940 127.795 160.365 ;
        RECT 126.805 159.600 127.795 159.770 ;
        RECT 125.315 158.790 125.590 159.120 ;
        RECT 125.420 158.535 125.590 158.790 ;
        RECT 125.815 158.715 126.155 159.085 ;
        RECT 126.805 158.725 127.290 159.430 ;
        RECT 127.460 159.055 127.795 159.600 ;
        RECT 127.965 159.405 128.390 160.195 ;
        RECT 128.560 159.770 128.835 160.195 ;
        RECT 129.005 159.940 129.390 160.365 ;
        RECT 128.560 159.575 129.390 159.770 ;
        RECT 127.965 159.225 128.870 159.405 ;
        RECT 127.460 158.725 127.870 159.055 ;
        RECT 128.040 158.725 128.870 159.225 ;
        RECT 129.040 159.055 129.390 159.575 ;
        RECT 129.560 159.405 129.805 160.195 ;
        RECT 129.995 159.770 130.250 160.195 ;
        RECT 130.420 159.940 130.805 160.365 ;
        RECT 129.995 159.575 130.805 159.770 ;
        RECT 129.560 159.225 130.285 159.405 ;
        RECT 129.040 158.725 129.465 159.055 ;
        RECT 129.635 158.725 130.285 159.225 ;
        RECT 130.455 159.055 130.805 159.575 ;
        RECT 130.975 159.225 131.235 160.195 ;
        RECT 131.405 159.275 132.615 160.365 ;
        RECT 130.455 158.725 130.880 159.055 ;
        RECT 127.460 158.555 127.795 158.725 ;
        RECT 128.040 158.555 128.390 158.725 ;
        RECT 129.040 158.555 129.390 158.725 ;
        RECT 129.635 158.555 129.805 158.725 ;
        RECT 130.455 158.555 130.805 158.725 ;
        RECT 131.050 158.555 131.235 159.225 ;
        RECT 124.965 157.985 125.225 158.490 ;
        RECT 125.420 158.365 126.085 158.535 ;
        RECT 125.405 157.815 125.735 158.195 ;
        RECT 125.915 157.985 126.085 158.365 ;
        RECT 126.345 157.815 126.635 158.540 ;
        RECT 126.805 158.385 127.795 158.555 ;
        RECT 126.805 157.985 127.240 158.385 ;
        RECT 127.410 157.815 127.795 158.215 ;
        RECT 127.965 157.985 128.390 158.555 ;
        RECT 128.580 158.385 129.390 158.555 ;
        RECT 128.580 157.985 128.835 158.385 ;
        RECT 129.005 157.815 129.390 158.215 ;
        RECT 129.560 157.985 129.805 158.555 ;
        RECT 129.995 158.385 130.805 158.555 ;
        RECT 129.995 157.985 130.250 158.385 ;
        RECT 130.420 157.815 130.805 158.215 ;
        RECT 130.975 157.985 131.235 158.555 ;
        RECT 131.405 158.565 131.925 159.105 ;
        RECT 132.095 158.735 132.615 159.275 ;
        RECT 132.990 159.395 133.320 160.195 ;
        RECT 133.490 159.565 133.820 160.365 ;
        RECT 134.120 159.395 134.450 160.195 ;
        RECT 135.095 159.565 135.345 160.365 ;
        RECT 132.990 159.225 135.425 159.395 ;
        RECT 135.615 159.225 135.785 160.365 ;
        RECT 135.955 159.225 136.295 160.195 ;
        RECT 136.670 159.395 137.000 160.195 ;
        RECT 137.170 159.565 137.500 160.365 ;
        RECT 137.800 159.395 138.130 160.195 ;
        RECT 138.775 159.565 139.025 160.365 ;
        RECT 136.670 159.225 139.105 159.395 ;
        RECT 139.295 159.225 139.465 160.365 ;
        RECT 139.635 159.225 139.975 160.195 ;
        RECT 132.785 158.805 133.135 159.055 ;
        RECT 133.320 158.595 133.490 159.225 ;
        RECT 133.660 158.805 133.990 159.005 ;
        RECT 134.160 158.805 134.490 159.005 ;
        RECT 134.660 158.805 135.080 159.005 ;
        RECT 135.255 158.975 135.425 159.225 ;
        RECT 135.255 158.805 135.950 158.975 ;
        RECT 136.120 158.665 136.295 159.225 ;
        RECT 136.465 158.805 136.815 159.055 ;
        RECT 131.405 157.815 132.615 158.565 ;
        RECT 132.990 157.985 133.490 158.595 ;
        RECT 134.120 158.465 135.345 158.635 ;
        RECT 136.065 158.615 136.295 158.665 ;
        RECT 134.120 157.985 134.450 158.465 ;
        RECT 134.620 157.815 134.845 158.275 ;
        RECT 135.015 157.985 135.345 158.465 ;
        RECT 135.535 157.815 135.785 158.615 ;
        RECT 135.955 157.985 136.295 158.615 ;
        RECT 137.000 158.595 137.170 159.225 ;
        RECT 137.340 158.805 137.670 159.005 ;
        RECT 137.840 158.805 138.170 159.005 ;
        RECT 138.340 158.805 138.760 159.005 ;
        RECT 138.935 158.975 139.105 159.225 ;
        RECT 138.935 158.805 139.630 158.975 ;
        RECT 136.670 157.985 137.170 158.595 ;
        RECT 137.800 158.465 139.025 158.635 ;
        RECT 139.800 158.615 139.975 159.225 ;
        RECT 137.800 157.985 138.130 158.465 ;
        RECT 138.300 157.815 138.525 158.275 ;
        RECT 138.695 157.985 139.025 158.465 ;
        RECT 139.215 157.815 139.465 158.615 ;
        RECT 139.635 157.985 139.975 158.615 ;
        RECT 140.145 159.290 140.415 160.195 ;
        RECT 140.585 159.605 140.915 160.365 ;
        RECT 141.095 159.435 141.275 160.195 ;
        RECT 140.145 158.490 140.325 159.290 ;
        RECT 140.600 159.265 141.275 159.435 ;
        RECT 141.525 159.290 141.795 160.195 ;
        RECT 141.965 159.605 142.295 160.365 ;
        RECT 142.475 159.435 142.655 160.195 ;
        RECT 142.910 159.940 143.245 160.365 ;
        RECT 143.415 159.760 143.600 160.165 ;
        RECT 140.600 159.120 140.770 159.265 ;
        RECT 140.495 158.790 140.770 159.120 ;
        RECT 140.600 158.535 140.770 158.790 ;
        RECT 140.995 158.715 141.335 159.085 ;
        RECT 140.145 157.985 140.405 158.490 ;
        RECT 140.600 158.365 141.265 158.535 ;
        RECT 140.585 157.815 140.915 158.195 ;
        RECT 141.095 157.985 141.265 158.365 ;
        RECT 141.525 158.490 141.705 159.290 ;
        RECT 141.980 159.265 142.655 159.435 ;
        RECT 142.935 159.585 143.600 159.760 ;
        RECT 143.805 159.585 144.135 160.365 ;
        RECT 141.980 159.120 142.150 159.265 ;
        RECT 141.875 158.790 142.150 159.120 ;
        RECT 141.980 158.535 142.150 158.790 ;
        RECT 142.375 158.715 142.715 159.085 ;
        RECT 142.935 158.555 143.275 159.585 ;
        RECT 144.305 159.395 144.575 160.165 ;
        RECT 143.445 159.225 144.575 159.395 ;
        RECT 143.445 158.725 143.695 159.225 ;
        RECT 141.525 157.985 141.785 158.490 ;
        RECT 141.980 158.365 142.645 158.535 ;
        RECT 142.935 158.385 143.620 158.555 ;
        RECT 143.875 158.475 144.235 159.055 ;
        RECT 141.965 157.815 142.295 158.195 ;
        RECT 142.475 157.985 142.645 158.365 ;
        RECT 142.910 157.815 143.245 158.215 ;
        RECT 143.415 157.985 143.620 158.385 ;
        RECT 144.405 158.315 144.575 159.225 ;
        RECT 143.830 157.815 144.105 158.295 ;
        RECT 144.315 157.985 144.575 158.315 ;
        RECT 144.745 159.290 145.015 160.195 ;
        RECT 145.185 159.605 145.515 160.365 ;
        RECT 145.695 159.435 145.875 160.195 ;
        RECT 144.745 158.490 144.925 159.290 ;
        RECT 145.200 159.265 145.875 159.435 ;
        RECT 146.125 159.290 146.395 160.195 ;
        RECT 146.565 159.605 146.895 160.365 ;
        RECT 147.075 159.435 147.255 160.195 ;
        RECT 145.200 159.120 145.370 159.265 ;
        RECT 145.095 158.790 145.370 159.120 ;
        RECT 145.200 158.535 145.370 158.790 ;
        RECT 145.595 158.715 145.935 159.085 ;
        RECT 144.745 157.985 145.005 158.490 ;
        RECT 145.200 158.365 145.865 158.535 ;
        RECT 145.185 157.815 145.515 158.195 ;
        RECT 145.695 157.985 145.865 158.365 ;
        RECT 146.125 158.490 146.305 159.290 ;
        RECT 146.580 159.265 147.255 159.435 ;
        RECT 147.505 159.275 148.715 160.365 ;
        RECT 146.580 159.120 146.750 159.265 ;
        RECT 146.475 158.790 146.750 159.120 ;
        RECT 146.580 158.535 146.750 158.790 ;
        RECT 146.975 158.715 147.315 159.085 ;
        RECT 147.505 158.565 148.025 159.105 ;
        RECT 148.195 158.735 148.715 159.275 ;
        RECT 148.885 159.275 150.095 160.365 ;
        RECT 148.885 158.735 149.405 159.275 ;
        RECT 149.575 158.565 150.095 159.105 ;
        RECT 146.125 157.985 146.385 158.490 ;
        RECT 146.580 158.365 147.245 158.535 ;
        RECT 146.565 157.815 146.895 158.195 ;
        RECT 147.075 157.985 147.245 158.365 ;
        RECT 147.505 157.815 148.715 158.565 ;
        RECT 148.885 157.815 150.095 158.565 ;
        RECT 36.100 157.645 150.180 157.815 ;
        RECT 36.185 156.895 37.395 157.645 ;
        RECT 38.115 157.095 38.285 157.385 ;
        RECT 38.455 157.265 38.785 157.645 ;
        RECT 38.115 156.925 38.780 157.095 ;
        RECT 36.185 156.355 36.705 156.895 ;
        RECT 36.875 156.185 37.395 156.725 ;
        RECT 36.185 155.095 37.395 156.185 ;
        RECT 38.030 156.105 38.380 156.755 ;
        RECT 38.550 155.935 38.780 156.925 ;
        RECT 38.115 155.765 38.780 155.935 ;
        RECT 38.115 155.265 38.285 155.765 ;
        RECT 38.455 155.095 38.785 155.595 ;
        RECT 38.955 155.265 39.140 157.385 ;
        RECT 39.395 157.185 39.645 157.645 ;
        RECT 39.815 157.195 40.150 157.365 ;
        RECT 40.345 157.195 41.020 157.365 ;
        RECT 39.815 157.055 39.985 157.195 ;
        RECT 39.310 156.065 39.590 157.015 ;
        RECT 39.760 156.925 39.985 157.055 ;
        RECT 39.760 155.820 39.930 156.925 ;
        RECT 40.155 156.775 40.680 156.995 ;
        RECT 40.100 156.010 40.340 156.605 ;
        RECT 40.510 156.075 40.680 156.775 ;
        RECT 40.850 156.415 41.020 157.195 ;
        RECT 41.340 157.145 41.710 157.645 ;
        RECT 41.890 157.195 42.295 157.365 ;
        RECT 42.465 157.195 43.250 157.365 ;
        RECT 41.890 156.965 42.060 157.195 ;
        RECT 41.230 156.665 42.060 156.965 ;
        RECT 42.445 156.695 42.910 157.025 ;
        RECT 41.230 156.635 41.430 156.665 ;
        RECT 41.550 156.415 41.720 156.485 ;
        RECT 40.850 156.245 41.720 156.415 ;
        RECT 41.210 156.155 41.720 156.245 ;
        RECT 39.760 155.690 40.065 155.820 ;
        RECT 40.510 155.710 41.040 156.075 ;
        RECT 39.380 155.095 39.645 155.555 ;
        RECT 39.815 155.265 40.065 155.690 ;
        RECT 41.210 155.540 41.380 156.155 ;
        RECT 40.275 155.370 41.380 155.540 ;
        RECT 41.550 155.095 41.720 155.895 ;
        RECT 41.890 155.595 42.060 156.665 ;
        RECT 42.230 155.765 42.420 156.485 ;
        RECT 42.590 155.735 42.910 156.695 ;
        RECT 43.080 156.735 43.250 157.195 ;
        RECT 43.525 157.115 43.735 157.645 ;
        RECT 43.995 156.905 44.325 157.430 ;
        RECT 44.495 157.035 44.665 157.645 ;
        RECT 44.835 156.990 45.165 157.425 ;
        RECT 44.835 156.905 45.215 156.990 ;
        RECT 44.125 156.735 44.325 156.905 ;
        RECT 44.990 156.865 45.215 156.905 ;
        RECT 43.080 156.405 43.955 156.735 ;
        RECT 44.125 156.405 44.875 156.735 ;
        RECT 41.890 155.265 42.140 155.595 ;
        RECT 43.080 155.565 43.250 156.405 ;
        RECT 44.125 156.200 44.315 156.405 ;
        RECT 45.045 156.285 45.215 156.865 ;
        RECT 45.385 156.895 46.595 157.645 ;
        RECT 46.765 157.145 47.025 157.475 ;
        RECT 47.235 157.165 47.510 157.645 ;
        RECT 45.385 156.355 45.905 156.895 ;
        RECT 45.000 156.235 45.215 156.285 ;
        RECT 43.420 155.825 44.315 156.200 ;
        RECT 44.825 156.155 45.215 156.235 ;
        RECT 46.075 156.185 46.595 156.725 ;
        RECT 42.365 155.395 43.250 155.565 ;
        RECT 43.430 155.095 43.745 155.595 ;
        RECT 43.975 155.265 44.315 155.825 ;
        RECT 44.485 155.095 44.655 156.105 ;
        RECT 44.825 155.310 45.155 156.155 ;
        RECT 45.385 155.095 46.595 156.185 ;
        RECT 46.765 156.235 46.935 157.145 ;
        RECT 47.720 157.075 47.925 157.475 ;
        RECT 48.095 157.245 48.430 157.645 ;
        RECT 47.105 156.405 47.465 156.985 ;
        RECT 47.720 156.905 48.405 157.075 ;
        RECT 47.645 156.235 47.895 156.735 ;
        RECT 46.765 156.065 47.895 156.235 ;
        RECT 46.765 155.295 47.035 156.065 ;
        RECT 48.065 155.875 48.405 156.905 ;
        RECT 48.605 156.875 51.195 157.645 ;
        RECT 51.415 156.990 51.745 157.425 ;
        RECT 51.915 157.035 52.085 157.645 ;
        RECT 51.365 156.905 51.745 156.990 ;
        RECT 52.255 156.905 52.585 157.430 ;
        RECT 52.845 157.115 53.055 157.645 ;
        RECT 53.330 157.195 54.115 157.365 ;
        RECT 54.285 157.195 54.690 157.365 ;
        RECT 48.605 156.355 49.815 156.875 ;
        RECT 51.365 156.865 51.590 156.905 ;
        RECT 49.985 156.185 51.195 156.705 ;
        RECT 47.205 155.095 47.535 155.875 ;
        RECT 47.740 155.700 48.405 155.875 ;
        RECT 47.740 155.295 47.925 155.700 ;
        RECT 48.095 155.095 48.430 155.520 ;
        RECT 48.605 155.095 51.195 156.185 ;
        RECT 51.365 156.285 51.535 156.865 ;
        RECT 52.255 156.735 52.455 156.905 ;
        RECT 53.330 156.735 53.500 157.195 ;
        RECT 51.705 156.405 52.455 156.735 ;
        RECT 52.625 156.405 53.500 156.735 ;
        RECT 51.365 156.235 51.580 156.285 ;
        RECT 51.365 156.155 51.755 156.235 ;
        RECT 51.425 155.310 51.755 156.155 ;
        RECT 52.265 156.200 52.455 156.405 ;
        RECT 51.925 155.095 52.095 156.105 ;
        RECT 52.265 155.825 53.160 156.200 ;
        RECT 52.265 155.265 52.605 155.825 ;
        RECT 52.835 155.095 53.150 155.595 ;
        RECT 53.330 155.565 53.500 156.405 ;
        RECT 53.670 156.695 54.135 157.025 ;
        RECT 54.520 156.965 54.690 157.195 ;
        RECT 54.870 157.145 55.240 157.645 ;
        RECT 55.560 157.195 56.235 157.365 ;
        RECT 56.430 157.195 56.765 157.365 ;
        RECT 53.670 155.735 53.990 156.695 ;
        RECT 54.520 156.665 55.350 156.965 ;
        RECT 54.160 155.765 54.350 156.485 ;
        RECT 54.520 155.595 54.690 156.665 ;
        RECT 55.150 156.635 55.350 156.665 ;
        RECT 54.860 156.415 55.030 156.485 ;
        RECT 55.560 156.415 55.730 157.195 ;
        RECT 56.595 157.055 56.765 157.195 ;
        RECT 56.935 157.185 57.185 157.645 ;
        RECT 54.860 156.245 55.730 156.415 ;
        RECT 55.900 156.775 56.425 156.995 ;
        RECT 56.595 156.925 56.820 157.055 ;
        RECT 54.860 156.155 55.370 156.245 ;
        RECT 53.330 155.395 54.215 155.565 ;
        RECT 54.440 155.265 54.690 155.595 ;
        RECT 54.860 155.095 55.030 155.895 ;
        RECT 55.200 155.540 55.370 156.155 ;
        RECT 55.900 156.075 56.070 156.775 ;
        RECT 55.540 155.710 56.070 156.075 ;
        RECT 56.240 156.010 56.480 156.605 ;
        RECT 56.650 155.820 56.820 156.925 ;
        RECT 56.990 156.065 57.270 157.015 ;
        RECT 56.515 155.690 56.820 155.820 ;
        RECT 55.200 155.370 56.305 155.540 ;
        RECT 56.515 155.265 56.765 155.690 ;
        RECT 56.935 155.095 57.200 155.555 ;
        RECT 57.440 155.265 57.625 157.385 ;
        RECT 57.795 157.265 58.125 157.645 ;
        RECT 58.295 157.095 58.465 157.385 ;
        RECT 57.800 156.925 58.465 157.095 ;
        RECT 57.800 155.935 58.030 156.925 ;
        RECT 58.725 156.905 59.045 157.385 ;
        RECT 59.215 157.075 59.445 157.475 ;
        RECT 59.615 157.255 59.965 157.645 ;
        RECT 59.215 156.995 59.725 157.075 ;
        RECT 60.135 156.995 60.465 157.475 ;
        RECT 59.215 156.905 60.465 156.995 ;
        RECT 58.200 156.105 58.550 156.755 ;
        RECT 58.725 155.975 58.895 156.905 ;
        RECT 59.555 156.825 60.465 156.905 ;
        RECT 60.635 156.825 60.805 157.645 ;
        RECT 61.310 156.905 61.775 157.450 ;
        RECT 61.945 156.920 62.235 157.645 ;
        RECT 63.605 157.015 63.985 157.465 ;
        RECT 59.065 156.315 59.235 156.735 ;
        RECT 59.465 156.485 60.065 156.655 ;
        RECT 59.065 156.145 59.725 156.315 ;
        RECT 57.800 155.765 58.465 155.935 ;
        RECT 58.725 155.775 59.385 155.975 ;
        RECT 59.555 155.945 59.725 156.145 ;
        RECT 59.895 156.285 60.065 156.485 ;
        RECT 60.235 156.455 60.930 156.655 ;
        RECT 61.190 156.285 61.435 156.735 ;
        RECT 59.895 156.115 61.435 156.285 ;
        RECT 61.605 155.945 61.775 156.905 ;
        RECT 59.555 155.775 61.775 155.945 ;
        RECT 57.795 155.095 58.125 155.595 ;
        RECT 58.295 155.265 58.465 155.765 ;
        RECT 59.215 155.605 59.385 155.775 ;
        RECT 58.745 155.095 59.045 155.605 ;
        RECT 59.215 155.435 59.595 155.605 ;
        RECT 60.175 155.095 60.805 155.605 ;
        RECT 60.975 155.265 61.305 155.775 ;
        RECT 61.475 155.095 61.775 155.605 ;
        RECT 61.945 155.095 62.235 156.260 ;
        RECT 63.345 156.065 63.575 156.755 ;
        RECT 63.755 156.565 63.985 157.015 ;
        RECT 64.165 156.865 64.395 157.645 ;
        RECT 64.575 156.935 65.005 157.465 ;
        RECT 64.575 156.685 64.820 156.935 ;
        RECT 65.185 156.735 65.395 157.355 ;
        RECT 65.565 156.915 65.895 157.645 ;
        RECT 63.755 155.885 64.095 156.565 ;
        RECT 63.335 155.685 64.095 155.885 ;
        RECT 64.285 156.385 64.820 156.685 ;
        RECT 65.000 156.385 65.395 156.735 ;
        RECT 65.590 156.385 65.880 156.735 ;
        RECT 66.085 156.700 66.425 157.475 ;
        RECT 66.595 157.185 66.765 157.645 ;
        RECT 67.005 157.210 67.365 157.475 ;
        RECT 67.005 157.205 67.360 157.210 ;
        RECT 67.005 157.195 67.355 157.205 ;
        RECT 67.005 157.190 67.350 157.195 ;
        RECT 67.005 157.180 67.345 157.190 ;
        RECT 67.995 157.185 68.165 157.645 ;
        RECT 67.005 157.175 67.340 157.180 ;
        RECT 67.005 157.165 67.330 157.175 ;
        RECT 67.005 157.155 67.320 157.165 ;
        RECT 67.005 157.015 67.305 157.155 ;
        RECT 66.595 156.825 67.305 157.015 ;
        RECT 67.495 157.015 67.825 157.095 ;
        RECT 68.335 157.015 68.675 157.475 ;
        RECT 67.495 156.825 68.675 157.015 ;
        RECT 68.845 156.875 71.435 157.645 ;
        RECT 71.695 157.095 71.865 157.475 ;
        RECT 72.045 157.265 72.375 157.645 ;
        RECT 71.695 156.925 72.360 157.095 ;
        RECT 72.555 156.970 72.815 157.475 ;
        RECT 63.335 155.295 63.595 155.685 ;
        RECT 63.765 155.095 64.095 155.505 ;
        RECT 64.285 155.275 64.615 156.385 ;
        RECT 64.785 156.005 65.825 156.205 ;
        RECT 64.785 155.275 64.975 156.005 ;
        RECT 65.145 155.095 65.475 155.825 ;
        RECT 65.655 155.275 65.825 156.005 ;
        RECT 66.085 155.265 66.365 156.700 ;
        RECT 66.595 156.255 66.880 156.825 ;
        RECT 67.065 156.425 67.535 156.655 ;
        RECT 67.705 156.635 68.035 156.655 ;
        RECT 67.705 156.455 68.155 156.635 ;
        RECT 68.345 156.455 68.675 156.655 ;
        RECT 66.595 156.040 67.745 156.255 ;
        RECT 66.535 155.095 67.245 155.870 ;
        RECT 67.415 155.265 67.745 156.040 ;
        RECT 67.940 155.340 68.155 156.455 ;
        RECT 68.445 156.115 68.675 156.455 ;
        RECT 68.845 156.355 70.055 156.875 ;
        RECT 70.225 156.185 71.435 156.705 ;
        RECT 71.625 156.375 71.965 156.745 ;
        RECT 72.190 156.670 72.360 156.925 ;
        RECT 72.190 156.340 72.465 156.670 ;
        RECT 72.190 156.195 72.360 156.340 ;
        RECT 68.335 155.095 68.665 155.815 ;
        RECT 68.845 155.095 71.435 156.185 ;
        RECT 71.685 156.025 72.360 156.195 ;
        RECT 72.635 156.170 72.815 156.970 ;
        RECT 72.995 156.835 73.265 157.645 ;
        RECT 73.435 156.835 73.765 157.475 ;
        RECT 73.935 156.835 74.175 157.645 ;
        RECT 74.455 157.095 74.625 157.475 ;
        RECT 74.805 157.265 75.135 157.645 ;
        RECT 74.455 156.925 75.120 157.095 ;
        RECT 75.315 156.970 75.575 157.475 ;
        RECT 76.075 157.245 76.405 157.645 ;
        RECT 76.575 157.075 76.905 157.415 ;
        RECT 77.955 157.245 78.285 157.645 ;
        RECT 72.985 156.405 73.335 156.655 ;
        RECT 73.505 156.235 73.675 156.835 ;
        RECT 73.845 156.405 74.195 156.655 ;
        RECT 74.385 156.375 74.725 156.745 ;
        RECT 74.950 156.670 75.120 156.925 ;
        RECT 74.950 156.340 75.225 156.670 ;
        RECT 71.685 155.265 71.865 156.025 ;
        RECT 72.045 155.095 72.375 155.855 ;
        RECT 72.545 155.265 72.815 156.170 ;
        RECT 72.995 155.095 73.325 156.235 ;
        RECT 73.505 156.065 74.185 156.235 ;
        RECT 74.950 156.195 75.120 156.340 ;
        RECT 73.855 155.280 74.185 156.065 ;
        RECT 74.445 156.025 75.120 156.195 ;
        RECT 75.395 156.170 75.575 156.970 ;
        RECT 74.445 155.265 74.625 156.025 ;
        RECT 74.805 155.095 75.135 155.855 ;
        RECT 75.305 155.265 75.575 156.170 ;
        RECT 75.920 156.905 78.285 157.075 ;
        RECT 78.455 156.920 78.785 157.430 ;
        RECT 75.920 155.905 76.090 156.905 ;
        RECT 78.115 156.735 78.285 156.905 ;
        RECT 76.260 156.075 76.505 156.735 ;
        RECT 76.720 156.075 76.985 156.735 ;
        RECT 77.180 156.075 77.465 156.735 ;
        RECT 77.640 156.405 77.945 156.735 ;
        RECT 78.115 156.405 78.425 156.735 ;
        RECT 77.640 156.075 77.855 156.405 ;
        RECT 75.920 155.735 76.375 155.905 ;
        RECT 76.045 155.305 76.375 155.735 ;
        RECT 76.555 155.735 77.845 155.905 ;
        RECT 76.555 155.315 76.805 155.735 ;
        RECT 77.035 155.095 77.365 155.565 ;
        RECT 77.595 155.315 77.845 155.735 ;
        RECT 78.035 155.095 78.285 156.235 ;
        RECT 78.595 156.155 78.785 156.920 ;
        RECT 78.455 155.305 78.785 156.155 ;
        RECT 78.980 155.275 79.260 157.465 ;
        RECT 79.460 157.275 80.190 157.645 ;
        RECT 80.770 157.105 81.200 157.465 ;
        RECT 79.460 156.915 81.200 157.105 ;
        RECT 79.460 156.405 79.720 156.915 ;
        RECT 79.450 155.095 79.735 156.235 ;
        RECT 79.930 156.115 80.190 156.735 ;
        RECT 80.385 156.115 80.810 156.735 ;
        RECT 80.980 156.685 81.200 156.915 ;
        RECT 81.370 156.865 81.615 157.645 ;
        RECT 80.980 156.385 81.525 156.685 ;
        RECT 81.815 156.565 82.045 157.465 ;
        RECT 80.000 155.745 81.025 155.945 ;
        RECT 80.000 155.275 80.170 155.745 ;
        RECT 80.345 155.095 80.675 155.575 ;
        RECT 80.845 155.275 81.025 155.745 ;
        RECT 81.195 155.275 81.525 156.385 ;
        RECT 81.705 155.885 82.045 156.565 ;
        RECT 82.225 156.065 82.455 157.405 ;
        RECT 82.645 156.920 82.985 157.645 ;
        RECT 83.155 156.735 83.360 157.335 ;
        RECT 83.590 157.130 84.540 157.315 ;
        RECT 82.670 156.105 82.925 156.735 ;
        RECT 83.155 156.105 83.535 156.735 ;
        RECT 83.795 156.405 84.015 157.130 ;
        RECT 84.710 156.995 85.125 157.430 ;
        RECT 85.315 157.165 85.645 157.645 ;
        RECT 85.815 157.170 86.155 157.430 ;
        RECT 84.710 156.920 85.725 156.995 ;
        RECT 84.905 156.825 85.725 156.920 ;
        RECT 84.325 156.405 84.705 156.735 ;
        RECT 84.405 156.285 84.705 156.405 ;
        RECT 84.405 156.115 84.715 156.285 ;
        RECT 84.405 156.110 84.705 156.115 ;
        RECT 84.905 156.095 85.235 156.655 ;
        RECT 81.705 155.685 82.455 155.885 ;
        RECT 81.695 155.095 82.045 155.505 ;
        RECT 82.215 155.295 82.455 155.685 ;
        RECT 82.735 155.765 84.705 155.935 ;
        RECT 85.555 155.905 85.725 156.825 ;
        RECT 82.735 155.265 82.905 155.765 ;
        RECT 83.145 155.095 83.395 155.555 ;
        RECT 83.695 155.265 83.865 155.765 ;
        RECT 84.075 155.095 84.325 155.555 ;
        RECT 84.535 155.265 84.705 155.765 ;
        RECT 84.875 155.735 85.725 155.905 ;
        RECT 84.875 155.305 85.205 155.735 ;
        RECT 85.895 155.565 86.155 157.170 ;
        RECT 86.325 156.845 87.020 157.475 ;
        RECT 87.225 156.845 87.535 157.645 ;
        RECT 87.705 156.920 87.995 157.645 ;
        RECT 89.105 156.955 89.345 157.475 ;
        RECT 89.515 157.150 89.910 157.645 ;
        RECT 90.475 157.315 90.645 157.460 ;
        RECT 90.270 157.120 90.645 157.315 ;
        RECT 86.345 156.405 86.680 156.655 ;
        RECT 86.850 156.245 87.020 156.845 ;
        RECT 87.190 156.405 87.525 156.675 ;
        RECT 85.395 155.095 85.645 155.555 ;
        RECT 85.815 155.305 86.155 155.565 ;
        RECT 86.325 155.095 86.585 156.235 ;
        RECT 86.755 155.265 87.085 156.245 ;
        RECT 87.255 155.095 87.535 156.235 ;
        RECT 87.705 155.095 87.995 156.260 ;
        RECT 89.105 156.150 89.280 156.955 ;
        RECT 90.270 156.785 90.440 157.120 ;
        RECT 90.925 157.075 91.165 157.450 ;
        RECT 91.335 157.140 91.670 157.645 ;
        RECT 90.925 156.925 91.145 157.075 ;
        RECT 92.305 156.995 92.565 157.475 ;
        RECT 92.735 157.105 92.985 157.645 ;
        RECT 89.455 156.425 90.440 156.785 ;
        RECT 90.610 156.595 91.145 156.925 ;
        RECT 89.455 156.405 90.740 156.425 ;
        RECT 89.880 156.255 90.740 156.405 ;
        RECT 89.105 155.365 89.410 156.150 ;
        RECT 89.585 155.775 90.280 156.085 ;
        RECT 89.590 155.095 90.275 155.565 ;
        RECT 90.455 155.310 90.740 156.255 ;
        RECT 90.910 155.945 91.145 156.595 ;
        RECT 91.315 156.115 91.615 156.965 ;
        RECT 92.305 155.965 92.475 156.995 ;
        RECT 93.155 156.940 93.375 157.425 ;
        RECT 92.645 156.345 92.875 156.740 ;
        RECT 93.045 156.515 93.375 156.940 ;
        RECT 93.545 157.265 94.435 157.435 ;
        RECT 93.545 156.540 93.715 157.265 ;
        RECT 94.695 157.095 94.865 157.475 ;
        RECT 95.045 157.265 95.375 157.645 ;
        RECT 93.885 156.710 94.435 157.095 ;
        RECT 94.695 156.925 95.360 157.095 ;
        RECT 95.555 156.970 95.815 157.475 ;
        RECT 93.545 156.470 94.435 156.540 ;
        RECT 93.540 156.445 94.435 156.470 ;
        RECT 93.530 156.430 94.435 156.445 ;
        RECT 93.525 156.415 94.435 156.430 ;
        RECT 93.515 156.410 94.435 156.415 ;
        RECT 93.510 156.400 94.435 156.410 ;
        RECT 93.505 156.390 94.435 156.400 ;
        RECT 93.495 156.385 94.435 156.390 ;
        RECT 93.485 156.375 94.435 156.385 ;
        RECT 94.625 156.375 94.965 156.745 ;
        RECT 95.190 156.670 95.360 156.925 ;
        RECT 93.475 156.370 94.435 156.375 ;
        RECT 93.475 156.365 93.810 156.370 ;
        RECT 93.460 156.360 93.810 156.365 ;
        RECT 93.445 156.350 93.810 156.360 ;
        RECT 93.420 156.345 93.810 156.350 ;
        RECT 92.645 156.340 93.810 156.345 ;
        RECT 92.645 156.305 93.780 156.340 ;
        RECT 92.645 156.280 93.745 156.305 ;
        RECT 92.645 156.250 93.715 156.280 ;
        RECT 92.645 156.220 93.695 156.250 ;
        RECT 92.645 156.190 93.675 156.220 ;
        RECT 92.645 156.180 93.605 156.190 ;
        RECT 92.645 156.170 93.580 156.180 ;
        RECT 92.645 156.155 93.560 156.170 ;
        RECT 92.645 156.140 93.540 156.155 ;
        RECT 92.750 156.130 93.535 156.140 ;
        RECT 92.750 156.095 93.520 156.130 ;
        RECT 90.910 155.715 91.585 155.945 ;
        RECT 90.915 155.095 91.245 155.545 ;
        RECT 91.415 155.285 91.585 155.715 ;
        RECT 92.305 155.265 92.580 155.965 ;
        RECT 92.750 155.845 93.505 156.095 ;
        RECT 93.675 155.775 94.005 156.020 ;
        RECT 94.175 155.920 94.435 156.370 ;
        RECT 95.190 156.340 95.465 156.670 ;
        RECT 95.190 156.195 95.360 156.340 ;
        RECT 94.685 156.025 95.360 156.195 ;
        RECT 95.635 156.170 95.815 156.970 ;
        RECT 95.985 156.875 98.575 157.645 ;
        RECT 95.985 156.355 97.195 156.875 ;
        RECT 97.365 156.185 98.575 156.705 ;
        RECT 93.820 155.750 94.005 155.775 ;
        RECT 93.820 155.650 94.435 155.750 ;
        RECT 92.750 155.095 93.005 155.640 ;
        RECT 93.175 155.265 93.655 155.605 ;
        RECT 93.830 155.095 94.435 155.650 ;
        RECT 94.685 155.265 94.865 156.025 ;
        RECT 95.045 155.095 95.375 155.855 ;
        RECT 95.545 155.265 95.815 156.170 ;
        RECT 95.985 155.095 98.575 156.185 ;
        RECT 98.745 155.265 99.025 157.365 ;
        RECT 99.255 157.185 99.425 157.645 ;
        RECT 99.695 157.255 100.945 157.435 ;
        RECT 100.080 157.015 100.445 157.085 ;
        RECT 99.195 156.835 100.445 157.015 ;
        RECT 100.615 157.035 100.945 157.255 ;
        RECT 101.115 157.205 101.285 157.645 ;
        RECT 101.455 157.035 101.795 157.450 ;
        RECT 100.615 156.865 101.795 157.035 ;
        RECT 101.965 156.845 102.275 157.645 ;
        RECT 102.480 156.845 103.175 157.475 ;
        RECT 103.345 157.100 108.690 157.645 ;
        RECT 99.195 156.235 99.470 156.835 ;
        RECT 99.640 156.405 99.995 156.655 ;
        RECT 100.190 156.625 100.655 156.655 ;
        RECT 100.185 156.455 100.655 156.625 ;
        RECT 100.190 156.405 100.655 156.455 ;
        RECT 100.825 156.405 101.155 156.655 ;
        RECT 101.330 156.455 101.795 156.655 ;
        RECT 101.975 156.405 102.310 156.675 ;
        RECT 100.975 156.285 101.155 156.405 ;
        RECT 99.195 156.025 100.805 156.235 ;
        RECT 100.975 156.115 101.305 156.285 ;
        RECT 100.395 155.925 100.805 156.025 ;
        RECT 99.215 155.095 100.000 155.855 ;
        RECT 100.395 155.265 100.780 155.925 ;
        RECT 101.105 155.325 101.305 156.115 ;
        RECT 101.475 155.095 101.795 156.275 ;
        RECT 102.480 156.245 102.650 156.845 ;
        RECT 102.820 156.405 103.155 156.655 ;
        RECT 104.930 156.270 105.270 157.100 ;
        RECT 109.070 156.865 109.570 157.475 ;
        RECT 101.965 155.095 102.245 156.235 ;
        RECT 102.415 155.265 102.745 156.245 ;
        RECT 102.915 155.095 103.175 156.235 ;
        RECT 106.750 155.530 107.100 156.780 ;
        RECT 108.865 156.405 109.215 156.655 ;
        RECT 109.400 156.235 109.570 156.865 ;
        RECT 110.200 156.995 110.530 157.475 ;
        RECT 110.700 157.185 110.925 157.645 ;
        RECT 111.095 156.995 111.425 157.475 ;
        RECT 110.200 156.825 111.425 156.995 ;
        RECT 111.615 156.845 111.865 157.645 ;
        RECT 112.035 156.845 112.375 157.475 ;
        RECT 113.465 156.920 113.755 157.645 ;
        RECT 113.925 156.845 114.620 157.475 ;
        RECT 114.825 156.845 115.135 157.645 ;
        RECT 115.305 156.875 118.815 157.645 ;
        RECT 109.740 156.455 110.070 156.655 ;
        RECT 110.240 156.455 110.570 156.655 ;
        RECT 110.740 156.455 111.160 156.655 ;
        RECT 111.335 156.485 112.030 156.655 ;
        RECT 111.335 156.235 111.505 156.485 ;
        RECT 112.200 156.235 112.375 156.845 ;
        RECT 113.945 156.405 114.280 156.655 ;
        RECT 109.070 156.065 111.505 156.235 ;
        RECT 103.345 155.095 108.690 155.530 ;
        RECT 109.070 155.265 109.400 156.065 ;
        RECT 109.570 155.095 109.900 155.895 ;
        RECT 110.200 155.265 110.530 156.065 ;
        RECT 111.175 155.095 111.425 155.895 ;
        RECT 111.695 155.095 111.865 156.235 ;
        RECT 112.035 155.265 112.375 156.235 ;
        RECT 113.465 155.095 113.755 156.260 ;
        RECT 114.450 156.245 114.620 156.845 ;
        RECT 114.790 156.405 115.125 156.675 ;
        RECT 115.305 156.355 116.955 156.875 ;
        RECT 119.925 156.835 120.165 157.645 ;
        RECT 120.335 156.835 120.665 157.475 ;
        RECT 120.835 156.835 121.105 157.645 ;
        RECT 121.285 156.875 122.955 157.645 ;
        RECT 113.925 155.095 114.185 156.235 ;
        RECT 114.355 155.265 114.685 156.245 ;
        RECT 114.855 155.095 115.135 156.235 ;
        RECT 117.125 156.185 118.815 156.705 ;
        RECT 119.905 156.405 120.255 156.655 ;
        RECT 120.425 156.235 120.595 156.835 ;
        RECT 120.765 156.405 121.115 156.655 ;
        RECT 121.285 156.355 122.035 156.875 ;
        RECT 123.185 156.825 123.395 157.645 ;
        RECT 123.565 156.845 123.895 157.475 ;
        RECT 115.305 155.095 118.815 156.185 ;
        RECT 119.915 156.065 120.595 156.235 ;
        RECT 119.915 155.280 120.245 156.065 ;
        RECT 120.775 155.095 121.105 156.235 ;
        RECT 122.205 156.185 122.955 156.705 ;
        RECT 123.565 156.245 123.815 156.845 ;
        RECT 124.065 156.825 124.295 157.645 ;
        RECT 124.595 157.095 124.765 157.475 ;
        RECT 124.945 157.265 125.275 157.645 ;
        RECT 124.595 156.925 125.260 157.095 ;
        RECT 125.455 156.970 125.715 157.475 ;
        RECT 123.985 156.405 124.315 156.655 ;
        RECT 124.525 156.375 124.865 156.745 ;
        RECT 125.090 156.670 125.260 156.925 ;
        RECT 125.090 156.340 125.365 156.670 ;
        RECT 121.285 155.095 122.955 156.185 ;
        RECT 123.185 155.095 123.395 156.235 ;
        RECT 123.565 155.265 123.895 156.245 ;
        RECT 124.065 155.095 124.295 156.235 ;
        RECT 125.090 156.195 125.260 156.340 ;
        RECT 124.585 156.025 125.260 156.195 ;
        RECT 125.535 156.170 125.715 156.970 ;
        RECT 125.945 156.825 126.155 157.645 ;
        RECT 126.325 156.845 126.655 157.475 ;
        RECT 126.325 156.245 126.575 156.845 ;
        RECT 126.825 156.825 127.055 157.645 ;
        RECT 128.185 157.265 129.075 157.435 ;
        RECT 128.185 156.710 128.735 157.095 ;
        RECT 126.745 156.405 127.075 156.655 ;
        RECT 128.905 156.540 129.075 157.265 ;
        RECT 128.185 156.470 129.075 156.540 ;
        RECT 129.245 156.940 129.465 157.425 ;
        RECT 129.635 157.105 129.885 157.645 ;
        RECT 130.055 156.995 130.315 157.475 ;
        RECT 131.570 157.135 131.810 157.645 ;
        RECT 131.990 157.135 132.270 157.465 ;
        RECT 132.500 157.135 132.715 157.645 ;
        RECT 129.245 156.515 129.575 156.940 ;
        RECT 128.185 156.445 129.080 156.470 ;
        RECT 128.185 156.430 129.090 156.445 ;
        RECT 128.185 156.415 129.095 156.430 ;
        RECT 128.185 156.410 129.105 156.415 ;
        RECT 128.185 156.400 129.110 156.410 ;
        RECT 128.185 156.390 129.115 156.400 ;
        RECT 128.185 156.385 129.125 156.390 ;
        RECT 128.185 156.375 129.135 156.385 ;
        RECT 128.185 156.370 129.145 156.375 ;
        RECT 124.585 155.265 124.765 156.025 ;
        RECT 124.945 155.095 125.275 155.855 ;
        RECT 125.445 155.265 125.715 156.170 ;
        RECT 125.945 155.095 126.155 156.235 ;
        RECT 126.325 155.265 126.655 156.245 ;
        RECT 126.825 155.095 127.055 156.235 ;
        RECT 128.185 155.920 128.445 156.370 ;
        RECT 128.810 156.365 129.145 156.370 ;
        RECT 128.810 156.360 129.160 156.365 ;
        RECT 128.810 156.350 129.175 156.360 ;
        RECT 128.810 156.345 129.200 156.350 ;
        RECT 129.745 156.345 129.975 156.740 ;
        RECT 128.810 156.340 129.975 156.345 ;
        RECT 128.840 156.305 129.975 156.340 ;
        RECT 128.875 156.280 129.975 156.305 ;
        RECT 128.905 156.250 129.975 156.280 ;
        RECT 128.925 156.220 129.975 156.250 ;
        RECT 128.945 156.190 129.975 156.220 ;
        RECT 129.015 156.180 129.975 156.190 ;
        RECT 129.040 156.170 129.975 156.180 ;
        RECT 129.060 156.155 129.975 156.170 ;
        RECT 129.080 156.140 129.975 156.155 ;
        RECT 129.085 156.130 129.870 156.140 ;
        RECT 129.100 156.095 129.870 156.130 ;
        RECT 128.615 155.775 128.945 156.020 ;
        RECT 129.115 155.845 129.870 156.095 ;
        RECT 130.145 155.965 130.315 156.995 ;
        RECT 131.465 156.405 131.820 156.965 ;
        RECT 131.990 156.235 132.160 157.135 ;
        RECT 132.330 156.405 132.595 156.965 ;
        RECT 132.885 156.905 133.500 157.475 ;
        RECT 132.845 156.235 133.015 156.735 ;
        RECT 128.615 155.750 128.800 155.775 ;
        RECT 128.185 155.650 128.800 155.750 ;
        RECT 128.185 155.095 128.790 155.650 ;
        RECT 128.965 155.265 129.445 155.605 ;
        RECT 129.615 155.095 129.870 155.640 ;
        RECT 130.040 155.265 130.315 155.965 ;
        RECT 131.590 156.065 133.015 156.235 ;
        RECT 131.590 155.890 131.980 156.065 ;
        RECT 132.465 155.095 132.795 155.895 ;
        RECT 133.185 155.885 133.500 156.905 ;
        RECT 132.965 155.265 133.500 155.885 ;
        RECT 133.705 156.970 133.965 157.475 ;
        RECT 134.145 157.265 134.475 157.645 ;
        RECT 134.655 157.095 134.825 157.475 ;
        RECT 133.705 156.170 133.885 156.970 ;
        RECT 134.160 156.925 134.825 157.095 ;
        RECT 134.160 156.670 134.330 156.925 ;
        RECT 135.085 156.875 138.595 157.645 ;
        RECT 139.225 156.920 139.515 157.645 ;
        RECT 139.775 157.095 139.945 157.385 ;
        RECT 140.115 157.265 140.445 157.645 ;
        RECT 139.775 156.925 140.440 157.095 ;
        RECT 134.055 156.340 134.330 156.670 ;
        RECT 134.555 156.375 134.895 156.745 ;
        RECT 135.085 156.355 136.735 156.875 ;
        RECT 134.160 156.195 134.330 156.340 ;
        RECT 133.705 155.265 133.975 156.170 ;
        RECT 134.160 156.025 134.835 156.195 ;
        RECT 136.905 156.185 138.595 156.705 ;
        RECT 134.145 155.095 134.475 155.855 ;
        RECT 134.655 155.265 134.835 156.025 ;
        RECT 135.085 155.095 138.595 156.185 ;
        RECT 139.225 155.095 139.515 156.260 ;
        RECT 139.690 156.105 140.040 156.755 ;
        RECT 140.210 155.935 140.440 156.925 ;
        RECT 139.775 155.765 140.440 155.935 ;
        RECT 139.775 155.265 139.945 155.765 ;
        RECT 140.115 155.095 140.445 155.595 ;
        RECT 140.615 155.265 140.800 157.385 ;
        RECT 141.055 157.185 141.305 157.645 ;
        RECT 141.475 157.195 141.810 157.365 ;
        RECT 142.005 157.195 142.680 157.365 ;
        RECT 141.475 157.055 141.645 157.195 ;
        RECT 140.970 156.065 141.250 157.015 ;
        RECT 141.420 156.925 141.645 157.055 ;
        RECT 141.420 155.820 141.590 156.925 ;
        RECT 141.815 156.775 142.340 156.995 ;
        RECT 141.760 156.010 142.000 156.605 ;
        RECT 142.170 156.075 142.340 156.775 ;
        RECT 142.510 156.415 142.680 157.195 ;
        RECT 143.000 157.145 143.370 157.645 ;
        RECT 143.550 157.195 143.955 157.365 ;
        RECT 144.125 157.195 144.910 157.365 ;
        RECT 143.550 156.965 143.720 157.195 ;
        RECT 142.890 156.665 143.720 156.965 ;
        RECT 144.105 156.695 144.570 157.025 ;
        RECT 142.890 156.635 143.090 156.665 ;
        RECT 143.210 156.415 143.380 156.485 ;
        RECT 142.510 156.245 143.380 156.415 ;
        RECT 142.870 156.155 143.380 156.245 ;
        RECT 141.420 155.690 141.725 155.820 ;
        RECT 142.170 155.710 142.700 156.075 ;
        RECT 141.040 155.095 141.305 155.555 ;
        RECT 141.475 155.265 141.725 155.690 ;
        RECT 142.870 155.540 143.040 156.155 ;
        RECT 141.935 155.370 143.040 155.540 ;
        RECT 143.210 155.095 143.380 155.895 ;
        RECT 143.550 155.595 143.720 156.665 ;
        RECT 143.890 155.765 144.080 156.485 ;
        RECT 144.250 155.735 144.570 156.695 ;
        RECT 144.740 156.735 144.910 157.195 ;
        RECT 145.185 157.115 145.395 157.645 ;
        RECT 145.655 156.905 145.985 157.430 ;
        RECT 146.155 157.035 146.325 157.645 ;
        RECT 146.495 156.990 146.825 157.425 ;
        RECT 146.495 156.905 146.875 156.990 ;
        RECT 145.785 156.735 145.985 156.905 ;
        RECT 146.650 156.865 146.875 156.905 ;
        RECT 144.740 156.405 145.615 156.735 ;
        RECT 145.785 156.405 146.535 156.735 ;
        RECT 143.550 155.265 143.800 155.595 ;
        RECT 144.740 155.565 144.910 156.405 ;
        RECT 145.785 156.200 145.975 156.405 ;
        RECT 146.705 156.285 146.875 156.865 ;
        RECT 147.045 156.875 148.715 157.645 ;
        RECT 148.885 156.895 150.095 157.645 ;
        RECT 147.045 156.355 147.795 156.875 ;
        RECT 146.660 156.235 146.875 156.285 ;
        RECT 145.080 155.825 145.975 156.200 ;
        RECT 146.485 156.155 146.875 156.235 ;
        RECT 147.965 156.185 148.715 156.705 ;
        RECT 144.025 155.395 144.910 155.565 ;
        RECT 145.090 155.095 145.405 155.595 ;
        RECT 145.635 155.265 145.975 155.825 ;
        RECT 146.145 155.095 146.315 156.105 ;
        RECT 146.485 155.310 146.815 156.155 ;
        RECT 147.045 155.095 148.715 156.185 ;
        RECT 148.885 156.185 149.405 156.725 ;
        RECT 149.575 156.355 150.095 156.895 ;
        RECT 148.885 155.095 150.095 156.185 ;
        RECT 36.100 154.925 150.180 155.095 ;
        RECT 36.185 153.835 37.395 154.925 ;
        RECT 37.565 153.835 40.155 154.925 ;
        RECT 36.185 153.125 36.705 153.665 ;
        RECT 36.875 153.295 37.395 153.835 ;
        RECT 37.565 153.145 38.775 153.665 ;
        RECT 38.945 153.315 40.155 153.835 ;
        RECT 40.325 153.850 40.595 154.755 ;
        RECT 40.765 154.165 41.095 154.925 ;
        RECT 41.275 153.995 41.445 154.755 ;
        RECT 36.185 152.375 37.395 153.125 ;
        RECT 37.565 152.375 40.155 153.145 ;
        RECT 40.325 153.050 40.495 153.850 ;
        RECT 40.780 153.825 41.445 153.995 ;
        RECT 42.165 153.850 42.435 154.755 ;
        RECT 42.605 154.165 42.935 154.925 ;
        RECT 43.115 153.995 43.285 154.755 ;
        RECT 40.780 153.680 40.950 153.825 ;
        RECT 40.665 153.350 40.950 153.680 ;
        RECT 40.780 153.095 40.950 153.350 ;
        RECT 41.185 153.275 41.515 153.645 ;
        RECT 40.325 152.545 40.585 153.050 ;
        RECT 40.780 152.925 41.445 153.095 ;
        RECT 40.765 152.375 41.095 152.755 ;
        RECT 41.275 152.545 41.445 152.925 ;
        RECT 42.165 153.050 42.335 153.850 ;
        RECT 42.620 153.825 43.285 153.995 ;
        RECT 43.545 153.835 44.755 154.925 ;
        RECT 42.620 153.680 42.790 153.825 ;
        RECT 42.505 153.350 42.790 153.680 ;
        RECT 42.620 153.095 42.790 153.350 ;
        RECT 43.025 153.275 43.355 153.645 ;
        RECT 43.545 153.125 44.065 153.665 ;
        RECT 44.235 153.295 44.755 153.835 ;
        RECT 44.925 153.785 45.185 154.925 ;
        RECT 45.355 153.775 45.685 154.755 ;
        RECT 45.855 153.785 46.135 154.925 ;
        RECT 46.305 154.055 46.580 154.755 ;
        RECT 46.750 154.380 47.005 154.925 ;
        RECT 47.175 154.415 47.655 154.755 ;
        RECT 47.830 154.370 48.435 154.925 ;
        RECT 47.820 154.270 48.435 154.370 ;
        RECT 47.820 154.245 48.005 154.270 ;
        RECT 44.945 153.365 45.280 153.615 ;
        RECT 45.450 153.175 45.620 153.775 ;
        RECT 45.790 153.345 46.125 153.615 ;
        RECT 42.165 152.545 42.425 153.050 ;
        RECT 42.620 152.925 43.285 153.095 ;
        RECT 42.605 152.375 42.935 152.755 ;
        RECT 43.115 152.545 43.285 152.925 ;
        RECT 43.545 152.375 44.755 153.125 ;
        RECT 44.925 152.545 45.620 153.175 ;
        RECT 45.825 152.375 46.135 153.175 ;
        RECT 46.305 153.025 46.475 154.055 ;
        RECT 46.750 153.925 47.505 154.175 ;
        RECT 47.675 154.000 48.005 154.245 ;
        RECT 46.750 153.890 47.520 153.925 ;
        RECT 46.750 153.880 47.535 153.890 ;
        RECT 46.645 153.865 47.540 153.880 ;
        RECT 46.645 153.850 47.560 153.865 ;
        RECT 46.645 153.840 47.580 153.850 ;
        RECT 46.645 153.830 47.605 153.840 ;
        RECT 46.645 153.800 47.675 153.830 ;
        RECT 46.645 153.770 47.695 153.800 ;
        RECT 46.645 153.740 47.715 153.770 ;
        RECT 46.645 153.715 47.745 153.740 ;
        RECT 46.645 153.680 47.780 153.715 ;
        RECT 46.645 153.675 47.810 153.680 ;
        RECT 46.645 153.280 46.875 153.675 ;
        RECT 47.420 153.670 47.810 153.675 ;
        RECT 47.445 153.660 47.810 153.670 ;
        RECT 47.460 153.655 47.810 153.660 ;
        RECT 47.475 153.650 47.810 153.655 ;
        RECT 48.175 153.650 48.435 154.100 ;
        RECT 49.065 153.760 49.355 154.925 ;
        RECT 49.560 154.135 50.095 154.755 ;
        RECT 47.475 153.645 48.435 153.650 ;
        RECT 47.485 153.635 48.435 153.645 ;
        RECT 47.495 153.630 48.435 153.635 ;
        RECT 47.505 153.620 48.435 153.630 ;
        RECT 47.510 153.610 48.435 153.620 ;
        RECT 47.515 153.605 48.435 153.610 ;
        RECT 47.525 153.590 48.435 153.605 ;
        RECT 47.530 153.575 48.435 153.590 ;
        RECT 47.540 153.550 48.435 153.575 ;
        RECT 47.045 153.080 47.375 153.505 ;
        RECT 46.305 152.545 46.565 153.025 ;
        RECT 46.735 152.375 46.985 152.915 ;
        RECT 47.155 152.595 47.375 153.080 ;
        RECT 47.545 153.480 48.435 153.550 ;
        RECT 47.545 152.755 47.715 153.480 ;
        RECT 47.885 152.925 48.435 153.310 ;
        RECT 49.560 153.115 49.875 154.135 ;
        RECT 50.265 154.125 50.595 154.925 ;
        RECT 51.825 154.490 57.170 154.925 ;
        RECT 57.345 154.490 62.690 154.925 ;
        RECT 51.080 153.955 51.470 154.130 ;
        RECT 50.045 153.785 51.470 153.955 ;
        RECT 50.045 153.285 50.215 153.785 ;
        RECT 47.545 152.585 48.435 152.755 ;
        RECT 49.065 152.375 49.355 153.100 ;
        RECT 49.560 152.545 50.175 153.115 ;
        RECT 50.465 153.055 50.730 153.615 ;
        RECT 50.900 152.885 51.070 153.785 ;
        RECT 51.240 153.055 51.595 153.615 ;
        RECT 53.410 152.920 53.750 153.750 ;
        RECT 55.230 153.240 55.580 154.490 ;
        RECT 58.930 152.920 59.270 153.750 ;
        RECT 60.750 153.240 61.100 154.490 ;
        RECT 62.865 153.835 64.535 154.925 ;
        RECT 62.865 153.145 63.615 153.665 ;
        RECT 63.785 153.315 64.535 153.835 ;
        RECT 65.165 154.055 65.440 154.755 ;
        RECT 65.650 154.380 65.865 154.925 ;
        RECT 66.035 154.415 66.510 154.755 ;
        RECT 66.680 154.420 67.295 154.925 ;
        RECT 66.680 154.245 66.875 154.420 ;
        RECT 50.345 152.375 50.560 152.885 ;
        RECT 50.790 152.555 51.070 152.885 ;
        RECT 51.250 152.375 51.490 152.885 ;
        RECT 51.825 152.375 57.170 152.920 ;
        RECT 57.345 152.375 62.690 152.920 ;
        RECT 62.865 152.375 64.535 153.145 ;
        RECT 65.165 153.025 65.335 154.055 ;
        RECT 65.610 153.885 66.325 154.180 ;
        RECT 66.545 154.055 66.875 154.245 ;
        RECT 67.045 153.885 67.295 154.250 ;
        RECT 65.505 153.715 67.295 153.885 ;
        RECT 65.505 153.285 65.735 153.715 ;
        RECT 65.165 152.545 65.425 153.025 ;
        RECT 65.905 153.015 66.315 153.535 ;
        RECT 65.595 152.375 65.925 152.835 ;
        RECT 66.115 152.595 66.315 153.015 ;
        RECT 66.485 152.860 66.740 153.715 ;
        RECT 67.535 153.535 67.705 154.755 ;
        RECT 67.955 154.415 68.215 154.925 ;
        RECT 66.910 153.285 67.705 153.535 ;
        RECT 67.875 153.365 68.215 154.245 ;
        RECT 68.385 153.835 70.055 154.925 ;
        RECT 67.455 153.195 67.705 153.285 ;
        RECT 66.485 152.595 67.275 152.860 ;
        RECT 67.455 152.775 67.785 153.195 ;
        RECT 67.955 152.375 68.215 153.195 ;
        RECT 68.385 153.145 69.135 153.665 ;
        RECT 69.305 153.315 70.055 153.835 ;
        RECT 70.720 154.135 71.255 154.755 ;
        RECT 68.385 152.375 70.055 153.145 ;
        RECT 70.720 153.115 71.035 154.135 ;
        RECT 71.425 154.125 71.755 154.925 ;
        RECT 72.240 153.955 72.630 154.130 ;
        RECT 71.205 153.785 72.630 153.955 ;
        RECT 72.985 153.835 74.655 154.925 ;
        RECT 71.205 153.285 71.375 153.785 ;
        RECT 70.720 152.545 71.335 153.115 ;
        RECT 71.625 153.055 71.890 153.615 ;
        RECT 72.060 152.885 72.230 153.785 ;
        RECT 72.400 153.055 72.755 153.615 ;
        RECT 72.985 153.145 73.735 153.665 ;
        RECT 73.905 153.315 74.655 153.835 ;
        RECT 74.825 153.760 75.115 154.925 ;
        RECT 75.285 153.835 77.875 154.925 ;
        RECT 75.285 153.145 76.495 153.665 ;
        RECT 76.665 153.315 77.875 153.835 ;
        RECT 78.125 153.995 78.305 154.755 ;
        RECT 78.485 154.165 78.815 154.925 ;
        RECT 78.125 153.825 78.800 153.995 ;
        RECT 78.985 153.850 79.255 154.755 ;
        RECT 78.630 153.680 78.800 153.825 ;
        RECT 78.065 153.275 78.405 153.645 ;
        RECT 78.630 153.350 78.905 153.680 ;
        RECT 71.505 152.375 71.720 152.885 ;
        RECT 71.950 152.555 72.230 152.885 ;
        RECT 72.410 152.375 72.650 152.885 ;
        RECT 72.985 152.375 74.655 153.145 ;
        RECT 74.825 152.375 75.115 153.100 ;
        RECT 75.285 152.375 77.875 153.145 ;
        RECT 78.630 153.095 78.800 153.350 ;
        RECT 78.135 152.925 78.800 153.095 ;
        RECT 79.075 153.050 79.255 153.850 ;
        RECT 79.465 153.975 79.755 154.745 ;
        RECT 80.325 154.385 80.585 154.745 ;
        RECT 80.755 154.555 81.085 154.925 ;
        RECT 81.255 154.385 81.515 154.745 ;
        RECT 80.325 154.155 81.515 154.385 ;
        RECT 81.705 154.205 82.035 154.925 ;
        RECT 82.205 153.975 82.470 154.745 ;
        RECT 79.465 153.795 81.960 153.975 ;
        RECT 79.435 153.285 79.705 153.615 ;
        RECT 79.885 153.285 80.320 153.615 ;
        RECT 80.500 153.285 81.075 153.615 ;
        RECT 81.255 153.285 81.535 153.615 ;
        RECT 81.735 153.105 81.960 153.795 ;
        RECT 78.135 152.545 78.305 152.925 ;
        RECT 78.485 152.375 78.815 152.755 ;
        RECT 78.995 152.545 79.255 153.050 ;
        RECT 79.475 152.915 81.960 153.105 ;
        RECT 79.475 152.555 79.700 152.915 ;
        RECT 79.880 152.375 80.210 152.745 ;
        RECT 80.390 152.555 80.645 152.915 ;
        RECT 81.210 152.375 81.955 152.745 ;
        RECT 82.135 152.555 82.470 153.975 ;
        RECT 83.290 153.955 83.680 154.130 ;
        RECT 84.165 154.125 84.495 154.925 ;
        RECT 84.665 154.135 85.200 154.755 ;
        RECT 85.865 154.330 86.300 154.755 ;
        RECT 86.470 154.500 86.855 154.925 ;
        RECT 85.865 154.160 86.855 154.330 ;
        RECT 83.290 153.785 84.715 153.955 ;
        RECT 83.165 153.055 83.520 153.615 ;
        RECT 83.690 152.885 83.860 153.785 ;
        RECT 84.030 153.055 84.295 153.615 ;
        RECT 84.545 153.285 84.715 153.785 ;
        RECT 84.885 153.115 85.200 154.135 ;
        RECT 85.865 153.285 86.350 153.990 ;
        RECT 86.520 153.615 86.855 154.160 ;
        RECT 87.025 153.965 87.450 154.755 ;
        RECT 87.620 154.330 87.895 154.755 ;
        RECT 88.065 154.500 88.450 154.925 ;
        RECT 87.620 154.135 88.450 154.330 ;
        RECT 87.025 153.785 87.930 153.965 ;
        RECT 86.520 153.285 86.930 153.615 ;
        RECT 87.100 153.285 87.930 153.785 ;
        RECT 88.100 153.615 88.450 154.135 ;
        RECT 88.620 153.965 88.865 154.755 ;
        RECT 89.055 154.330 89.310 154.755 ;
        RECT 89.480 154.500 89.865 154.925 ;
        RECT 89.055 154.135 89.865 154.330 ;
        RECT 88.620 153.785 89.345 153.965 ;
        RECT 88.100 153.285 88.525 153.615 ;
        RECT 88.695 153.285 89.345 153.785 ;
        RECT 89.515 153.615 89.865 154.135 ;
        RECT 90.035 153.785 90.295 154.755 ;
        RECT 90.465 154.490 95.810 154.925 ;
        RECT 89.515 153.285 89.940 153.615 ;
        RECT 86.520 153.115 86.855 153.285 ;
        RECT 87.100 153.115 87.450 153.285 ;
        RECT 88.100 153.115 88.450 153.285 ;
        RECT 88.695 153.115 88.865 153.285 ;
        RECT 89.515 153.115 89.865 153.285 ;
        RECT 90.110 153.115 90.295 153.785 ;
        RECT 83.270 152.375 83.510 152.885 ;
        RECT 83.690 152.555 83.970 152.885 ;
        RECT 84.200 152.375 84.415 152.885 ;
        RECT 84.585 152.545 85.200 153.115 ;
        RECT 85.865 152.945 86.855 153.115 ;
        RECT 85.865 152.545 86.300 152.945 ;
        RECT 86.470 152.375 86.855 152.775 ;
        RECT 87.025 152.545 87.450 153.115 ;
        RECT 87.640 152.945 88.450 153.115 ;
        RECT 87.640 152.545 87.895 152.945 ;
        RECT 88.065 152.375 88.450 152.775 ;
        RECT 88.620 152.545 88.865 153.115 ;
        RECT 89.055 152.945 89.865 153.115 ;
        RECT 89.055 152.545 89.310 152.945 ;
        RECT 89.480 152.375 89.865 152.775 ;
        RECT 90.035 152.545 90.295 153.115 ;
        RECT 92.050 152.920 92.390 153.750 ;
        RECT 93.870 153.240 94.220 154.490 ;
        RECT 96.905 153.850 97.175 154.755 ;
        RECT 97.345 154.165 97.675 154.925 ;
        RECT 97.855 153.995 98.035 154.755 ;
        RECT 96.905 153.050 97.085 153.850 ;
        RECT 97.360 153.825 98.035 153.995 ;
        RECT 98.470 153.955 98.860 154.130 ;
        RECT 99.345 154.125 99.675 154.925 ;
        RECT 99.845 154.135 100.380 154.755 ;
        RECT 97.360 153.680 97.530 153.825 ;
        RECT 98.470 153.785 99.895 153.955 ;
        RECT 97.255 153.350 97.530 153.680 ;
        RECT 97.360 153.095 97.530 153.350 ;
        RECT 97.755 153.275 98.095 153.645 ;
        RECT 90.465 152.375 95.810 152.920 ;
        RECT 96.905 152.545 97.165 153.050 ;
        RECT 97.360 152.925 98.025 153.095 ;
        RECT 98.345 153.055 98.700 153.615 ;
        RECT 97.345 152.375 97.675 152.755 ;
        RECT 97.855 152.545 98.025 152.925 ;
        RECT 98.870 152.885 99.040 153.785 ;
        RECT 99.210 153.055 99.475 153.615 ;
        RECT 99.725 153.285 99.895 153.785 ;
        RECT 100.065 153.115 100.380 154.135 ;
        RECT 100.585 153.760 100.875 154.925 ;
        RECT 101.345 154.285 101.675 154.715 ;
        RECT 101.220 154.115 101.675 154.285 ;
        RECT 101.855 154.285 102.105 154.705 ;
        RECT 102.335 154.455 102.665 154.925 ;
        RECT 102.895 154.285 103.145 154.705 ;
        RECT 101.855 154.115 103.145 154.285 ;
        RECT 98.450 152.375 98.690 152.885 ;
        RECT 98.870 152.555 99.150 152.885 ;
        RECT 99.380 152.375 99.595 152.885 ;
        RECT 99.765 152.545 100.380 153.115 ;
        RECT 101.220 153.115 101.390 154.115 ;
        RECT 101.560 153.285 101.805 153.945 ;
        RECT 102.020 153.285 102.285 153.945 ;
        RECT 102.480 153.285 102.765 153.945 ;
        RECT 102.940 153.615 103.155 153.945 ;
        RECT 103.335 153.785 103.585 154.925 ;
        RECT 103.755 153.865 104.085 154.715 ;
        RECT 102.940 153.285 103.245 153.615 ;
        RECT 103.415 153.285 103.725 153.615 ;
        RECT 103.415 153.115 103.585 153.285 ;
        RECT 100.585 152.375 100.875 153.100 ;
        RECT 101.220 152.945 103.585 153.115 ;
        RECT 103.895 153.100 104.085 153.865 ;
        RECT 101.375 152.375 101.705 152.775 ;
        RECT 101.875 152.605 102.205 152.945 ;
        RECT 103.255 152.375 103.585 152.775 ;
        RECT 103.755 152.590 104.085 153.100 ;
        RECT 104.275 153.865 104.605 154.715 ;
        RECT 104.275 153.100 104.465 153.865 ;
        RECT 104.775 153.785 105.025 154.925 ;
        RECT 105.215 154.285 105.465 154.705 ;
        RECT 105.695 154.455 106.025 154.925 ;
        RECT 106.255 154.285 106.505 154.705 ;
        RECT 105.215 154.115 106.505 154.285 ;
        RECT 106.685 154.285 107.015 154.715 ;
        RECT 106.685 154.115 107.140 154.285 ;
        RECT 105.205 153.615 105.420 153.945 ;
        RECT 104.635 153.285 104.945 153.615 ;
        RECT 105.115 153.285 105.420 153.615 ;
        RECT 105.595 153.285 105.880 153.945 ;
        RECT 106.075 153.285 106.340 153.945 ;
        RECT 106.555 153.285 106.800 153.945 ;
        RECT 104.775 153.115 104.945 153.285 ;
        RECT 106.970 153.115 107.140 154.115 ;
        RECT 107.670 153.955 108.060 154.130 ;
        RECT 108.545 154.125 108.875 154.925 ;
        RECT 109.045 154.135 109.580 154.755 ;
        RECT 107.670 153.785 109.095 153.955 ;
        RECT 104.275 152.590 104.605 153.100 ;
        RECT 104.775 152.945 107.140 153.115 ;
        RECT 107.545 153.055 107.900 153.615 ;
        RECT 104.775 152.375 105.105 152.775 ;
        RECT 106.155 152.605 106.485 152.945 ;
        RECT 108.070 152.885 108.240 153.785 ;
        RECT 108.410 153.055 108.675 153.615 ;
        RECT 108.925 153.285 109.095 153.785 ;
        RECT 109.265 153.115 109.580 154.135 ;
        RECT 106.655 152.375 106.985 152.775 ;
        RECT 107.650 152.375 107.890 152.885 ;
        RECT 108.070 152.555 108.350 152.885 ;
        RECT 108.580 152.375 108.795 152.885 ;
        RECT 108.965 152.545 109.580 153.115 ;
        RECT 109.795 153.865 110.125 154.715 ;
        RECT 109.795 153.100 109.985 153.865 ;
        RECT 110.295 153.785 110.545 154.925 ;
        RECT 110.735 154.285 110.985 154.705 ;
        RECT 111.215 154.455 111.545 154.925 ;
        RECT 111.775 154.285 112.025 154.705 ;
        RECT 110.735 154.115 112.025 154.285 ;
        RECT 112.205 154.285 112.535 154.715 ;
        RECT 112.205 154.115 112.660 154.285 ;
        RECT 110.725 153.615 110.940 153.945 ;
        RECT 110.155 153.285 110.465 153.615 ;
        RECT 110.635 153.285 110.940 153.615 ;
        RECT 111.115 153.285 111.400 153.945 ;
        RECT 111.595 153.285 111.860 153.945 ;
        RECT 112.075 153.285 112.320 153.945 ;
        RECT 110.295 153.115 110.465 153.285 ;
        RECT 112.490 153.115 112.660 154.115 ;
        RECT 109.795 152.590 110.125 153.100 ;
        RECT 110.295 152.945 112.660 153.115 ;
        RECT 113.015 153.865 113.345 154.715 ;
        RECT 113.015 153.100 113.205 153.865 ;
        RECT 113.515 153.785 113.765 154.925 ;
        RECT 113.955 154.285 114.205 154.705 ;
        RECT 114.435 154.455 114.765 154.925 ;
        RECT 114.995 154.285 115.245 154.705 ;
        RECT 113.955 154.115 115.245 154.285 ;
        RECT 115.425 154.285 115.755 154.715 ;
        RECT 115.425 154.115 115.880 154.285 ;
        RECT 113.945 153.615 114.160 153.945 ;
        RECT 113.375 153.285 113.685 153.615 ;
        RECT 113.855 153.285 114.160 153.615 ;
        RECT 114.335 153.285 114.620 153.945 ;
        RECT 114.815 153.285 115.080 153.945 ;
        RECT 115.295 153.285 115.540 153.945 ;
        RECT 113.515 153.115 113.685 153.285 ;
        RECT 115.710 153.115 115.880 154.115 ;
        RECT 116.235 153.860 116.545 154.925 ;
        RECT 116.715 154.255 116.950 154.755 ;
        RECT 117.120 154.465 117.450 154.925 ;
        RECT 117.645 154.585 118.755 154.755 ;
        RECT 117.645 154.425 117.835 154.585 ;
        RECT 118.065 154.255 118.365 154.415 ;
        RECT 116.715 154.075 118.365 154.255 ;
        RECT 118.535 154.075 118.755 154.585 ;
        RECT 118.925 154.075 119.255 154.925 ;
        RECT 119.445 154.490 124.790 154.925 ;
        RECT 110.295 152.375 110.625 152.775 ;
        RECT 111.675 152.605 112.005 152.945 ;
        RECT 112.175 152.375 112.505 152.775 ;
        RECT 113.015 152.590 113.345 153.100 ;
        RECT 113.515 152.945 115.880 153.115 ;
        RECT 116.230 153.055 116.545 153.690 ;
        RECT 113.515 152.375 113.845 152.775 ;
        RECT 114.895 152.605 115.225 152.945 ;
        RECT 116.715 152.885 116.925 154.075 ;
        RECT 117.265 153.735 119.240 153.905 ;
        RECT 117.265 153.365 117.760 153.735 ;
        RECT 117.940 153.365 118.740 153.565 ;
        RECT 118.910 153.345 119.240 153.735 ;
        RECT 117.095 153.005 119.255 153.175 ;
        RECT 115.395 152.375 115.725 152.775 ;
        RECT 116.235 152.715 116.545 152.885 ;
        RECT 117.095 152.715 117.425 153.005 ;
        RECT 116.235 152.545 117.425 152.715 ;
        RECT 117.665 152.375 117.835 152.835 ;
        RECT 118.065 152.545 118.395 153.005 ;
        RECT 118.575 152.375 118.745 152.835 ;
        RECT 118.925 152.545 119.255 153.005 ;
        RECT 121.030 152.920 121.370 153.750 ;
        RECT 122.850 153.240 123.200 154.490 ;
        RECT 124.965 153.835 126.175 154.925 ;
        RECT 124.965 153.125 125.485 153.665 ;
        RECT 125.655 153.295 126.175 153.835 ;
        RECT 126.345 153.760 126.635 154.925 ;
        RECT 126.810 153.955 127.085 154.755 ;
        RECT 127.255 154.125 127.585 154.925 ;
        RECT 127.755 154.585 128.895 154.755 ;
        RECT 127.755 153.955 127.925 154.585 ;
        RECT 126.810 153.745 127.925 153.955 ;
        RECT 128.095 153.955 128.425 154.415 ;
        RECT 128.595 154.125 128.895 154.585 ;
        RECT 130.025 154.415 130.285 154.925 ;
        RECT 128.095 153.735 128.855 153.955 ;
        RECT 126.810 153.365 127.530 153.565 ;
        RECT 127.700 153.365 128.470 153.565 ;
        RECT 128.640 153.195 128.855 153.735 ;
        RECT 130.025 153.365 130.365 154.245 ;
        RECT 130.535 153.535 130.705 154.755 ;
        RECT 130.945 154.420 131.560 154.925 ;
        RECT 130.945 153.885 131.195 154.250 ;
        RECT 131.365 154.245 131.560 154.420 ;
        RECT 131.730 154.415 132.205 154.755 ;
        RECT 132.375 154.380 132.590 154.925 ;
        RECT 131.365 154.055 131.695 154.245 ;
        RECT 131.915 153.885 132.630 154.180 ;
        RECT 132.800 154.055 133.075 154.755 ;
        RECT 130.945 153.715 132.735 153.885 ;
        RECT 130.535 153.285 131.330 153.535 ;
        RECT 130.535 153.195 130.785 153.285 ;
        RECT 119.445 152.375 124.790 152.920 ;
        RECT 124.965 152.375 126.175 153.125 ;
        RECT 126.345 152.375 126.635 153.100 ;
        RECT 126.810 152.375 127.085 153.195 ;
        RECT 127.255 153.025 128.855 153.195 ;
        RECT 127.255 153.015 128.425 153.025 ;
        RECT 127.255 152.545 127.585 153.015 ;
        RECT 127.755 152.375 127.925 152.845 ;
        RECT 128.095 152.545 128.425 153.015 ;
        RECT 128.595 152.375 128.885 152.845 ;
        RECT 130.025 152.375 130.285 153.195 ;
        RECT 130.455 152.775 130.785 153.195 ;
        RECT 131.500 152.860 131.755 153.715 ;
        RECT 130.965 152.595 131.755 152.860 ;
        RECT 131.925 153.015 132.335 153.535 ;
        RECT 132.505 153.285 132.735 153.715 ;
        RECT 132.905 153.025 133.075 154.055 ;
        RECT 131.925 152.595 132.125 153.015 ;
        RECT 132.315 152.375 132.645 152.835 ;
        RECT 132.815 152.545 133.075 153.025 ;
        RECT 133.280 154.135 133.815 154.755 ;
        RECT 133.280 153.115 133.595 154.135 ;
        RECT 133.985 154.125 134.315 154.925 ;
        RECT 134.800 153.955 135.190 154.130 ;
        RECT 133.765 153.785 135.190 153.955 ;
        RECT 135.545 153.835 138.135 154.925 ;
        RECT 133.765 153.285 133.935 153.785 ;
        RECT 133.280 152.545 133.895 153.115 ;
        RECT 134.185 153.055 134.450 153.615 ;
        RECT 134.620 152.885 134.790 153.785 ;
        RECT 134.960 153.055 135.315 153.615 ;
        RECT 135.545 153.145 136.755 153.665 ;
        RECT 136.925 153.315 138.135 153.835 ;
        RECT 138.855 153.995 139.025 154.755 ;
        RECT 139.205 154.165 139.535 154.925 ;
        RECT 138.855 153.825 139.520 153.995 ;
        RECT 139.705 153.850 139.975 154.755 ;
        RECT 140.145 154.490 145.490 154.925 ;
        RECT 139.350 153.680 139.520 153.825 ;
        RECT 138.785 153.275 139.115 153.645 ;
        RECT 139.350 153.350 139.635 153.680 ;
        RECT 134.065 152.375 134.280 152.885 ;
        RECT 134.510 152.555 134.790 152.885 ;
        RECT 134.970 152.375 135.210 152.885 ;
        RECT 135.545 152.375 138.135 153.145 ;
        RECT 139.350 153.095 139.520 153.350 ;
        RECT 138.855 152.925 139.520 153.095 ;
        RECT 139.805 153.050 139.975 153.850 ;
        RECT 138.855 152.545 139.025 152.925 ;
        RECT 139.205 152.375 139.535 152.755 ;
        RECT 139.715 152.545 139.975 153.050 ;
        RECT 141.730 152.920 142.070 153.750 ;
        RECT 143.550 153.240 143.900 154.490 ;
        RECT 145.665 153.835 148.255 154.925 ;
        RECT 145.665 153.145 146.875 153.665 ;
        RECT 147.045 153.315 148.255 153.835 ;
        RECT 148.885 153.835 150.095 154.925 ;
        RECT 148.885 153.295 149.405 153.835 ;
        RECT 140.145 152.375 145.490 152.920 ;
        RECT 145.665 152.375 148.255 153.145 ;
        RECT 149.575 153.125 150.095 153.665 ;
        RECT 148.885 152.375 150.095 153.125 ;
        RECT 36.100 152.205 150.180 152.375 ;
        RECT 36.185 151.455 37.395 152.205 ;
        RECT 37.565 151.455 38.775 152.205 ;
        RECT 39.035 151.655 39.205 151.945 ;
        RECT 39.375 151.825 39.705 152.205 ;
        RECT 39.035 151.485 39.700 151.655 ;
        RECT 36.185 150.915 36.705 151.455 ;
        RECT 36.875 150.745 37.395 151.285 ;
        RECT 37.565 150.915 38.085 151.455 ;
        RECT 38.255 150.745 38.775 151.285 ;
        RECT 36.185 149.655 37.395 150.745 ;
        RECT 37.565 149.655 38.775 150.745 ;
        RECT 38.950 150.665 39.300 151.315 ;
        RECT 39.470 150.495 39.700 151.485 ;
        RECT 39.035 150.325 39.700 150.495 ;
        RECT 39.035 149.825 39.205 150.325 ;
        RECT 39.375 149.655 39.705 150.155 ;
        RECT 39.875 149.825 40.060 151.945 ;
        RECT 40.315 151.745 40.565 152.205 ;
        RECT 40.735 151.755 41.070 151.925 ;
        RECT 41.265 151.755 41.940 151.925 ;
        RECT 40.735 151.615 40.905 151.755 ;
        RECT 40.230 150.625 40.510 151.575 ;
        RECT 40.680 151.485 40.905 151.615 ;
        RECT 40.680 150.380 40.850 151.485 ;
        RECT 41.075 151.335 41.600 151.555 ;
        RECT 41.020 150.570 41.260 151.165 ;
        RECT 41.430 150.635 41.600 151.335 ;
        RECT 41.770 150.975 41.940 151.755 ;
        RECT 42.260 151.705 42.630 152.205 ;
        RECT 42.810 151.755 43.215 151.925 ;
        RECT 43.385 151.755 44.170 151.925 ;
        RECT 42.810 151.525 42.980 151.755 ;
        RECT 42.150 151.225 42.980 151.525 ;
        RECT 43.365 151.255 43.830 151.585 ;
        RECT 42.150 151.195 42.350 151.225 ;
        RECT 42.470 150.975 42.640 151.045 ;
        RECT 41.770 150.805 42.640 150.975 ;
        RECT 42.130 150.715 42.640 150.805 ;
        RECT 40.680 150.250 40.985 150.380 ;
        RECT 41.430 150.270 41.960 150.635 ;
        RECT 40.300 149.655 40.565 150.115 ;
        RECT 40.735 149.825 40.985 150.250 ;
        RECT 42.130 150.100 42.300 150.715 ;
        RECT 41.195 149.930 42.300 150.100 ;
        RECT 42.470 149.655 42.640 150.455 ;
        RECT 42.810 150.155 42.980 151.225 ;
        RECT 43.150 150.325 43.340 151.045 ;
        RECT 43.510 150.295 43.830 151.255 ;
        RECT 44.000 151.295 44.170 151.755 ;
        RECT 44.445 151.675 44.655 152.205 ;
        RECT 44.915 151.465 45.245 151.990 ;
        RECT 45.415 151.595 45.585 152.205 ;
        RECT 45.755 151.550 46.085 151.985 ;
        RECT 46.255 151.690 46.425 152.205 ;
        RECT 47.685 151.635 48.120 152.035 ;
        RECT 48.290 151.805 48.675 152.205 ;
        RECT 45.755 151.465 46.135 151.550 ;
        RECT 47.685 151.465 48.675 151.635 ;
        RECT 48.845 151.465 49.270 152.035 ;
        RECT 49.460 151.635 49.715 152.035 ;
        RECT 49.885 151.805 50.270 152.205 ;
        RECT 49.460 151.465 50.270 151.635 ;
        RECT 50.440 151.465 50.685 152.035 ;
        RECT 50.875 151.635 51.130 152.035 ;
        RECT 51.300 151.805 51.685 152.205 ;
        RECT 50.875 151.465 51.685 151.635 ;
        RECT 51.855 151.465 52.115 152.035 ;
        RECT 45.045 151.295 45.245 151.465 ;
        RECT 45.910 151.425 46.135 151.465 ;
        RECT 44.000 150.965 44.875 151.295 ;
        RECT 45.045 150.965 45.795 151.295 ;
        RECT 42.810 149.825 43.060 150.155 ;
        RECT 44.000 150.125 44.170 150.965 ;
        RECT 45.045 150.760 45.235 150.965 ;
        RECT 45.965 150.845 46.135 151.425 ;
        RECT 48.340 151.295 48.675 151.465 ;
        RECT 48.920 151.295 49.270 151.465 ;
        RECT 49.920 151.295 50.270 151.465 ;
        RECT 50.515 151.295 50.685 151.465 ;
        RECT 51.335 151.295 51.685 151.465 ;
        RECT 45.920 150.795 46.135 150.845 ;
        RECT 44.340 150.385 45.235 150.760 ;
        RECT 45.745 150.715 46.135 150.795 ;
        RECT 43.285 149.955 44.170 150.125 ;
        RECT 44.350 149.655 44.665 150.155 ;
        RECT 44.895 149.825 45.235 150.385 ;
        RECT 45.405 149.655 45.575 150.665 ;
        RECT 45.745 149.870 46.075 150.715 ;
        RECT 47.685 150.590 48.170 151.295 ;
        RECT 48.340 150.965 48.750 151.295 ;
        RECT 46.245 149.655 46.415 150.570 ;
        RECT 48.340 150.420 48.675 150.965 ;
        RECT 48.920 150.795 49.750 151.295 ;
        RECT 47.685 150.250 48.675 150.420 ;
        RECT 48.845 150.615 49.750 150.795 ;
        RECT 49.920 150.965 50.345 151.295 ;
        RECT 47.685 149.825 48.120 150.250 ;
        RECT 48.290 149.655 48.675 150.080 ;
        RECT 48.845 149.825 49.270 150.615 ;
        RECT 49.920 150.445 50.270 150.965 ;
        RECT 50.515 150.795 51.165 151.295 ;
        RECT 49.440 150.250 50.270 150.445 ;
        RECT 50.440 150.615 51.165 150.795 ;
        RECT 51.335 150.965 51.760 151.295 ;
        RECT 49.440 149.825 49.715 150.250 ;
        RECT 49.885 149.655 50.270 150.080 ;
        RECT 50.440 149.825 50.685 150.615 ;
        RECT 51.335 150.445 51.685 150.965 ;
        RECT 51.930 150.795 52.115 151.465 ;
        RECT 50.875 150.250 51.685 150.445 ;
        RECT 50.875 149.825 51.130 150.250 ;
        RECT 51.300 149.655 51.685 150.080 ;
        RECT 51.855 149.825 52.115 150.795 ;
        RECT 52.285 151.530 52.545 152.035 ;
        RECT 52.725 151.825 53.055 152.205 ;
        RECT 53.235 151.655 53.405 152.035 ;
        RECT 52.285 150.730 52.455 151.530 ;
        RECT 52.740 151.485 53.405 151.655 ;
        RECT 52.740 151.230 52.910 151.485 ;
        RECT 53.665 151.435 55.335 152.205 ;
        RECT 55.505 151.635 55.940 152.035 ;
        RECT 56.110 151.805 56.495 152.205 ;
        RECT 55.505 151.465 56.495 151.635 ;
        RECT 56.665 151.465 57.090 152.035 ;
        RECT 57.280 151.635 57.535 152.035 ;
        RECT 57.705 151.805 58.090 152.205 ;
        RECT 57.280 151.465 58.090 151.635 ;
        RECT 58.260 151.465 58.505 152.035 ;
        RECT 58.695 151.635 58.950 152.035 ;
        RECT 59.120 151.805 59.505 152.205 ;
        RECT 58.695 151.465 59.505 151.635 ;
        RECT 59.675 151.465 59.935 152.035 ;
        RECT 52.625 150.900 52.910 151.230 ;
        RECT 53.145 150.935 53.475 151.305 ;
        RECT 53.665 150.915 54.415 151.435 ;
        RECT 56.160 151.295 56.495 151.465 ;
        RECT 56.740 151.295 57.090 151.465 ;
        RECT 57.740 151.295 58.090 151.465 ;
        RECT 58.335 151.295 58.505 151.465 ;
        RECT 59.155 151.295 59.505 151.465 ;
        RECT 52.740 150.755 52.910 150.900 ;
        RECT 52.285 149.825 52.555 150.730 ;
        RECT 52.740 150.585 53.405 150.755 ;
        RECT 54.585 150.745 55.335 151.265 ;
        RECT 52.725 149.655 53.055 150.415 ;
        RECT 53.235 149.825 53.405 150.585 ;
        RECT 53.665 149.655 55.335 150.745 ;
        RECT 55.505 150.590 55.990 151.295 ;
        RECT 56.160 150.965 56.570 151.295 ;
        RECT 56.160 150.420 56.495 150.965 ;
        RECT 56.740 150.795 57.570 151.295 ;
        RECT 55.505 150.250 56.495 150.420 ;
        RECT 56.665 150.615 57.570 150.795 ;
        RECT 57.740 150.965 58.165 151.295 ;
        RECT 55.505 149.825 55.940 150.250 ;
        RECT 56.110 149.655 56.495 150.080 ;
        RECT 56.665 149.825 57.090 150.615 ;
        RECT 57.740 150.445 58.090 150.965 ;
        RECT 58.335 150.795 58.985 151.295 ;
        RECT 57.260 150.250 58.090 150.445 ;
        RECT 58.260 150.615 58.985 150.795 ;
        RECT 59.155 150.965 59.580 151.295 ;
        RECT 57.260 149.825 57.535 150.250 ;
        RECT 57.705 149.655 58.090 150.080 ;
        RECT 58.260 149.825 58.505 150.615 ;
        RECT 59.155 150.445 59.505 150.965 ;
        RECT 59.750 150.795 59.935 151.465 ;
        RECT 60.105 151.435 61.775 152.205 ;
        RECT 61.945 151.480 62.235 152.205 ;
        RECT 62.405 151.660 67.750 152.205 ;
        RECT 67.925 151.660 73.270 152.205 ;
        RECT 73.445 151.660 78.790 152.205 ;
        RECT 60.105 150.915 60.855 151.435 ;
        RECT 58.695 150.250 59.505 150.445 ;
        RECT 58.695 149.825 58.950 150.250 ;
        RECT 59.120 149.655 59.505 150.080 ;
        RECT 59.675 149.825 59.935 150.795 ;
        RECT 61.025 150.745 61.775 151.265 ;
        RECT 63.990 150.830 64.330 151.660 ;
        RECT 60.105 149.655 61.775 150.745 ;
        RECT 61.945 149.655 62.235 150.820 ;
        RECT 65.810 150.090 66.160 151.340 ;
        RECT 69.510 150.830 69.850 151.660 ;
        RECT 71.330 150.090 71.680 151.340 ;
        RECT 75.030 150.830 75.370 151.660 ;
        RECT 78.965 151.435 80.635 152.205 ;
        RECT 80.810 151.715 81.065 152.205 ;
        RECT 81.235 151.695 82.465 152.035 ;
        RECT 76.850 150.090 77.200 151.340 ;
        RECT 78.965 150.915 79.715 151.435 ;
        RECT 79.885 150.745 80.635 151.265 ;
        RECT 80.830 150.965 81.050 151.545 ;
        RECT 81.235 150.795 81.415 151.695 ;
        RECT 81.585 150.965 81.960 151.525 ;
        RECT 82.135 151.465 82.465 151.695 ;
        RECT 83.105 151.405 83.415 152.205 ;
        RECT 83.620 151.405 84.315 152.035 ;
        RECT 82.165 150.965 82.475 151.295 ;
        RECT 83.115 150.965 83.450 151.235 ;
        RECT 83.620 150.805 83.790 151.405 ;
        RECT 84.525 151.385 84.755 152.205 ;
        RECT 84.925 151.405 85.255 152.035 ;
        RECT 83.960 150.965 84.295 151.215 ;
        RECT 84.505 150.965 84.835 151.215 ;
        RECT 85.005 150.805 85.255 151.405 ;
        RECT 85.425 151.385 85.635 152.205 ;
        RECT 85.865 151.435 87.535 152.205 ;
        RECT 87.705 151.480 87.995 152.205 ;
        RECT 88.495 151.805 88.825 152.205 ;
        RECT 88.995 151.635 89.325 151.975 ;
        RECT 90.375 151.805 90.705 152.205 ;
        RECT 88.340 151.465 90.705 151.635 ;
        RECT 90.875 151.480 91.205 151.990 ;
        RECT 85.865 150.915 86.615 151.435 ;
        RECT 62.405 149.655 67.750 150.090 ;
        RECT 67.925 149.655 73.270 150.090 ;
        RECT 73.445 149.655 78.790 150.090 ;
        RECT 78.965 149.655 80.635 150.745 ;
        RECT 80.810 149.655 81.065 150.795 ;
        RECT 81.235 150.625 82.465 150.795 ;
        RECT 81.235 149.825 81.565 150.625 ;
        RECT 81.735 149.655 81.965 150.455 ;
        RECT 82.135 149.825 82.465 150.625 ;
        RECT 83.105 149.655 83.385 150.795 ;
        RECT 83.555 149.825 83.885 150.805 ;
        RECT 84.055 149.655 84.315 150.795 ;
        RECT 84.525 149.655 84.755 150.795 ;
        RECT 84.925 149.825 85.255 150.805 ;
        RECT 85.425 149.655 85.635 150.795 ;
        RECT 86.785 150.745 87.535 151.265 ;
        RECT 85.865 149.655 87.535 150.745 ;
        RECT 87.705 149.655 87.995 150.820 ;
        RECT 88.340 150.465 88.510 151.465 ;
        RECT 90.535 151.295 90.705 151.465 ;
        RECT 88.680 150.635 88.925 151.295 ;
        RECT 89.140 150.635 89.405 151.295 ;
        RECT 89.600 150.635 89.885 151.295 ;
        RECT 90.060 150.965 90.365 151.295 ;
        RECT 90.535 150.965 90.845 151.295 ;
        RECT 90.060 150.635 90.275 150.965 ;
        RECT 88.340 150.295 88.795 150.465 ;
        RECT 88.465 149.865 88.795 150.295 ;
        RECT 88.975 150.295 90.265 150.465 ;
        RECT 88.975 149.875 89.225 150.295 ;
        RECT 89.455 149.655 89.785 150.125 ;
        RECT 90.015 149.875 90.265 150.295 ;
        RECT 90.455 149.655 90.705 150.795 ;
        RECT 91.015 150.715 91.205 151.480 ;
        RECT 91.385 151.635 91.820 152.035 ;
        RECT 91.990 151.805 92.375 152.205 ;
        RECT 91.385 151.465 92.375 151.635 ;
        RECT 92.545 151.465 92.970 152.035 ;
        RECT 93.160 151.635 93.415 152.035 ;
        RECT 93.585 151.805 93.970 152.205 ;
        RECT 93.160 151.465 93.970 151.635 ;
        RECT 94.140 151.465 94.385 152.035 ;
        RECT 94.575 151.635 94.830 152.035 ;
        RECT 95.000 151.805 95.385 152.205 ;
        RECT 94.575 151.465 95.385 151.635 ;
        RECT 95.555 151.465 95.815 152.035 ;
        RECT 92.040 151.295 92.375 151.465 ;
        RECT 92.620 151.295 92.970 151.465 ;
        RECT 93.620 151.295 93.970 151.465 ;
        RECT 94.215 151.295 94.385 151.465 ;
        RECT 95.035 151.295 95.385 151.465 ;
        RECT 90.875 149.865 91.205 150.715 ;
        RECT 91.385 150.590 91.870 151.295 ;
        RECT 92.040 150.965 92.450 151.295 ;
        RECT 92.040 150.420 92.375 150.965 ;
        RECT 92.620 150.795 93.450 151.295 ;
        RECT 91.385 150.250 92.375 150.420 ;
        RECT 92.545 150.615 93.450 150.795 ;
        RECT 93.620 150.965 94.045 151.295 ;
        RECT 91.385 149.825 91.820 150.250 ;
        RECT 91.990 149.655 92.375 150.080 ;
        RECT 92.545 149.825 92.970 150.615 ;
        RECT 93.620 150.445 93.970 150.965 ;
        RECT 94.215 150.795 94.865 151.295 ;
        RECT 93.140 150.250 93.970 150.445 ;
        RECT 94.140 150.615 94.865 150.795 ;
        RECT 95.035 150.965 95.460 151.295 ;
        RECT 93.140 149.825 93.415 150.250 ;
        RECT 93.585 149.655 93.970 150.080 ;
        RECT 94.140 149.825 94.385 150.615 ;
        RECT 95.035 150.445 95.385 150.965 ;
        RECT 95.630 150.795 95.815 151.465 ;
        RECT 95.985 151.435 97.655 152.205 ;
        RECT 98.285 151.530 98.545 152.035 ;
        RECT 98.725 151.825 99.055 152.205 ;
        RECT 99.235 151.655 99.405 152.035 ;
        RECT 95.985 150.915 96.735 151.435 ;
        RECT 94.575 150.250 95.385 150.445 ;
        RECT 94.575 149.825 94.830 150.250 ;
        RECT 95.000 149.655 95.385 150.080 ;
        RECT 95.555 149.825 95.815 150.795 ;
        RECT 96.905 150.745 97.655 151.265 ;
        RECT 95.985 149.655 97.655 150.745 ;
        RECT 98.285 150.730 98.465 151.530 ;
        RECT 98.740 151.485 99.405 151.655 ;
        RECT 98.740 151.230 98.910 151.485 ;
        RECT 99.665 151.455 100.875 152.205 ;
        RECT 101.050 151.700 101.385 152.205 ;
        RECT 101.555 151.635 101.795 152.010 ;
        RECT 102.075 151.875 102.245 152.020 ;
        RECT 102.075 151.680 102.450 151.875 ;
        RECT 102.810 151.710 103.205 152.205 ;
        RECT 98.635 150.900 98.910 151.230 ;
        RECT 99.135 150.935 99.475 151.305 ;
        RECT 99.665 150.915 100.185 151.455 ;
        RECT 98.740 150.755 98.910 150.900 ;
        RECT 98.285 149.825 98.555 150.730 ;
        RECT 98.740 150.585 99.415 150.755 ;
        RECT 100.355 150.745 100.875 151.285 ;
        RECT 98.725 149.655 99.055 150.415 ;
        RECT 99.235 149.825 99.415 150.585 ;
        RECT 99.665 149.655 100.875 150.745 ;
        RECT 101.105 150.675 101.405 151.525 ;
        RECT 101.575 151.485 101.795 151.635 ;
        RECT 101.575 151.155 102.110 151.485 ;
        RECT 102.280 151.345 102.450 151.680 ;
        RECT 103.375 151.515 103.615 152.035 ;
        RECT 101.575 150.505 101.810 151.155 ;
        RECT 102.280 150.985 103.265 151.345 ;
        RECT 101.135 150.275 101.810 150.505 ;
        RECT 101.980 150.965 103.265 150.985 ;
        RECT 101.980 150.815 102.840 150.965 ;
        RECT 103.440 150.845 103.615 151.515 ;
        RECT 101.135 149.845 101.305 150.275 ;
        RECT 101.475 149.655 101.805 150.105 ;
        RECT 101.980 149.870 102.265 150.815 ;
        RECT 103.405 150.710 103.615 150.845 ;
        RECT 102.440 150.335 103.135 150.645 ;
        RECT 102.445 149.655 103.130 150.125 ;
        RECT 103.310 149.925 103.615 150.710 ;
        RECT 103.805 151.530 104.065 152.035 ;
        RECT 104.245 151.825 104.575 152.205 ;
        RECT 104.755 151.655 104.925 152.035 ;
        RECT 105.185 151.660 110.530 152.205 ;
        RECT 103.805 150.730 103.985 151.530 ;
        RECT 104.260 151.485 104.925 151.655 ;
        RECT 104.260 151.230 104.430 151.485 ;
        RECT 104.155 150.900 104.430 151.230 ;
        RECT 104.655 150.935 104.995 151.305 ;
        RECT 104.260 150.755 104.430 150.900 ;
        RECT 106.770 150.830 107.110 151.660 ;
        RECT 110.705 151.435 113.295 152.205 ;
        RECT 113.465 151.480 113.755 152.205 ;
        RECT 103.805 149.825 104.075 150.730 ;
        RECT 104.260 150.585 104.935 150.755 ;
        RECT 104.245 149.655 104.575 150.415 ;
        RECT 104.755 149.825 104.935 150.585 ;
        RECT 108.590 150.090 108.940 151.340 ;
        RECT 110.705 150.915 111.915 151.435 ;
        RECT 112.085 150.745 113.295 151.265 ;
        RECT 113.925 151.220 114.195 152.035 ;
        RECT 114.365 151.465 115.035 152.205 ;
        RECT 115.205 151.635 115.500 151.980 ;
        RECT 115.680 151.805 116.055 152.205 ;
        RECT 116.270 151.635 116.600 151.980 ;
        RECT 115.205 151.465 116.600 151.635 ;
        RECT 116.850 151.465 117.435 152.035 ;
        RECT 117.605 151.660 122.950 152.205 ;
        RECT 105.185 149.655 110.530 150.090 ;
        RECT 110.705 149.655 113.295 150.745 ;
        RECT 113.465 149.655 113.755 150.820 ;
        RECT 113.925 149.825 114.275 151.220 ;
        RECT 114.445 150.795 114.615 151.295 ;
        RECT 114.785 150.965 115.120 151.295 ;
        RECT 115.290 150.965 115.630 151.295 ;
        RECT 114.445 150.625 115.190 150.795 ;
        RECT 114.445 149.655 114.850 150.455 ;
        RECT 115.020 149.995 115.190 150.625 ;
        RECT 115.360 150.220 115.630 150.965 ;
        RECT 115.820 150.965 116.110 151.295 ;
        RECT 116.280 150.965 116.680 151.295 ;
        RECT 115.820 150.220 116.055 150.965 ;
        RECT 116.850 150.795 117.020 151.465 ;
        RECT 117.190 150.965 117.435 151.295 ;
        RECT 119.190 150.830 119.530 151.660 ;
        RECT 123.125 151.455 124.335 152.205 ;
        RECT 116.225 150.625 117.435 150.795 ;
        RECT 116.225 149.995 116.555 150.625 ;
        RECT 115.020 149.825 116.555 149.995 ;
        RECT 116.740 149.655 116.975 150.455 ;
        RECT 117.145 149.825 117.435 150.625 ;
        RECT 121.010 150.090 121.360 151.340 ;
        RECT 123.125 150.915 123.645 151.455 ;
        RECT 124.545 151.385 124.775 152.205 ;
        RECT 124.945 151.405 125.275 152.035 ;
        RECT 123.815 150.745 124.335 151.285 ;
        RECT 124.525 150.965 124.855 151.215 ;
        RECT 125.025 150.805 125.275 151.405 ;
        RECT 125.445 151.385 125.655 152.205 ;
        RECT 125.885 151.435 127.555 152.205 ;
        RECT 127.925 151.575 128.255 151.935 ;
        RECT 128.875 151.745 129.125 152.205 ;
        RECT 129.295 151.745 129.855 152.035 ;
        RECT 125.885 150.915 126.635 151.435 ;
        RECT 127.925 151.385 129.315 151.575 ;
        RECT 129.145 151.295 129.315 151.385 ;
        RECT 117.605 149.655 122.950 150.090 ;
        RECT 123.125 149.655 124.335 150.745 ;
        RECT 124.545 149.655 124.775 150.795 ;
        RECT 124.945 149.825 125.275 150.805 ;
        RECT 125.445 149.655 125.655 150.795 ;
        RECT 126.805 150.745 127.555 151.265 ;
        RECT 125.885 149.655 127.555 150.745 ;
        RECT 127.740 150.965 128.415 151.215 ;
        RECT 128.635 150.965 128.975 151.215 ;
        RECT 129.145 150.965 129.435 151.295 ;
        RECT 127.740 150.605 128.005 150.965 ;
        RECT 129.145 150.715 129.315 150.965 ;
        RECT 128.375 150.545 129.315 150.715 ;
        RECT 127.925 149.655 128.205 150.325 ;
        RECT 128.375 149.995 128.675 150.545 ;
        RECT 129.605 150.375 129.855 151.745 ;
        RECT 130.030 151.675 130.320 152.025 ;
        RECT 130.515 151.845 130.845 152.205 ;
        RECT 131.015 151.675 131.245 151.980 ;
        RECT 130.030 151.505 131.245 151.675 ;
        RECT 131.435 151.525 131.605 151.900 ;
        RECT 131.435 151.355 131.635 151.525 ;
        RECT 131.875 151.395 132.145 152.205 ;
        RECT 132.315 151.395 132.645 152.035 ;
        RECT 132.815 151.395 133.055 152.205 ;
        RECT 133.245 151.660 138.590 152.205 ;
        RECT 131.435 151.335 131.605 151.355 ;
        RECT 130.090 151.185 130.350 151.295 ;
        RECT 130.085 151.015 130.350 151.185 ;
        RECT 130.090 150.965 130.350 151.015 ;
        RECT 130.530 150.965 130.915 151.295 ;
        RECT 131.085 151.165 131.605 151.335 ;
        RECT 128.875 149.655 129.205 150.375 ;
        RECT 129.395 149.825 129.855 150.375 ;
        RECT 130.030 149.655 130.350 150.795 ;
        RECT 130.530 149.915 130.725 150.965 ;
        RECT 131.085 150.785 131.255 151.165 ;
        RECT 130.905 150.505 131.255 150.785 ;
        RECT 131.445 150.635 131.690 150.995 ;
        RECT 131.865 150.965 132.215 151.215 ;
        RECT 132.385 150.795 132.555 151.395 ;
        RECT 132.725 150.965 133.075 151.215 ;
        RECT 134.830 150.830 135.170 151.660 ;
        RECT 139.225 151.480 139.515 152.205 ;
        RECT 140.695 151.655 140.865 151.945 ;
        RECT 141.035 151.825 141.365 152.205 ;
        RECT 140.695 151.485 141.360 151.655 ;
        RECT 130.905 149.825 131.235 150.505 ;
        RECT 131.435 149.655 131.690 150.455 ;
        RECT 131.875 149.655 132.205 150.795 ;
        RECT 132.385 150.625 133.065 150.795 ;
        RECT 132.735 149.840 133.065 150.625 ;
        RECT 136.650 150.090 137.000 151.340 ;
        RECT 133.245 149.655 138.590 150.090 ;
        RECT 139.225 149.655 139.515 150.820 ;
        RECT 140.610 150.665 140.960 151.315 ;
        RECT 141.130 150.495 141.360 151.485 ;
        RECT 140.695 150.325 141.360 150.495 ;
        RECT 140.695 149.825 140.865 150.325 ;
        RECT 141.035 149.655 141.365 150.155 ;
        RECT 141.535 149.825 141.720 151.945 ;
        RECT 141.975 151.745 142.225 152.205 ;
        RECT 142.395 151.755 142.730 151.925 ;
        RECT 142.925 151.755 143.600 151.925 ;
        RECT 142.395 151.615 142.565 151.755 ;
        RECT 141.890 150.625 142.170 151.575 ;
        RECT 142.340 151.485 142.565 151.615 ;
        RECT 142.340 150.380 142.510 151.485 ;
        RECT 142.735 151.335 143.260 151.555 ;
        RECT 142.680 150.570 142.920 151.165 ;
        RECT 143.090 150.635 143.260 151.335 ;
        RECT 143.430 150.975 143.600 151.755 ;
        RECT 143.920 151.705 144.290 152.205 ;
        RECT 144.470 151.755 144.875 151.925 ;
        RECT 145.045 151.755 145.830 151.925 ;
        RECT 144.470 151.525 144.640 151.755 ;
        RECT 143.810 151.225 144.640 151.525 ;
        RECT 145.025 151.255 145.490 151.585 ;
        RECT 143.810 151.195 144.010 151.225 ;
        RECT 144.130 150.975 144.300 151.045 ;
        RECT 143.430 150.805 144.300 150.975 ;
        RECT 143.790 150.715 144.300 150.805 ;
        RECT 142.340 150.250 142.645 150.380 ;
        RECT 143.090 150.270 143.620 150.635 ;
        RECT 141.960 149.655 142.225 150.115 ;
        RECT 142.395 149.825 142.645 150.250 ;
        RECT 143.790 150.100 143.960 150.715 ;
        RECT 142.855 149.930 143.960 150.100 ;
        RECT 144.130 149.655 144.300 150.455 ;
        RECT 144.470 150.155 144.640 151.225 ;
        RECT 144.810 150.325 145.000 151.045 ;
        RECT 145.170 150.295 145.490 151.255 ;
        RECT 145.660 151.295 145.830 151.755 ;
        RECT 146.105 151.675 146.315 152.205 ;
        RECT 146.575 151.465 146.905 151.990 ;
        RECT 147.075 151.595 147.245 152.205 ;
        RECT 147.415 151.550 147.745 151.985 ;
        RECT 147.415 151.465 147.795 151.550 ;
        RECT 146.705 151.295 146.905 151.465 ;
        RECT 147.570 151.425 147.795 151.465 ;
        RECT 148.885 151.455 150.095 152.205 ;
        RECT 145.660 150.965 146.535 151.295 ;
        RECT 146.705 150.965 147.455 151.295 ;
        RECT 144.470 149.825 144.720 150.155 ;
        RECT 145.660 150.125 145.830 150.965 ;
        RECT 146.705 150.760 146.895 150.965 ;
        RECT 147.625 150.845 147.795 151.425 ;
        RECT 147.580 150.795 147.795 150.845 ;
        RECT 146.000 150.385 146.895 150.760 ;
        RECT 147.405 150.715 147.795 150.795 ;
        RECT 148.885 150.745 149.405 151.285 ;
        RECT 149.575 150.915 150.095 151.455 ;
        RECT 144.945 149.955 145.830 150.125 ;
        RECT 146.010 149.655 146.325 150.155 ;
        RECT 146.555 149.825 146.895 150.385 ;
        RECT 147.065 149.655 147.235 150.665 ;
        RECT 147.405 149.870 147.735 150.715 ;
        RECT 148.885 149.655 150.095 150.745 ;
        RECT 36.100 149.485 150.180 149.655 ;
        RECT 36.185 148.395 37.395 149.485 ;
        RECT 37.565 148.395 40.155 149.485 ;
        RECT 36.185 147.685 36.705 148.225 ;
        RECT 36.875 147.855 37.395 148.395 ;
        RECT 37.565 147.705 38.775 148.225 ;
        RECT 38.945 147.875 40.155 148.395 ;
        RECT 40.325 148.410 40.595 149.315 ;
        RECT 40.765 148.725 41.095 149.485 ;
        RECT 41.275 148.555 41.445 149.315 ;
        RECT 36.185 146.935 37.395 147.685 ;
        RECT 37.565 146.935 40.155 147.705 ;
        RECT 40.325 147.610 40.495 148.410 ;
        RECT 40.780 148.385 41.445 148.555 ;
        RECT 41.705 148.410 41.975 149.315 ;
        RECT 42.145 148.725 42.475 149.485 ;
        RECT 42.655 148.555 42.825 149.315 ;
        RECT 43.085 149.050 48.430 149.485 ;
        RECT 40.780 148.240 40.950 148.385 ;
        RECT 40.665 147.910 40.950 148.240 ;
        RECT 40.780 147.655 40.950 147.910 ;
        RECT 41.185 147.835 41.515 148.205 ;
        RECT 40.325 147.105 40.585 147.610 ;
        RECT 40.780 147.485 41.445 147.655 ;
        RECT 40.765 146.935 41.095 147.315 ;
        RECT 41.275 147.105 41.445 147.485 ;
        RECT 41.705 147.610 41.875 148.410 ;
        RECT 42.160 148.385 42.825 148.555 ;
        RECT 42.160 148.240 42.330 148.385 ;
        RECT 42.045 147.910 42.330 148.240 ;
        RECT 42.160 147.655 42.330 147.910 ;
        RECT 42.565 147.835 42.895 148.205 ;
        RECT 41.705 147.105 41.965 147.610 ;
        RECT 42.160 147.485 42.825 147.655 ;
        RECT 42.145 146.935 42.475 147.315 ;
        RECT 42.655 147.105 42.825 147.485 ;
        RECT 44.670 147.480 45.010 148.310 ;
        RECT 46.490 147.800 46.840 149.050 ;
        RECT 49.065 148.320 49.355 149.485 ;
        RECT 49.525 148.395 52.115 149.485 ;
        RECT 52.485 148.815 52.765 149.485 ;
        RECT 52.935 148.595 53.235 149.145 ;
        RECT 53.435 148.765 53.765 149.485 ;
        RECT 53.955 148.765 54.415 149.315 ;
        RECT 49.525 147.705 50.735 148.225 ;
        RECT 50.905 147.875 52.115 148.395 ;
        RECT 52.300 148.175 52.565 148.535 ;
        RECT 52.935 148.425 53.875 148.595 ;
        RECT 53.705 148.175 53.875 148.425 ;
        RECT 52.300 147.925 52.975 148.175 ;
        RECT 53.195 147.925 53.535 148.175 ;
        RECT 53.705 147.845 53.995 148.175 ;
        RECT 53.705 147.755 53.875 147.845 ;
        RECT 43.085 146.935 48.430 147.480 ;
        RECT 49.065 146.935 49.355 147.660 ;
        RECT 49.525 146.935 52.115 147.705 ;
        RECT 52.485 147.565 53.875 147.755 ;
        RECT 52.485 147.205 52.815 147.565 ;
        RECT 54.165 147.395 54.415 148.765 ;
        RECT 54.605 148.595 54.865 149.305 ;
        RECT 55.035 148.775 55.365 149.485 ;
        RECT 55.535 148.595 55.765 149.305 ;
        RECT 54.605 148.355 55.765 148.595 ;
        RECT 55.945 148.575 56.215 149.305 ;
        RECT 56.395 148.755 56.735 149.485 ;
        RECT 55.945 148.355 56.715 148.575 ;
        RECT 54.595 147.845 54.895 148.175 ;
        RECT 55.075 147.865 55.600 148.175 ;
        RECT 55.780 147.865 56.245 148.175 ;
        RECT 53.435 146.935 53.685 147.395 ;
        RECT 53.855 147.105 54.415 147.395 ;
        RECT 54.605 146.935 54.895 147.665 ;
        RECT 55.075 147.225 55.305 147.865 ;
        RECT 56.425 147.685 56.715 148.355 ;
        RECT 55.485 147.485 56.715 147.685 ;
        RECT 55.485 147.115 55.795 147.485 ;
        RECT 55.975 146.935 56.645 147.305 ;
        RECT 56.905 147.115 57.165 149.305 ;
        RECT 57.345 148.635 57.725 149.315 ;
        RECT 58.315 148.635 58.485 149.485 ;
        RECT 58.655 148.805 58.985 149.315 ;
        RECT 59.155 148.975 59.325 149.485 ;
        RECT 59.495 148.805 59.895 149.315 ;
        RECT 58.655 148.635 59.895 148.805 ;
        RECT 57.345 147.675 57.515 148.635 ;
        RECT 57.685 148.295 58.990 148.465 ;
        RECT 60.075 148.385 60.395 149.315 ;
        RECT 60.655 149.145 61.815 149.315 ;
        RECT 60.655 148.645 60.825 149.145 ;
        RECT 61.085 148.515 61.255 148.975 ;
        RECT 61.485 148.895 61.815 149.145 ;
        RECT 62.040 149.065 62.370 149.485 ;
        RECT 62.625 148.895 62.910 149.315 ;
        RECT 61.485 148.725 62.910 148.895 ;
        RECT 63.155 148.685 63.485 149.485 ;
        RECT 63.735 148.765 64.070 149.275 ;
        RECT 57.685 147.845 57.930 148.295 ;
        RECT 58.100 147.925 58.650 148.125 ;
        RECT 58.820 148.095 58.990 148.295 ;
        RECT 59.765 148.215 60.395 148.385 ;
        RECT 58.820 147.925 59.195 148.095 ;
        RECT 59.365 147.675 59.595 148.175 ;
        RECT 57.345 147.505 59.595 147.675 ;
        RECT 57.395 146.935 57.725 147.325 ;
        RECT 57.895 147.185 58.065 147.505 ;
        RECT 59.765 147.335 59.935 148.215 ;
        RECT 60.630 148.175 60.835 148.465 ;
        RECT 61.085 148.345 63.455 148.515 ;
        RECT 63.285 148.175 63.455 148.345 ;
        RECT 60.630 148.125 60.980 148.175 ;
        RECT 60.625 147.955 60.980 148.125 ;
        RECT 60.630 147.845 60.980 147.955 ;
        RECT 58.235 146.935 58.565 147.325 ;
        RECT 58.980 147.165 59.935 147.335 ;
        RECT 60.105 146.935 60.395 147.770 ;
        RECT 60.575 146.935 60.905 147.655 ;
        RECT 61.290 147.510 61.710 148.175 ;
        RECT 61.880 147.785 62.170 148.175 ;
        RECT 62.360 147.785 62.630 148.175 ;
        RECT 62.840 148.125 63.090 148.175 ;
        RECT 62.840 147.955 63.095 148.125 ;
        RECT 62.840 147.845 63.090 147.955 ;
        RECT 63.285 147.845 63.590 148.175 ;
        RECT 61.880 147.615 62.175 147.785 ;
        RECT 62.360 147.615 62.635 147.785 ;
        RECT 63.285 147.675 63.455 147.845 ;
        RECT 61.880 147.515 62.170 147.615 ;
        RECT 62.360 147.515 62.630 147.615 ;
        RECT 62.895 147.505 63.455 147.675 ;
        RECT 62.895 147.335 63.065 147.505 ;
        RECT 63.815 147.410 64.070 148.765 ;
        RECT 64.245 148.395 65.915 149.485 ;
        RECT 61.450 147.165 63.065 147.335 ;
        RECT 63.235 146.935 63.565 147.335 ;
        RECT 63.735 147.150 64.070 147.410 ;
        RECT 64.245 147.705 64.995 148.225 ;
        RECT 65.165 147.875 65.915 148.395 ;
        RECT 66.165 148.555 66.345 149.315 ;
        RECT 66.525 148.725 66.855 149.485 ;
        RECT 66.165 148.385 66.840 148.555 ;
        RECT 67.025 148.410 67.295 149.315 ;
        RECT 66.670 148.240 66.840 148.385 ;
        RECT 66.105 147.835 66.445 148.205 ;
        RECT 66.670 147.910 66.945 148.240 ;
        RECT 64.245 146.935 65.915 147.705 ;
        RECT 66.670 147.655 66.840 147.910 ;
        RECT 66.175 147.485 66.840 147.655 ;
        RECT 67.115 147.610 67.295 148.410 ;
        RECT 67.465 148.395 68.675 149.485 ;
        RECT 66.175 147.105 66.345 147.485 ;
        RECT 66.525 146.935 66.855 147.315 ;
        RECT 67.035 147.105 67.295 147.610 ;
        RECT 67.465 147.685 67.985 148.225 ;
        RECT 68.155 147.855 68.675 148.395 ;
        RECT 68.845 148.345 69.125 149.485 ;
        RECT 69.295 148.335 69.625 149.315 ;
        RECT 69.795 148.345 70.055 149.485 ;
        RECT 70.225 148.345 70.505 149.485 ;
        RECT 70.675 148.335 71.005 149.315 ;
        RECT 71.175 148.345 71.435 149.485 ;
        RECT 71.905 148.845 72.235 149.275 ;
        RECT 71.780 148.675 72.235 148.845 ;
        RECT 72.415 148.845 72.665 149.265 ;
        RECT 72.895 149.015 73.225 149.485 ;
        RECT 73.455 148.845 73.705 149.265 ;
        RECT 72.415 148.675 73.705 148.845 ;
        RECT 68.855 147.905 69.190 148.175 ;
        RECT 69.360 147.735 69.530 148.335 ;
        RECT 70.740 148.295 70.915 148.335 ;
        RECT 69.700 147.925 70.035 148.175 ;
        RECT 70.235 147.905 70.570 148.175 ;
        RECT 70.740 147.735 70.910 148.295 ;
        RECT 71.080 147.925 71.415 148.175 ;
        RECT 67.465 146.935 68.675 147.685 ;
        RECT 68.845 146.935 69.155 147.735 ;
        RECT 69.360 147.105 70.055 147.735 ;
        RECT 70.225 146.935 70.535 147.735 ;
        RECT 70.740 147.105 71.435 147.735 ;
        RECT 71.780 147.675 71.950 148.675 ;
        RECT 72.120 147.845 72.365 148.505 ;
        RECT 72.580 147.845 72.845 148.505 ;
        RECT 73.040 147.845 73.325 148.505 ;
        RECT 73.500 148.175 73.715 148.505 ;
        RECT 73.895 148.345 74.145 149.485 ;
        RECT 74.315 148.425 74.645 149.275 ;
        RECT 73.500 147.845 73.805 148.175 ;
        RECT 73.975 147.845 74.285 148.175 ;
        RECT 73.975 147.675 74.145 147.845 ;
        RECT 71.780 147.505 74.145 147.675 ;
        RECT 74.455 147.660 74.645 148.425 ;
        RECT 74.825 148.320 75.115 149.485 ;
        RECT 75.585 148.845 75.915 149.275 ;
        RECT 75.460 148.675 75.915 148.845 ;
        RECT 76.095 148.845 76.345 149.265 ;
        RECT 76.575 149.015 76.905 149.485 ;
        RECT 77.135 148.845 77.385 149.265 ;
        RECT 76.095 148.675 77.385 148.845 ;
        RECT 75.460 147.675 75.630 148.675 ;
        RECT 75.800 147.845 76.045 148.505 ;
        RECT 76.260 147.845 76.525 148.505 ;
        RECT 76.720 147.845 77.005 148.505 ;
        RECT 77.180 148.175 77.395 148.505 ;
        RECT 77.575 148.345 77.825 149.485 ;
        RECT 77.995 148.425 78.325 149.275 ;
        RECT 78.705 148.815 78.985 149.485 ;
        RECT 79.155 148.595 79.455 149.145 ;
        RECT 79.655 148.765 79.985 149.485 ;
        RECT 80.175 148.765 80.635 149.315 ;
        RECT 77.180 147.845 77.485 148.175 ;
        RECT 77.655 147.845 77.965 148.175 ;
        RECT 77.655 147.675 77.825 147.845 ;
        RECT 71.935 146.935 72.265 147.335 ;
        RECT 72.435 147.165 72.765 147.505 ;
        RECT 73.815 146.935 74.145 147.335 ;
        RECT 74.315 147.150 74.645 147.660 ;
        RECT 74.825 146.935 75.115 147.660 ;
        RECT 75.460 147.505 77.825 147.675 ;
        RECT 78.135 147.660 78.325 148.425 ;
        RECT 78.520 148.175 78.785 148.535 ;
        RECT 79.155 148.425 80.095 148.595 ;
        RECT 79.925 148.175 80.095 148.425 ;
        RECT 78.520 147.925 79.195 148.175 ;
        RECT 79.415 147.925 79.755 148.175 ;
        RECT 79.925 147.845 80.215 148.175 ;
        RECT 79.925 147.755 80.095 147.845 ;
        RECT 75.615 146.935 75.945 147.335 ;
        RECT 76.115 147.165 76.445 147.505 ;
        RECT 77.495 146.935 77.825 147.335 ;
        RECT 77.995 147.150 78.325 147.660 ;
        RECT 78.705 147.565 80.095 147.755 ;
        RECT 78.705 147.205 79.035 147.565 ;
        RECT 80.385 147.395 80.635 148.765 ;
        RECT 81.450 148.515 81.840 148.690 ;
        RECT 82.325 148.685 82.655 149.485 ;
        RECT 82.825 148.695 83.360 149.315 ;
        RECT 81.450 148.345 82.875 148.515 ;
        RECT 81.325 147.615 81.680 148.175 ;
        RECT 81.850 147.445 82.020 148.345 ;
        RECT 82.190 147.615 82.455 148.175 ;
        RECT 82.705 147.845 82.875 148.345 ;
        RECT 83.045 147.675 83.360 148.695 ;
        RECT 79.655 146.935 79.905 147.395 ;
        RECT 80.075 147.105 80.635 147.395 ;
        RECT 81.430 146.935 81.670 147.445 ;
        RECT 81.850 147.115 82.130 147.445 ;
        RECT 82.360 146.935 82.575 147.445 ;
        RECT 82.745 147.105 83.360 147.675 ;
        RECT 84.495 148.425 84.825 149.275 ;
        RECT 84.495 147.660 84.685 148.425 ;
        RECT 84.995 148.345 85.245 149.485 ;
        RECT 85.435 148.845 85.685 149.265 ;
        RECT 85.915 149.015 86.245 149.485 ;
        RECT 86.475 148.845 86.725 149.265 ;
        RECT 85.435 148.675 86.725 148.845 ;
        RECT 86.905 148.845 87.235 149.275 ;
        RECT 86.905 148.675 87.360 148.845 ;
        RECT 85.425 148.175 85.640 148.505 ;
        RECT 84.855 147.845 85.165 148.175 ;
        RECT 85.335 147.845 85.640 148.175 ;
        RECT 85.815 147.845 86.100 148.505 ;
        RECT 86.295 147.845 86.560 148.505 ;
        RECT 86.775 147.845 87.020 148.505 ;
        RECT 84.995 147.675 85.165 147.845 ;
        RECT 87.190 147.675 87.360 148.675 ;
        RECT 84.495 147.150 84.825 147.660 ;
        RECT 84.995 147.505 87.360 147.675 ;
        RECT 87.705 148.345 88.045 149.315 ;
        RECT 88.215 148.345 88.385 149.485 ;
        RECT 88.655 148.685 88.905 149.485 ;
        RECT 89.550 148.515 89.880 149.315 ;
        RECT 90.180 148.685 90.510 149.485 ;
        RECT 90.680 148.515 91.010 149.315 ;
        RECT 88.575 148.345 91.010 148.515 ;
        RECT 91.385 148.395 93.975 149.485 ;
        RECT 87.705 147.735 87.880 148.345 ;
        RECT 88.575 148.095 88.745 148.345 ;
        RECT 88.050 147.925 88.745 148.095 ;
        RECT 88.920 147.925 89.340 148.125 ;
        RECT 89.510 147.925 89.840 148.125 ;
        RECT 90.010 147.925 90.340 148.125 ;
        RECT 84.995 146.935 85.325 147.335 ;
        RECT 86.375 147.165 86.705 147.505 ;
        RECT 86.875 146.935 87.205 147.335 ;
        RECT 87.705 147.105 88.045 147.735 ;
        RECT 88.215 146.935 88.465 147.735 ;
        RECT 88.655 147.585 89.880 147.755 ;
        RECT 88.655 147.105 88.985 147.585 ;
        RECT 89.155 146.935 89.380 147.395 ;
        RECT 89.550 147.105 89.880 147.585 ;
        RECT 90.510 147.715 90.680 148.345 ;
        RECT 90.865 147.925 91.215 148.175 ;
        RECT 90.510 147.105 91.010 147.715 ;
        RECT 91.385 147.705 92.595 148.225 ;
        RECT 92.765 147.875 93.975 148.395 ;
        RECT 94.605 148.345 94.885 149.485 ;
        RECT 95.055 148.335 95.385 149.315 ;
        RECT 95.555 148.345 95.815 149.485 ;
        RECT 95.985 148.395 98.575 149.485 ;
        RECT 98.750 149.060 99.085 149.485 ;
        RECT 99.255 148.880 99.440 149.285 ;
        RECT 95.120 148.295 95.295 148.335 ;
        RECT 94.615 147.905 94.950 148.175 ;
        RECT 95.120 147.735 95.290 148.295 ;
        RECT 95.460 147.925 95.795 148.175 ;
        RECT 91.385 146.935 93.975 147.705 ;
        RECT 94.605 146.935 94.915 147.735 ;
        RECT 95.120 147.105 95.815 147.735 ;
        RECT 95.985 147.705 97.195 148.225 ;
        RECT 97.365 147.875 98.575 148.395 ;
        RECT 98.775 148.705 99.440 148.880 ;
        RECT 99.645 148.705 99.975 149.485 ;
        RECT 95.985 146.935 98.575 147.705 ;
        RECT 98.775 147.675 99.115 148.705 ;
        RECT 100.145 148.515 100.415 149.285 ;
        RECT 99.285 148.345 100.415 148.515 ;
        RECT 99.285 147.845 99.535 148.345 ;
        RECT 98.775 147.505 99.460 147.675 ;
        RECT 99.715 147.595 100.075 148.175 ;
        RECT 98.750 146.935 99.085 147.335 ;
        RECT 99.255 147.105 99.460 147.505 ;
        RECT 100.245 147.435 100.415 148.345 ;
        RECT 100.585 148.320 100.875 149.485 ;
        RECT 101.050 149.060 101.385 149.485 ;
        RECT 101.555 148.880 101.740 149.285 ;
        RECT 101.075 148.705 101.740 148.880 ;
        RECT 101.945 148.705 102.275 149.485 ;
        RECT 101.075 147.675 101.415 148.705 ;
        RECT 102.445 148.515 102.715 149.285 ;
        RECT 101.585 148.345 102.715 148.515 ;
        RECT 102.885 148.395 105.475 149.485 ;
        RECT 101.585 147.845 101.835 148.345 ;
        RECT 99.670 146.935 99.945 147.415 ;
        RECT 100.155 147.105 100.415 147.435 ;
        RECT 100.585 146.935 100.875 147.660 ;
        RECT 101.075 147.505 101.760 147.675 ;
        RECT 102.015 147.595 102.375 148.175 ;
        RECT 101.050 146.935 101.385 147.335 ;
        RECT 101.555 147.105 101.760 147.505 ;
        RECT 102.545 147.435 102.715 148.345 ;
        RECT 101.970 146.935 102.245 147.415 ;
        RECT 102.455 147.105 102.715 147.435 ;
        RECT 102.885 147.705 104.095 148.225 ;
        RECT 104.265 147.875 105.475 148.395 ;
        RECT 105.645 148.515 105.915 149.285 ;
        RECT 106.085 148.705 106.415 149.485 ;
        RECT 106.620 148.880 106.805 149.285 ;
        RECT 106.975 149.060 107.310 149.485 ;
        RECT 106.620 148.705 107.285 148.880 ;
        RECT 105.645 148.345 106.775 148.515 ;
        RECT 102.885 146.935 105.475 147.705 ;
        RECT 105.645 147.435 105.815 148.345 ;
        RECT 105.985 147.595 106.345 148.175 ;
        RECT 106.525 147.845 106.775 148.345 ;
        RECT 106.945 147.675 107.285 148.705 ;
        RECT 107.485 148.395 110.075 149.485 ;
        RECT 106.600 147.505 107.285 147.675 ;
        RECT 107.485 147.705 108.695 148.225 ;
        RECT 108.865 147.875 110.075 148.395 ;
        RECT 110.245 148.345 110.585 149.315 ;
        RECT 110.755 148.345 110.925 149.485 ;
        RECT 111.195 148.685 111.445 149.485 ;
        RECT 112.090 148.515 112.420 149.315 ;
        RECT 112.720 148.685 113.050 149.485 ;
        RECT 113.220 148.515 113.550 149.315 ;
        RECT 114.225 148.845 114.555 149.275 ;
        RECT 111.115 148.345 113.550 148.515 ;
        RECT 114.100 148.675 114.555 148.845 ;
        RECT 114.735 148.845 114.985 149.265 ;
        RECT 115.215 149.015 115.545 149.485 ;
        RECT 115.775 148.845 116.025 149.265 ;
        RECT 114.735 148.675 116.025 148.845 ;
        RECT 110.245 147.735 110.420 148.345 ;
        RECT 111.115 148.095 111.285 148.345 ;
        RECT 110.590 147.925 111.285 148.095 ;
        RECT 111.460 147.925 111.880 148.125 ;
        RECT 112.050 147.925 112.380 148.125 ;
        RECT 112.550 147.925 112.880 148.125 ;
        RECT 105.645 147.105 105.905 147.435 ;
        RECT 106.115 146.935 106.390 147.415 ;
        RECT 106.600 147.105 106.805 147.505 ;
        RECT 106.975 146.935 107.310 147.335 ;
        RECT 107.485 146.935 110.075 147.705 ;
        RECT 110.245 147.105 110.585 147.735 ;
        RECT 110.755 146.935 111.005 147.735 ;
        RECT 111.195 147.585 112.420 147.755 ;
        RECT 111.195 147.105 111.525 147.585 ;
        RECT 111.695 146.935 111.920 147.395 ;
        RECT 112.090 147.105 112.420 147.585 ;
        RECT 113.050 147.715 113.220 148.345 ;
        RECT 113.405 147.925 113.755 148.175 ;
        RECT 113.050 147.105 113.550 147.715 ;
        RECT 114.100 147.675 114.270 148.675 ;
        RECT 114.440 147.845 114.685 148.505 ;
        RECT 114.900 147.845 115.165 148.505 ;
        RECT 115.360 147.845 115.645 148.505 ;
        RECT 115.820 148.175 116.035 148.505 ;
        RECT 116.215 148.345 116.465 149.485 ;
        RECT 116.635 148.425 116.965 149.275 ;
        RECT 115.820 147.845 116.125 148.175 ;
        RECT 116.295 147.845 116.605 148.175 ;
        RECT 116.295 147.675 116.465 147.845 ;
        RECT 114.100 147.505 116.465 147.675 ;
        RECT 116.775 147.660 116.965 148.425 ;
        RECT 114.255 146.935 114.585 147.335 ;
        RECT 114.755 147.165 115.085 147.505 ;
        RECT 116.135 146.935 116.465 147.335 ;
        RECT 116.635 147.150 116.965 147.660 ;
        RECT 118.100 148.695 118.635 149.315 ;
        RECT 118.100 147.675 118.415 148.695 ;
        RECT 118.805 148.685 119.135 149.485 ;
        RECT 119.620 148.515 120.010 148.690 ;
        RECT 118.585 148.345 120.010 148.515 ;
        RECT 120.365 148.345 120.625 149.485 ;
        RECT 118.585 147.845 118.755 148.345 ;
        RECT 118.100 147.105 118.715 147.675 ;
        RECT 119.005 147.615 119.270 148.175 ;
        RECT 119.440 147.445 119.610 148.345 ;
        RECT 120.795 148.335 121.125 149.315 ;
        RECT 121.295 148.345 121.575 149.485 ;
        RECT 122.685 148.635 123.015 149.485 ;
        RECT 123.185 149.145 124.295 149.315 ;
        RECT 123.185 148.635 123.405 149.145 ;
        RECT 124.105 148.985 124.295 149.145 ;
        RECT 124.490 149.025 124.820 149.485 ;
        RECT 123.575 148.815 123.875 148.975 ;
        RECT 124.990 148.815 125.225 149.315 ;
        RECT 123.575 148.635 125.225 148.815 ;
        RECT 119.780 147.615 120.135 148.175 ;
        RECT 120.385 147.925 120.720 148.175 ;
        RECT 120.890 147.735 121.060 148.335 ;
        RECT 122.700 148.295 124.675 148.465 ;
        RECT 121.230 147.905 121.565 148.175 ;
        RECT 122.700 147.905 123.030 148.295 ;
        RECT 123.200 147.925 124.000 148.125 ;
        RECT 124.180 147.925 124.675 148.295 ;
        RECT 118.885 146.935 119.100 147.445 ;
        RECT 119.330 147.115 119.610 147.445 ;
        RECT 119.790 146.935 120.030 147.445 ;
        RECT 120.365 147.105 121.060 147.735 ;
        RECT 121.265 146.935 121.575 147.735 ;
        RECT 122.685 147.565 124.845 147.735 ;
        RECT 122.685 147.105 123.015 147.565 ;
        RECT 123.195 146.935 123.365 147.395 ;
        RECT 123.545 147.105 123.875 147.565 ;
        RECT 124.105 146.935 124.275 147.395 ;
        RECT 124.515 147.275 124.845 147.565 ;
        RECT 125.015 147.445 125.225 148.635 ;
        RECT 125.395 148.420 125.705 149.485 ;
        RECT 126.345 148.320 126.635 149.485 ;
        RECT 126.805 148.345 127.075 149.315 ;
        RECT 127.285 148.685 127.565 149.485 ;
        RECT 127.745 148.935 128.940 149.265 ;
        RECT 128.070 148.515 128.490 148.765 ;
        RECT 127.245 148.345 128.490 148.515 ;
        RECT 125.395 147.615 125.710 148.250 ;
        RECT 125.395 147.275 125.705 147.445 ;
        RECT 124.515 147.105 125.705 147.275 ;
        RECT 126.345 146.935 126.635 147.660 ;
        RECT 126.805 147.610 126.975 148.345 ;
        RECT 127.245 148.175 127.415 148.345 ;
        RECT 128.715 148.175 128.885 148.735 ;
        RECT 129.135 148.345 129.390 149.485 ;
        RECT 129.565 149.050 134.910 149.485 ;
        RECT 127.185 147.845 127.415 148.175 ;
        RECT 128.145 147.845 128.885 148.175 ;
        RECT 129.055 147.925 129.390 148.175 ;
        RECT 127.245 147.675 127.415 147.845 ;
        RECT 128.635 147.755 128.885 147.845 ;
        RECT 126.805 147.265 127.075 147.610 ;
        RECT 127.245 147.505 127.985 147.675 ;
        RECT 128.635 147.585 129.370 147.755 ;
        RECT 127.265 146.935 127.645 147.335 ;
        RECT 127.815 147.155 127.985 147.505 ;
        RECT 128.155 146.935 128.890 147.415 ;
        RECT 129.060 147.115 129.370 147.585 ;
        RECT 131.150 147.480 131.490 148.310 ;
        RECT 132.970 147.800 133.320 149.050 ;
        RECT 135.085 148.395 136.755 149.485 ;
        RECT 135.085 147.705 135.835 148.225 ;
        RECT 136.005 147.875 136.755 148.395 ;
        RECT 129.565 146.935 134.910 147.480 ;
        RECT 135.085 146.935 136.755 147.705 ;
        RECT 136.935 147.115 137.195 149.305 ;
        RECT 137.365 148.755 137.705 149.485 ;
        RECT 137.885 148.575 138.155 149.305 ;
        RECT 137.385 148.355 138.155 148.575 ;
        RECT 138.335 148.595 138.565 149.305 ;
        RECT 138.735 148.775 139.065 149.485 ;
        RECT 139.235 148.595 139.495 149.305 ;
        RECT 138.335 148.355 139.495 148.595 ;
        RECT 139.685 148.765 140.145 149.315 ;
        RECT 140.335 148.765 140.665 149.485 ;
        RECT 137.385 147.685 137.675 148.355 ;
        RECT 137.855 147.865 138.320 148.175 ;
        RECT 138.500 147.865 139.025 148.175 ;
        RECT 137.385 147.485 138.615 147.685 ;
        RECT 137.455 146.935 138.125 147.305 ;
        RECT 138.305 147.115 138.615 147.485 ;
        RECT 138.795 147.225 139.025 147.865 ;
        RECT 139.205 147.845 139.505 148.175 ;
        RECT 139.205 146.935 139.495 147.665 ;
        RECT 139.685 147.395 139.935 148.765 ;
        RECT 140.865 148.595 141.165 149.145 ;
        RECT 141.335 148.815 141.615 149.485 ;
        RECT 140.225 148.425 141.165 148.595 ;
        RECT 140.225 148.175 140.395 148.425 ;
        RECT 141.535 148.175 141.800 148.535 ;
        RECT 140.105 147.845 140.395 148.175 ;
        RECT 140.565 147.925 140.905 148.175 ;
        RECT 141.125 147.925 141.800 148.175 ;
        RECT 141.985 148.410 142.255 149.315 ;
        RECT 142.425 148.725 142.755 149.485 ;
        RECT 142.935 148.555 143.115 149.315 ;
        RECT 140.225 147.755 140.395 147.845 ;
        RECT 140.225 147.565 141.615 147.755 ;
        RECT 139.685 147.105 140.245 147.395 ;
        RECT 140.415 146.935 140.665 147.395 ;
        RECT 141.285 147.205 141.615 147.565 ;
        RECT 141.985 147.610 142.165 148.410 ;
        RECT 142.440 148.385 143.115 148.555 ;
        RECT 142.440 148.240 142.610 148.385 ;
        RECT 143.425 148.345 143.635 149.485 ;
        RECT 142.335 147.910 142.610 148.240 ;
        RECT 143.805 148.335 144.135 149.315 ;
        RECT 144.305 148.345 144.535 149.485 ;
        RECT 144.745 148.395 148.255 149.485 ;
        RECT 142.440 147.655 142.610 147.910 ;
        RECT 142.835 147.835 143.175 148.205 ;
        RECT 141.985 147.105 142.245 147.610 ;
        RECT 142.440 147.485 143.105 147.655 ;
        RECT 142.425 146.935 142.755 147.315 ;
        RECT 142.935 147.105 143.105 147.485 ;
        RECT 143.425 146.935 143.635 147.755 ;
        RECT 143.805 147.735 144.055 148.335 ;
        RECT 144.225 147.925 144.555 148.175 ;
        RECT 143.805 147.105 144.135 147.735 ;
        RECT 144.305 146.935 144.535 147.755 ;
        RECT 144.745 147.705 146.395 148.225 ;
        RECT 146.565 147.875 148.255 148.395 ;
        RECT 148.885 148.395 150.095 149.485 ;
        RECT 148.885 147.855 149.405 148.395 ;
        RECT 144.745 146.935 148.255 147.705 ;
        RECT 149.575 147.685 150.095 148.225 ;
        RECT 148.885 146.935 150.095 147.685 ;
        RECT 36.100 146.765 150.180 146.935 ;
        RECT 36.185 146.015 37.395 146.765 ;
        RECT 37.625 146.285 37.905 146.765 ;
        RECT 38.075 146.115 38.335 146.505 ;
        RECT 38.510 146.285 38.765 146.765 ;
        RECT 38.935 146.115 39.230 146.505 ;
        RECT 39.410 146.285 39.685 146.765 ;
        RECT 39.855 146.265 40.155 146.595 ;
        RECT 41.305 146.285 41.585 146.765 ;
        RECT 36.185 145.475 36.705 146.015 ;
        RECT 37.580 145.945 39.230 146.115 ;
        RECT 36.875 145.305 37.395 145.845 ;
        RECT 36.185 144.215 37.395 145.305 ;
        RECT 37.580 145.435 37.985 145.945 ;
        RECT 38.155 145.605 39.295 145.775 ;
        RECT 37.580 145.265 38.335 145.435 ;
        RECT 37.620 144.215 37.905 145.085 ;
        RECT 38.075 145.015 38.335 145.265 ;
        RECT 39.125 145.355 39.295 145.605 ;
        RECT 39.465 145.525 39.815 146.095 ;
        RECT 39.985 145.355 40.155 146.265 ;
        RECT 41.755 146.115 42.015 146.505 ;
        RECT 42.190 146.285 42.445 146.765 ;
        RECT 42.615 146.115 42.910 146.505 ;
        RECT 43.090 146.285 43.365 146.765 ;
        RECT 43.535 146.265 43.835 146.595 ;
        RECT 39.125 145.185 40.155 145.355 ;
        RECT 41.260 145.945 42.910 146.115 ;
        RECT 41.260 145.435 41.665 145.945 ;
        RECT 41.835 145.605 42.975 145.775 ;
        RECT 41.260 145.265 42.015 145.435 ;
        RECT 38.075 144.845 39.195 145.015 ;
        RECT 38.075 144.385 38.335 144.845 ;
        RECT 38.510 144.215 38.765 144.675 ;
        RECT 38.935 144.385 39.195 144.845 ;
        RECT 39.365 144.215 39.675 145.015 ;
        RECT 39.845 144.385 40.155 145.185 ;
        RECT 41.300 144.215 41.585 145.085 ;
        RECT 41.755 145.015 42.015 145.265 ;
        RECT 42.805 145.355 42.975 145.605 ;
        RECT 43.145 145.525 43.495 146.095 ;
        RECT 43.665 145.355 43.835 146.265 ;
        RECT 44.555 146.215 44.725 146.505 ;
        RECT 44.895 146.385 45.225 146.765 ;
        RECT 44.555 146.045 45.220 146.215 ;
        RECT 42.805 145.185 43.835 145.355 ;
        RECT 44.470 145.225 44.820 145.875 ;
        RECT 42.225 145.015 42.395 145.065 ;
        RECT 41.755 144.845 42.875 145.015 ;
        RECT 41.755 144.385 42.015 144.845 ;
        RECT 42.190 144.215 42.445 144.675 ;
        RECT 42.615 144.385 42.875 144.845 ;
        RECT 43.045 144.215 43.355 145.015 ;
        RECT 43.525 144.385 43.835 145.185 ;
        RECT 44.990 145.055 45.220 146.045 ;
        RECT 44.555 144.885 45.220 145.055 ;
        RECT 44.555 144.385 44.725 144.885 ;
        RECT 44.895 144.215 45.225 144.715 ;
        RECT 45.395 144.385 45.580 146.505 ;
        RECT 45.835 146.305 46.085 146.765 ;
        RECT 46.255 146.315 46.590 146.485 ;
        RECT 46.785 146.315 47.460 146.485 ;
        RECT 46.255 146.175 46.425 146.315 ;
        RECT 45.750 145.185 46.030 146.135 ;
        RECT 46.200 146.045 46.425 146.175 ;
        RECT 46.200 144.940 46.370 146.045 ;
        RECT 46.595 145.895 47.120 146.115 ;
        RECT 46.540 145.130 46.780 145.725 ;
        RECT 46.950 145.195 47.120 145.895 ;
        RECT 47.290 145.535 47.460 146.315 ;
        RECT 47.780 146.265 48.150 146.765 ;
        RECT 48.330 146.315 48.735 146.485 ;
        RECT 48.905 146.315 49.690 146.485 ;
        RECT 48.330 146.085 48.500 146.315 ;
        RECT 47.670 145.785 48.500 146.085 ;
        RECT 48.885 145.815 49.350 146.145 ;
        RECT 47.670 145.755 47.870 145.785 ;
        RECT 47.990 145.535 48.160 145.605 ;
        RECT 47.290 145.365 48.160 145.535 ;
        RECT 47.650 145.275 48.160 145.365 ;
        RECT 46.200 144.810 46.505 144.940 ;
        RECT 46.950 144.830 47.480 145.195 ;
        RECT 45.820 144.215 46.085 144.675 ;
        RECT 46.255 144.385 46.505 144.810 ;
        RECT 47.650 144.660 47.820 145.275 ;
        RECT 46.715 144.490 47.820 144.660 ;
        RECT 47.990 144.215 48.160 145.015 ;
        RECT 48.330 144.715 48.500 145.785 ;
        RECT 48.670 144.885 48.860 145.605 ;
        RECT 49.030 144.855 49.350 145.815 ;
        RECT 49.520 145.855 49.690 146.315 ;
        RECT 49.965 146.235 50.175 146.765 ;
        RECT 50.435 146.025 50.765 146.550 ;
        RECT 50.935 146.155 51.105 146.765 ;
        RECT 51.275 146.110 51.605 146.545 ;
        RECT 51.875 146.375 52.205 146.765 ;
        RECT 52.375 146.195 52.545 146.515 ;
        RECT 52.715 146.375 53.045 146.765 ;
        RECT 53.460 146.365 54.415 146.535 ;
        RECT 51.275 146.025 51.655 146.110 ;
        RECT 50.565 145.855 50.765 146.025 ;
        RECT 51.430 145.985 51.655 146.025 ;
        RECT 49.520 145.525 50.395 145.855 ;
        RECT 50.565 145.525 51.315 145.855 ;
        RECT 48.330 144.385 48.580 144.715 ;
        RECT 49.520 144.685 49.690 145.525 ;
        RECT 50.565 145.320 50.755 145.525 ;
        RECT 51.485 145.405 51.655 145.985 ;
        RECT 51.440 145.355 51.655 145.405 ;
        RECT 49.860 144.945 50.755 145.320 ;
        RECT 51.265 145.275 51.655 145.355 ;
        RECT 51.825 146.025 54.075 146.195 ;
        RECT 48.805 144.515 49.690 144.685 ;
        RECT 49.870 144.215 50.185 144.715 ;
        RECT 50.415 144.385 50.755 144.945 ;
        RECT 50.925 144.215 51.095 145.225 ;
        RECT 51.265 144.430 51.595 145.275 ;
        RECT 51.825 145.065 51.995 146.025 ;
        RECT 52.165 145.405 52.410 145.855 ;
        RECT 52.580 145.575 53.130 145.775 ;
        RECT 53.300 145.605 53.675 145.775 ;
        RECT 53.300 145.405 53.470 145.605 ;
        RECT 53.845 145.525 54.075 146.025 ;
        RECT 52.165 145.235 53.470 145.405 ;
        RECT 54.245 145.485 54.415 146.365 ;
        RECT 54.585 145.930 54.875 146.765 ;
        RECT 55.135 146.215 55.305 146.595 ;
        RECT 55.485 146.385 55.815 146.765 ;
        RECT 55.135 146.045 55.800 146.215 ;
        RECT 55.995 146.090 56.255 146.595 ;
        RECT 55.065 145.495 55.405 145.865 ;
        RECT 55.630 145.790 55.800 146.045 ;
        RECT 54.245 145.315 54.875 145.485 ;
        RECT 55.630 145.460 55.905 145.790 ;
        RECT 55.630 145.315 55.800 145.460 ;
        RECT 51.825 144.385 52.205 145.065 ;
        RECT 52.795 144.215 52.965 145.065 ;
        RECT 53.135 144.895 54.375 145.065 ;
        RECT 53.135 144.385 53.465 144.895 ;
        RECT 53.635 144.215 53.805 144.725 ;
        RECT 53.975 144.385 54.375 144.895 ;
        RECT 54.555 144.385 54.875 145.315 ;
        RECT 55.125 145.145 55.800 145.315 ;
        RECT 56.075 145.290 56.255 146.090 ;
        RECT 55.125 144.385 55.305 145.145 ;
        RECT 55.485 144.215 55.815 144.975 ;
        RECT 55.985 144.385 56.255 145.290 ;
        RECT 57.345 146.025 57.810 146.570 ;
        RECT 57.345 145.065 57.515 146.025 ;
        RECT 58.315 145.945 58.485 146.765 ;
        RECT 58.655 146.115 58.985 146.595 ;
        RECT 59.155 146.375 59.505 146.765 ;
        RECT 59.675 146.195 59.905 146.595 ;
        RECT 59.395 146.115 59.905 146.195 ;
        RECT 58.655 146.025 59.905 146.115 ;
        RECT 60.075 146.025 60.395 146.505 ;
        RECT 58.655 145.945 59.565 146.025 ;
        RECT 57.685 145.405 57.930 145.855 ;
        RECT 58.190 145.575 58.885 145.775 ;
        RECT 59.055 145.605 59.655 145.775 ;
        RECT 59.055 145.405 59.225 145.605 ;
        RECT 59.885 145.435 60.055 145.855 ;
        RECT 57.685 145.235 59.225 145.405 ;
        RECT 59.395 145.265 60.055 145.435 ;
        RECT 59.395 145.065 59.565 145.265 ;
        RECT 60.225 145.095 60.395 146.025 ;
        RECT 60.565 146.015 61.775 146.765 ;
        RECT 61.945 146.040 62.235 146.765 ;
        RECT 60.565 145.475 61.085 146.015 ;
        RECT 62.405 145.995 64.075 146.765 ;
        RECT 64.905 146.135 65.235 146.495 ;
        RECT 65.855 146.305 66.105 146.765 ;
        RECT 66.275 146.305 66.835 146.595 ;
        RECT 61.255 145.305 61.775 145.845 ;
        RECT 62.405 145.475 63.155 145.995 ;
        RECT 64.905 145.945 66.295 146.135 ;
        RECT 66.125 145.855 66.295 145.945 ;
        RECT 57.345 144.895 59.565 145.065 ;
        RECT 59.735 144.895 60.395 145.095 ;
        RECT 57.345 144.215 57.645 144.725 ;
        RECT 57.815 144.385 58.145 144.895 ;
        RECT 59.735 144.725 59.905 144.895 ;
        RECT 58.315 144.215 58.945 144.725 ;
        RECT 59.525 144.555 59.905 144.725 ;
        RECT 60.075 144.215 60.375 144.725 ;
        RECT 60.565 144.215 61.775 145.305 ;
        RECT 61.945 144.215 62.235 145.380 ;
        RECT 63.325 145.305 64.075 145.825 ;
        RECT 62.405 144.215 64.075 145.305 ;
        RECT 64.720 145.525 65.395 145.775 ;
        RECT 65.615 145.525 65.955 145.775 ;
        RECT 66.125 145.525 66.415 145.855 ;
        RECT 64.720 145.165 64.985 145.525 ;
        RECT 66.125 145.275 66.295 145.525 ;
        RECT 65.355 145.105 66.295 145.275 ;
        RECT 64.905 144.215 65.185 144.885 ;
        RECT 65.355 144.555 65.655 145.105 ;
        RECT 66.585 144.935 66.835 146.305 ;
        RECT 67.935 145.955 68.205 146.765 ;
        RECT 68.375 145.955 68.705 146.595 ;
        RECT 68.875 145.955 69.115 146.765 ;
        RECT 69.315 145.955 69.585 146.765 ;
        RECT 69.755 145.955 70.085 146.595 ;
        RECT 70.255 145.955 70.495 146.765 ;
        RECT 70.685 146.015 71.895 146.765 ;
        RECT 72.065 146.025 72.505 146.585 ;
        RECT 72.675 146.025 73.125 146.765 ;
        RECT 73.295 146.195 73.465 146.595 ;
        RECT 73.635 146.365 74.055 146.765 ;
        RECT 74.225 146.195 74.455 146.595 ;
        RECT 73.295 146.025 74.455 146.195 ;
        RECT 74.625 146.025 75.115 146.595 ;
        RECT 67.925 145.525 68.275 145.775 ;
        RECT 68.445 145.355 68.615 145.955 ;
        RECT 68.785 145.525 69.135 145.775 ;
        RECT 69.305 145.525 69.655 145.775 ;
        RECT 69.825 145.355 69.995 145.955 ;
        RECT 70.165 145.525 70.515 145.775 ;
        RECT 70.685 145.475 71.205 146.015 ;
        RECT 65.855 144.215 66.185 144.935 ;
        RECT 66.375 144.385 66.835 144.935 ;
        RECT 67.935 144.215 68.265 145.355 ;
        RECT 68.445 145.185 69.125 145.355 ;
        RECT 68.795 144.400 69.125 145.185 ;
        RECT 69.315 144.215 69.645 145.355 ;
        RECT 69.825 145.185 70.505 145.355 ;
        RECT 71.375 145.305 71.895 145.845 ;
        RECT 70.175 144.400 70.505 145.185 ;
        RECT 70.685 144.215 71.895 145.305 ;
        RECT 72.065 145.015 72.375 146.025 ;
        RECT 72.545 145.405 72.715 145.855 ;
        RECT 72.885 145.575 73.275 145.855 ;
        RECT 73.460 145.525 73.705 145.855 ;
        RECT 72.545 145.235 73.335 145.405 ;
        RECT 72.065 144.385 72.505 145.015 ;
        RECT 72.680 144.215 72.995 145.065 ;
        RECT 73.165 144.555 73.335 145.235 ;
        RECT 73.505 144.725 73.705 145.525 ;
        RECT 73.905 144.725 74.155 145.855 ;
        RECT 74.370 145.525 74.775 145.855 ;
        RECT 74.945 145.355 75.115 146.025 ;
        RECT 74.345 145.185 75.115 145.355 ;
        RECT 75.285 145.820 75.625 146.595 ;
        RECT 75.795 146.305 75.965 146.765 ;
        RECT 76.205 146.330 76.565 146.595 ;
        RECT 76.205 146.325 76.560 146.330 ;
        RECT 76.205 146.315 76.555 146.325 ;
        RECT 76.205 146.310 76.550 146.315 ;
        RECT 76.205 146.300 76.545 146.310 ;
        RECT 77.195 146.305 77.365 146.765 ;
        RECT 76.205 146.295 76.540 146.300 ;
        RECT 76.205 146.285 76.530 146.295 ;
        RECT 76.205 146.275 76.520 146.285 ;
        RECT 76.205 146.135 76.505 146.275 ;
        RECT 75.795 145.945 76.505 146.135 ;
        RECT 76.695 146.135 77.025 146.215 ;
        RECT 77.535 146.135 77.875 146.595 ;
        RECT 76.695 145.945 77.875 146.135 ;
        RECT 74.345 144.555 74.595 145.185 ;
        RECT 73.165 144.385 74.595 144.555 ;
        RECT 74.775 144.215 75.105 145.015 ;
        RECT 75.285 144.385 75.565 145.820 ;
        RECT 75.795 145.375 76.080 145.945 ;
        RECT 78.505 145.820 78.845 146.595 ;
        RECT 79.015 146.305 79.185 146.765 ;
        RECT 79.425 146.330 79.785 146.595 ;
        RECT 79.425 146.325 79.780 146.330 ;
        RECT 79.425 146.315 79.775 146.325 ;
        RECT 79.425 146.310 79.770 146.315 ;
        RECT 79.425 146.300 79.765 146.310 ;
        RECT 80.415 146.305 80.585 146.765 ;
        RECT 79.425 146.295 79.760 146.300 ;
        RECT 79.425 146.285 79.750 146.295 ;
        RECT 79.425 146.275 79.740 146.285 ;
        RECT 79.425 146.135 79.725 146.275 ;
        RECT 79.015 145.945 79.725 146.135 ;
        RECT 79.915 146.135 80.245 146.215 ;
        RECT 80.755 146.135 81.095 146.595 ;
        RECT 79.915 145.945 81.095 146.135 ;
        RECT 76.265 145.545 76.735 145.775 ;
        RECT 76.905 145.755 77.235 145.775 ;
        RECT 76.905 145.575 77.355 145.755 ;
        RECT 77.545 145.575 77.875 145.775 ;
        RECT 75.795 145.160 76.945 145.375 ;
        RECT 75.735 144.215 76.445 144.990 ;
        RECT 76.615 144.385 76.945 145.160 ;
        RECT 77.140 144.460 77.355 145.575 ;
        RECT 77.645 145.235 77.875 145.575 ;
        RECT 77.535 144.215 77.865 144.935 ;
        RECT 78.505 144.385 78.785 145.820 ;
        RECT 79.015 145.375 79.300 145.945 ;
        RECT 82.185 145.820 82.525 146.595 ;
        RECT 82.695 146.305 82.865 146.765 ;
        RECT 83.105 146.330 83.465 146.595 ;
        RECT 83.105 146.325 83.460 146.330 ;
        RECT 83.105 146.315 83.455 146.325 ;
        RECT 83.105 146.310 83.450 146.315 ;
        RECT 83.105 146.300 83.445 146.310 ;
        RECT 84.095 146.305 84.265 146.765 ;
        RECT 83.105 146.295 83.440 146.300 ;
        RECT 83.105 146.285 83.430 146.295 ;
        RECT 83.105 146.275 83.420 146.285 ;
        RECT 83.105 146.135 83.405 146.275 ;
        RECT 82.695 145.945 83.405 146.135 ;
        RECT 83.595 146.135 83.925 146.215 ;
        RECT 84.435 146.135 84.775 146.595 ;
        RECT 83.595 145.945 84.775 146.135 ;
        RECT 84.945 146.135 85.285 146.595 ;
        RECT 85.455 146.305 85.625 146.765 ;
        RECT 86.255 146.330 86.615 146.595 ;
        RECT 86.260 146.325 86.615 146.330 ;
        RECT 86.265 146.315 86.615 146.325 ;
        RECT 86.270 146.310 86.615 146.315 ;
        RECT 86.275 146.300 86.615 146.310 ;
        RECT 86.855 146.305 87.025 146.765 ;
        RECT 86.280 146.295 86.615 146.300 ;
        RECT 86.290 146.285 86.615 146.295 ;
        RECT 86.300 146.275 86.615 146.285 ;
        RECT 85.795 146.135 86.125 146.215 ;
        RECT 84.945 145.945 86.125 146.135 ;
        RECT 86.315 146.135 86.615 146.275 ;
        RECT 86.315 145.945 87.025 146.135 ;
        RECT 79.485 145.545 79.955 145.775 ;
        RECT 80.125 145.755 80.455 145.775 ;
        RECT 80.125 145.575 80.575 145.755 ;
        RECT 80.765 145.575 81.095 145.775 ;
        RECT 79.015 145.160 80.165 145.375 ;
        RECT 78.955 144.215 79.665 144.990 ;
        RECT 79.835 144.385 80.165 145.160 ;
        RECT 80.360 144.460 80.575 145.575 ;
        RECT 80.865 145.235 81.095 145.575 ;
        RECT 80.755 144.215 81.085 144.935 ;
        RECT 82.185 144.385 82.465 145.820 ;
        RECT 82.695 145.375 82.980 145.945 ;
        RECT 83.165 145.545 83.635 145.775 ;
        RECT 83.805 145.755 84.135 145.775 ;
        RECT 83.805 145.575 84.255 145.755 ;
        RECT 84.445 145.575 84.775 145.775 ;
        RECT 82.695 145.160 83.845 145.375 ;
        RECT 82.635 144.215 83.345 144.990 ;
        RECT 83.515 144.385 83.845 145.160 ;
        RECT 84.040 144.460 84.255 145.575 ;
        RECT 84.545 145.235 84.775 145.575 ;
        RECT 84.945 145.575 85.275 145.775 ;
        RECT 85.585 145.755 85.915 145.775 ;
        RECT 85.465 145.575 85.915 145.755 ;
        RECT 84.945 145.235 85.175 145.575 ;
        RECT 84.435 144.215 84.765 144.935 ;
        RECT 84.955 144.215 85.285 144.935 ;
        RECT 85.465 144.460 85.680 145.575 ;
        RECT 86.085 145.545 86.555 145.775 ;
        RECT 86.740 145.375 87.025 145.945 ;
        RECT 87.195 145.820 87.535 146.595 ;
        RECT 87.705 146.040 87.995 146.765 ;
        RECT 85.875 145.160 87.025 145.375 ;
        RECT 85.875 144.385 86.205 145.160 ;
        RECT 86.375 144.215 87.085 144.990 ;
        RECT 87.255 144.385 87.535 145.820 ;
        RECT 88.625 145.965 88.965 146.595 ;
        RECT 89.135 145.965 89.385 146.765 ;
        RECT 89.575 146.115 89.905 146.595 ;
        RECT 90.075 146.305 90.300 146.765 ;
        RECT 90.470 146.115 90.800 146.595 ;
        RECT 87.705 144.215 87.995 145.380 ;
        RECT 88.625 145.355 88.800 145.965 ;
        RECT 89.575 145.945 90.800 146.115 ;
        RECT 91.430 145.985 91.930 146.595 ;
        RECT 92.305 145.995 93.975 146.765 ;
        RECT 94.145 146.135 94.485 146.595 ;
        RECT 94.655 146.305 94.825 146.765 ;
        RECT 95.455 146.330 95.815 146.595 ;
        RECT 95.460 146.325 95.815 146.330 ;
        RECT 95.465 146.315 95.815 146.325 ;
        RECT 95.470 146.310 95.815 146.315 ;
        RECT 95.475 146.300 95.815 146.310 ;
        RECT 96.055 146.305 96.225 146.765 ;
        RECT 95.480 146.295 95.815 146.300 ;
        RECT 95.490 146.285 95.815 146.295 ;
        RECT 95.500 146.275 95.815 146.285 ;
        RECT 94.995 146.135 95.325 146.215 ;
        RECT 88.970 145.605 89.665 145.775 ;
        RECT 89.495 145.355 89.665 145.605 ;
        RECT 89.840 145.575 90.260 145.775 ;
        RECT 90.430 145.575 90.760 145.775 ;
        RECT 90.930 145.575 91.260 145.775 ;
        RECT 91.430 145.355 91.600 145.985 ;
        RECT 91.785 145.525 92.135 145.775 ;
        RECT 92.305 145.475 93.055 145.995 ;
        RECT 94.145 145.945 95.325 146.135 ;
        RECT 95.515 146.135 95.815 146.275 ;
        RECT 95.515 145.945 96.225 146.135 ;
        RECT 88.625 144.385 88.965 145.355 ;
        RECT 89.135 144.215 89.305 145.355 ;
        RECT 89.495 145.185 91.930 145.355 ;
        RECT 93.225 145.305 93.975 145.825 ;
        RECT 89.575 144.215 89.825 145.015 ;
        RECT 90.470 144.385 90.800 145.185 ;
        RECT 91.100 144.215 91.430 145.015 ;
        RECT 91.600 144.385 91.930 145.185 ;
        RECT 92.305 144.215 93.975 145.305 ;
        RECT 94.145 145.575 94.475 145.775 ;
        RECT 94.785 145.755 95.115 145.775 ;
        RECT 94.665 145.575 95.115 145.755 ;
        RECT 94.145 145.235 94.375 145.575 ;
        RECT 94.155 144.215 94.485 144.935 ;
        RECT 94.665 144.460 94.880 145.575 ;
        RECT 95.285 145.545 95.755 145.775 ;
        RECT 95.940 145.375 96.225 145.945 ;
        RECT 96.395 145.820 96.735 146.595 ;
        RECT 95.075 145.160 96.225 145.375 ;
        RECT 95.075 144.385 95.405 145.160 ;
        RECT 95.575 144.215 96.285 144.990 ;
        RECT 96.455 144.385 96.735 145.820 ;
        RECT 96.905 146.015 98.115 146.765 ;
        RECT 96.905 145.475 97.425 146.015 ;
        RECT 97.595 145.305 98.115 145.845 ;
        RECT 96.905 144.215 98.115 145.305 ;
        RECT 98.285 145.820 98.625 146.595 ;
        RECT 98.795 146.305 98.965 146.765 ;
        RECT 99.205 146.330 99.565 146.595 ;
        RECT 99.205 146.325 99.560 146.330 ;
        RECT 99.205 146.315 99.555 146.325 ;
        RECT 99.205 146.310 99.550 146.315 ;
        RECT 99.205 146.300 99.545 146.310 ;
        RECT 100.195 146.305 100.365 146.765 ;
        RECT 99.205 146.295 99.540 146.300 ;
        RECT 99.205 146.285 99.530 146.295 ;
        RECT 99.205 146.275 99.520 146.285 ;
        RECT 99.205 146.135 99.505 146.275 ;
        RECT 98.795 145.945 99.505 146.135 ;
        RECT 99.695 146.135 100.025 146.215 ;
        RECT 100.535 146.135 100.875 146.595 ;
        RECT 99.695 145.945 100.875 146.135 ;
        RECT 98.285 144.385 98.565 145.820 ;
        RECT 98.795 145.375 99.080 145.945 ;
        RECT 101.045 145.820 101.385 146.595 ;
        RECT 101.555 146.305 101.725 146.765 ;
        RECT 101.965 146.330 102.325 146.595 ;
        RECT 101.965 146.325 102.320 146.330 ;
        RECT 101.965 146.315 102.315 146.325 ;
        RECT 101.965 146.310 102.310 146.315 ;
        RECT 101.965 146.300 102.305 146.310 ;
        RECT 102.955 146.305 103.125 146.765 ;
        RECT 101.965 146.295 102.300 146.300 ;
        RECT 101.965 146.285 102.290 146.295 ;
        RECT 101.965 146.275 102.280 146.285 ;
        RECT 101.965 146.135 102.265 146.275 ;
        RECT 101.555 145.945 102.265 146.135 ;
        RECT 102.455 146.135 102.785 146.215 ;
        RECT 103.295 146.135 103.635 146.595 ;
        RECT 102.455 145.945 103.635 146.135 ;
        RECT 103.805 146.090 104.065 146.595 ;
        RECT 104.245 146.385 104.575 146.765 ;
        RECT 104.755 146.215 104.925 146.595 ;
        RECT 99.265 145.545 99.735 145.775 ;
        RECT 99.905 145.755 100.235 145.775 ;
        RECT 99.905 145.575 100.355 145.755 ;
        RECT 100.545 145.575 100.875 145.775 ;
        RECT 98.795 145.160 99.945 145.375 ;
        RECT 98.735 144.215 99.445 144.990 ;
        RECT 99.615 144.385 99.945 145.160 ;
        RECT 100.140 144.460 100.355 145.575 ;
        RECT 100.645 145.235 100.875 145.575 ;
        RECT 100.535 144.215 100.865 144.935 ;
        RECT 101.045 144.385 101.325 145.820 ;
        RECT 101.555 145.375 101.840 145.945 ;
        RECT 102.025 145.545 102.495 145.775 ;
        RECT 102.665 145.755 102.995 145.775 ;
        RECT 102.665 145.575 103.115 145.755 ;
        RECT 103.305 145.575 103.635 145.775 ;
        RECT 101.555 145.160 102.705 145.375 ;
        RECT 101.495 144.215 102.205 144.990 ;
        RECT 102.375 144.385 102.705 145.160 ;
        RECT 102.900 144.460 103.115 145.575 ;
        RECT 103.405 145.235 103.635 145.575 ;
        RECT 103.805 145.290 103.985 146.090 ;
        RECT 104.260 146.045 104.925 146.215 ;
        RECT 104.260 145.790 104.430 146.045 ;
        RECT 104.155 145.460 104.430 145.790 ;
        RECT 104.655 145.495 104.995 145.865 ;
        RECT 105.185 145.820 105.525 146.595 ;
        RECT 105.695 146.305 105.865 146.765 ;
        RECT 106.105 146.330 106.465 146.595 ;
        RECT 106.105 146.325 106.460 146.330 ;
        RECT 106.105 146.315 106.455 146.325 ;
        RECT 106.105 146.310 106.450 146.315 ;
        RECT 106.105 146.300 106.445 146.310 ;
        RECT 107.095 146.305 107.265 146.765 ;
        RECT 106.105 146.295 106.440 146.300 ;
        RECT 106.105 146.285 106.430 146.295 ;
        RECT 106.105 146.275 106.420 146.285 ;
        RECT 106.105 146.135 106.405 146.275 ;
        RECT 105.695 145.945 106.405 146.135 ;
        RECT 106.595 146.135 106.925 146.215 ;
        RECT 107.435 146.135 107.775 146.595 ;
        RECT 106.595 145.945 107.775 146.135 ;
        RECT 108.035 146.215 108.205 146.595 ;
        RECT 108.385 146.385 108.715 146.765 ;
        RECT 108.035 146.045 108.700 146.215 ;
        RECT 108.895 146.090 109.155 146.595 ;
        RECT 104.260 145.315 104.430 145.460 ;
        RECT 103.295 144.215 103.625 144.935 ;
        RECT 103.805 144.385 104.075 145.290 ;
        RECT 104.260 145.145 104.935 145.315 ;
        RECT 104.245 144.215 104.575 144.975 ;
        RECT 104.755 144.385 104.935 145.145 ;
        RECT 105.185 144.385 105.465 145.820 ;
        RECT 105.695 145.375 105.980 145.945 ;
        RECT 106.165 145.545 106.635 145.775 ;
        RECT 106.805 145.755 107.135 145.775 ;
        RECT 106.805 145.575 107.255 145.755 ;
        RECT 107.445 145.575 107.775 145.775 ;
        RECT 105.695 145.160 106.845 145.375 ;
        RECT 105.635 144.215 106.345 144.990 ;
        RECT 106.515 144.385 106.845 145.160 ;
        RECT 107.040 144.460 107.255 145.575 ;
        RECT 107.545 145.235 107.775 145.575 ;
        RECT 107.965 145.495 108.295 145.865 ;
        RECT 108.530 145.790 108.700 146.045 ;
        RECT 108.530 145.460 108.815 145.790 ;
        RECT 108.530 145.315 108.700 145.460 ;
        RECT 108.035 145.145 108.700 145.315 ;
        RECT 108.985 145.290 109.155 146.090 ;
        RECT 109.415 146.215 109.585 146.595 ;
        RECT 109.765 146.385 110.095 146.765 ;
        RECT 109.415 146.045 110.080 146.215 ;
        RECT 110.275 146.090 110.535 146.595 ;
        RECT 109.345 145.495 109.685 145.865 ;
        RECT 109.910 145.790 110.080 146.045 ;
        RECT 109.910 145.460 110.185 145.790 ;
        RECT 109.910 145.315 110.080 145.460 ;
        RECT 107.435 144.215 107.765 144.935 ;
        RECT 108.035 144.385 108.205 145.145 ;
        RECT 108.385 144.215 108.715 144.975 ;
        RECT 108.885 144.385 109.155 145.290 ;
        RECT 109.405 145.145 110.080 145.315 ;
        RECT 110.355 145.290 110.535 146.090 ;
        RECT 110.705 146.135 111.045 146.595 ;
        RECT 111.215 146.305 111.385 146.765 ;
        RECT 112.015 146.330 112.375 146.595 ;
        RECT 112.020 146.325 112.375 146.330 ;
        RECT 112.025 146.315 112.375 146.325 ;
        RECT 112.030 146.310 112.375 146.315 ;
        RECT 112.035 146.300 112.375 146.310 ;
        RECT 112.615 146.305 112.785 146.765 ;
        RECT 112.040 146.295 112.375 146.300 ;
        RECT 112.050 146.285 112.375 146.295 ;
        RECT 112.060 146.275 112.375 146.285 ;
        RECT 111.555 146.135 111.885 146.215 ;
        RECT 110.705 145.945 111.885 146.135 ;
        RECT 112.075 146.135 112.375 146.275 ;
        RECT 112.075 145.945 112.785 146.135 ;
        RECT 109.405 144.385 109.585 145.145 ;
        RECT 109.765 144.215 110.095 144.975 ;
        RECT 110.265 144.385 110.535 145.290 ;
        RECT 110.705 145.575 111.035 145.775 ;
        RECT 111.345 145.755 111.675 145.775 ;
        RECT 111.225 145.575 111.675 145.755 ;
        RECT 110.705 145.235 110.935 145.575 ;
        RECT 110.715 144.215 111.045 144.935 ;
        RECT 111.225 144.460 111.440 145.575 ;
        RECT 111.845 145.545 112.315 145.775 ;
        RECT 112.500 145.375 112.785 145.945 ;
        RECT 112.955 145.820 113.295 146.595 ;
        RECT 113.465 146.040 113.755 146.765 ;
        RECT 113.925 146.135 114.265 146.595 ;
        RECT 114.435 146.305 114.605 146.765 ;
        RECT 115.235 146.330 115.595 146.595 ;
        RECT 115.240 146.325 115.595 146.330 ;
        RECT 115.245 146.315 115.595 146.325 ;
        RECT 115.250 146.310 115.595 146.315 ;
        RECT 115.255 146.300 115.595 146.310 ;
        RECT 115.835 146.305 116.005 146.765 ;
        RECT 115.260 146.295 115.595 146.300 ;
        RECT 115.270 146.285 115.595 146.295 ;
        RECT 115.280 146.275 115.595 146.285 ;
        RECT 114.775 146.135 115.105 146.215 ;
        RECT 113.925 145.945 115.105 146.135 ;
        RECT 115.295 146.135 115.595 146.275 ;
        RECT 115.295 145.945 116.005 146.135 ;
        RECT 111.635 145.160 112.785 145.375 ;
        RECT 111.635 144.385 111.965 145.160 ;
        RECT 112.135 144.215 112.845 144.990 ;
        RECT 113.015 144.385 113.295 145.820 ;
        RECT 113.925 145.575 114.255 145.775 ;
        RECT 114.565 145.755 114.895 145.775 ;
        RECT 114.445 145.575 114.895 145.755 ;
        RECT 113.465 144.215 113.755 145.380 ;
        RECT 113.925 145.235 114.155 145.575 ;
        RECT 113.935 144.215 114.265 144.935 ;
        RECT 114.445 144.460 114.660 145.575 ;
        RECT 115.065 145.545 115.535 145.775 ;
        RECT 115.720 145.375 116.005 145.945 ;
        RECT 116.175 145.820 116.515 146.595 ;
        RECT 116.685 146.135 117.025 146.595 ;
        RECT 117.195 146.305 117.365 146.765 ;
        RECT 117.995 146.330 118.355 146.595 ;
        RECT 118.000 146.325 118.355 146.330 ;
        RECT 118.005 146.315 118.355 146.325 ;
        RECT 118.010 146.310 118.355 146.315 ;
        RECT 118.015 146.300 118.355 146.310 ;
        RECT 118.595 146.305 118.765 146.765 ;
        RECT 118.020 146.295 118.355 146.300 ;
        RECT 118.030 146.285 118.355 146.295 ;
        RECT 118.040 146.275 118.355 146.285 ;
        RECT 117.535 146.135 117.865 146.215 ;
        RECT 116.685 145.945 117.865 146.135 ;
        RECT 118.055 146.135 118.355 146.275 ;
        RECT 118.055 145.945 118.765 146.135 ;
        RECT 114.855 145.160 116.005 145.375 ;
        RECT 114.855 144.385 115.185 145.160 ;
        RECT 115.355 144.215 116.065 144.990 ;
        RECT 116.235 144.385 116.515 145.820 ;
        RECT 116.685 145.575 117.015 145.775 ;
        RECT 117.325 145.755 117.655 145.775 ;
        RECT 117.205 145.575 117.655 145.755 ;
        RECT 116.685 145.235 116.915 145.575 ;
        RECT 116.695 144.215 117.025 144.935 ;
        RECT 117.205 144.460 117.420 145.575 ;
        RECT 117.825 145.545 118.295 145.775 ;
        RECT 118.480 145.375 118.765 145.945 ;
        RECT 118.935 145.820 119.275 146.595 ;
        RECT 119.535 146.215 119.705 146.595 ;
        RECT 119.885 146.385 120.215 146.765 ;
        RECT 119.535 146.045 120.200 146.215 ;
        RECT 120.395 146.090 120.655 146.595 ;
        RECT 117.615 145.160 118.765 145.375 ;
        RECT 117.615 144.385 117.945 145.160 ;
        RECT 118.115 144.215 118.825 144.990 ;
        RECT 118.995 144.385 119.275 145.820 ;
        RECT 119.465 145.495 119.795 145.865 ;
        RECT 120.030 145.790 120.200 146.045 ;
        RECT 120.030 145.460 120.315 145.790 ;
        RECT 120.030 145.315 120.200 145.460 ;
        RECT 119.535 145.145 120.200 145.315 ;
        RECT 120.485 145.290 120.655 146.090 ;
        RECT 120.825 146.135 121.165 146.595 ;
        RECT 121.335 146.305 121.505 146.765 ;
        RECT 122.135 146.330 122.495 146.595 ;
        RECT 122.140 146.325 122.495 146.330 ;
        RECT 122.145 146.315 122.495 146.325 ;
        RECT 122.150 146.310 122.495 146.315 ;
        RECT 122.155 146.300 122.495 146.310 ;
        RECT 122.735 146.305 122.905 146.765 ;
        RECT 122.160 146.295 122.495 146.300 ;
        RECT 122.170 146.285 122.495 146.295 ;
        RECT 122.180 146.275 122.495 146.285 ;
        RECT 121.675 146.135 122.005 146.215 ;
        RECT 120.825 145.945 122.005 146.135 ;
        RECT 122.195 146.135 122.495 146.275 ;
        RECT 122.195 145.945 122.905 146.135 ;
        RECT 119.535 144.385 119.705 145.145 ;
        RECT 119.885 144.215 120.215 144.975 ;
        RECT 120.385 144.385 120.655 145.290 ;
        RECT 120.825 145.575 121.155 145.775 ;
        RECT 121.465 145.755 121.795 145.775 ;
        RECT 121.345 145.575 121.795 145.755 ;
        RECT 120.825 145.235 121.055 145.575 ;
        RECT 120.835 144.215 121.165 144.935 ;
        RECT 121.345 144.460 121.560 145.575 ;
        RECT 121.965 145.545 122.435 145.775 ;
        RECT 122.620 145.375 122.905 145.945 ;
        RECT 123.075 145.820 123.415 146.595 ;
        RECT 123.825 146.295 123.995 146.765 ;
        RECT 124.665 146.295 124.835 146.765 ;
        RECT 125.100 146.375 126.330 146.595 ;
        RECT 124.165 146.125 124.495 146.205 ;
        RECT 125.525 146.125 125.855 146.205 ;
        RECT 121.755 145.160 122.905 145.375 ;
        RECT 121.755 144.385 122.085 145.160 ;
        RECT 122.255 144.215 122.965 144.990 ;
        RECT 123.135 144.385 123.415 145.820 ;
        RECT 123.585 145.945 125.855 146.125 ;
        RECT 126.080 146.125 126.330 146.375 ;
        RECT 126.500 146.295 126.670 146.765 ;
        RECT 126.840 146.125 127.170 146.595 ;
        RECT 127.440 146.295 127.610 146.765 ;
        RECT 126.080 145.945 127.170 146.125 ;
        RECT 127.780 146.125 128.110 146.595 ;
        RECT 128.280 146.295 128.450 146.765 ;
        RECT 128.620 146.125 128.950 146.595 ;
        RECT 129.120 146.295 129.290 146.765 ;
        RECT 127.780 145.945 129.360 146.125 ;
        RECT 123.585 145.435 123.995 145.945 ;
        RECT 124.205 145.605 124.865 145.775 ;
        RECT 123.585 145.225 124.455 145.435 ;
        RECT 124.695 145.405 124.865 145.605 ;
        RECT 125.390 145.575 126.060 145.775 ;
        RECT 126.250 145.575 127.770 145.775 ;
        RECT 127.940 145.575 128.435 145.775 ;
        RECT 128.605 145.575 128.935 145.775 ;
        RECT 127.600 145.405 127.770 145.575 ;
        RECT 128.605 145.405 128.775 145.575 ;
        RECT 124.695 145.235 127.430 145.405 ;
        RECT 127.600 145.235 128.775 145.405 ;
        RECT 123.785 144.555 124.035 145.055 ;
        RECT 124.205 144.725 124.455 145.225 ;
        RECT 127.260 145.065 127.430 145.235 ;
        RECT 129.190 145.065 129.360 145.945 ;
        RECT 129.565 145.995 131.235 146.765 ;
        RECT 131.955 146.215 132.125 146.505 ;
        RECT 132.295 146.385 132.625 146.765 ;
        RECT 131.955 146.045 132.620 146.215 ;
        RECT 129.565 145.475 130.315 145.995 ;
        RECT 130.485 145.305 131.235 145.825 ;
        RECT 124.625 144.895 127.090 145.065 ;
        RECT 127.260 144.895 129.360 145.065 ;
        RECT 124.625 144.555 125.395 144.895 ;
        RECT 123.785 144.385 125.395 144.555 ;
        RECT 125.565 144.215 125.870 144.715 ;
        RECT 126.040 144.385 126.290 144.895 ;
        RECT 126.880 144.725 127.090 144.895 ;
        RECT 127.820 144.725 128.070 144.895 ;
        RECT 126.460 144.215 126.710 144.715 ;
        RECT 126.880 144.385 127.195 144.725 ;
        RECT 128.245 144.715 128.415 144.725 ;
        RECT 129.165 144.715 129.335 144.725 ;
        RECT 127.400 144.555 127.650 144.715 ;
        RECT 128.240 144.555 128.490 144.715 ;
        RECT 127.400 144.385 128.490 144.555 ;
        RECT 128.660 144.215 128.910 144.715 ;
        RECT 129.080 144.385 129.360 144.715 ;
        RECT 129.565 144.215 131.235 145.305 ;
        RECT 131.870 145.225 132.220 145.875 ;
        RECT 132.390 145.055 132.620 146.045 ;
        RECT 131.955 144.885 132.620 145.055 ;
        RECT 131.955 144.385 132.125 144.885 ;
        RECT 132.295 144.215 132.625 144.715 ;
        RECT 132.795 144.385 132.980 146.505 ;
        RECT 133.235 146.305 133.485 146.765 ;
        RECT 133.655 146.315 133.990 146.485 ;
        RECT 134.185 146.315 134.860 146.485 ;
        RECT 133.655 146.175 133.825 146.315 ;
        RECT 133.150 145.185 133.430 146.135 ;
        RECT 133.600 146.045 133.825 146.175 ;
        RECT 133.600 144.940 133.770 146.045 ;
        RECT 133.995 145.895 134.520 146.115 ;
        RECT 133.940 145.130 134.180 145.725 ;
        RECT 134.350 145.195 134.520 145.895 ;
        RECT 134.690 145.535 134.860 146.315 ;
        RECT 135.180 146.265 135.550 146.765 ;
        RECT 135.730 146.315 136.135 146.485 ;
        RECT 136.305 146.315 137.090 146.485 ;
        RECT 135.730 146.085 135.900 146.315 ;
        RECT 135.070 145.785 135.900 146.085 ;
        RECT 136.285 145.815 136.750 146.145 ;
        RECT 135.070 145.755 135.270 145.785 ;
        RECT 135.390 145.535 135.560 145.605 ;
        RECT 134.690 145.365 135.560 145.535 ;
        RECT 135.050 145.275 135.560 145.365 ;
        RECT 133.600 144.810 133.905 144.940 ;
        RECT 134.350 144.830 134.880 145.195 ;
        RECT 133.220 144.215 133.485 144.675 ;
        RECT 133.655 144.385 133.905 144.810 ;
        RECT 135.050 144.660 135.220 145.275 ;
        RECT 134.115 144.490 135.220 144.660 ;
        RECT 135.390 144.215 135.560 145.015 ;
        RECT 135.730 144.715 135.900 145.785 ;
        RECT 136.070 144.885 136.260 145.605 ;
        RECT 136.430 144.855 136.750 145.815 ;
        RECT 136.920 145.855 137.090 146.315 ;
        RECT 137.365 146.235 137.575 146.765 ;
        RECT 137.835 146.025 138.165 146.550 ;
        RECT 138.335 146.155 138.505 146.765 ;
        RECT 138.675 146.110 139.005 146.545 ;
        RECT 138.675 146.025 139.055 146.110 ;
        RECT 139.225 146.040 139.515 146.765 ;
        RECT 139.790 146.295 139.960 146.765 ;
        RECT 140.130 146.125 140.460 146.595 ;
        RECT 140.630 146.295 140.800 146.765 ;
        RECT 140.970 146.125 141.300 146.595 ;
        RECT 141.470 146.295 141.640 146.765 ;
        RECT 137.965 145.855 138.165 146.025 ;
        RECT 138.830 145.985 139.055 146.025 ;
        RECT 136.920 145.525 137.795 145.855 ;
        RECT 137.965 145.525 138.715 145.855 ;
        RECT 135.730 144.385 135.980 144.715 ;
        RECT 136.920 144.685 137.090 145.525 ;
        RECT 137.965 145.320 138.155 145.525 ;
        RECT 138.885 145.405 139.055 145.985 ;
        RECT 138.840 145.355 139.055 145.405 ;
        RECT 139.720 145.945 141.300 146.125 ;
        RECT 141.910 146.125 142.240 146.595 ;
        RECT 142.410 146.295 142.580 146.765 ;
        RECT 142.750 146.375 143.980 146.595 ;
        RECT 142.750 146.125 143.000 146.375 ;
        RECT 144.245 146.295 144.415 146.765 ;
        RECT 145.085 146.295 145.255 146.765 ;
        RECT 145.755 146.215 145.925 146.595 ;
        RECT 146.140 146.385 146.470 146.765 ;
        RECT 141.910 145.945 143.000 146.125 ;
        RECT 143.225 146.125 143.555 146.205 ;
        RECT 144.585 146.125 144.915 146.205 ;
        RECT 143.225 145.945 145.495 146.125 ;
        RECT 145.755 146.045 146.470 146.215 ;
        RECT 137.260 144.945 138.155 145.320 ;
        RECT 138.665 145.275 139.055 145.355 ;
        RECT 136.205 144.515 137.090 144.685 ;
        RECT 137.270 144.215 137.585 144.715 ;
        RECT 137.815 144.385 138.155 144.945 ;
        RECT 138.325 144.215 138.495 145.225 ;
        RECT 138.665 144.430 138.995 145.275 ;
        RECT 139.225 144.215 139.515 145.380 ;
        RECT 139.720 145.065 139.890 145.945 ;
        RECT 143.885 145.915 144.055 145.945 ;
        RECT 140.145 145.575 140.475 145.775 ;
        RECT 140.645 145.575 141.140 145.775 ;
        RECT 141.310 145.575 142.830 145.775 ;
        RECT 143.020 145.575 143.690 145.775 ;
        RECT 144.215 145.605 144.875 145.775 ;
        RECT 140.305 145.405 140.475 145.575 ;
        RECT 141.310 145.405 141.480 145.575 ;
        RECT 144.215 145.405 144.385 145.605 ;
        RECT 145.085 145.435 145.495 145.945 ;
        RECT 145.665 145.495 146.020 145.865 ;
        RECT 146.300 145.855 146.470 146.045 ;
        RECT 146.640 146.020 146.895 146.595 ;
        RECT 146.300 145.525 146.555 145.855 ;
        RECT 140.305 145.235 141.480 145.405 ;
        RECT 141.650 145.235 144.385 145.405 ;
        RECT 141.650 145.065 141.820 145.235 ;
        RECT 144.625 145.225 145.495 145.435 ;
        RECT 146.300 145.315 146.470 145.525 ;
        RECT 139.720 144.895 141.820 145.065 ;
        RECT 141.990 144.895 144.455 145.065 ;
        RECT 141.010 144.725 141.260 144.895 ;
        RECT 141.990 144.725 142.200 144.895 ;
        RECT 139.745 144.715 139.915 144.725 ;
        RECT 140.665 144.715 140.835 144.725 ;
        RECT 139.720 144.385 140.000 144.715 ;
        RECT 140.170 144.215 140.420 144.715 ;
        RECT 140.590 144.555 140.840 144.715 ;
        RECT 141.430 144.555 141.680 144.715 ;
        RECT 140.590 144.385 141.680 144.555 ;
        RECT 141.885 144.385 142.200 144.725 ;
        RECT 142.370 144.215 142.620 144.715 ;
        RECT 142.790 144.385 143.040 144.895 ;
        RECT 143.210 144.215 143.515 144.715 ;
        RECT 143.685 144.555 144.455 144.895 ;
        RECT 144.625 144.725 144.875 145.225 ;
        RECT 145.755 145.145 146.470 145.315 ;
        RECT 146.725 145.290 146.895 146.020 ;
        RECT 147.070 145.925 147.330 146.765 ;
        RECT 147.505 146.015 148.715 146.765 ;
        RECT 148.885 146.015 150.095 146.765 ;
        RECT 147.505 145.475 148.025 146.015 ;
        RECT 145.045 144.555 145.295 145.055 ;
        RECT 143.685 144.385 145.295 144.555 ;
        RECT 145.755 144.385 145.925 145.145 ;
        RECT 146.140 144.215 146.470 144.975 ;
        RECT 146.640 144.385 146.895 145.290 ;
        RECT 147.070 144.215 147.330 145.365 ;
        RECT 148.195 145.305 148.715 145.845 ;
        RECT 147.505 144.215 148.715 145.305 ;
        RECT 148.885 145.305 149.405 145.845 ;
        RECT 149.575 145.475 150.095 146.015 ;
        RECT 148.885 144.215 150.095 145.305 ;
        RECT 36.100 144.045 150.180 144.215 ;
        RECT 36.185 142.955 37.395 144.045 ;
        RECT 36.185 142.245 36.705 142.785 ;
        RECT 36.875 142.415 37.395 142.955 ;
        RECT 38.030 142.895 38.290 144.045 ;
        RECT 38.465 142.970 38.720 143.875 ;
        RECT 38.890 143.285 39.220 144.045 ;
        RECT 39.435 143.115 39.605 143.875 ;
        RECT 40.415 143.375 40.585 143.875 ;
        RECT 40.755 143.545 41.085 144.045 ;
        RECT 40.415 143.205 41.080 143.375 ;
        RECT 36.185 141.495 37.395 142.245 ;
        RECT 38.030 141.495 38.290 142.335 ;
        RECT 38.465 142.240 38.635 142.970 ;
        RECT 38.890 142.945 39.605 143.115 ;
        RECT 38.890 142.735 39.060 142.945 ;
        RECT 38.805 142.405 39.060 142.735 ;
        RECT 38.465 141.665 38.720 142.240 ;
        RECT 38.890 142.215 39.060 142.405 ;
        RECT 39.340 142.395 39.695 142.765 ;
        RECT 40.330 142.385 40.680 143.035 ;
        RECT 40.850 142.215 41.080 143.205 ;
        RECT 38.890 142.045 39.605 142.215 ;
        RECT 38.890 141.495 39.220 141.875 ;
        RECT 39.435 141.665 39.605 142.045 ;
        RECT 40.415 142.045 41.080 142.215 ;
        RECT 40.415 141.755 40.585 142.045 ;
        RECT 40.755 141.495 41.085 141.875 ;
        RECT 41.255 141.755 41.440 143.875 ;
        RECT 41.680 143.585 41.945 144.045 ;
        RECT 42.115 143.450 42.365 143.875 ;
        RECT 42.575 143.600 43.680 143.770 ;
        RECT 42.060 143.320 42.365 143.450 ;
        RECT 41.610 142.125 41.890 143.075 ;
        RECT 42.060 142.215 42.230 143.320 ;
        RECT 42.400 142.535 42.640 143.130 ;
        RECT 42.810 143.065 43.340 143.430 ;
        RECT 42.810 142.365 42.980 143.065 ;
        RECT 43.510 142.985 43.680 143.600 ;
        RECT 43.850 143.245 44.020 144.045 ;
        RECT 44.190 143.545 44.440 143.875 ;
        RECT 44.665 143.575 45.550 143.745 ;
        RECT 43.510 142.895 44.020 142.985 ;
        RECT 42.060 142.085 42.285 142.215 ;
        RECT 42.455 142.145 42.980 142.365 ;
        RECT 43.150 142.725 44.020 142.895 ;
        RECT 41.695 141.495 41.945 141.955 ;
        RECT 42.115 141.945 42.285 142.085 ;
        RECT 43.150 141.945 43.320 142.725 ;
        RECT 43.850 142.655 44.020 142.725 ;
        RECT 43.530 142.475 43.730 142.505 ;
        RECT 44.190 142.475 44.360 143.545 ;
        RECT 44.530 142.655 44.720 143.375 ;
        RECT 43.530 142.175 44.360 142.475 ;
        RECT 44.890 142.445 45.210 143.405 ;
        RECT 42.115 141.775 42.450 141.945 ;
        RECT 42.645 141.775 43.320 141.945 ;
        RECT 43.640 141.495 44.010 141.995 ;
        RECT 44.190 141.945 44.360 142.175 ;
        RECT 44.745 142.115 45.210 142.445 ;
        RECT 45.380 142.735 45.550 143.575 ;
        RECT 45.730 143.545 46.045 144.045 ;
        RECT 46.275 143.315 46.615 143.875 ;
        RECT 45.720 142.940 46.615 143.315 ;
        RECT 46.785 143.035 46.955 144.045 ;
        RECT 46.425 142.735 46.615 142.940 ;
        RECT 47.125 142.985 47.455 143.830 ;
        RECT 47.125 142.905 47.515 142.985 ;
        RECT 47.685 142.955 48.895 144.045 ;
        RECT 47.300 142.855 47.515 142.905 ;
        RECT 45.380 142.405 46.255 142.735 ;
        RECT 46.425 142.405 47.175 142.735 ;
        RECT 45.380 141.945 45.550 142.405 ;
        RECT 46.425 142.235 46.625 142.405 ;
        RECT 47.345 142.275 47.515 142.855 ;
        RECT 47.290 142.235 47.515 142.275 ;
        RECT 44.190 141.775 44.595 141.945 ;
        RECT 44.765 141.775 45.550 141.945 ;
        RECT 45.825 141.495 46.035 142.025 ;
        RECT 46.295 141.710 46.625 142.235 ;
        RECT 47.135 142.150 47.515 142.235 ;
        RECT 47.685 142.245 48.205 142.785 ;
        RECT 48.375 142.415 48.895 142.955 ;
        RECT 49.065 142.880 49.355 144.045 ;
        RECT 49.530 142.895 49.790 144.045 ;
        RECT 49.965 142.970 50.220 143.875 ;
        RECT 50.390 143.285 50.720 144.045 ;
        RECT 50.935 143.115 51.105 143.875 ;
        RECT 51.420 143.175 51.705 144.045 ;
        RECT 51.875 143.415 52.135 143.875 ;
        RECT 52.310 143.585 52.565 144.045 ;
        RECT 52.735 143.415 52.995 143.875 ;
        RECT 51.875 143.245 52.995 143.415 ;
        RECT 53.165 143.245 53.475 144.045 ;
        RECT 46.795 141.495 46.965 142.105 ;
        RECT 47.135 141.715 47.465 142.150 ;
        RECT 47.685 141.495 48.895 142.245 ;
        RECT 49.065 141.495 49.355 142.220 ;
        RECT 49.530 141.495 49.790 142.335 ;
        RECT 49.965 142.240 50.135 142.970 ;
        RECT 50.390 142.945 51.105 143.115 ;
        RECT 51.875 142.995 52.135 143.245 ;
        RECT 53.645 143.075 53.955 143.875 ;
        RECT 50.390 142.735 50.560 142.945 ;
        RECT 51.380 142.825 52.135 142.995 ;
        RECT 52.925 142.905 53.955 143.075 ;
        RECT 50.305 142.405 50.560 142.735 ;
        RECT 49.965 141.665 50.220 142.240 ;
        RECT 50.390 142.215 50.560 142.405 ;
        RECT 50.840 142.395 51.195 142.765 ;
        RECT 51.380 142.315 51.785 142.825 ;
        RECT 52.925 142.655 53.095 142.905 ;
        RECT 51.955 142.485 53.095 142.655 ;
        RECT 50.390 142.045 51.105 142.215 ;
        RECT 51.380 142.145 53.030 142.315 ;
        RECT 53.265 142.165 53.615 142.735 ;
        RECT 50.390 141.495 50.720 141.875 ;
        RECT 50.935 141.665 51.105 142.045 ;
        RECT 51.425 141.495 51.705 141.975 ;
        RECT 51.875 141.755 52.135 142.145 ;
        RECT 52.310 141.495 52.565 141.975 ;
        RECT 52.735 141.755 53.030 142.145 ;
        RECT 53.785 141.995 53.955 142.905 ;
        RECT 54.590 142.895 54.850 144.045 ;
        RECT 55.025 142.970 55.280 143.875 ;
        RECT 55.450 143.285 55.780 144.045 ;
        RECT 55.995 143.115 56.165 143.875 ;
        RECT 53.210 141.495 53.485 141.975 ;
        RECT 53.655 141.665 53.955 141.995 ;
        RECT 54.590 141.495 54.850 142.335 ;
        RECT 55.025 142.240 55.195 142.970 ;
        RECT 55.450 142.945 56.165 143.115 ;
        RECT 56.425 142.955 58.095 144.045 ;
        RECT 55.450 142.735 55.620 142.945 ;
        RECT 55.365 142.405 55.620 142.735 ;
        RECT 55.025 141.665 55.280 142.240 ;
        RECT 55.450 142.215 55.620 142.405 ;
        RECT 55.900 142.395 56.255 142.765 ;
        RECT 56.425 142.265 57.175 142.785 ;
        RECT 57.345 142.435 58.095 142.955 ;
        RECT 58.730 142.895 58.990 144.045 ;
        RECT 59.165 142.970 59.420 143.875 ;
        RECT 59.590 143.285 59.920 144.045 ;
        RECT 60.135 143.115 60.305 143.875 ;
        RECT 55.450 142.045 56.165 142.215 ;
        RECT 55.450 141.495 55.780 141.875 ;
        RECT 55.995 141.665 56.165 142.045 ;
        RECT 56.425 141.495 58.095 142.265 ;
        RECT 58.730 141.495 58.990 142.335 ;
        RECT 59.165 142.240 59.335 142.970 ;
        RECT 59.590 142.945 60.305 143.115 ;
        RECT 60.565 142.955 61.775 144.045 ;
        RECT 59.590 142.735 59.760 142.945 ;
        RECT 59.505 142.405 59.760 142.735 ;
        RECT 59.165 141.665 59.420 142.240 ;
        RECT 59.590 142.215 59.760 142.405 ;
        RECT 60.040 142.395 60.395 142.765 ;
        RECT 60.565 142.245 61.085 142.785 ;
        RECT 61.255 142.415 61.775 142.955 ;
        RECT 61.945 142.880 62.235 144.045 ;
        RECT 62.870 142.895 63.130 144.045 ;
        RECT 63.305 142.970 63.560 143.875 ;
        RECT 63.730 143.285 64.060 144.045 ;
        RECT 64.275 143.115 64.445 143.875 ;
        RECT 64.705 143.610 70.050 144.045 ;
        RECT 59.590 142.045 60.305 142.215 ;
        RECT 59.590 141.495 59.920 141.875 ;
        RECT 60.135 141.665 60.305 142.045 ;
        RECT 60.565 141.495 61.775 142.245 ;
        RECT 61.945 141.495 62.235 142.220 ;
        RECT 62.870 141.495 63.130 142.335 ;
        RECT 63.305 142.240 63.475 142.970 ;
        RECT 63.730 142.945 64.445 143.115 ;
        RECT 63.730 142.735 63.900 142.945 ;
        RECT 63.645 142.405 63.900 142.735 ;
        RECT 63.305 141.665 63.560 142.240 ;
        RECT 63.730 142.215 63.900 142.405 ;
        RECT 64.180 142.395 64.535 142.765 ;
        RECT 63.730 142.045 64.445 142.215 ;
        RECT 63.730 141.495 64.060 141.875 ;
        RECT 64.275 141.665 64.445 142.045 ;
        RECT 66.290 142.040 66.630 142.870 ;
        RECT 68.110 142.360 68.460 143.610 ;
        RECT 70.225 142.955 73.735 144.045 ;
        RECT 70.225 142.265 71.875 142.785 ;
        RECT 72.045 142.435 73.735 142.955 ;
        RECT 74.825 142.880 75.115 144.045 ;
        RECT 75.290 142.895 75.550 144.045 ;
        RECT 75.725 142.970 75.980 143.875 ;
        RECT 76.150 143.285 76.480 144.045 ;
        RECT 76.695 143.115 76.865 143.875 ;
        RECT 64.705 141.495 70.050 142.040 ;
        RECT 70.225 141.495 73.735 142.265 ;
        RECT 74.825 141.495 75.115 142.220 ;
        RECT 75.290 141.495 75.550 142.335 ;
        RECT 75.725 142.240 75.895 142.970 ;
        RECT 76.150 142.945 76.865 143.115 ;
        RECT 77.675 143.115 77.845 143.875 ;
        RECT 78.025 143.285 78.355 144.045 ;
        RECT 77.675 142.945 78.340 143.115 ;
        RECT 78.525 142.970 78.795 143.875 ;
        RECT 76.150 142.735 76.320 142.945 ;
        RECT 78.170 142.800 78.340 142.945 ;
        RECT 76.065 142.405 76.320 142.735 ;
        RECT 75.725 141.665 75.980 142.240 ;
        RECT 76.150 142.215 76.320 142.405 ;
        RECT 76.600 142.395 76.955 142.765 ;
        RECT 77.605 142.395 77.935 142.765 ;
        RECT 78.170 142.470 78.455 142.800 ;
        RECT 78.170 142.215 78.340 142.470 ;
        RECT 76.150 142.045 76.865 142.215 ;
        RECT 76.150 141.495 76.480 141.875 ;
        RECT 76.695 141.665 76.865 142.045 ;
        RECT 77.675 142.045 78.340 142.215 ;
        RECT 78.625 142.170 78.795 142.970 ;
        RECT 79.515 143.115 79.685 143.875 ;
        RECT 79.900 143.285 80.230 144.045 ;
        RECT 79.515 142.945 80.230 143.115 ;
        RECT 80.400 142.970 80.655 143.875 ;
        RECT 79.425 142.395 79.780 142.765 ;
        RECT 80.060 142.735 80.230 142.945 ;
        RECT 80.060 142.405 80.315 142.735 ;
        RECT 80.060 142.215 80.230 142.405 ;
        RECT 80.485 142.240 80.655 142.970 ;
        RECT 80.830 142.895 81.090 144.045 ;
        RECT 81.265 142.970 81.535 143.875 ;
        RECT 81.705 143.285 82.035 144.045 ;
        RECT 82.215 143.115 82.385 143.875 ;
        RECT 77.675 141.665 77.845 142.045 ;
        RECT 78.025 141.495 78.355 141.875 ;
        RECT 78.535 141.665 78.795 142.170 ;
        RECT 79.515 142.045 80.230 142.215 ;
        RECT 79.515 141.665 79.685 142.045 ;
        RECT 79.900 141.495 80.230 141.875 ;
        RECT 80.400 141.665 80.655 142.240 ;
        RECT 80.830 141.495 81.090 142.335 ;
        RECT 81.265 142.170 81.435 142.970 ;
        RECT 81.720 142.945 82.385 143.115 ;
        RECT 83.655 143.115 83.825 143.875 ;
        RECT 84.040 143.285 84.370 144.045 ;
        RECT 83.655 142.945 84.370 143.115 ;
        RECT 84.540 142.970 84.795 143.875 ;
        RECT 81.720 142.800 81.890 142.945 ;
        RECT 81.605 142.470 81.890 142.800 ;
        RECT 81.720 142.215 81.890 142.470 ;
        RECT 82.125 142.395 82.455 142.765 ;
        RECT 83.565 142.395 83.920 142.765 ;
        RECT 84.200 142.735 84.370 142.945 ;
        RECT 84.200 142.405 84.455 142.735 ;
        RECT 84.200 142.215 84.370 142.405 ;
        RECT 84.625 142.240 84.795 142.970 ;
        RECT 84.970 142.895 85.230 144.045 ;
        RECT 85.405 142.955 87.075 144.045 ;
        RECT 81.265 141.665 81.525 142.170 ;
        RECT 81.720 142.045 82.385 142.215 ;
        RECT 81.705 141.495 82.035 141.875 ;
        RECT 82.215 141.665 82.385 142.045 ;
        RECT 83.655 142.045 84.370 142.215 ;
        RECT 83.655 141.665 83.825 142.045 ;
        RECT 84.040 141.495 84.370 141.875 ;
        RECT 84.540 141.665 84.795 142.240 ;
        RECT 84.970 141.495 85.230 142.335 ;
        RECT 85.405 142.265 86.155 142.785 ;
        RECT 86.325 142.435 87.075 142.955 ;
        RECT 87.705 142.880 87.995 144.045 ;
        RECT 88.165 143.075 88.475 143.875 ;
        RECT 88.645 143.245 88.955 144.045 ;
        RECT 89.125 143.415 89.385 143.875 ;
        RECT 89.555 143.585 89.810 144.045 ;
        RECT 89.985 143.415 90.245 143.875 ;
        RECT 89.125 143.245 90.245 143.415 ;
        RECT 88.165 142.905 89.195 143.075 ;
        RECT 85.405 141.495 87.075 142.265 ;
        RECT 87.705 141.495 87.995 142.220 ;
        RECT 88.165 141.995 88.335 142.905 ;
        RECT 88.505 142.165 88.855 142.735 ;
        RECT 89.025 142.655 89.195 142.905 ;
        RECT 89.985 142.995 90.245 143.245 ;
        RECT 90.415 143.175 90.700 144.045 ;
        RECT 91.395 143.325 91.725 144.045 ;
        RECT 89.985 142.825 90.740 142.995 ;
        RECT 89.025 142.485 90.165 142.655 ;
        RECT 90.335 142.315 90.740 142.825 ;
        RECT 91.385 142.685 91.615 143.025 ;
        RECT 91.905 142.685 92.120 143.800 ;
        RECT 92.315 143.100 92.645 143.875 ;
        RECT 92.815 143.270 93.525 144.045 ;
        RECT 92.315 142.885 93.465 143.100 ;
        RECT 91.385 142.485 91.715 142.685 ;
        RECT 91.905 142.505 92.355 142.685 ;
        RECT 92.025 142.485 92.355 142.505 ;
        RECT 92.525 142.485 92.995 142.715 ;
        RECT 93.180 142.315 93.465 142.885 ;
        RECT 93.695 142.440 93.975 143.875 ;
        RECT 94.235 143.115 94.405 143.875 ;
        RECT 94.620 143.285 94.950 144.045 ;
        RECT 94.235 142.945 94.950 143.115 ;
        RECT 95.120 142.970 95.375 143.875 ;
        RECT 89.090 142.145 90.740 142.315 ;
        RECT 88.165 141.665 88.465 141.995 ;
        RECT 88.635 141.495 88.910 141.975 ;
        RECT 89.090 141.755 89.385 142.145 ;
        RECT 89.555 141.495 89.810 141.975 ;
        RECT 89.985 141.755 90.245 142.145 ;
        RECT 91.385 142.125 92.565 142.315 ;
        RECT 90.415 141.495 90.695 141.975 ;
        RECT 91.385 141.665 91.725 142.125 ;
        RECT 92.235 142.045 92.565 142.125 ;
        RECT 92.755 142.125 93.465 142.315 ;
        RECT 92.755 141.985 93.055 142.125 ;
        RECT 92.740 141.975 93.055 141.985 ;
        RECT 92.730 141.965 93.055 141.975 ;
        RECT 92.720 141.960 93.055 141.965 ;
        RECT 91.895 141.495 92.065 141.955 ;
        RECT 92.715 141.950 93.055 141.960 ;
        RECT 92.710 141.945 93.055 141.950 ;
        RECT 92.705 141.935 93.055 141.945 ;
        RECT 92.700 141.930 93.055 141.935 ;
        RECT 92.695 141.665 93.055 141.930 ;
        RECT 93.295 141.495 93.465 141.955 ;
        RECT 93.635 141.665 93.975 142.440 ;
        RECT 94.145 142.395 94.500 142.765 ;
        RECT 94.780 142.735 94.950 142.945 ;
        RECT 94.780 142.405 95.035 142.735 ;
        RECT 94.780 142.215 94.950 142.405 ;
        RECT 95.205 142.240 95.375 142.970 ;
        RECT 95.550 142.895 95.810 144.045 ;
        RECT 95.990 142.895 96.250 144.045 ;
        RECT 96.425 142.970 96.680 143.875 ;
        RECT 96.850 143.285 97.180 144.045 ;
        RECT 97.395 143.115 97.565 143.875 ;
        RECT 94.235 142.045 94.950 142.215 ;
        RECT 94.235 141.665 94.405 142.045 ;
        RECT 94.620 141.495 94.950 141.875 ;
        RECT 95.120 141.665 95.375 142.240 ;
        RECT 95.550 141.495 95.810 142.335 ;
        RECT 95.990 141.495 96.250 142.335 ;
        RECT 96.425 142.240 96.595 142.970 ;
        RECT 96.850 142.945 97.565 143.115 ;
        RECT 97.825 142.955 100.415 144.045 ;
        RECT 96.850 142.735 97.020 142.945 ;
        RECT 96.765 142.405 97.020 142.735 ;
        RECT 96.425 141.665 96.680 142.240 ;
        RECT 96.850 142.215 97.020 142.405 ;
        RECT 97.300 142.395 97.655 142.765 ;
        RECT 97.825 142.265 99.035 142.785 ;
        RECT 99.205 142.435 100.415 142.955 ;
        RECT 100.585 142.880 100.875 144.045 ;
        RECT 101.135 143.115 101.305 143.875 ;
        RECT 101.520 143.285 101.850 144.045 ;
        RECT 101.135 142.945 101.850 143.115 ;
        RECT 102.020 142.970 102.275 143.875 ;
        RECT 101.045 142.395 101.400 142.765 ;
        RECT 101.680 142.735 101.850 142.945 ;
        RECT 101.680 142.405 101.935 142.735 ;
        RECT 96.850 142.045 97.565 142.215 ;
        RECT 96.850 141.495 97.180 141.875 ;
        RECT 97.395 141.665 97.565 142.045 ;
        RECT 97.825 141.495 100.415 142.265 ;
        RECT 100.585 141.495 100.875 142.220 ;
        RECT 101.680 142.215 101.850 142.405 ;
        RECT 102.105 142.240 102.275 142.970 ;
        RECT 102.450 142.895 102.710 144.045 ;
        RECT 102.885 142.955 104.095 144.045 ;
        RECT 101.135 142.045 101.850 142.215 ;
        RECT 101.135 141.665 101.305 142.045 ;
        RECT 101.520 141.495 101.850 141.875 ;
        RECT 102.020 141.665 102.275 142.240 ;
        RECT 102.450 141.495 102.710 142.335 ;
        RECT 102.885 142.245 103.405 142.785 ;
        RECT 103.575 142.415 104.095 142.955 ;
        RECT 104.270 142.895 104.530 144.045 ;
        RECT 104.705 142.970 104.960 143.875 ;
        RECT 105.130 143.285 105.460 144.045 ;
        RECT 105.675 143.115 105.845 143.875 ;
        RECT 106.105 143.610 111.450 144.045 ;
        RECT 102.885 141.495 104.095 142.245 ;
        RECT 104.270 141.495 104.530 142.335 ;
        RECT 104.705 142.240 104.875 142.970 ;
        RECT 105.130 142.945 105.845 143.115 ;
        RECT 105.130 142.735 105.300 142.945 ;
        RECT 105.045 142.405 105.300 142.735 ;
        RECT 104.705 141.665 104.960 142.240 ;
        RECT 105.130 142.215 105.300 142.405 ;
        RECT 105.580 142.395 105.935 142.765 ;
        RECT 105.130 142.045 105.845 142.215 ;
        RECT 105.130 141.495 105.460 141.875 ;
        RECT 105.675 141.665 105.845 142.045 ;
        RECT 107.690 142.040 108.030 142.870 ;
        RECT 109.510 142.360 109.860 143.610 ;
        RECT 111.625 142.955 113.295 144.045 ;
        RECT 111.625 142.265 112.375 142.785 ;
        RECT 112.545 142.435 113.295 142.955 ;
        RECT 113.465 142.880 113.755 144.045 ;
        RECT 113.935 143.325 114.265 144.045 ;
        RECT 113.925 142.685 114.155 143.025 ;
        RECT 114.445 142.685 114.660 143.800 ;
        RECT 114.855 143.100 115.185 143.875 ;
        RECT 115.355 143.270 116.065 144.045 ;
        RECT 114.855 142.885 116.005 143.100 ;
        RECT 113.925 142.485 114.255 142.685 ;
        RECT 114.445 142.505 114.895 142.685 ;
        RECT 114.565 142.485 114.895 142.505 ;
        RECT 115.065 142.485 115.535 142.715 ;
        RECT 115.720 142.315 116.005 142.885 ;
        RECT 116.235 142.440 116.515 143.875 ;
        RECT 116.775 143.115 116.945 143.875 ;
        RECT 117.160 143.285 117.490 144.045 ;
        RECT 116.775 142.945 117.490 143.115 ;
        RECT 117.660 142.970 117.915 143.875 ;
        RECT 106.105 141.495 111.450 142.040 ;
        RECT 111.625 141.495 113.295 142.265 ;
        RECT 113.465 141.495 113.755 142.220 ;
        RECT 113.925 142.125 115.105 142.315 ;
        RECT 113.925 141.665 114.265 142.125 ;
        RECT 114.775 142.045 115.105 142.125 ;
        RECT 115.295 142.125 116.005 142.315 ;
        RECT 115.295 141.985 115.595 142.125 ;
        RECT 115.280 141.975 115.595 141.985 ;
        RECT 115.270 141.965 115.595 141.975 ;
        RECT 115.260 141.960 115.595 141.965 ;
        RECT 114.435 141.495 114.605 141.955 ;
        RECT 115.255 141.950 115.595 141.960 ;
        RECT 115.250 141.945 115.595 141.950 ;
        RECT 115.245 141.935 115.595 141.945 ;
        RECT 115.240 141.930 115.595 141.935 ;
        RECT 115.235 141.665 115.595 141.930 ;
        RECT 115.835 141.495 116.005 141.955 ;
        RECT 116.175 141.665 116.515 142.440 ;
        RECT 116.685 142.395 117.040 142.765 ;
        RECT 117.320 142.735 117.490 142.945 ;
        RECT 117.320 142.405 117.575 142.735 ;
        RECT 117.320 142.215 117.490 142.405 ;
        RECT 117.745 142.240 117.915 142.970 ;
        RECT 118.090 142.895 118.350 144.045 ;
        RECT 118.525 142.955 120.195 144.045 ;
        RECT 116.775 142.045 117.490 142.215 ;
        RECT 116.775 141.665 116.945 142.045 ;
        RECT 117.160 141.495 117.490 141.875 ;
        RECT 117.660 141.665 117.915 142.240 ;
        RECT 118.090 141.495 118.350 142.335 ;
        RECT 118.525 142.265 119.275 142.785 ;
        RECT 119.445 142.435 120.195 142.955 ;
        RECT 120.915 143.115 121.085 143.875 ;
        RECT 121.300 143.285 121.630 144.045 ;
        RECT 120.915 142.945 121.630 143.115 ;
        RECT 121.800 142.970 122.055 143.875 ;
        RECT 120.825 142.395 121.180 142.765 ;
        RECT 121.460 142.735 121.630 142.945 ;
        RECT 121.460 142.405 121.715 142.735 ;
        RECT 118.525 141.495 120.195 142.265 ;
        RECT 121.460 142.215 121.630 142.405 ;
        RECT 121.885 142.240 122.055 142.970 ;
        RECT 122.230 142.895 122.490 144.045 ;
        RECT 122.665 142.955 124.335 144.045 ;
        RECT 120.915 142.045 121.630 142.215 ;
        RECT 120.915 141.665 121.085 142.045 ;
        RECT 121.300 141.495 121.630 141.875 ;
        RECT 121.800 141.665 122.055 142.240 ;
        RECT 122.230 141.495 122.490 142.335 ;
        RECT 122.665 142.265 123.415 142.785 ;
        RECT 123.585 142.435 124.335 142.955 ;
        RECT 124.595 143.115 124.765 143.875 ;
        RECT 124.980 143.285 125.310 144.045 ;
        RECT 124.595 142.945 125.310 143.115 ;
        RECT 125.480 142.970 125.735 143.875 ;
        RECT 124.505 142.395 124.860 142.765 ;
        RECT 125.140 142.735 125.310 142.945 ;
        RECT 125.140 142.405 125.395 142.735 ;
        RECT 122.665 141.495 124.335 142.265 ;
        RECT 125.140 142.215 125.310 142.405 ;
        RECT 125.565 142.240 125.735 142.970 ;
        RECT 125.910 142.895 126.170 144.045 ;
        RECT 126.345 142.880 126.635 144.045 ;
        RECT 126.815 143.325 127.145 144.045 ;
        RECT 126.805 142.685 127.035 143.025 ;
        RECT 127.325 142.685 127.540 143.800 ;
        RECT 127.735 143.100 128.065 143.875 ;
        RECT 128.235 143.270 128.945 144.045 ;
        RECT 127.735 142.885 128.885 143.100 ;
        RECT 126.805 142.485 127.135 142.685 ;
        RECT 127.325 142.505 127.775 142.685 ;
        RECT 127.445 142.485 127.775 142.505 ;
        RECT 127.945 142.485 128.415 142.715 ;
        RECT 124.595 142.045 125.310 142.215 ;
        RECT 124.595 141.665 124.765 142.045 ;
        RECT 124.980 141.495 125.310 141.875 ;
        RECT 125.480 141.665 125.735 142.240 ;
        RECT 125.910 141.495 126.170 142.335 ;
        RECT 128.600 142.315 128.885 142.885 ;
        RECT 129.115 142.440 129.395 143.875 ;
        RECT 126.345 141.495 126.635 142.220 ;
        RECT 126.805 142.125 127.985 142.315 ;
        RECT 126.805 141.665 127.145 142.125 ;
        RECT 127.655 142.045 127.985 142.125 ;
        RECT 128.175 142.125 128.885 142.315 ;
        RECT 128.175 141.985 128.475 142.125 ;
        RECT 128.160 141.975 128.475 141.985 ;
        RECT 128.150 141.965 128.475 141.975 ;
        RECT 128.140 141.960 128.475 141.965 ;
        RECT 127.315 141.495 127.485 141.955 ;
        RECT 128.135 141.950 128.475 141.960 ;
        RECT 128.130 141.945 128.475 141.950 ;
        RECT 128.125 141.935 128.475 141.945 ;
        RECT 128.120 141.930 128.475 141.935 ;
        RECT 128.115 141.665 128.475 141.930 ;
        RECT 128.715 141.495 128.885 141.955 ;
        RECT 129.055 141.665 129.395 142.440 ;
        RECT 129.565 143.075 129.875 143.875 ;
        RECT 130.045 143.245 130.355 144.045 ;
        RECT 130.525 143.415 130.785 143.875 ;
        RECT 130.955 143.585 131.210 144.045 ;
        RECT 131.385 143.415 131.645 143.875 ;
        RECT 130.525 143.245 131.645 143.415 ;
        RECT 129.565 142.905 130.595 143.075 ;
        RECT 129.565 141.995 129.735 142.905 ;
        RECT 129.905 142.165 130.255 142.735 ;
        RECT 130.425 142.655 130.595 142.905 ;
        RECT 131.385 142.995 131.645 143.245 ;
        RECT 131.815 143.175 132.100 144.045 ;
        RECT 133.335 143.115 133.505 143.875 ;
        RECT 133.720 143.285 134.050 144.045 ;
        RECT 131.385 142.825 132.140 142.995 ;
        RECT 133.335 142.945 134.050 143.115 ;
        RECT 134.220 142.970 134.475 143.875 ;
        RECT 130.425 142.485 131.565 142.655 ;
        RECT 131.735 142.315 132.140 142.825 ;
        RECT 133.245 142.395 133.600 142.765 ;
        RECT 133.880 142.735 134.050 142.945 ;
        RECT 133.880 142.405 134.135 142.735 ;
        RECT 130.490 142.145 132.140 142.315 ;
        RECT 133.880 142.215 134.050 142.405 ;
        RECT 134.305 142.240 134.475 142.970 ;
        RECT 134.650 142.895 134.910 144.045 ;
        RECT 135.085 142.955 136.755 144.045 ;
        RECT 129.565 141.665 129.865 141.995 ;
        RECT 130.035 141.495 130.310 141.975 ;
        RECT 130.490 141.755 130.785 142.145 ;
        RECT 130.955 141.495 131.210 141.975 ;
        RECT 131.385 141.755 131.645 142.145 ;
        RECT 133.335 142.045 134.050 142.215 ;
        RECT 131.815 141.495 132.095 141.975 ;
        RECT 133.335 141.665 133.505 142.045 ;
        RECT 133.720 141.495 134.050 141.875 ;
        RECT 134.220 141.665 134.475 142.240 ;
        RECT 134.650 141.495 134.910 142.335 ;
        RECT 135.085 142.265 135.835 142.785 ;
        RECT 136.005 142.435 136.755 142.955 ;
        RECT 137.475 143.115 137.645 143.875 ;
        RECT 137.860 143.285 138.190 144.045 ;
        RECT 137.475 142.945 138.190 143.115 ;
        RECT 138.360 142.970 138.615 143.875 ;
        RECT 137.385 142.395 137.740 142.765 ;
        RECT 138.020 142.735 138.190 142.945 ;
        RECT 138.020 142.405 138.275 142.735 ;
        RECT 135.085 141.495 136.755 142.265 ;
        RECT 138.020 142.215 138.190 142.405 ;
        RECT 138.445 142.240 138.615 142.970 ;
        RECT 138.790 142.895 139.050 144.045 ;
        RECT 139.225 142.880 139.515 144.045 ;
        RECT 140.145 143.205 140.575 144.045 ;
        RECT 141.165 143.545 141.415 144.045 ;
        RECT 141.685 143.705 142.810 143.875 ;
        RECT 141.685 143.545 141.935 143.705 ;
        RECT 142.485 143.535 142.810 143.705 ;
        RECT 142.980 143.545 143.230 144.045 ;
        RECT 143.400 143.535 143.650 143.875 ;
        RECT 140.745 143.375 140.995 143.535 ;
        RECT 142.105 143.375 142.315 143.535 ;
        RECT 140.745 143.205 142.315 143.375 ;
        RECT 143.960 143.375 144.210 143.875 ;
        RECT 144.380 143.545 144.630 144.045 ;
        RECT 144.800 143.375 145.050 143.875 ;
        RECT 145.220 143.545 145.470 144.045 ;
        RECT 145.640 143.375 145.955 143.875 ;
        RECT 143.960 143.365 145.955 143.375 ;
        RECT 140.745 143.035 140.995 143.205 ;
        RECT 142.560 143.195 145.955 143.365 ;
        RECT 142.560 143.035 142.730 143.195 ;
        RECT 140.145 142.825 140.995 143.035 ;
        RECT 141.235 142.865 142.730 143.035 ;
        RECT 137.475 142.045 138.190 142.215 ;
        RECT 137.475 141.665 137.645 142.045 ;
        RECT 137.860 141.495 138.190 141.875 ;
        RECT 138.360 141.665 138.615 142.240 ;
        RECT 138.790 141.495 139.050 142.335 ;
        RECT 139.225 141.495 139.515 142.220 ;
        RECT 140.145 141.885 140.535 142.825 ;
        RECT 141.235 142.655 141.405 142.865 ;
        RECT 142.940 142.855 145.250 143.025 ;
        RECT 142.940 142.695 143.110 142.855 ;
        RECT 140.745 142.485 141.405 142.655 ;
        RECT 142.085 142.485 143.110 142.695 ;
        RECT 145.080 142.695 145.250 142.855 ;
        RECT 143.335 142.485 144.785 142.685 ;
        RECT 145.080 142.485 145.555 142.695 ;
        RECT 140.705 142.135 143.270 142.315 ;
        RECT 140.705 142.055 141.035 142.135 ;
        RECT 140.145 141.715 141.455 141.885 ;
        RECT 141.725 141.495 141.895 141.965 ;
        RECT 142.065 141.665 142.430 142.135 ;
        RECT 142.600 141.495 142.770 141.965 ;
        RECT 142.940 141.665 143.270 142.135 ;
        RECT 143.440 141.495 143.610 142.315 ;
        RECT 143.920 142.135 145.010 142.315 ;
        RECT 145.725 142.305 145.955 143.195 ;
        RECT 146.215 143.115 146.385 143.875 ;
        RECT 146.600 143.285 146.930 144.045 ;
        RECT 146.215 142.945 146.930 143.115 ;
        RECT 147.100 142.970 147.355 143.875 ;
        RECT 146.125 142.395 146.480 142.765 ;
        RECT 146.760 142.735 146.930 142.945 ;
        RECT 146.760 142.405 147.015 142.735 ;
        RECT 143.920 141.665 144.250 142.135 ;
        RECT 144.420 141.495 144.590 141.965 ;
        RECT 144.760 141.885 145.010 142.135 ;
        RECT 145.180 142.055 145.955 142.305 ;
        RECT 146.760 142.215 146.930 142.405 ;
        RECT 147.185 142.240 147.355 142.970 ;
        RECT 147.530 142.895 147.790 144.045 ;
        RECT 148.885 142.955 150.095 144.045 ;
        RECT 148.885 142.415 149.405 142.955 ;
        RECT 146.215 142.045 146.930 142.215 ;
        RECT 144.760 141.665 145.935 141.885 ;
        RECT 146.215 141.665 146.385 142.045 ;
        RECT 146.600 141.495 146.930 141.875 ;
        RECT 147.100 141.665 147.355 142.240 ;
        RECT 147.530 141.495 147.790 142.335 ;
        RECT 149.575 142.245 150.095 142.785 ;
        RECT 148.885 141.495 150.095 142.245 ;
        RECT 36.100 141.325 150.180 141.495 ;
        RECT 34.110 128.480 36.100 128.650 ;
        RECT 34.110 104.970 34.280 128.480 ;
        RECT 34.760 125.840 35.450 128.000 ;
        RECT 35.930 104.970 36.100 128.480 ;
        RECT 38.110 128.480 40.100 128.650 ;
        RECT 38.110 104.970 38.280 128.480 ;
        RECT 38.760 125.840 39.450 128.000 ;
        RECT 39.930 104.970 40.100 128.480 ;
        RECT 42.110 128.480 44.100 128.650 ;
        RECT 42.110 104.970 42.280 128.480 ;
        RECT 42.760 125.840 43.450 128.000 ;
        RECT 43.930 104.970 44.100 128.480 ;
        RECT 46.110 128.480 48.100 128.650 ;
        RECT 46.110 104.970 46.280 128.480 ;
        RECT 46.760 125.840 47.450 128.000 ;
        RECT 47.930 104.970 48.100 128.480 ;
        RECT 50.110 128.480 52.100 128.650 ;
        RECT 50.110 104.970 50.280 128.480 ;
        RECT 50.760 125.840 51.450 128.000 ;
        RECT 51.930 104.970 52.100 128.480 ;
        RECT 54.110 128.480 56.100 128.650 ;
        RECT 54.110 104.970 54.280 128.480 ;
        RECT 54.760 125.840 55.450 128.000 ;
        RECT 55.930 104.970 56.100 128.480 ;
        RECT 58.110 128.480 60.100 128.650 ;
        RECT 58.110 104.970 58.280 128.480 ;
        RECT 58.760 125.840 59.450 128.000 ;
        RECT 59.930 104.970 60.100 128.480 ;
        RECT 62.110 128.480 64.100 128.650 ;
        RECT 62.110 104.970 62.280 128.480 ;
        RECT 62.760 125.840 63.450 128.000 ;
        RECT 63.930 104.970 64.100 128.480 ;
        RECT 75.110 128.480 77.100 128.650 ;
        RECT 75.110 104.970 75.280 128.480 ;
        RECT 75.760 125.840 76.450 128.000 ;
        RECT 76.930 104.970 77.100 128.480 ;
        RECT 79.110 128.480 81.100 128.650 ;
        RECT 79.110 104.970 79.280 128.480 ;
        RECT 79.760 125.840 80.450 128.000 ;
        RECT 80.930 104.970 81.100 128.480 ;
        RECT 83.110 128.480 85.100 128.650 ;
        RECT 83.110 104.970 83.280 128.480 ;
        RECT 83.760 125.840 84.450 128.000 ;
        RECT 84.930 104.970 85.100 128.480 ;
        RECT 87.110 128.480 89.100 128.650 ;
        RECT 87.110 104.970 87.280 128.480 ;
        RECT 87.760 125.840 88.450 128.000 ;
        RECT 88.930 104.970 89.100 128.480 ;
        RECT 91.110 128.480 93.100 128.650 ;
        RECT 91.110 104.970 91.280 128.480 ;
        RECT 91.760 125.840 92.450 128.000 ;
        RECT 92.930 104.970 93.100 128.480 ;
        RECT 95.110 128.480 97.100 128.650 ;
        RECT 95.110 104.970 95.280 128.480 ;
        RECT 95.760 125.840 96.450 128.000 ;
        RECT 96.930 104.970 97.100 128.480 ;
        RECT 99.110 128.480 101.100 128.650 ;
        RECT 99.110 104.970 99.280 128.480 ;
        RECT 99.760 125.840 100.450 128.000 ;
        RECT 100.930 104.970 101.100 128.480 ;
        RECT 103.110 128.480 105.100 128.650 ;
        RECT 103.110 104.970 103.280 128.480 ;
        RECT 103.760 125.840 104.450 128.000 ;
        RECT 104.930 104.970 105.100 128.480 ;
        RECT 116.110 128.480 118.100 128.650 ;
        RECT 116.110 104.970 116.280 128.480 ;
        RECT 116.760 125.840 117.450 128.000 ;
        RECT 117.930 104.970 118.100 128.480 ;
        RECT 120.110 128.480 122.100 128.650 ;
        RECT 120.110 104.970 120.280 128.480 ;
        RECT 120.760 125.840 121.450 128.000 ;
        RECT 121.930 104.970 122.100 128.480 ;
        RECT 124.110 128.480 126.100 128.650 ;
        RECT 124.110 104.970 124.280 128.480 ;
        RECT 124.760 125.840 125.450 128.000 ;
        RECT 125.930 104.970 126.100 128.480 ;
        RECT 128.110 128.480 130.100 128.650 ;
        RECT 128.110 104.970 128.280 128.480 ;
        RECT 128.760 125.840 129.450 128.000 ;
        RECT 129.930 104.970 130.100 128.480 ;
        RECT 132.110 128.480 134.100 128.650 ;
        RECT 132.110 104.970 132.280 128.480 ;
        RECT 132.760 125.840 133.450 128.000 ;
        RECT 133.930 104.970 134.100 128.480 ;
        RECT 136.110 128.480 138.100 128.650 ;
        RECT 136.110 104.970 136.280 128.480 ;
        RECT 136.760 125.840 137.450 128.000 ;
        RECT 137.930 104.970 138.100 128.480 ;
        RECT 140.110 128.480 142.100 128.650 ;
        RECT 140.110 104.970 140.280 128.480 ;
        RECT 140.760 125.840 141.450 128.000 ;
        RECT 141.930 104.970 142.100 128.480 ;
        RECT 144.110 128.480 146.100 128.650 ;
        RECT 144.110 104.970 144.280 128.480 ;
        RECT 144.760 125.840 145.450 128.000 ;
        RECT 145.930 104.970 146.100 128.480 ;
        RECT 34.030 104.170 34.370 104.970 ;
        RECT 35.830 104.170 36.170 104.970 ;
        RECT 38.030 104.170 38.370 104.970 ;
        RECT 39.830 104.170 40.170 104.970 ;
        RECT 42.030 104.170 42.370 104.970 ;
        RECT 43.830 104.170 44.170 104.970 ;
        RECT 46.030 104.170 46.370 104.970 ;
        RECT 47.830 104.170 48.170 104.970 ;
        RECT 50.030 104.170 50.370 104.970 ;
        RECT 51.830 104.170 52.170 104.970 ;
        RECT 54.030 104.170 54.370 104.970 ;
        RECT 55.830 104.170 56.170 104.970 ;
        RECT 58.030 104.170 58.370 104.970 ;
        RECT 59.830 104.170 60.170 104.970 ;
        RECT 62.030 104.170 62.370 104.970 ;
        RECT 63.830 104.170 64.170 104.970 ;
        RECT 75.030 104.170 75.370 104.970 ;
        RECT 76.830 104.170 77.170 104.970 ;
        RECT 79.030 104.170 79.370 104.970 ;
        RECT 80.830 104.170 81.170 104.970 ;
        RECT 83.030 104.170 83.370 104.970 ;
        RECT 84.830 104.170 85.170 104.970 ;
        RECT 87.030 104.170 87.370 104.970 ;
        RECT 88.830 104.170 89.170 104.970 ;
        RECT 91.030 104.170 91.370 104.970 ;
        RECT 92.830 104.170 93.170 104.970 ;
        RECT 95.030 104.170 95.370 104.970 ;
        RECT 96.830 104.170 97.170 104.970 ;
        RECT 99.030 104.170 99.370 104.970 ;
        RECT 100.830 104.170 101.170 104.970 ;
        RECT 103.030 104.170 103.370 104.970 ;
        RECT 104.830 104.170 105.170 104.970 ;
        RECT 116.030 104.170 116.370 104.970 ;
        RECT 117.830 104.170 118.170 104.970 ;
        RECT 120.030 104.170 120.370 104.970 ;
        RECT 121.830 104.170 122.170 104.970 ;
        RECT 124.030 104.170 124.370 104.970 ;
        RECT 125.830 104.170 126.170 104.970 ;
        RECT 128.030 104.170 128.370 104.970 ;
        RECT 129.830 104.170 130.170 104.970 ;
        RECT 132.030 104.170 132.370 104.970 ;
        RECT 133.830 104.170 134.170 104.970 ;
        RECT 136.030 104.170 136.370 104.970 ;
        RECT 137.830 104.170 138.170 104.970 ;
        RECT 140.030 104.170 140.370 104.970 ;
        RECT 141.830 104.170 142.170 104.970 ;
        RECT 144.030 104.170 144.370 104.970 ;
        RECT 145.830 104.170 146.170 104.970 ;
        RECT 34.110 83.460 34.280 104.170 ;
        RECT 34.760 83.940 35.450 86.100 ;
        RECT 35.930 83.460 36.100 104.170 ;
        RECT 34.110 83.290 36.100 83.460 ;
        RECT 38.110 83.460 38.280 104.170 ;
        RECT 38.760 83.940 39.450 86.100 ;
        RECT 39.930 83.460 40.100 104.170 ;
        RECT 38.110 83.290 40.100 83.460 ;
        RECT 42.110 83.460 42.280 104.170 ;
        RECT 42.760 83.940 43.450 86.100 ;
        RECT 43.930 83.460 44.100 104.170 ;
        RECT 42.110 83.290 44.100 83.460 ;
        RECT 46.110 83.460 46.280 104.170 ;
        RECT 46.760 83.940 47.450 86.100 ;
        RECT 47.930 83.460 48.100 104.170 ;
        RECT 46.110 83.290 48.100 83.460 ;
        RECT 50.110 83.460 50.280 104.170 ;
        RECT 50.760 83.940 51.450 86.100 ;
        RECT 51.930 83.460 52.100 104.170 ;
        RECT 50.110 83.290 52.100 83.460 ;
        RECT 54.110 83.460 54.280 104.170 ;
        RECT 54.760 83.940 55.450 86.100 ;
        RECT 55.930 83.460 56.100 104.170 ;
        RECT 54.110 83.290 56.100 83.460 ;
        RECT 58.110 83.460 58.280 104.170 ;
        RECT 58.760 83.940 59.450 86.100 ;
        RECT 59.930 83.460 60.100 104.170 ;
        RECT 58.110 83.290 60.100 83.460 ;
        RECT 62.110 83.460 62.280 104.170 ;
        RECT 62.760 83.940 63.450 86.100 ;
        RECT 63.930 83.460 64.100 104.170 ;
        RECT 62.110 83.290 64.100 83.460 ;
        RECT 75.110 83.460 75.280 104.170 ;
        RECT 75.760 83.940 76.450 86.100 ;
        RECT 76.930 83.460 77.100 104.170 ;
        RECT 75.110 83.290 77.100 83.460 ;
        RECT 79.110 83.460 79.280 104.170 ;
        RECT 79.760 83.940 80.450 86.100 ;
        RECT 80.930 83.460 81.100 104.170 ;
        RECT 79.110 83.290 81.100 83.460 ;
        RECT 83.110 83.460 83.280 104.170 ;
        RECT 83.760 83.940 84.450 86.100 ;
        RECT 84.930 83.460 85.100 104.170 ;
        RECT 83.110 83.290 85.100 83.460 ;
        RECT 87.110 83.460 87.280 104.170 ;
        RECT 87.760 83.940 88.450 86.100 ;
        RECT 88.930 83.460 89.100 104.170 ;
        RECT 87.110 83.290 89.100 83.460 ;
        RECT 91.110 83.460 91.280 104.170 ;
        RECT 91.760 83.940 92.450 86.100 ;
        RECT 92.930 83.460 93.100 104.170 ;
        RECT 91.110 83.290 93.100 83.460 ;
        RECT 95.110 83.460 95.280 104.170 ;
        RECT 95.760 83.940 96.450 86.100 ;
        RECT 96.930 83.460 97.100 104.170 ;
        RECT 95.110 83.290 97.100 83.460 ;
        RECT 99.110 83.460 99.280 104.170 ;
        RECT 99.760 83.940 100.450 86.100 ;
        RECT 100.930 83.460 101.100 104.170 ;
        RECT 99.110 83.290 101.100 83.460 ;
        RECT 103.110 83.460 103.280 104.170 ;
        RECT 103.760 83.940 104.450 86.100 ;
        RECT 104.930 83.460 105.100 104.170 ;
        RECT 103.110 83.290 105.100 83.460 ;
        RECT 116.110 83.460 116.280 104.170 ;
        RECT 116.760 83.940 117.450 86.100 ;
        RECT 117.930 83.460 118.100 104.170 ;
        RECT 116.110 83.290 118.100 83.460 ;
        RECT 120.110 83.460 120.280 104.170 ;
        RECT 120.760 83.940 121.450 86.100 ;
        RECT 121.930 83.460 122.100 104.170 ;
        RECT 120.110 83.290 122.100 83.460 ;
        RECT 124.110 83.460 124.280 104.170 ;
        RECT 124.760 83.940 125.450 86.100 ;
        RECT 125.930 83.460 126.100 104.170 ;
        RECT 124.110 83.290 126.100 83.460 ;
        RECT 128.110 83.460 128.280 104.170 ;
        RECT 128.760 83.940 129.450 86.100 ;
        RECT 129.930 83.460 130.100 104.170 ;
        RECT 128.110 83.290 130.100 83.460 ;
        RECT 132.110 83.460 132.280 104.170 ;
        RECT 132.760 83.940 133.450 86.100 ;
        RECT 133.930 83.460 134.100 104.170 ;
        RECT 132.110 83.290 134.100 83.460 ;
        RECT 136.110 83.460 136.280 104.170 ;
        RECT 136.760 83.940 137.450 86.100 ;
        RECT 137.930 83.460 138.100 104.170 ;
        RECT 136.110 83.290 138.100 83.460 ;
        RECT 140.110 83.460 140.280 104.170 ;
        RECT 140.760 83.940 141.450 86.100 ;
        RECT 141.930 83.460 142.100 104.170 ;
        RECT 140.110 83.290 142.100 83.460 ;
        RECT 144.110 83.460 144.280 104.170 ;
        RECT 144.760 83.940 145.450 86.100 ;
        RECT 145.930 83.460 146.100 104.170 ;
        RECT 144.110 83.290 146.100 83.460 ;
        RECT 34.110 80.480 36.100 80.650 ;
        RECT 34.110 55.810 34.280 80.480 ;
        RECT 34.760 77.840 35.450 80.000 ;
        RECT 34.760 56.290 35.450 58.450 ;
        RECT 34.480 55.810 35.740 55.900 ;
        RECT 35.930 55.810 36.100 80.480 ;
        RECT 34.110 55.640 36.100 55.810 ;
        RECT 38.110 80.480 40.100 80.650 ;
        RECT 38.110 55.810 38.280 80.480 ;
        RECT 38.760 77.840 39.450 80.000 ;
        RECT 38.760 56.290 39.450 58.450 ;
        RECT 38.480 55.810 39.740 55.900 ;
        RECT 39.930 55.810 40.100 80.480 ;
        RECT 38.110 55.640 40.100 55.810 ;
        RECT 42.110 80.480 44.100 80.650 ;
        RECT 42.110 55.810 42.280 80.480 ;
        RECT 42.760 77.840 43.450 80.000 ;
        RECT 42.760 56.290 43.450 58.450 ;
        RECT 42.480 55.810 43.740 55.900 ;
        RECT 43.930 55.810 44.100 80.480 ;
        RECT 42.110 55.640 44.100 55.810 ;
        RECT 46.110 80.480 48.100 80.650 ;
        RECT 46.110 55.810 46.280 80.480 ;
        RECT 46.760 77.840 47.450 80.000 ;
        RECT 46.760 56.290 47.450 58.450 ;
        RECT 46.480 55.810 47.740 55.900 ;
        RECT 47.930 55.810 48.100 80.480 ;
        RECT 46.110 55.640 48.100 55.810 ;
        RECT 50.110 80.480 52.100 80.650 ;
        RECT 50.110 55.810 50.280 80.480 ;
        RECT 50.760 77.840 51.450 80.000 ;
        RECT 50.760 56.290 51.450 58.450 ;
        RECT 50.480 55.810 51.740 55.900 ;
        RECT 51.930 55.810 52.100 80.480 ;
        RECT 50.110 55.640 52.100 55.810 ;
        RECT 54.110 80.480 56.100 80.650 ;
        RECT 54.110 55.810 54.280 80.480 ;
        RECT 54.760 77.840 55.450 80.000 ;
        RECT 54.760 56.290 55.450 58.450 ;
        RECT 54.480 55.810 55.740 55.900 ;
        RECT 55.930 55.810 56.100 80.480 ;
        RECT 54.110 55.640 56.100 55.810 ;
        RECT 58.110 80.480 60.100 80.650 ;
        RECT 58.110 55.810 58.280 80.480 ;
        RECT 58.760 77.840 59.450 80.000 ;
        RECT 58.760 56.290 59.450 58.450 ;
        RECT 58.480 55.810 59.740 55.900 ;
        RECT 59.930 55.810 60.100 80.480 ;
        RECT 58.110 55.640 60.100 55.810 ;
        RECT 62.110 80.480 64.100 80.650 ;
        RECT 62.110 55.810 62.280 80.480 ;
        RECT 62.760 77.840 63.450 80.000 ;
        RECT 62.760 56.290 63.450 58.450 ;
        RECT 62.480 55.810 63.740 55.900 ;
        RECT 63.930 55.810 64.100 80.480 ;
        RECT 62.110 55.640 64.100 55.810 ;
        RECT 75.110 80.480 77.100 80.650 ;
        RECT 75.110 55.810 75.280 80.480 ;
        RECT 75.760 77.840 76.450 80.000 ;
        RECT 75.760 56.290 76.450 58.450 ;
        RECT 75.480 55.810 76.740 55.900 ;
        RECT 76.930 55.810 77.100 80.480 ;
        RECT 75.110 55.640 77.100 55.810 ;
        RECT 79.110 80.480 81.100 80.650 ;
        RECT 79.110 55.810 79.280 80.480 ;
        RECT 79.760 77.840 80.450 80.000 ;
        RECT 79.760 56.290 80.450 58.450 ;
        RECT 79.480 55.810 80.740 55.900 ;
        RECT 80.930 55.810 81.100 80.480 ;
        RECT 79.110 55.640 81.100 55.810 ;
        RECT 83.110 80.480 85.100 80.650 ;
        RECT 83.110 55.810 83.280 80.480 ;
        RECT 83.760 77.840 84.450 80.000 ;
        RECT 83.760 56.290 84.450 58.450 ;
        RECT 83.480 55.810 84.740 55.900 ;
        RECT 84.930 55.810 85.100 80.480 ;
        RECT 83.110 55.640 85.100 55.810 ;
        RECT 87.110 80.480 89.100 80.650 ;
        RECT 87.110 55.810 87.280 80.480 ;
        RECT 87.760 77.840 88.450 80.000 ;
        RECT 87.760 56.290 88.450 58.450 ;
        RECT 87.480 55.810 88.740 55.900 ;
        RECT 88.930 55.810 89.100 80.480 ;
        RECT 87.110 55.640 89.100 55.810 ;
        RECT 91.110 80.480 93.100 80.650 ;
        RECT 91.110 55.810 91.280 80.480 ;
        RECT 91.760 77.840 92.450 80.000 ;
        RECT 91.760 56.290 92.450 58.450 ;
        RECT 91.480 55.810 92.740 55.900 ;
        RECT 92.930 55.810 93.100 80.480 ;
        RECT 91.110 55.640 93.100 55.810 ;
        RECT 95.110 80.480 97.100 80.650 ;
        RECT 95.110 55.810 95.280 80.480 ;
        RECT 95.760 77.840 96.450 80.000 ;
        RECT 95.760 56.290 96.450 58.450 ;
        RECT 95.480 55.810 96.740 55.900 ;
        RECT 96.930 55.810 97.100 80.480 ;
        RECT 95.110 55.640 97.100 55.810 ;
        RECT 99.110 80.480 101.100 80.650 ;
        RECT 99.110 55.810 99.280 80.480 ;
        RECT 99.760 77.840 100.450 80.000 ;
        RECT 99.760 56.290 100.450 58.450 ;
        RECT 99.480 55.810 100.740 55.900 ;
        RECT 100.930 55.810 101.100 80.480 ;
        RECT 99.110 55.640 101.100 55.810 ;
        RECT 103.110 80.480 105.100 80.650 ;
        RECT 103.110 55.810 103.280 80.480 ;
        RECT 103.760 77.840 104.450 80.000 ;
        RECT 103.760 56.290 104.450 58.450 ;
        RECT 103.480 55.810 104.740 55.900 ;
        RECT 104.930 55.810 105.100 80.480 ;
        RECT 103.110 55.640 105.100 55.810 ;
        RECT 116.110 80.480 118.100 80.650 ;
        RECT 116.110 55.810 116.280 80.480 ;
        RECT 116.760 77.840 117.450 80.000 ;
        RECT 116.760 56.290 117.450 58.450 ;
        RECT 116.480 55.810 117.740 55.900 ;
        RECT 117.930 55.810 118.100 80.480 ;
        RECT 116.110 55.640 118.100 55.810 ;
        RECT 120.110 80.480 122.100 80.650 ;
        RECT 120.110 55.810 120.280 80.480 ;
        RECT 120.760 77.840 121.450 80.000 ;
        RECT 120.760 56.290 121.450 58.450 ;
        RECT 120.480 55.810 121.740 55.900 ;
        RECT 121.930 55.810 122.100 80.480 ;
        RECT 120.110 55.640 122.100 55.810 ;
        RECT 124.110 80.480 126.100 80.650 ;
        RECT 124.110 55.810 124.280 80.480 ;
        RECT 124.760 77.840 125.450 80.000 ;
        RECT 124.760 56.290 125.450 58.450 ;
        RECT 124.480 55.810 125.740 55.900 ;
        RECT 125.930 55.810 126.100 80.480 ;
        RECT 124.110 55.640 126.100 55.810 ;
        RECT 128.110 80.480 130.100 80.650 ;
        RECT 128.110 55.810 128.280 80.480 ;
        RECT 128.760 77.840 129.450 80.000 ;
        RECT 128.760 56.290 129.450 58.450 ;
        RECT 128.480 55.810 129.740 55.900 ;
        RECT 129.930 55.810 130.100 80.480 ;
        RECT 128.110 55.640 130.100 55.810 ;
        RECT 132.110 80.480 134.100 80.650 ;
        RECT 132.110 55.810 132.280 80.480 ;
        RECT 132.760 77.840 133.450 80.000 ;
        RECT 132.760 56.290 133.450 58.450 ;
        RECT 132.480 55.810 133.740 55.900 ;
        RECT 133.930 55.810 134.100 80.480 ;
        RECT 132.110 55.640 134.100 55.810 ;
        RECT 136.110 80.480 138.100 80.650 ;
        RECT 136.110 55.810 136.280 80.480 ;
        RECT 136.760 77.840 137.450 80.000 ;
        RECT 136.760 56.290 137.450 58.450 ;
        RECT 136.480 55.810 137.740 55.900 ;
        RECT 137.930 55.810 138.100 80.480 ;
        RECT 136.110 55.640 138.100 55.810 ;
        RECT 140.110 80.480 142.100 80.650 ;
        RECT 140.110 55.810 140.280 80.480 ;
        RECT 140.760 77.840 141.450 80.000 ;
        RECT 140.760 56.290 141.450 58.450 ;
        RECT 140.480 55.810 141.740 55.900 ;
        RECT 141.930 55.810 142.100 80.480 ;
        RECT 140.110 55.640 142.100 55.810 ;
        RECT 144.110 80.480 146.100 80.650 ;
        RECT 144.110 55.810 144.280 80.480 ;
        RECT 144.760 77.840 145.450 80.000 ;
        RECT 144.760 56.290 145.450 58.450 ;
        RECT 144.480 55.810 145.740 55.900 ;
        RECT 145.930 55.810 146.100 80.480 ;
        RECT 144.110 55.640 146.100 55.810 ;
        RECT 34.480 55.540 35.740 55.640 ;
        RECT 38.480 55.540 39.740 55.640 ;
        RECT 42.480 55.540 43.740 55.640 ;
        RECT 46.480 55.540 47.740 55.640 ;
        RECT 50.480 55.540 51.740 55.640 ;
        RECT 54.480 55.540 55.740 55.640 ;
        RECT 58.480 55.540 59.740 55.640 ;
        RECT 62.480 55.540 63.740 55.640 ;
        RECT 75.480 55.540 76.740 55.640 ;
        RECT 79.480 55.540 80.740 55.640 ;
        RECT 83.480 55.540 84.740 55.640 ;
        RECT 87.480 55.540 88.740 55.640 ;
        RECT 91.480 55.540 92.740 55.640 ;
        RECT 95.480 55.540 96.740 55.640 ;
        RECT 99.480 55.540 100.740 55.640 ;
        RECT 103.480 55.540 104.740 55.640 ;
        RECT 116.480 55.540 117.740 55.640 ;
        RECT 120.480 55.540 121.740 55.640 ;
        RECT 124.480 55.540 125.740 55.640 ;
        RECT 128.480 55.540 129.740 55.640 ;
        RECT 132.480 55.540 133.740 55.640 ;
        RECT 136.480 55.540 137.740 55.640 ;
        RECT 140.480 55.540 141.740 55.640 ;
        RECT 144.480 55.540 145.740 55.640 ;
        RECT 26.865 20.640 28.615 20.810 ;
        RECT 26.865 16.465 27.035 20.640 ;
        RECT 27.575 20.130 27.905 20.300 ;
        RECT 26.800 15.765 27.100 16.465 ;
        RECT 26.865 11.150 27.035 15.765 ;
        RECT 27.435 11.875 27.605 19.915 ;
        RECT 27.875 11.875 28.045 19.915 ;
        RECT 27.575 11.490 27.905 11.660 ;
        RECT 28.445 11.150 28.615 20.640 ;
        RECT 29.680 18.615 31.430 18.785 ;
        RECT 29.680 13.215 29.850 18.615 ;
        RECT 30.390 18.105 30.720 18.275 ;
        RECT 30.250 13.895 30.420 17.935 ;
        RECT 30.690 13.895 30.860 17.935 ;
        RECT 31.260 17.665 31.430 18.615 ;
        RECT 31.200 16.865 31.500 17.665 ;
        RECT 30.390 13.555 30.720 13.725 ;
        RECT 31.260 13.215 31.430 16.865 ;
        RECT 29.680 13.045 31.430 13.215 ;
        RECT 26.865 10.980 28.615 11.150 ;
      LAYER mcon ;
        RECT 36.245 214.765 36.415 214.935 ;
        RECT 36.705 214.765 36.875 214.935 ;
        RECT 37.165 214.765 37.335 214.935 ;
        RECT 37.625 214.765 37.795 214.935 ;
        RECT 38.085 214.765 38.255 214.935 ;
        RECT 38.545 214.765 38.715 214.935 ;
        RECT 39.005 214.765 39.175 214.935 ;
        RECT 39.465 214.765 39.635 214.935 ;
        RECT 39.925 214.765 40.095 214.935 ;
        RECT 40.385 214.765 40.555 214.935 ;
        RECT 40.845 214.765 41.015 214.935 ;
        RECT 41.305 214.765 41.475 214.935 ;
        RECT 41.765 214.765 41.935 214.935 ;
        RECT 42.225 214.765 42.395 214.935 ;
        RECT 42.685 214.765 42.855 214.935 ;
        RECT 43.145 214.765 43.315 214.935 ;
        RECT 43.605 214.765 43.775 214.935 ;
        RECT 44.065 214.765 44.235 214.935 ;
        RECT 44.525 214.765 44.695 214.935 ;
        RECT 44.985 214.765 45.155 214.935 ;
        RECT 45.445 214.765 45.615 214.935 ;
        RECT 45.905 214.765 46.075 214.935 ;
        RECT 46.365 214.765 46.535 214.935 ;
        RECT 46.825 214.765 46.995 214.935 ;
        RECT 47.285 214.765 47.455 214.935 ;
        RECT 47.745 214.765 47.915 214.935 ;
        RECT 48.205 214.765 48.375 214.935 ;
        RECT 48.665 214.765 48.835 214.935 ;
        RECT 49.125 214.765 49.295 214.935 ;
        RECT 49.585 214.765 49.755 214.935 ;
        RECT 50.045 214.765 50.215 214.935 ;
        RECT 50.505 214.765 50.675 214.935 ;
        RECT 50.965 214.765 51.135 214.935 ;
        RECT 51.425 214.765 51.595 214.935 ;
        RECT 51.885 214.765 52.055 214.935 ;
        RECT 52.345 214.765 52.515 214.935 ;
        RECT 52.805 214.765 52.975 214.935 ;
        RECT 53.265 214.765 53.435 214.935 ;
        RECT 53.725 214.765 53.895 214.935 ;
        RECT 54.185 214.765 54.355 214.935 ;
        RECT 54.645 214.765 54.815 214.935 ;
        RECT 55.105 214.765 55.275 214.935 ;
        RECT 55.565 214.765 55.735 214.935 ;
        RECT 56.025 214.765 56.195 214.935 ;
        RECT 56.485 214.765 56.655 214.935 ;
        RECT 56.945 214.765 57.115 214.935 ;
        RECT 57.405 214.765 57.575 214.935 ;
        RECT 57.865 214.765 58.035 214.935 ;
        RECT 58.325 214.765 58.495 214.935 ;
        RECT 58.785 214.765 58.955 214.935 ;
        RECT 59.245 214.765 59.415 214.935 ;
        RECT 59.705 214.765 59.875 214.935 ;
        RECT 60.165 214.765 60.335 214.935 ;
        RECT 60.625 214.765 60.795 214.935 ;
        RECT 61.085 214.765 61.255 214.935 ;
        RECT 61.545 214.765 61.715 214.935 ;
        RECT 62.005 214.765 62.175 214.935 ;
        RECT 62.465 214.765 62.635 214.935 ;
        RECT 62.925 214.765 63.095 214.935 ;
        RECT 63.385 214.765 63.555 214.935 ;
        RECT 63.845 214.765 64.015 214.935 ;
        RECT 64.305 214.765 64.475 214.935 ;
        RECT 64.765 214.765 64.935 214.935 ;
        RECT 65.225 214.765 65.395 214.935 ;
        RECT 65.685 214.765 65.855 214.935 ;
        RECT 66.145 214.765 66.315 214.935 ;
        RECT 66.605 214.765 66.775 214.935 ;
        RECT 67.065 214.765 67.235 214.935 ;
        RECT 67.525 214.765 67.695 214.935 ;
        RECT 67.985 214.765 68.155 214.935 ;
        RECT 68.445 214.765 68.615 214.935 ;
        RECT 68.905 214.765 69.075 214.935 ;
        RECT 69.365 214.765 69.535 214.935 ;
        RECT 69.825 214.765 69.995 214.935 ;
        RECT 70.285 214.765 70.455 214.935 ;
        RECT 70.745 214.765 70.915 214.935 ;
        RECT 71.205 214.765 71.375 214.935 ;
        RECT 71.665 214.765 71.835 214.935 ;
        RECT 72.125 214.765 72.295 214.935 ;
        RECT 72.585 214.765 72.755 214.935 ;
        RECT 73.045 214.765 73.215 214.935 ;
        RECT 73.505 214.765 73.675 214.935 ;
        RECT 73.965 214.765 74.135 214.935 ;
        RECT 74.425 214.765 74.595 214.935 ;
        RECT 74.885 214.765 75.055 214.935 ;
        RECT 75.345 214.765 75.515 214.935 ;
        RECT 75.805 214.765 75.975 214.935 ;
        RECT 76.265 214.765 76.435 214.935 ;
        RECT 76.725 214.765 76.895 214.935 ;
        RECT 77.185 214.765 77.355 214.935 ;
        RECT 77.645 214.765 77.815 214.935 ;
        RECT 78.105 214.765 78.275 214.935 ;
        RECT 78.565 214.765 78.735 214.935 ;
        RECT 79.025 214.765 79.195 214.935 ;
        RECT 79.485 214.765 79.655 214.935 ;
        RECT 79.945 214.765 80.115 214.935 ;
        RECT 80.405 214.765 80.575 214.935 ;
        RECT 80.865 214.765 81.035 214.935 ;
        RECT 81.325 214.765 81.495 214.935 ;
        RECT 81.785 214.765 81.955 214.935 ;
        RECT 82.245 214.765 82.415 214.935 ;
        RECT 82.705 214.765 82.875 214.935 ;
        RECT 83.165 214.765 83.335 214.935 ;
        RECT 83.625 214.765 83.795 214.935 ;
        RECT 84.085 214.765 84.255 214.935 ;
        RECT 84.545 214.765 84.715 214.935 ;
        RECT 85.005 214.765 85.175 214.935 ;
        RECT 85.465 214.765 85.635 214.935 ;
        RECT 85.925 214.765 86.095 214.935 ;
        RECT 86.385 214.765 86.555 214.935 ;
        RECT 86.845 214.765 87.015 214.935 ;
        RECT 87.305 214.765 87.475 214.935 ;
        RECT 87.765 214.765 87.935 214.935 ;
        RECT 88.225 214.765 88.395 214.935 ;
        RECT 88.685 214.765 88.855 214.935 ;
        RECT 89.145 214.765 89.315 214.935 ;
        RECT 89.605 214.765 89.775 214.935 ;
        RECT 90.065 214.765 90.235 214.935 ;
        RECT 90.525 214.765 90.695 214.935 ;
        RECT 90.985 214.765 91.155 214.935 ;
        RECT 91.445 214.765 91.615 214.935 ;
        RECT 91.905 214.765 92.075 214.935 ;
        RECT 92.365 214.765 92.535 214.935 ;
        RECT 92.825 214.765 92.995 214.935 ;
        RECT 93.285 214.765 93.455 214.935 ;
        RECT 93.745 214.765 93.915 214.935 ;
        RECT 94.205 214.765 94.375 214.935 ;
        RECT 94.665 214.765 94.835 214.935 ;
        RECT 95.125 214.765 95.295 214.935 ;
        RECT 95.585 214.765 95.755 214.935 ;
        RECT 96.045 214.765 96.215 214.935 ;
        RECT 96.505 214.765 96.675 214.935 ;
        RECT 96.965 214.765 97.135 214.935 ;
        RECT 97.425 214.765 97.595 214.935 ;
        RECT 97.885 214.765 98.055 214.935 ;
        RECT 98.345 214.765 98.515 214.935 ;
        RECT 98.805 214.765 98.975 214.935 ;
        RECT 99.265 214.765 99.435 214.935 ;
        RECT 99.725 214.765 99.895 214.935 ;
        RECT 100.185 214.765 100.355 214.935 ;
        RECT 100.645 214.765 100.815 214.935 ;
        RECT 101.105 214.765 101.275 214.935 ;
        RECT 101.565 214.765 101.735 214.935 ;
        RECT 102.025 214.765 102.195 214.935 ;
        RECT 102.485 214.765 102.655 214.935 ;
        RECT 102.945 214.765 103.115 214.935 ;
        RECT 103.405 214.765 103.575 214.935 ;
        RECT 103.865 214.765 104.035 214.935 ;
        RECT 104.325 214.765 104.495 214.935 ;
        RECT 104.785 214.765 104.955 214.935 ;
        RECT 105.245 214.765 105.415 214.935 ;
        RECT 105.705 214.765 105.875 214.935 ;
        RECT 106.165 214.765 106.335 214.935 ;
        RECT 106.625 214.765 106.795 214.935 ;
        RECT 107.085 214.765 107.255 214.935 ;
        RECT 107.545 214.765 107.715 214.935 ;
        RECT 108.005 214.765 108.175 214.935 ;
        RECT 108.465 214.765 108.635 214.935 ;
        RECT 108.925 214.765 109.095 214.935 ;
        RECT 109.385 214.765 109.555 214.935 ;
        RECT 109.845 214.765 110.015 214.935 ;
        RECT 110.305 214.765 110.475 214.935 ;
        RECT 110.765 214.765 110.935 214.935 ;
        RECT 111.225 214.765 111.395 214.935 ;
        RECT 111.685 214.765 111.855 214.935 ;
        RECT 112.145 214.765 112.315 214.935 ;
        RECT 112.605 214.765 112.775 214.935 ;
        RECT 113.065 214.765 113.235 214.935 ;
        RECT 113.525 214.765 113.695 214.935 ;
        RECT 113.985 214.765 114.155 214.935 ;
        RECT 114.445 214.765 114.615 214.935 ;
        RECT 114.905 214.765 115.075 214.935 ;
        RECT 115.365 214.765 115.535 214.935 ;
        RECT 115.825 214.765 115.995 214.935 ;
        RECT 116.285 214.765 116.455 214.935 ;
        RECT 116.745 214.765 116.915 214.935 ;
        RECT 117.205 214.765 117.375 214.935 ;
        RECT 117.665 214.765 117.835 214.935 ;
        RECT 118.125 214.765 118.295 214.935 ;
        RECT 118.585 214.765 118.755 214.935 ;
        RECT 119.045 214.765 119.215 214.935 ;
        RECT 119.505 214.765 119.675 214.935 ;
        RECT 119.965 214.765 120.135 214.935 ;
        RECT 120.425 214.765 120.595 214.935 ;
        RECT 120.885 214.765 121.055 214.935 ;
        RECT 121.345 214.765 121.515 214.935 ;
        RECT 121.805 214.765 121.975 214.935 ;
        RECT 122.265 214.765 122.435 214.935 ;
        RECT 122.725 214.765 122.895 214.935 ;
        RECT 123.185 214.765 123.355 214.935 ;
        RECT 123.645 214.765 123.815 214.935 ;
        RECT 124.105 214.765 124.275 214.935 ;
        RECT 124.565 214.765 124.735 214.935 ;
        RECT 125.025 214.765 125.195 214.935 ;
        RECT 125.485 214.765 125.655 214.935 ;
        RECT 125.945 214.765 126.115 214.935 ;
        RECT 126.405 214.765 126.575 214.935 ;
        RECT 126.865 214.765 127.035 214.935 ;
        RECT 127.325 214.765 127.495 214.935 ;
        RECT 127.785 214.765 127.955 214.935 ;
        RECT 128.245 214.765 128.415 214.935 ;
        RECT 128.705 214.765 128.875 214.935 ;
        RECT 129.165 214.765 129.335 214.935 ;
        RECT 129.625 214.765 129.795 214.935 ;
        RECT 130.085 214.765 130.255 214.935 ;
        RECT 130.545 214.765 130.715 214.935 ;
        RECT 131.005 214.765 131.175 214.935 ;
        RECT 131.465 214.765 131.635 214.935 ;
        RECT 131.925 214.765 132.095 214.935 ;
        RECT 132.385 214.765 132.555 214.935 ;
        RECT 132.845 214.765 133.015 214.935 ;
        RECT 133.305 214.765 133.475 214.935 ;
        RECT 133.765 214.765 133.935 214.935 ;
        RECT 134.225 214.765 134.395 214.935 ;
        RECT 134.685 214.765 134.855 214.935 ;
        RECT 135.145 214.765 135.315 214.935 ;
        RECT 135.605 214.765 135.775 214.935 ;
        RECT 136.065 214.765 136.235 214.935 ;
        RECT 136.525 214.765 136.695 214.935 ;
        RECT 136.985 214.765 137.155 214.935 ;
        RECT 137.445 214.765 137.615 214.935 ;
        RECT 137.905 214.765 138.075 214.935 ;
        RECT 138.365 214.765 138.535 214.935 ;
        RECT 138.825 214.765 138.995 214.935 ;
        RECT 139.285 214.765 139.455 214.935 ;
        RECT 139.745 214.765 139.915 214.935 ;
        RECT 140.205 214.765 140.375 214.935 ;
        RECT 140.665 214.765 140.835 214.935 ;
        RECT 141.125 214.765 141.295 214.935 ;
        RECT 141.585 214.765 141.755 214.935 ;
        RECT 142.045 214.765 142.215 214.935 ;
        RECT 142.505 214.765 142.675 214.935 ;
        RECT 142.965 214.765 143.135 214.935 ;
        RECT 143.425 214.765 143.595 214.935 ;
        RECT 143.885 214.765 144.055 214.935 ;
        RECT 144.345 214.765 144.515 214.935 ;
        RECT 144.805 214.765 144.975 214.935 ;
        RECT 145.265 214.765 145.435 214.935 ;
        RECT 145.725 214.765 145.895 214.935 ;
        RECT 146.185 214.765 146.355 214.935 ;
        RECT 146.645 214.765 146.815 214.935 ;
        RECT 147.105 214.765 147.275 214.935 ;
        RECT 147.565 214.765 147.735 214.935 ;
        RECT 148.025 214.765 148.195 214.935 ;
        RECT 148.485 214.765 148.655 214.935 ;
        RECT 148.945 214.765 149.115 214.935 ;
        RECT 149.405 214.765 149.575 214.935 ;
        RECT 149.865 214.765 150.035 214.935 ;
        RECT 44.985 213.235 45.155 213.405 ;
        RECT 48.205 212.555 48.375 212.725 ;
        RECT 56.485 214.255 56.655 214.425 ;
        RECT 59.245 214.255 59.415 214.425 ;
        RECT 57.405 213.235 57.575 213.405 ;
        RECT 60.625 212.895 60.795 213.065 ;
        RECT 64.305 214.255 64.475 214.425 ;
        RECT 63.385 213.235 63.555 213.405 ;
        RECT 66.605 214.255 66.775 214.425 ;
        RECT 67.985 212.895 68.155 213.065 ;
        RECT 71.205 214.255 71.375 214.425 ;
        RECT 72.125 213.235 72.295 213.405 ;
        RECT 72.585 213.235 72.755 213.405 ;
        RECT 75.805 214.255 75.975 214.425 ;
        RECT 79.025 214.255 79.195 214.425 ;
        RECT 73.505 213.235 73.675 213.405 ;
        RECT 73.045 212.555 73.215 212.725 ;
        RECT 77.185 212.895 77.355 213.065 ;
        RECT 78.105 213.235 78.275 213.405 ;
        RECT 81.325 214.255 81.495 214.425 ;
        RECT 82.705 212.895 82.875 213.065 ;
        RECT 85.925 214.255 86.095 214.425 ;
        RECT 88.685 214.255 88.855 214.425 ;
        RECT 86.845 213.235 87.015 213.405 ;
        RECT 90.065 212.895 90.235 213.065 ;
        RECT 99.265 213.235 99.435 213.405 ;
        RECT 101.105 213.235 101.275 213.405 ;
        RECT 102.485 213.235 102.655 213.405 ;
        RECT 98.805 212.555 98.975 212.725 ;
        RECT 113.985 213.915 114.155 214.085 ;
        RECT 116.285 213.575 116.455 213.745 ;
        RECT 116.745 213.575 116.915 213.745 ;
        RECT 122.265 213.235 122.435 213.405 ;
        RECT 123.185 212.555 123.355 212.725 ;
        RECT 126.865 213.235 127.035 213.405 ;
        RECT 127.785 212.555 127.955 212.725 ;
        RECT 130.545 213.235 130.715 213.405 ;
        RECT 129.625 212.555 129.795 212.725 ;
        RECT 133.765 213.235 133.935 213.405 ;
        RECT 132.845 212.555 133.015 212.725 ;
        RECT 135.145 213.235 135.315 213.405 ;
        RECT 134.225 212.555 134.395 212.725 ;
        RECT 139.745 213.915 139.915 214.085 ;
        RECT 140.665 214.255 140.835 214.425 ;
        RECT 137.905 213.235 138.075 213.405 ;
        RECT 136.985 212.555 137.155 212.725 ;
        RECT 142.045 213.235 142.215 213.405 ;
        RECT 144.345 213.915 144.515 214.085 ;
        RECT 143.425 213.235 143.595 213.405 ;
        RECT 142.505 212.555 142.675 212.725 ;
        RECT 145.265 213.235 145.435 213.405 ;
        RECT 147.565 213.915 147.735 214.085 ;
        RECT 148.485 213.235 148.655 213.405 ;
        RECT 36.245 212.045 36.415 212.215 ;
        RECT 36.705 212.045 36.875 212.215 ;
        RECT 37.165 212.045 37.335 212.215 ;
        RECT 37.625 212.045 37.795 212.215 ;
        RECT 38.085 212.045 38.255 212.215 ;
        RECT 38.545 212.045 38.715 212.215 ;
        RECT 39.005 212.045 39.175 212.215 ;
        RECT 39.465 212.045 39.635 212.215 ;
        RECT 39.925 212.045 40.095 212.215 ;
        RECT 40.385 212.045 40.555 212.215 ;
        RECT 40.845 212.045 41.015 212.215 ;
        RECT 41.305 212.045 41.475 212.215 ;
        RECT 41.765 212.045 41.935 212.215 ;
        RECT 42.225 212.045 42.395 212.215 ;
        RECT 42.685 212.045 42.855 212.215 ;
        RECT 43.145 212.045 43.315 212.215 ;
        RECT 43.605 212.045 43.775 212.215 ;
        RECT 44.065 212.045 44.235 212.215 ;
        RECT 44.525 212.045 44.695 212.215 ;
        RECT 44.985 212.045 45.155 212.215 ;
        RECT 45.445 212.045 45.615 212.215 ;
        RECT 45.905 212.045 46.075 212.215 ;
        RECT 46.365 212.045 46.535 212.215 ;
        RECT 46.825 212.045 46.995 212.215 ;
        RECT 47.285 212.045 47.455 212.215 ;
        RECT 47.745 212.045 47.915 212.215 ;
        RECT 48.205 212.045 48.375 212.215 ;
        RECT 48.665 212.045 48.835 212.215 ;
        RECT 49.125 212.045 49.295 212.215 ;
        RECT 49.585 212.045 49.755 212.215 ;
        RECT 50.045 212.045 50.215 212.215 ;
        RECT 50.505 212.045 50.675 212.215 ;
        RECT 50.965 212.045 51.135 212.215 ;
        RECT 51.425 212.045 51.595 212.215 ;
        RECT 51.885 212.045 52.055 212.215 ;
        RECT 52.345 212.045 52.515 212.215 ;
        RECT 52.805 212.045 52.975 212.215 ;
        RECT 53.265 212.045 53.435 212.215 ;
        RECT 53.725 212.045 53.895 212.215 ;
        RECT 54.185 212.045 54.355 212.215 ;
        RECT 54.645 212.045 54.815 212.215 ;
        RECT 55.105 212.045 55.275 212.215 ;
        RECT 55.565 212.045 55.735 212.215 ;
        RECT 56.025 212.045 56.195 212.215 ;
        RECT 56.485 212.045 56.655 212.215 ;
        RECT 56.945 212.045 57.115 212.215 ;
        RECT 57.405 212.045 57.575 212.215 ;
        RECT 57.865 212.045 58.035 212.215 ;
        RECT 58.325 212.045 58.495 212.215 ;
        RECT 58.785 212.045 58.955 212.215 ;
        RECT 59.245 212.045 59.415 212.215 ;
        RECT 59.705 212.045 59.875 212.215 ;
        RECT 60.165 212.045 60.335 212.215 ;
        RECT 60.625 212.045 60.795 212.215 ;
        RECT 61.085 212.045 61.255 212.215 ;
        RECT 61.545 212.045 61.715 212.215 ;
        RECT 62.005 212.045 62.175 212.215 ;
        RECT 62.465 212.045 62.635 212.215 ;
        RECT 62.925 212.045 63.095 212.215 ;
        RECT 63.385 212.045 63.555 212.215 ;
        RECT 63.845 212.045 64.015 212.215 ;
        RECT 64.305 212.045 64.475 212.215 ;
        RECT 64.765 212.045 64.935 212.215 ;
        RECT 65.225 212.045 65.395 212.215 ;
        RECT 65.685 212.045 65.855 212.215 ;
        RECT 66.145 212.045 66.315 212.215 ;
        RECT 66.605 212.045 66.775 212.215 ;
        RECT 67.065 212.045 67.235 212.215 ;
        RECT 67.525 212.045 67.695 212.215 ;
        RECT 67.985 212.045 68.155 212.215 ;
        RECT 68.445 212.045 68.615 212.215 ;
        RECT 68.905 212.045 69.075 212.215 ;
        RECT 69.365 212.045 69.535 212.215 ;
        RECT 69.825 212.045 69.995 212.215 ;
        RECT 70.285 212.045 70.455 212.215 ;
        RECT 70.745 212.045 70.915 212.215 ;
        RECT 71.205 212.045 71.375 212.215 ;
        RECT 71.665 212.045 71.835 212.215 ;
        RECT 72.125 212.045 72.295 212.215 ;
        RECT 72.585 212.045 72.755 212.215 ;
        RECT 73.045 212.045 73.215 212.215 ;
        RECT 73.505 212.045 73.675 212.215 ;
        RECT 73.965 212.045 74.135 212.215 ;
        RECT 74.425 212.045 74.595 212.215 ;
        RECT 74.885 212.045 75.055 212.215 ;
        RECT 75.345 212.045 75.515 212.215 ;
        RECT 75.805 212.045 75.975 212.215 ;
        RECT 76.265 212.045 76.435 212.215 ;
        RECT 76.725 212.045 76.895 212.215 ;
        RECT 77.185 212.045 77.355 212.215 ;
        RECT 77.645 212.045 77.815 212.215 ;
        RECT 78.105 212.045 78.275 212.215 ;
        RECT 78.565 212.045 78.735 212.215 ;
        RECT 79.025 212.045 79.195 212.215 ;
        RECT 79.485 212.045 79.655 212.215 ;
        RECT 79.945 212.045 80.115 212.215 ;
        RECT 80.405 212.045 80.575 212.215 ;
        RECT 80.865 212.045 81.035 212.215 ;
        RECT 81.325 212.045 81.495 212.215 ;
        RECT 81.785 212.045 81.955 212.215 ;
        RECT 82.245 212.045 82.415 212.215 ;
        RECT 82.705 212.045 82.875 212.215 ;
        RECT 83.165 212.045 83.335 212.215 ;
        RECT 83.625 212.045 83.795 212.215 ;
        RECT 84.085 212.045 84.255 212.215 ;
        RECT 84.545 212.045 84.715 212.215 ;
        RECT 85.005 212.045 85.175 212.215 ;
        RECT 85.465 212.045 85.635 212.215 ;
        RECT 85.925 212.045 86.095 212.215 ;
        RECT 86.385 212.045 86.555 212.215 ;
        RECT 86.845 212.045 87.015 212.215 ;
        RECT 87.305 212.045 87.475 212.215 ;
        RECT 87.765 212.045 87.935 212.215 ;
        RECT 88.225 212.045 88.395 212.215 ;
        RECT 88.685 212.045 88.855 212.215 ;
        RECT 89.145 212.045 89.315 212.215 ;
        RECT 89.605 212.045 89.775 212.215 ;
        RECT 90.065 212.045 90.235 212.215 ;
        RECT 90.525 212.045 90.695 212.215 ;
        RECT 90.985 212.045 91.155 212.215 ;
        RECT 91.445 212.045 91.615 212.215 ;
        RECT 91.905 212.045 92.075 212.215 ;
        RECT 92.365 212.045 92.535 212.215 ;
        RECT 92.825 212.045 92.995 212.215 ;
        RECT 93.285 212.045 93.455 212.215 ;
        RECT 93.745 212.045 93.915 212.215 ;
        RECT 94.205 212.045 94.375 212.215 ;
        RECT 94.665 212.045 94.835 212.215 ;
        RECT 95.125 212.045 95.295 212.215 ;
        RECT 95.585 212.045 95.755 212.215 ;
        RECT 96.045 212.045 96.215 212.215 ;
        RECT 96.505 212.045 96.675 212.215 ;
        RECT 96.965 212.045 97.135 212.215 ;
        RECT 97.425 212.045 97.595 212.215 ;
        RECT 97.885 212.045 98.055 212.215 ;
        RECT 98.345 212.045 98.515 212.215 ;
        RECT 98.805 212.045 98.975 212.215 ;
        RECT 99.265 212.045 99.435 212.215 ;
        RECT 99.725 212.045 99.895 212.215 ;
        RECT 100.185 212.045 100.355 212.215 ;
        RECT 100.645 212.045 100.815 212.215 ;
        RECT 101.105 212.045 101.275 212.215 ;
        RECT 101.565 212.045 101.735 212.215 ;
        RECT 102.025 212.045 102.195 212.215 ;
        RECT 102.485 212.045 102.655 212.215 ;
        RECT 102.945 212.045 103.115 212.215 ;
        RECT 103.405 212.045 103.575 212.215 ;
        RECT 103.865 212.045 104.035 212.215 ;
        RECT 104.325 212.045 104.495 212.215 ;
        RECT 104.785 212.045 104.955 212.215 ;
        RECT 105.245 212.045 105.415 212.215 ;
        RECT 105.705 212.045 105.875 212.215 ;
        RECT 106.165 212.045 106.335 212.215 ;
        RECT 106.625 212.045 106.795 212.215 ;
        RECT 107.085 212.045 107.255 212.215 ;
        RECT 107.545 212.045 107.715 212.215 ;
        RECT 108.005 212.045 108.175 212.215 ;
        RECT 108.465 212.045 108.635 212.215 ;
        RECT 108.925 212.045 109.095 212.215 ;
        RECT 109.385 212.045 109.555 212.215 ;
        RECT 109.845 212.045 110.015 212.215 ;
        RECT 110.305 212.045 110.475 212.215 ;
        RECT 110.765 212.045 110.935 212.215 ;
        RECT 111.225 212.045 111.395 212.215 ;
        RECT 111.685 212.045 111.855 212.215 ;
        RECT 112.145 212.045 112.315 212.215 ;
        RECT 112.605 212.045 112.775 212.215 ;
        RECT 113.065 212.045 113.235 212.215 ;
        RECT 113.525 212.045 113.695 212.215 ;
        RECT 113.985 212.045 114.155 212.215 ;
        RECT 114.445 212.045 114.615 212.215 ;
        RECT 114.905 212.045 115.075 212.215 ;
        RECT 115.365 212.045 115.535 212.215 ;
        RECT 115.825 212.045 115.995 212.215 ;
        RECT 116.285 212.045 116.455 212.215 ;
        RECT 116.745 212.045 116.915 212.215 ;
        RECT 117.205 212.045 117.375 212.215 ;
        RECT 117.665 212.045 117.835 212.215 ;
        RECT 118.125 212.045 118.295 212.215 ;
        RECT 118.585 212.045 118.755 212.215 ;
        RECT 119.045 212.045 119.215 212.215 ;
        RECT 119.505 212.045 119.675 212.215 ;
        RECT 119.965 212.045 120.135 212.215 ;
        RECT 120.425 212.045 120.595 212.215 ;
        RECT 120.885 212.045 121.055 212.215 ;
        RECT 121.345 212.045 121.515 212.215 ;
        RECT 121.805 212.045 121.975 212.215 ;
        RECT 122.265 212.045 122.435 212.215 ;
        RECT 122.725 212.045 122.895 212.215 ;
        RECT 123.185 212.045 123.355 212.215 ;
        RECT 123.645 212.045 123.815 212.215 ;
        RECT 124.105 212.045 124.275 212.215 ;
        RECT 124.565 212.045 124.735 212.215 ;
        RECT 125.025 212.045 125.195 212.215 ;
        RECT 125.485 212.045 125.655 212.215 ;
        RECT 125.945 212.045 126.115 212.215 ;
        RECT 126.405 212.045 126.575 212.215 ;
        RECT 126.865 212.045 127.035 212.215 ;
        RECT 127.325 212.045 127.495 212.215 ;
        RECT 127.785 212.045 127.955 212.215 ;
        RECT 128.245 212.045 128.415 212.215 ;
        RECT 128.705 212.045 128.875 212.215 ;
        RECT 129.165 212.045 129.335 212.215 ;
        RECT 129.625 212.045 129.795 212.215 ;
        RECT 130.085 212.045 130.255 212.215 ;
        RECT 130.545 212.045 130.715 212.215 ;
        RECT 131.005 212.045 131.175 212.215 ;
        RECT 131.465 212.045 131.635 212.215 ;
        RECT 131.925 212.045 132.095 212.215 ;
        RECT 132.385 212.045 132.555 212.215 ;
        RECT 132.845 212.045 133.015 212.215 ;
        RECT 133.305 212.045 133.475 212.215 ;
        RECT 133.765 212.045 133.935 212.215 ;
        RECT 134.225 212.045 134.395 212.215 ;
        RECT 134.685 212.045 134.855 212.215 ;
        RECT 135.145 212.045 135.315 212.215 ;
        RECT 135.605 212.045 135.775 212.215 ;
        RECT 136.065 212.045 136.235 212.215 ;
        RECT 136.525 212.045 136.695 212.215 ;
        RECT 136.985 212.045 137.155 212.215 ;
        RECT 137.445 212.045 137.615 212.215 ;
        RECT 137.905 212.045 138.075 212.215 ;
        RECT 138.365 212.045 138.535 212.215 ;
        RECT 138.825 212.045 138.995 212.215 ;
        RECT 139.285 212.045 139.455 212.215 ;
        RECT 139.745 212.045 139.915 212.215 ;
        RECT 140.205 212.045 140.375 212.215 ;
        RECT 140.665 212.045 140.835 212.215 ;
        RECT 141.125 212.045 141.295 212.215 ;
        RECT 141.585 212.045 141.755 212.215 ;
        RECT 142.045 212.045 142.215 212.215 ;
        RECT 142.505 212.045 142.675 212.215 ;
        RECT 142.965 212.045 143.135 212.215 ;
        RECT 143.425 212.045 143.595 212.215 ;
        RECT 143.885 212.045 144.055 212.215 ;
        RECT 144.345 212.045 144.515 212.215 ;
        RECT 144.805 212.045 144.975 212.215 ;
        RECT 145.265 212.045 145.435 212.215 ;
        RECT 145.725 212.045 145.895 212.215 ;
        RECT 146.185 212.045 146.355 212.215 ;
        RECT 146.645 212.045 146.815 212.215 ;
        RECT 147.105 212.045 147.275 212.215 ;
        RECT 147.565 212.045 147.735 212.215 ;
        RECT 148.025 212.045 148.195 212.215 ;
        RECT 148.485 212.045 148.655 212.215 ;
        RECT 148.945 212.045 149.115 212.215 ;
        RECT 149.405 212.045 149.575 212.215 ;
        RECT 149.865 212.045 150.035 212.215 ;
        RECT 37.625 210.515 37.795 210.685 ;
        RECT 38.110 210.175 38.280 210.345 ;
        RECT 38.505 210.515 38.675 210.685 ;
        RECT 38.960 210.855 39.130 211.025 ;
        RECT 39.695 210.515 39.865 210.685 ;
        RECT 40.210 210.175 40.380 210.345 ;
        RECT 41.780 210.175 41.950 210.345 ;
        RECT 42.215 210.515 42.385 210.685 ;
        RECT 44.525 211.535 44.695 211.705 ;
        RECT 45.445 211.535 45.615 211.705 ;
        RECT 45.905 210.855 46.075 211.025 ;
        RECT 46.365 210.855 46.535 211.025 ;
        RECT 46.850 210.175 47.020 210.345 ;
        RECT 47.245 210.515 47.415 210.685 ;
        RECT 47.700 210.855 47.870 211.025 ;
        RECT 48.435 210.515 48.605 210.685 ;
        RECT 48.950 210.175 49.120 210.345 ;
        RECT 50.520 210.175 50.690 210.345 ;
        RECT 50.955 210.515 51.125 210.685 ;
        RECT 54.645 210.855 54.815 211.025 ;
        RECT 53.265 209.835 53.435 210.005 ;
        RECT 55.130 210.175 55.300 210.345 ;
        RECT 55.525 210.515 55.695 210.685 ;
        RECT 55.980 210.855 56.150 211.025 ;
        RECT 56.715 210.515 56.885 210.685 ;
        RECT 57.230 210.175 57.400 210.345 ;
        RECT 58.800 210.175 58.970 210.345 ;
        RECT 59.235 210.515 59.405 210.685 ;
        RECT 61.545 211.535 61.715 211.705 ;
        RECT 64.305 211.535 64.475 211.705 ;
        RECT 63.845 211.195 64.015 211.365 ;
        RECT 67.065 211.535 67.235 211.705 ;
        RECT 66.145 210.855 66.315 211.025 ;
        RECT 66.605 210.855 66.775 211.025 ;
        RECT 67.525 210.855 67.695 211.025 ;
        RECT 65.225 209.835 65.395 210.005 ;
        RECT 68.905 210.855 69.075 211.025 ;
        RECT 67.985 210.175 68.155 210.345 ;
        RECT 71.205 210.855 71.375 211.025 ;
        RECT 71.665 210.515 71.835 210.685 ;
        RECT 73.045 210.175 73.215 210.345 ;
        RECT 74.425 210.855 74.595 211.025 ;
        RECT 73.965 210.515 74.135 210.685 ;
        RECT 75.805 209.835 75.975 210.005 ;
        RECT 80.865 210.855 81.035 211.025 ;
        RECT 79.945 210.515 80.115 210.685 ;
        RECT 81.785 210.515 81.955 210.685 ;
        RECT 84.545 211.535 84.715 211.705 ;
        RECT 85.465 211.535 85.635 211.705 ;
        RECT 85.005 210.855 85.175 211.025 ;
        RECT 86.385 210.855 86.555 211.025 ;
        RECT 83.625 210.175 83.795 210.345 ;
        RECT 88.685 211.535 88.855 211.705 ;
        RECT 88.225 211.195 88.395 211.365 ;
        RECT 87.305 209.835 87.475 210.005 ;
        RECT 90.065 210.515 90.235 210.685 ;
        RECT 93.745 210.855 93.915 211.025 ;
        RECT 89.605 209.835 89.775 210.005 ;
        RECT 90.065 209.835 90.235 210.005 ;
        RECT 95.125 210.855 95.295 211.025 ;
        RECT 94.665 210.175 94.835 210.345 ;
        RECT 95.610 210.175 95.780 210.345 ;
        RECT 96.005 210.515 96.175 210.685 ;
        RECT 96.405 210.855 96.575 211.025 ;
        RECT 97.195 210.515 97.365 210.685 ;
        RECT 97.710 210.175 97.880 210.345 ;
        RECT 99.280 210.175 99.450 210.345 ;
        RECT 99.715 210.515 99.885 210.685 ;
        RECT 102.485 210.855 102.655 211.025 ;
        RECT 102.025 209.835 102.195 210.005 ;
        RECT 102.970 210.175 103.140 210.345 ;
        RECT 103.365 210.515 103.535 210.685 ;
        RECT 103.820 210.855 103.990 211.025 ;
        RECT 104.555 210.515 104.725 210.685 ;
        RECT 105.070 210.175 105.240 210.345 ;
        RECT 106.640 210.175 106.810 210.345 ;
        RECT 107.075 210.515 107.245 210.685 ;
        RECT 109.385 209.835 109.555 210.005 ;
        RECT 110.765 210.515 110.935 210.685 ;
        RECT 111.685 210.855 111.855 211.025 ;
        RECT 112.605 210.175 112.775 210.345 ;
        RECT 113.985 209.835 114.155 210.005 ;
        RECT 116.285 211.535 116.455 211.705 ;
        RECT 118.125 211.535 118.295 211.705 ;
        RECT 117.205 210.515 117.375 210.685 ;
        RECT 123.645 211.535 123.815 211.705 ;
        RECT 119.045 210.855 119.215 211.025 ;
        RECT 121.805 210.855 121.975 211.025 ;
        RECT 119.965 209.835 120.135 210.005 ;
        RECT 120.885 210.175 121.055 210.345 ;
        RECT 122.725 209.835 122.895 210.005 ;
        RECT 125.945 210.515 126.115 210.685 ;
        RECT 126.865 210.515 127.035 210.685 ;
        RECT 129.165 210.855 129.335 211.025 ;
        RECT 128.245 210.515 128.415 210.685 ;
        RECT 129.625 210.855 129.795 211.025 ;
        RECT 131.925 210.855 132.095 211.025 ;
        RECT 131.465 209.835 131.635 210.005 ;
        RECT 132.410 210.175 132.580 210.345 ;
        RECT 132.805 210.515 132.975 210.685 ;
        RECT 133.260 210.855 133.430 211.025 ;
        RECT 133.995 210.515 134.165 210.685 ;
        RECT 134.510 210.175 134.680 210.345 ;
        RECT 136.080 210.175 136.250 210.345 ;
        RECT 136.515 210.515 136.685 210.685 ;
        RECT 138.825 211.535 138.995 211.705 ;
        RECT 141.125 211.535 141.295 211.705 ;
        RECT 140.205 210.855 140.375 211.025 ;
        RECT 141.585 210.855 141.755 211.025 ;
        RECT 142.070 210.175 142.240 210.345 ;
        RECT 142.465 210.515 142.635 210.685 ;
        RECT 142.810 211.195 142.980 211.365 ;
        RECT 143.655 210.515 143.825 210.685 ;
        RECT 144.170 210.175 144.340 210.345 ;
        RECT 145.740 210.175 145.910 210.345 ;
        RECT 146.175 210.515 146.345 210.685 ;
        RECT 148.485 211.535 148.655 211.705 ;
        RECT 36.245 209.325 36.415 209.495 ;
        RECT 36.705 209.325 36.875 209.495 ;
        RECT 37.165 209.325 37.335 209.495 ;
        RECT 37.625 209.325 37.795 209.495 ;
        RECT 38.085 209.325 38.255 209.495 ;
        RECT 38.545 209.325 38.715 209.495 ;
        RECT 39.005 209.325 39.175 209.495 ;
        RECT 39.465 209.325 39.635 209.495 ;
        RECT 39.925 209.325 40.095 209.495 ;
        RECT 40.385 209.325 40.555 209.495 ;
        RECT 40.845 209.325 41.015 209.495 ;
        RECT 41.305 209.325 41.475 209.495 ;
        RECT 41.765 209.325 41.935 209.495 ;
        RECT 42.225 209.325 42.395 209.495 ;
        RECT 42.685 209.325 42.855 209.495 ;
        RECT 43.145 209.325 43.315 209.495 ;
        RECT 43.605 209.325 43.775 209.495 ;
        RECT 44.065 209.325 44.235 209.495 ;
        RECT 44.525 209.325 44.695 209.495 ;
        RECT 44.985 209.325 45.155 209.495 ;
        RECT 45.445 209.325 45.615 209.495 ;
        RECT 45.905 209.325 46.075 209.495 ;
        RECT 46.365 209.325 46.535 209.495 ;
        RECT 46.825 209.325 46.995 209.495 ;
        RECT 47.285 209.325 47.455 209.495 ;
        RECT 47.745 209.325 47.915 209.495 ;
        RECT 48.205 209.325 48.375 209.495 ;
        RECT 48.665 209.325 48.835 209.495 ;
        RECT 49.125 209.325 49.295 209.495 ;
        RECT 49.585 209.325 49.755 209.495 ;
        RECT 50.045 209.325 50.215 209.495 ;
        RECT 50.505 209.325 50.675 209.495 ;
        RECT 50.965 209.325 51.135 209.495 ;
        RECT 51.425 209.325 51.595 209.495 ;
        RECT 51.885 209.325 52.055 209.495 ;
        RECT 52.345 209.325 52.515 209.495 ;
        RECT 52.805 209.325 52.975 209.495 ;
        RECT 53.265 209.325 53.435 209.495 ;
        RECT 53.725 209.325 53.895 209.495 ;
        RECT 54.185 209.325 54.355 209.495 ;
        RECT 54.645 209.325 54.815 209.495 ;
        RECT 55.105 209.325 55.275 209.495 ;
        RECT 55.565 209.325 55.735 209.495 ;
        RECT 56.025 209.325 56.195 209.495 ;
        RECT 56.485 209.325 56.655 209.495 ;
        RECT 56.945 209.325 57.115 209.495 ;
        RECT 57.405 209.325 57.575 209.495 ;
        RECT 57.865 209.325 58.035 209.495 ;
        RECT 58.325 209.325 58.495 209.495 ;
        RECT 58.785 209.325 58.955 209.495 ;
        RECT 59.245 209.325 59.415 209.495 ;
        RECT 59.705 209.325 59.875 209.495 ;
        RECT 60.165 209.325 60.335 209.495 ;
        RECT 60.625 209.325 60.795 209.495 ;
        RECT 61.085 209.325 61.255 209.495 ;
        RECT 61.545 209.325 61.715 209.495 ;
        RECT 62.005 209.325 62.175 209.495 ;
        RECT 62.465 209.325 62.635 209.495 ;
        RECT 62.925 209.325 63.095 209.495 ;
        RECT 63.385 209.325 63.555 209.495 ;
        RECT 63.845 209.325 64.015 209.495 ;
        RECT 64.305 209.325 64.475 209.495 ;
        RECT 64.765 209.325 64.935 209.495 ;
        RECT 65.225 209.325 65.395 209.495 ;
        RECT 65.685 209.325 65.855 209.495 ;
        RECT 66.145 209.325 66.315 209.495 ;
        RECT 66.605 209.325 66.775 209.495 ;
        RECT 67.065 209.325 67.235 209.495 ;
        RECT 67.525 209.325 67.695 209.495 ;
        RECT 67.985 209.325 68.155 209.495 ;
        RECT 68.445 209.325 68.615 209.495 ;
        RECT 68.905 209.325 69.075 209.495 ;
        RECT 69.365 209.325 69.535 209.495 ;
        RECT 69.825 209.325 69.995 209.495 ;
        RECT 70.285 209.325 70.455 209.495 ;
        RECT 70.745 209.325 70.915 209.495 ;
        RECT 71.205 209.325 71.375 209.495 ;
        RECT 71.665 209.325 71.835 209.495 ;
        RECT 72.125 209.325 72.295 209.495 ;
        RECT 72.585 209.325 72.755 209.495 ;
        RECT 73.045 209.325 73.215 209.495 ;
        RECT 73.505 209.325 73.675 209.495 ;
        RECT 73.965 209.325 74.135 209.495 ;
        RECT 74.425 209.325 74.595 209.495 ;
        RECT 74.885 209.325 75.055 209.495 ;
        RECT 75.345 209.325 75.515 209.495 ;
        RECT 75.805 209.325 75.975 209.495 ;
        RECT 76.265 209.325 76.435 209.495 ;
        RECT 76.725 209.325 76.895 209.495 ;
        RECT 77.185 209.325 77.355 209.495 ;
        RECT 77.645 209.325 77.815 209.495 ;
        RECT 78.105 209.325 78.275 209.495 ;
        RECT 78.565 209.325 78.735 209.495 ;
        RECT 79.025 209.325 79.195 209.495 ;
        RECT 79.485 209.325 79.655 209.495 ;
        RECT 79.945 209.325 80.115 209.495 ;
        RECT 80.405 209.325 80.575 209.495 ;
        RECT 80.865 209.325 81.035 209.495 ;
        RECT 81.325 209.325 81.495 209.495 ;
        RECT 81.785 209.325 81.955 209.495 ;
        RECT 82.245 209.325 82.415 209.495 ;
        RECT 82.705 209.325 82.875 209.495 ;
        RECT 83.165 209.325 83.335 209.495 ;
        RECT 83.625 209.325 83.795 209.495 ;
        RECT 84.085 209.325 84.255 209.495 ;
        RECT 84.545 209.325 84.715 209.495 ;
        RECT 85.005 209.325 85.175 209.495 ;
        RECT 85.465 209.325 85.635 209.495 ;
        RECT 85.925 209.325 86.095 209.495 ;
        RECT 86.385 209.325 86.555 209.495 ;
        RECT 86.845 209.325 87.015 209.495 ;
        RECT 87.305 209.325 87.475 209.495 ;
        RECT 87.765 209.325 87.935 209.495 ;
        RECT 88.225 209.325 88.395 209.495 ;
        RECT 88.685 209.325 88.855 209.495 ;
        RECT 89.145 209.325 89.315 209.495 ;
        RECT 89.605 209.325 89.775 209.495 ;
        RECT 90.065 209.325 90.235 209.495 ;
        RECT 90.525 209.325 90.695 209.495 ;
        RECT 90.985 209.325 91.155 209.495 ;
        RECT 91.445 209.325 91.615 209.495 ;
        RECT 91.905 209.325 92.075 209.495 ;
        RECT 92.365 209.325 92.535 209.495 ;
        RECT 92.825 209.325 92.995 209.495 ;
        RECT 93.285 209.325 93.455 209.495 ;
        RECT 93.745 209.325 93.915 209.495 ;
        RECT 94.205 209.325 94.375 209.495 ;
        RECT 94.665 209.325 94.835 209.495 ;
        RECT 95.125 209.325 95.295 209.495 ;
        RECT 95.585 209.325 95.755 209.495 ;
        RECT 96.045 209.325 96.215 209.495 ;
        RECT 96.505 209.325 96.675 209.495 ;
        RECT 96.965 209.325 97.135 209.495 ;
        RECT 97.425 209.325 97.595 209.495 ;
        RECT 97.885 209.325 98.055 209.495 ;
        RECT 98.345 209.325 98.515 209.495 ;
        RECT 98.805 209.325 98.975 209.495 ;
        RECT 99.265 209.325 99.435 209.495 ;
        RECT 99.725 209.325 99.895 209.495 ;
        RECT 100.185 209.325 100.355 209.495 ;
        RECT 100.645 209.325 100.815 209.495 ;
        RECT 101.105 209.325 101.275 209.495 ;
        RECT 101.565 209.325 101.735 209.495 ;
        RECT 102.025 209.325 102.195 209.495 ;
        RECT 102.485 209.325 102.655 209.495 ;
        RECT 102.945 209.325 103.115 209.495 ;
        RECT 103.405 209.325 103.575 209.495 ;
        RECT 103.865 209.325 104.035 209.495 ;
        RECT 104.325 209.325 104.495 209.495 ;
        RECT 104.785 209.325 104.955 209.495 ;
        RECT 105.245 209.325 105.415 209.495 ;
        RECT 105.705 209.325 105.875 209.495 ;
        RECT 106.165 209.325 106.335 209.495 ;
        RECT 106.625 209.325 106.795 209.495 ;
        RECT 107.085 209.325 107.255 209.495 ;
        RECT 107.545 209.325 107.715 209.495 ;
        RECT 108.005 209.325 108.175 209.495 ;
        RECT 108.465 209.325 108.635 209.495 ;
        RECT 108.925 209.325 109.095 209.495 ;
        RECT 109.385 209.325 109.555 209.495 ;
        RECT 109.845 209.325 110.015 209.495 ;
        RECT 110.305 209.325 110.475 209.495 ;
        RECT 110.765 209.325 110.935 209.495 ;
        RECT 111.225 209.325 111.395 209.495 ;
        RECT 111.685 209.325 111.855 209.495 ;
        RECT 112.145 209.325 112.315 209.495 ;
        RECT 112.605 209.325 112.775 209.495 ;
        RECT 113.065 209.325 113.235 209.495 ;
        RECT 113.525 209.325 113.695 209.495 ;
        RECT 113.985 209.325 114.155 209.495 ;
        RECT 114.445 209.325 114.615 209.495 ;
        RECT 114.905 209.325 115.075 209.495 ;
        RECT 115.365 209.325 115.535 209.495 ;
        RECT 115.825 209.325 115.995 209.495 ;
        RECT 116.285 209.325 116.455 209.495 ;
        RECT 116.745 209.325 116.915 209.495 ;
        RECT 117.205 209.325 117.375 209.495 ;
        RECT 117.665 209.325 117.835 209.495 ;
        RECT 118.125 209.325 118.295 209.495 ;
        RECT 118.585 209.325 118.755 209.495 ;
        RECT 119.045 209.325 119.215 209.495 ;
        RECT 119.505 209.325 119.675 209.495 ;
        RECT 119.965 209.325 120.135 209.495 ;
        RECT 120.425 209.325 120.595 209.495 ;
        RECT 120.885 209.325 121.055 209.495 ;
        RECT 121.345 209.325 121.515 209.495 ;
        RECT 121.805 209.325 121.975 209.495 ;
        RECT 122.265 209.325 122.435 209.495 ;
        RECT 122.725 209.325 122.895 209.495 ;
        RECT 123.185 209.325 123.355 209.495 ;
        RECT 123.645 209.325 123.815 209.495 ;
        RECT 124.105 209.325 124.275 209.495 ;
        RECT 124.565 209.325 124.735 209.495 ;
        RECT 125.025 209.325 125.195 209.495 ;
        RECT 125.485 209.325 125.655 209.495 ;
        RECT 125.945 209.325 126.115 209.495 ;
        RECT 126.405 209.325 126.575 209.495 ;
        RECT 126.865 209.325 127.035 209.495 ;
        RECT 127.325 209.325 127.495 209.495 ;
        RECT 127.785 209.325 127.955 209.495 ;
        RECT 128.245 209.325 128.415 209.495 ;
        RECT 128.705 209.325 128.875 209.495 ;
        RECT 129.165 209.325 129.335 209.495 ;
        RECT 129.625 209.325 129.795 209.495 ;
        RECT 130.085 209.325 130.255 209.495 ;
        RECT 130.545 209.325 130.715 209.495 ;
        RECT 131.005 209.325 131.175 209.495 ;
        RECT 131.465 209.325 131.635 209.495 ;
        RECT 131.925 209.325 132.095 209.495 ;
        RECT 132.385 209.325 132.555 209.495 ;
        RECT 132.845 209.325 133.015 209.495 ;
        RECT 133.305 209.325 133.475 209.495 ;
        RECT 133.765 209.325 133.935 209.495 ;
        RECT 134.225 209.325 134.395 209.495 ;
        RECT 134.685 209.325 134.855 209.495 ;
        RECT 135.145 209.325 135.315 209.495 ;
        RECT 135.605 209.325 135.775 209.495 ;
        RECT 136.065 209.325 136.235 209.495 ;
        RECT 136.525 209.325 136.695 209.495 ;
        RECT 136.985 209.325 137.155 209.495 ;
        RECT 137.445 209.325 137.615 209.495 ;
        RECT 137.905 209.325 138.075 209.495 ;
        RECT 138.365 209.325 138.535 209.495 ;
        RECT 138.825 209.325 138.995 209.495 ;
        RECT 139.285 209.325 139.455 209.495 ;
        RECT 139.745 209.325 139.915 209.495 ;
        RECT 140.205 209.325 140.375 209.495 ;
        RECT 140.665 209.325 140.835 209.495 ;
        RECT 141.125 209.325 141.295 209.495 ;
        RECT 141.585 209.325 141.755 209.495 ;
        RECT 142.045 209.325 142.215 209.495 ;
        RECT 142.505 209.325 142.675 209.495 ;
        RECT 142.965 209.325 143.135 209.495 ;
        RECT 143.425 209.325 143.595 209.495 ;
        RECT 143.885 209.325 144.055 209.495 ;
        RECT 144.345 209.325 144.515 209.495 ;
        RECT 144.805 209.325 144.975 209.495 ;
        RECT 145.265 209.325 145.435 209.495 ;
        RECT 145.725 209.325 145.895 209.495 ;
        RECT 146.185 209.325 146.355 209.495 ;
        RECT 146.645 209.325 146.815 209.495 ;
        RECT 147.105 209.325 147.275 209.495 ;
        RECT 147.565 209.325 147.735 209.495 ;
        RECT 148.025 209.325 148.195 209.495 ;
        RECT 148.485 209.325 148.655 209.495 ;
        RECT 148.945 209.325 149.115 209.495 ;
        RECT 149.405 209.325 149.575 209.495 ;
        RECT 149.865 209.325 150.035 209.495 ;
        RECT 42.685 208.815 42.855 208.985 ;
        RECT 42.685 207.795 42.855 207.965 ;
        RECT 43.605 207.795 43.775 207.965 ;
        RECT 44.065 207.795 44.235 207.965 ;
        RECT 44.985 207.795 45.155 207.965 ;
        RECT 47.745 208.815 47.915 208.985 ;
        RECT 46.825 207.795 46.995 207.965 ;
        RECT 45.905 207.115 46.075 207.285 ;
        RECT 57.865 207.115 58.035 207.285 ;
        RECT 60.175 208.135 60.345 208.305 ;
        RECT 60.610 208.475 60.780 208.645 ;
        RECT 62.180 208.475 62.350 208.645 ;
        RECT 62.695 208.135 62.865 208.305 ;
        RECT 63.540 207.455 63.710 207.625 ;
        RECT 63.885 208.135 64.055 208.305 ;
        RECT 64.280 208.475 64.450 208.645 ;
        RECT 65.225 208.475 65.395 208.645 ;
        RECT 64.765 207.795 64.935 207.965 ;
        RECT 66.145 207.455 66.315 207.625 ;
        RECT 72.585 208.815 72.755 208.985 ;
        RECT 72.585 207.795 72.755 207.965 ;
        RECT 75.805 208.815 75.975 208.985 ;
        RECT 73.505 207.795 73.675 207.965 ;
        RECT 75.345 207.795 75.515 207.965 ;
        RECT 76.725 207.795 76.895 207.965 ;
        RECT 77.645 208.135 77.815 208.305 ;
        RECT 78.565 208.815 78.735 208.985 ;
        RECT 82.245 208.815 82.415 208.985 ;
        RECT 78.105 207.795 78.275 207.965 ;
        RECT 81.325 207.455 81.495 207.625 ;
        RECT 85.005 208.135 85.175 208.305 ;
        RECT 84.545 207.795 84.715 207.965 ;
        RECT 86.385 208.475 86.555 208.645 ;
        RECT 88.225 208.815 88.395 208.985 ;
        RECT 86.845 207.795 87.015 207.965 ;
        RECT 87.765 207.795 87.935 207.965 ;
        RECT 88.685 208.135 88.855 208.305 ;
        RECT 90.525 208.475 90.695 208.645 ;
        RECT 89.145 207.795 89.315 207.965 ;
        RECT 90.985 207.795 91.155 207.965 ;
        RECT 91.905 207.795 92.075 207.965 ;
        RECT 91.445 207.115 91.615 207.285 ;
        RECT 98.805 207.795 98.975 207.965 ;
        RECT 102.025 208.475 102.195 208.645 ;
        RECT 99.265 207.795 99.435 207.965 ;
        RECT 99.725 207.795 99.895 207.965 ;
        RECT 102.485 207.795 102.655 207.965 ;
        RECT 103.405 207.795 103.575 207.965 ;
        RECT 106.165 208.815 106.335 208.985 ;
        RECT 107.085 207.795 107.255 207.965 ;
        RECT 110.305 208.135 110.475 208.305 ;
        RECT 111.685 208.135 111.855 208.305 ;
        RECT 114.905 208.815 115.075 208.985 ;
        RECT 117.205 208.135 117.375 208.305 ;
        RECT 118.125 208.135 118.295 208.305 ;
        RECT 121.345 208.815 121.515 208.985 ;
        RECT 119.965 207.795 120.135 207.965 ;
        RECT 120.425 207.795 120.595 207.965 ;
        RECT 119.045 207.115 119.215 207.285 ;
        RECT 122.725 207.795 122.895 207.965 ;
        RECT 124.565 208.815 124.735 208.985 ;
        RECT 125.025 208.135 125.195 208.305 ;
        RECT 127.785 208.815 127.955 208.985 ;
        RECT 123.645 207.795 123.815 207.965 ;
        RECT 127.785 207.795 127.955 207.965 ;
        RECT 128.705 207.795 128.875 207.965 ;
        RECT 130.545 208.135 130.715 208.305 ;
        RECT 131.465 208.135 131.635 208.305 ;
        RECT 126.865 207.115 127.035 207.285 ;
        RECT 131.925 207.795 132.095 207.965 ;
        RECT 133.765 208.815 133.935 208.985 ;
        RECT 136.525 208.135 136.695 208.305 ;
        RECT 137.445 207.795 137.615 207.965 ;
        RECT 36.245 206.605 36.415 206.775 ;
        RECT 36.705 206.605 36.875 206.775 ;
        RECT 37.165 206.605 37.335 206.775 ;
        RECT 37.625 206.605 37.795 206.775 ;
        RECT 38.085 206.605 38.255 206.775 ;
        RECT 38.545 206.605 38.715 206.775 ;
        RECT 39.005 206.605 39.175 206.775 ;
        RECT 39.465 206.605 39.635 206.775 ;
        RECT 39.925 206.605 40.095 206.775 ;
        RECT 40.385 206.605 40.555 206.775 ;
        RECT 40.845 206.605 41.015 206.775 ;
        RECT 41.305 206.605 41.475 206.775 ;
        RECT 41.765 206.605 41.935 206.775 ;
        RECT 42.225 206.605 42.395 206.775 ;
        RECT 42.685 206.605 42.855 206.775 ;
        RECT 43.145 206.605 43.315 206.775 ;
        RECT 43.605 206.605 43.775 206.775 ;
        RECT 44.065 206.605 44.235 206.775 ;
        RECT 44.525 206.605 44.695 206.775 ;
        RECT 44.985 206.605 45.155 206.775 ;
        RECT 45.445 206.605 45.615 206.775 ;
        RECT 45.905 206.605 46.075 206.775 ;
        RECT 46.365 206.605 46.535 206.775 ;
        RECT 46.825 206.605 46.995 206.775 ;
        RECT 47.285 206.605 47.455 206.775 ;
        RECT 47.745 206.605 47.915 206.775 ;
        RECT 48.205 206.605 48.375 206.775 ;
        RECT 48.665 206.605 48.835 206.775 ;
        RECT 49.125 206.605 49.295 206.775 ;
        RECT 49.585 206.605 49.755 206.775 ;
        RECT 50.045 206.605 50.215 206.775 ;
        RECT 50.505 206.605 50.675 206.775 ;
        RECT 50.965 206.605 51.135 206.775 ;
        RECT 51.425 206.605 51.595 206.775 ;
        RECT 51.885 206.605 52.055 206.775 ;
        RECT 52.345 206.605 52.515 206.775 ;
        RECT 52.805 206.605 52.975 206.775 ;
        RECT 53.265 206.605 53.435 206.775 ;
        RECT 53.725 206.605 53.895 206.775 ;
        RECT 54.185 206.605 54.355 206.775 ;
        RECT 54.645 206.605 54.815 206.775 ;
        RECT 55.105 206.605 55.275 206.775 ;
        RECT 55.565 206.605 55.735 206.775 ;
        RECT 56.025 206.605 56.195 206.775 ;
        RECT 56.485 206.605 56.655 206.775 ;
        RECT 56.945 206.605 57.115 206.775 ;
        RECT 57.405 206.605 57.575 206.775 ;
        RECT 57.865 206.605 58.035 206.775 ;
        RECT 58.325 206.605 58.495 206.775 ;
        RECT 58.785 206.605 58.955 206.775 ;
        RECT 59.245 206.605 59.415 206.775 ;
        RECT 59.705 206.605 59.875 206.775 ;
        RECT 60.165 206.605 60.335 206.775 ;
        RECT 60.625 206.605 60.795 206.775 ;
        RECT 61.085 206.605 61.255 206.775 ;
        RECT 61.545 206.605 61.715 206.775 ;
        RECT 62.005 206.605 62.175 206.775 ;
        RECT 62.465 206.605 62.635 206.775 ;
        RECT 62.925 206.605 63.095 206.775 ;
        RECT 63.385 206.605 63.555 206.775 ;
        RECT 63.845 206.605 64.015 206.775 ;
        RECT 64.305 206.605 64.475 206.775 ;
        RECT 64.765 206.605 64.935 206.775 ;
        RECT 65.225 206.605 65.395 206.775 ;
        RECT 65.685 206.605 65.855 206.775 ;
        RECT 66.145 206.605 66.315 206.775 ;
        RECT 66.605 206.605 66.775 206.775 ;
        RECT 67.065 206.605 67.235 206.775 ;
        RECT 67.525 206.605 67.695 206.775 ;
        RECT 67.985 206.605 68.155 206.775 ;
        RECT 68.445 206.605 68.615 206.775 ;
        RECT 68.905 206.605 69.075 206.775 ;
        RECT 69.365 206.605 69.535 206.775 ;
        RECT 69.825 206.605 69.995 206.775 ;
        RECT 70.285 206.605 70.455 206.775 ;
        RECT 70.745 206.605 70.915 206.775 ;
        RECT 71.205 206.605 71.375 206.775 ;
        RECT 71.665 206.605 71.835 206.775 ;
        RECT 72.125 206.605 72.295 206.775 ;
        RECT 72.585 206.605 72.755 206.775 ;
        RECT 73.045 206.605 73.215 206.775 ;
        RECT 73.505 206.605 73.675 206.775 ;
        RECT 73.965 206.605 74.135 206.775 ;
        RECT 74.425 206.605 74.595 206.775 ;
        RECT 74.885 206.605 75.055 206.775 ;
        RECT 75.345 206.605 75.515 206.775 ;
        RECT 75.805 206.605 75.975 206.775 ;
        RECT 76.265 206.605 76.435 206.775 ;
        RECT 76.725 206.605 76.895 206.775 ;
        RECT 77.185 206.605 77.355 206.775 ;
        RECT 77.645 206.605 77.815 206.775 ;
        RECT 78.105 206.605 78.275 206.775 ;
        RECT 78.565 206.605 78.735 206.775 ;
        RECT 79.025 206.605 79.195 206.775 ;
        RECT 79.485 206.605 79.655 206.775 ;
        RECT 79.945 206.605 80.115 206.775 ;
        RECT 80.405 206.605 80.575 206.775 ;
        RECT 80.865 206.605 81.035 206.775 ;
        RECT 81.325 206.605 81.495 206.775 ;
        RECT 81.785 206.605 81.955 206.775 ;
        RECT 82.245 206.605 82.415 206.775 ;
        RECT 82.705 206.605 82.875 206.775 ;
        RECT 83.165 206.605 83.335 206.775 ;
        RECT 83.625 206.605 83.795 206.775 ;
        RECT 84.085 206.605 84.255 206.775 ;
        RECT 84.545 206.605 84.715 206.775 ;
        RECT 85.005 206.605 85.175 206.775 ;
        RECT 85.465 206.605 85.635 206.775 ;
        RECT 85.925 206.605 86.095 206.775 ;
        RECT 86.385 206.605 86.555 206.775 ;
        RECT 86.845 206.605 87.015 206.775 ;
        RECT 87.305 206.605 87.475 206.775 ;
        RECT 87.765 206.605 87.935 206.775 ;
        RECT 88.225 206.605 88.395 206.775 ;
        RECT 88.685 206.605 88.855 206.775 ;
        RECT 89.145 206.605 89.315 206.775 ;
        RECT 89.605 206.605 89.775 206.775 ;
        RECT 90.065 206.605 90.235 206.775 ;
        RECT 90.525 206.605 90.695 206.775 ;
        RECT 90.985 206.605 91.155 206.775 ;
        RECT 91.445 206.605 91.615 206.775 ;
        RECT 91.905 206.605 92.075 206.775 ;
        RECT 92.365 206.605 92.535 206.775 ;
        RECT 92.825 206.605 92.995 206.775 ;
        RECT 93.285 206.605 93.455 206.775 ;
        RECT 93.745 206.605 93.915 206.775 ;
        RECT 94.205 206.605 94.375 206.775 ;
        RECT 94.665 206.605 94.835 206.775 ;
        RECT 95.125 206.605 95.295 206.775 ;
        RECT 95.585 206.605 95.755 206.775 ;
        RECT 96.045 206.605 96.215 206.775 ;
        RECT 96.505 206.605 96.675 206.775 ;
        RECT 96.965 206.605 97.135 206.775 ;
        RECT 97.425 206.605 97.595 206.775 ;
        RECT 97.885 206.605 98.055 206.775 ;
        RECT 98.345 206.605 98.515 206.775 ;
        RECT 98.805 206.605 98.975 206.775 ;
        RECT 99.265 206.605 99.435 206.775 ;
        RECT 99.725 206.605 99.895 206.775 ;
        RECT 100.185 206.605 100.355 206.775 ;
        RECT 100.645 206.605 100.815 206.775 ;
        RECT 101.105 206.605 101.275 206.775 ;
        RECT 101.565 206.605 101.735 206.775 ;
        RECT 102.025 206.605 102.195 206.775 ;
        RECT 102.485 206.605 102.655 206.775 ;
        RECT 102.945 206.605 103.115 206.775 ;
        RECT 103.405 206.605 103.575 206.775 ;
        RECT 103.865 206.605 104.035 206.775 ;
        RECT 104.325 206.605 104.495 206.775 ;
        RECT 104.785 206.605 104.955 206.775 ;
        RECT 105.245 206.605 105.415 206.775 ;
        RECT 105.705 206.605 105.875 206.775 ;
        RECT 106.165 206.605 106.335 206.775 ;
        RECT 106.625 206.605 106.795 206.775 ;
        RECT 107.085 206.605 107.255 206.775 ;
        RECT 107.545 206.605 107.715 206.775 ;
        RECT 108.005 206.605 108.175 206.775 ;
        RECT 108.465 206.605 108.635 206.775 ;
        RECT 108.925 206.605 109.095 206.775 ;
        RECT 109.385 206.605 109.555 206.775 ;
        RECT 109.845 206.605 110.015 206.775 ;
        RECT 110.305 206.605 110.475 206.775 ;
        RECT 110.765 206.605 110.935 206.775 ;
        RECT 111.225 206.605 111.395 206.775 ;
        RECT 111.685 206.605 111.855 206.775 ;
        RECT 112.145 206.605 112.315 206.775 ;
        RECT 112.605 206.605 112.775 206.775 ;
        RECT 113.065 206.605 113.235 206.775 ;
        RECT 113.525 206.605 113.695 206.775 ;
        RECT 113.985 206.605 114.155 206.775 ;
        RECT 114.445 206.605 114.615 206.775 ;
        RECT 114.905 206.605 115.075 206.775 ;
        RECT 115.365 206.605 115.535 206.775 ;
        RECT 115.825 206.605 115.995 206.775 ;
        RECT 116.285 206.605 116.455 206.775 ;
        RECT 116.745 206.605 116.915 206.775 ;
        RECT 117.205 206.605 117.375 206.775 ;
        RECT 117.665 206.605 117.835 206.775 ;
        RECT 118.125 206.605 118.295 206.775 ;
        RECT 118.585 206.605 118.755 206.775 ;
        RECT 119.045 206.605 119.215 206.775 ;
        RECT 119.505 206.605 119.675 206.775 ;
        RECT 119.965 206.605 120.135 206.775 ;
        RECT 120.425 206.605 120.595 206.775 ;
        RECT 120.885 206.605 121.055 206.775 ;
        RECT 121.345 206.605 121.515 206.775 ;
        RECT 121.805 206.605 121.975 206.775 ;
        RECT 122.265 206.605 122.435 206.775 ;
        RECT 122.725 206.605 122.895 206.775 ;
        RECT 123.185 206.605 123.355 206.775 ;
        RECT 123.645 206.605 123.815 206.775 ;
        RECT 124.105 206.605 124.275 206.775 ;
        RECT 124.565 206.605 124.735 206.775 ;
        RECT 125.025 206.605 125.195 206.775 ;
        RECT 125.485 206.605 125.655 206.775 ;
        RECT 125.945 206.605 126.115 206.775 ;
        RECT 126.405 206.605 126.575 206.775 ;
        RECT 126.865 206.605 127.035 206.775 ;
        RECT 127.325 206.605 127.495 206.775 ;
        RECT 127.785 206.605 127.955 206.775 ;
        RECT 128.245 206.605 128.415 206.775 ;
        RECT 128.705 206.605 128.875 206.775 ;
        RECT 129.165 206.605 129.335 206.775 ;
        RECT 129.625 206.605 129.795 206.775 ;
        RECT 130.085 206.605 130.255 206.775 ;
        RECT 130.545 206.605 130.715 206.775 ;
        RECT 131.005 206.605 131.175 206.775 ;
        RECT 131.465 206.605 131.635 206.775 ;
        RECT 131.925 206.605 132.095 206.775 ;
        RECT 132.385 206.605 132.555 206.775 ;
        RECT 132.845 206.605 133.015 206.775 ;
        RECT 133.305 206.605 133.475 206.775 ;
        RECT 133.765 206.605 133.935 206.775 ;
        RECT 134.225 206.605 134.395 206.775 ;
        RECT 134.685 206.605 134.855 206.775 ;
        RECT 135.145 206.605 135.315 206.775 ;
        RECT 135.605 206.605 135.775 206.775 ;
        RECT 136.065 206.605 136.235 206.775 ;
        RECT 136.525 206.605 136.695 206.775 ;
        RECT 136.985 206.605 137.155 206.775 ;
        RECT 137.445 206.605 137.615 206.775 ;
        RECT 137.905 206.605 138.075 206.775 ;
        RECT 138.365 206.605 138.535 206.775 ;
        RECT 138.825 206.605 138.995 206.775 ;
        RECT 139.285 206.605 139.455 206.775 ;
        RECT 139.745 206.605 139.915 206.775 ;
        RECT 140.205 206.605 140.375 206.775 ;
        RECT 140.665 206.605 140.835 206.775 ;
        RECT 141.125 206.605 141.295 206.775 ;
        RECT 141.585 206.605 141.755 206.775 ;
        RECT 142.045 206.605 142.215 206.775 ;
        RECT 142.505 206.605 142.675 206.775 ;
        RECT 142.965 206.605 143.135 206.775 ;
        RECT 143.425 206.605 143.595 206.775 ;
        RECT 143.885 206.605 144.055 206.775 ;
        RECT 144.345 206.605 144.515 206.775 ;
        RECT 144.805 206.605 144.975 206.775 ;
        RECT 145.265 206.605 145.435 206.775 ;
        RECT 145.725 206.605 145.895 206.775 ;
        RECT 146.185 206.605 146.355 206.775 ;
        RECT 146.645 206.605 146.815 206.775 ;
        RECT 147.105 206.605 147.275 206.775 ;
        RECT 147.565 206.605 147.735 206.775 ;
        RECT 148.025 206.605 148.195 206.775 ;
        RECT 148.485 206.605 148.655 206.775 ;
        RECT 148.945 206.605 149.115 206.775 ;
        RECT 149.405 206.605 149.575 206.775 ;
        RECT 149.865 206.605 150.035 206.775 ;
        RECT 42.685 205.755 42.855 205.925 ;
        RECT 43.765 205.755 43.935 205.925 ;
        RECT 44.985 205.415 45.155 205.585 ;
        RECT 43.605 204.395 43.775 204.565 ;
        RECT 44.525 204.395 44.695 204.565 ;
        RECT 45.470 204.735 45.640 204.905 ;
        RECT 45.865 205.075 46.035 205.245 ;
        RECT 46.320 205.755 46.490 205.925 ;
        RECT 47.055 205.075 47.225 205.245 ;
        RECT 47.570 204.735 47.740 204.905 ;
        RECT 49.140 204.735 49.310 204.905 ;
        RECT 49.575 205.075 49.745 205.245 ;
        RECT 51.885 204.395 52.055 204.565 ;
        RECT 64.765 205.415 64.935 205.585 ;
        RECT 65.225 205.415 65.395 205.585 ;
        RECT 63.845 204.395 64.015 204.565 ;
        RECT 65.685 204.395 65.855 204.565 ;
        RECT 72.585 206.095 72.755 206.265 ;
        RECT 71.665 205.415 71.835 205.585 ;
        RECT 72.585 205.415 72.755 205.585 ;
        RECT 77.185 205.415 77.355 205.585 ;
        RECT 78.105 204.395 78.275 204.565 ;
        RECT 84.085 205.415 84.255 205.585 ;
        RECT 85.465 205.755 85.635 205.925 ;
        RECT 85.005 205.415 85.175 205.585 ;
        RECT 86.385 205.415 86.555 205.585 ;
        RECT 84.545 204.395 84.715 204.565 ;
        RECT 89.145 205.415 89.315 205.585 ;
        RECT 87.305 204.395 87.475 204.565 ;
        RECT 88.685 205.075 88.855 205.245 ;
        RECT 90.525 204.735 90.695 204.905 ;
        RECT 91.905 205.075 92.075 205.245 ;
        RECT 113.985 205.755 114.155 205.925 ;
        RECT 114.905 205.415 115.075 205.585 ;
        RECT 115.825 204.735 115.995 204.905 ;
        RECT 117.665 205.415 117.835 205.585 ;
        RECT 119.045 205.415 119.215 205.585 ;
        RECT 116.745 204.395 116.915 204.565 ;
        RECT 118.585 204.395 118.755 204.565 ;
        RECT 122.725 206.095 122.895 206.265 ;
        RECT 122.265 205.415 122.435 205.585 ;
        RECT 121.345 204.395 121.515 204.565 ;
        RECT 125.485 206.095 125.655 206.265 ;
        RECT 123.645 205.415 123.815 205.585 ;
        RECT 125.025 205.075 125.195 205.245 ;
        RECT 125.945 206.095 126.115 206.265 ;
        RECT 127.785 206.095 127.955 206.265 ;
        RECT 129.165 206.095 129.335 206.265 ;
        RECT 129.625 205.415 129.795 205.585 ;
        RECT 133.305 205.415 133.475 205.585 ;
        RECT 141.125 206.095 141.295 206.265 ;
        RECT 140.205 205.415 140.375 205.585 ;
        RECT 134.225 204.395 134.395 204.565 ;
        RECT 141.585 205.075 141.755 205.245 ;
        RECT 142.070 204.735 142.240 204.905 ;
        RECT 142.465 205.075 142.635 205.245 ;
        RECT 142.810 205.755 142.980 205.925 ;
        RECT 143.655 205.075 143.825 205.245 ;
        RECT 144.170 204.735 144.340 204.905 ;
        RECT 145.740 204.735 145.910 204.905 ;
        RECT 146.175 205.075 146.345 205.245 ;
        RECT 148.485 204.395 148.655 204.565 ;
        RECT 36.245 203.885 36.415 204.055 ;
        RECT 36.705 203.885 36.875 204.055 ;
        RECT 37.165 203.885 37.335 204.055 ;
        RECT 37.625 203.885 37.795 204.055 ;
        RECT 38.085 203.885 38.255 204.055 ;
        RECT 38.545 203.885 38.715 204.055 ;
        RECT 39.005 203.885 39.175 204.055 ;
        RECT 39.465 203.885 39.635 204.055 ;
        RECT 39.925 203.885 40.095 204.055 ;
        RECT 40.385 203.885 40.555 204.055 ;
        RECT 40.845 203.885 41.015 204.055 ;
        RECT 41.305 203.885 41.475 204.055 ;
        RECT 41.765 203.885 41.935 204.055 ;
        RECT 42.225 203.885 42.395 204.055 ;
        RECT 42.685 203.885 42.855 204.055 ;
        RECT 43.145 203.885 43.315 204.055 ;
        RECT 43.605 203.885 43.775 204.055 ;
        RECT 44.065 203.885 44.235 204.055 ;
        RECT 44.525 203.885 44.695 204.055 ;
        RECT 44.985 203.885 45.155 204.055 ;
        RECT 45.445 203.885 45.615 204.055 ;
        RECT 45.905 203.885 46.075 204.055 ;
        RECT 46.365 203.885 46.535 204.055 ;
        RECT 46.825 203.885 46.995 204.055 ;
        RECT 47.285 203.885 47.455 204.055 ;
        RECT 47.745 203.885 47.915 204.055 ;
        RECT 48.205 203.885 48.375 204.055 ;
        RECT 48.665 203.885 48.835 204.055 ;
        RECT 49.125 203.885 49.295 204.055 ;
        RECT 49.585 203.885 49.755 204.055 ;
        RECT 50.045 203.885 50.215 204.055 ;
        RECT 50.505 203.885 50.675 204.055 ;
        RECT 50.965 203.885 51.135 204.055 ;
        RECT 51.425 203.885 51.595 204.055 ;
        RECT 51.885 203.885 52.055 204.055 ;
        RECT 52.345 203.885 52.515 204.055 ;
        RECT 52.805 203.885 52.975 204.055 ;
        RECT 53.265 203.885 53.435 204.055 ;
        RECT 53.725 203.885 53.895 204.055 ;
        RECT 54.185 203.885 54.355 204.055 ;
        RECT 54.645 203.885 54.815 204.055 ;
        RECT 55.105 203.885 55.275 204.055 ;
        RECT 55.565 203.885 55.735 204.055 ;
        RECT 56.025 203.885 56.195 204.055 ;
        RECT 56.485 203.885 56.655 204.055 ;
        RECT 56.945 203.885 57.115 204.055 ;
        RECT 57.405 203.885 57.575 204.055 ;
        RECT 57.865 203.885 58.035 204.055 ;
        RECT 58.325 203.885 58.495 204.055 ;
        RECT 58.785 203.885 58.955 204.055 ;
        RECT 59.245 203.885 59.415 204.055 ;
        RECT 59.705 203.885 59.875 204.055 ;
        RECT 60.165 203.885 60.335 204.055 ;
        RECT 60.625 203.885 60.795 204.055 ;
        RECT 61.085 203.885 61.255 204.055 ;
        RECT 61.545 203.885 61.715 204.055 ;
        RECT 62.005 203.885 62.175 204.055 ;
        RECT 62.465 203.885 62.635 204.055 ;
        RECT 62.925 203.885 63.095 204.055 ;
        RECT 63.385 203.885 63.555 204.055 ;
        RECT 63.845 203.885 64.015 204.055 ;
        RECT 64.305 203.885 64.475 204.055 ;
        RECT 64.765 203.885 64.935 204.055 ;
        RECT 65.225 203.885 65.395 204.055 ;
        RECT 65.685 203.885 65.855 204.055 ;
        RECT 66.145 203.885 66.315 204.055 ;
        RECT 66.605 203.885 66.775 204.055 ;
        RECT 67.065 203.885 67.235 204.055 ;
        RECT 67.525 203.885 67.695 204.055 ;
        RECT 67.985 203.885 68.155 204.055 ;
        RECT 68.445 203.885 68.615 204.055 ;
        RECT 68.905 203.885 69.075 204.055 ;
        RECT 69.365 203.885 69.535 204.055 ;
        RECT 69.825 203.885 69.995 204.055 ;
        RECT 70.285 203.885 70.455 204.055 ;
        RECT 70.745 203.885 70.915 204.055 ;
        RECT 71.205 203.885 71.375 204.055 ;
        RECT 71.665 203.885 71.835 204.055 ;
        RECT 72.125 203.885 72.295 204.055 ;
        RECT 72.585 203.885 72.755 204.055 ;
        RECT 73.045 203.885 73.215 204.055 ;
        RECT 73.505 203.885 73.675 204.055 ;
        RECT 73.965 203.885 74.135 204.055 ;
        RECT 74.425 203.885 74.595 204.055 ;
        RECT 74.885 203.885 75.055 204.055 ;
        RECT 75.345 203.885 75.515 204.055 ;
        RECT 75.805 203.885 75.975 204.055 ;
        RECT 76.265 203.885 76.435 204.055 ;
        RECT 76.725 203.885 76.895 204.055 ;
        RECT 77.185 203.885 77.355 204.055 ;
        RECT 77.645 203.885 77.815 204.055 ;
        RECT 78.105 203.885 78.275 204.055 ;
        RECT 78.565 203.885 78.735 204.055 ;
        RECT 79.025 203.885 79.195 204.055 ;
        RECT 79.485 203.885 79.655 204.055 ;
        RECT 79.945 203.885 80.115 204.055 ;
        RECT 80.405 203.885 80.575 204.055 ;
        RECT 80.865 203.885 81.035 204.055 ;
        RECT 81.325 203.885 81.495 204.055 ;
        RECT 81.785 203.885 81.955 204.055 ;
        RECT 82.245 203.885 82.415 204.055 ;
        RECT 82.705 203.885 82.875 204.055 ;
        RECT 83.165 203.885 83.335 204.055 ;
        RECT 83.625 203.885 83.795 204.055 ;
        RECT 84.085 203.885 84.255 204.055 ;
        RECT 84.545 203.885 84.715 204.055 ;
        RECT 85.005 203.885 85.175 204.055 ;
        RECT 85.465 203.885 85.635 204.055 ;
        RECT 85.925 203.885 86.095 204.055 ;
        RECT 86.385 203.885 86.555 204.055 ;
        RECT 86.845 203.885 87.015 204.055 ;
        RECT 87.305 203.885 87.475 204.055 ;
        RECT 87.765 203.885 87.935 204.055 ;
        RECT 88.225 203.885 88.395 204.055 ;
        RECT 88.685 203.885 88.855 204.055 ;
        RECT 89.145 203.885 89.315 204.055 ;
        RECT 89.605 203.885 89.775 204.055 ;
        RECT 90.065 203.885 90.235 204.055 ;
        RECT 90.525 203.885 90.695 204.055 ;
        RECT 90.985 203.885 91.155 204.055 ;
        RECT 91.445 203.885 91.615 204.055 ;
        RECT 91.905 203.885 92.075 204.055 ;
        RECT 92.365 203.885 92.535 204.055 ;
        RECT 92.825 203.885 92.995 204.055 ;
        RECT 93.285 203.885 93.455 204.055 ;
        RECT 93.745 203.885 93.915 204.055 ;
        RECT 94.205 203.885 94.375 204.055 ;
        RECT 94.665 203.885 94.835 204.055 ;
        RECT 95.125 203.885 95.295 204.055 ;
        RECT 95.585 203.885 95.755 204.055 ;
        RECT 96.045 203.885 96.215 204.055 ;
        RECT 96.505 203.885 96.675 204.055 ;
        RECT 96.965 203.885 97.135 204.055 ;
        RECT 97.425 203.885 97.595 204.055 ;
        RECT 97.885 203.885 98.055 204.055 ;
        RECT 98.345 203.885 98.515 204.055 ;
        RECT 98.805 203.885 98.975 204.055 ;
        RECT 99.265 203.885 99.435 204.055 ;
        RECT 99.725 203.885 99.895 204.055 ;
        RECT 100.185 203.885 100.355 204.055 ;
        RECT 100.645 203.885 100.815 204.055 ;
        RECT 101.105 203.885 101.275 204.055 ;
        RECT 101.565 203.885 101.735 204.055 ;
        RECT 102.025 203.885 102.195 204.055 ;
        RECT 102.485 203.885 102.655 204.055 ;
        RECT 102.945 203.885 103.115 204.055 ;
        RECT 103.405 203.885 103.575 204.055 ;
        RECT 103.865 203.885 104.035 204.055 ;
        RECT 104.325 203.885 104.495 204.055 ;
        RECT 104.785 203.885 104.955 204.055 ;
        RECT 105.245 203.885 105.415 204.055 ;
        RECT 105.705 203.885 105.875 204.055 ;
        RECT 106.165 203.885 106.335 204.055 ;
        RECT 106.625 203.885 106.795 204.055 ;
        RECT 107.085 203.885 107.255 204.055 ;
        RECT 107.545 203.885 107.715 204.055 ;
        RECT 108.005 203.885 108.175 204.055 ;
        RECT 108.465 203.885 108.635 204.055 ;
        RECT 108.925 203.885 109.095 204.055 ;
        RECT 109.385 203.885 109.555 204.055 ;
        RECT 109.845 203.885 110.015 204.055 ;
        RECT 110.305 203.885 110.475 204.055 ;
        RECT 110.765 203.885 110.935 204.055 ;
        RECT 111.225 203.885 111.395 204.055 ;
        RECT 111.685 203.885 111.855 204.055 ;
        RECT 112.145 203.885 112.315 204.055 ;
        RECT 112.605 203.885 112.775 204.055 ;
        RECT 113.065 203.885 113.235 204.055 ;
        RECT 113.525 203.885 113.695 204.055 ;
        RECT 113.985 203.885 114.155 204.055 ;
        RECT 114.445 203.885 114.615 204.055 ;
        RECT 114.905 203.885 115.075 204.055 ;
        RECT 115.365 203.885 115.535 204.055 ;
        RECT 115.825 203.885 115.995 204.055 ;
        RECT 116.285 203.885 116.455 204.055 ;
        RECT 116.745 203.885 116.915 204.055 ;
        RECT 117.205 203.885 117.375 204.055 ;
        RECT 117.665 203.885 117.835 204.055 ;
        RECT 118.125 203.885 118.295 204.055 ;
        RECT 118.585 203.885 118.755 204.055 ;
        RECT 119.045 203.885 119.215 204.055 ;
        RECT 119.505 203.885 119.675 204.055 ;
        RECT 119.965 203.885 120.135 204.055 ;
        RECT 120.425 203.885 120.595 204.055 ;
        RECT 120.885 203.885 121.055 204.055 ;
        RECT 121.345 203.885 121.515 204.055 ;
        RECT 121.805 203.885 121.975 204.055 ;
        RECT 122.265 203.885 122.435 204.055 ;
        RECT 122.725 203.885 122.895 204.055 ;
        RECT 123.185 203.885 123.355 204.055 ;
        RECT 123.645 203.885 123.815 204.055 ;
        RECT 124.105 203.885 124.275 204.055 ;
        RECT 124.565 203.885 124.735 204.055 ;
        RECT 125.025 203.885 125.195 204.055 ;
        RECT 125.485 203.885 125.655 204.055 ;
        RECT 125.945 203.885 126.115 204.055 ;
        RECT 126.405 203.885 126.575 204.055 ;
        RECT 126.865 203.885 127.035 204.055 ;
        RECT 127.325 203.885 127.495 204.055 ;
        RECT 127.785 203.885 127.955 204.055 ;
        RECT 128.245 203.885 128.415 204.055 ;
        RECT 128.705 203.885 128.875 204.055 ;
        RECT 129.165 203.885 129.335 204.055 ;
        RECT 129.625 203.885 129.795 204.055 ;
        RECT 130.085 203.885 130.255 204.055 ;
        RECT 130.545 203.885 130.715 204.055 ;
        RECT 131.005 203.885 131.175 204.055 ;
        RECT 131.465 203.885 131.635 204.055 ;
        RECT 131.925 203.885 132.095 204.055 ;
        RECT 132.385 203.885 132.555 204.055 ;
        RECT 132.845 203.885 133.015 204.055 ;
        RECT 133.305 203.885 133.475 204.055 ;
        RECT 133.765 203.885 133.935 204.055 ;
        RECT 134.225 203.885 134.395 204.055 ;
        RECT 134.685 203.885 134.855 204.055 ;
        RECT 135.145 203.885 135.315 204.055 ;
        RECT 135.605 203.885 135.775 204.055 ;
        RECT 136.065 203.885 136.235 204.055 ;
        RECT 136.525 203.885 136.695 204.055 ;
        RECT 136.985 203.885 137.155 204.055 ;
        RECT 137.445 203.885 137.615 204.055 ;
        RECT 137.905 203.885 138.075 204.055 ;
        RECT 138.365 203.885 138.535 204.055 ;
        RECT 138.825 203.885 138.995 204.055 ;
        RECT 139.285 203.885 139.455 204.055 ;
        RECT 139.745 203.885 139.915 204.055 ;
        RECT 140.205 203.885 140.375 204.055 ;
        RECT 140.665 203.885 140.835 204.055 ;
        RECT 141.125 203.885 141.295 204.055 ;
        RECT 141.585 203.885 141.755 204.055 ;
        RECT 142.045 203.885 142.215 204.055 ;
        RECT 142.505 203.885 142.675 204.055 ;
        RECT 142.965 203.885 143.135 204.055 ;
        RECT 143.425 203.885 143.595 204.055 ;
        RECT 143.885 203.885 144.055 204.055 ;
        RECT 144.345 203.885 144.515 204.055 ;
        RECT 144.805 203.885 144.975 204.055 ;
        RECT 145.265 203.885 145.435 204.055 ;
        RECT 145.725 203.885 145.895 204.055 ;
        RECT 146.185 203.885 146.355 204.055 ;
        RECT 146.645 203.885 146.815 204.055 ;
        RECT 147.105 203.885 147.275 204.055 ;
        RECT 147.565 203.885 147.735 204.055 ;
        RECT 148.025 203.885 148.195 204.055 ;
        RECT 148.485 203.885 148.655 204.055 ;
        RECT 148.945 203.885 149.115 204.055 ;
        RECT 149.405 203.885 149.575 204.055 ;
        RECT 149.865 203.885 150.035 204.055 ;
        RECT 39.925 203.035 40.095 203.205 ;
        RECT 41.765 203.375 41.935 203.545 ;
        RECT 42.685 203.375 42.855 203.545 ;
        RECT 39.465 202.355 39.635 202.525 ;
        RECT 40.385 202.355 40.555 202.525 ;
        RECT 40.845 202.015 41.015 202.185 ;
        RECT 44.985 203.375 45.155 203.545 ;
        RECT 43.145 202.355 43.315 202.525 ;
        RECT 41.845 201.675 42.015 201.845 ;
        RECT 44.065 202.355 44.235 202.525 ;
        RECT 45.445 202.355 45.615 202.525 ;
        RECT 46.365 202.355 46.535 202.525 ;
        RECT 46.825 202.355 46.995 202.525 ;
        RECT 47.515 202.355 47.685 202.525 ;
        RECT 50.045 203.375 50.215 203.545 ;
        RECT 51.450 203.035 51.620 203.205 ;
        RECT 49.585 202.355 49.755 202.525 ;
        RECT 50.965 202.695 51.135 202.865 ;
        RECT 50.505 202.355 50.675 202.525 ;
        RECT 48.665 201.675 48.835 201.845 ;
        RECT 51.845 202.695 52.015 202.865 ;
        RECT 52.245 202.015 52.415 202.185 ;
        RECT 53.550 203.035 53.720 203.205 ;
        RECT 53.035 202.695 53.205 202.865 ;
        RECT 55.120 203.035 55.290 203.205 ;
        RECT 55.555 202.695 55.725 202.865 ;
        RECT 59.245 202.695 59.415 202.865 ;
        RECT 60.165 202.695 60.335 202.865 ;
        RECT 57.865 201.675 58.035 201.845 ;
        RECT 60.625 202.355 60.795 202.525 ;
        RECT 62.465 201.675 62.635 201.845 ;
        RECT 62.925 203.375 63.095 203.545 ;
        RECT 63.845 202.355 64.015 202.525 ;
        RECT 64.305 202.355 64.475 202.525 ;
        RECT 64.765 203.035 64.935 203.205 ;
        RECT 65.225 202.355 65.395 202.525 ;
        RECT 68.010 203.035 68.180 203.205 ;
        RECT 66.145 202.355 66.315 202.525 ;
        RECT 67.065 202.355 67.235 202.525 ;
        RECT 67.525 202.355 67.695 202.525 ;
        RECT 66.605 202.015 66.775 202.185 ;
        RECT 68.405 202.695 68.575 202.865 ;
        RECT 68.860 202.015 69.030 202.185 ;
        RECT 70.110 203.035 70.280 203.205 ;
        RECT 69.595 202.695 69.765 202.865 ;
        RECT 71.680 203.035 71.850 203.205 ;
        RECT 72.115 202.695 72.285 202.865 ;
        RECT 79.485 203.375 79.655 203.545 ;
        RECT 74.425 201.675 74.595 201.845 ;
        RECT 81.325 202.695 81.495 202.865 ;
        RECT 80.405 202.355 80.575 202.525 ;
        RECT 81.785 202.355 81.955 202.525 ;
        RECT 86.385 202.695 86.555 202.865 ;
        RECT 87.305 202.355 87.475 202.525 ;
        RECT 87.765 202.695 87.935 202.865 ;
        RECT 88.225 202.355 88.395 202.525 ;
        RECT 88.685 202.695 88.855 202.865 ;
        RECT 89.605 202.695 89.775 202.865 ;
        RECT 90.525 202.355 90.695 202.525 ;
        RECT 91.445 202.355 91.615 202.525 ;
        RECT 91.905 202.355 92.075 202.525 ;
        RECT 97.885 203.035 98.055 203.205 ;
        RECT 99.725 202.695 99.895 202.865 ;
        RECT 100.185 202.695 100.355 202.865 ;
        RECT 101.565 203.375 101.735 203.545 ;
        RECT 98.805 202.355 98.975 202.525 ;
        RECT 102.485 202.695 102.655 202.865 ;
        RECT 102.945 202.355 103.115 202.525 ;
        RECT 104.325 202.695 104.495 202.865 ;
        RECT 104.785 202.355 104.955 202.525 ;
        RECT 105.705 202.355 105.875 202.525 ;
        RECT 116.285 203.375 116.455 203.545 ;
        RECT 106.625 201.675 106.795 201.845 ;
        RECT 115.365 202.355 115.535 202.525 ;
        RECT 116.745 202.355 116.915 202.525 ;
        RECT 114.445 201.675 114.615 201.845 ;
        RECT 125.485 203.375 125.655 203.545 ;
        RECT 124.565 202.355 124.735 202.525 ;
        RECT 125.945 202.355 126.115 202.525 ;
        RECT 123.645 201.675 123.815 201.845 ;
        RECT 131.465 203.035 131.635 203.205 ;
        RECT 129.625 202.355 129.795 202.525 ;
        RECT 131.005 202.695 131.175 202.865 ;
        RECT 134.710 203.035 134.880 203.205 ;
        RECT 132.385 202.355 132.555 202.525 ;
        RECT 134.225 202.355 134.395 202.525 ;
        RECT 135.105 202.695 135.275 202.865 ;
        RECT 135.560 202.355 135.730 202.525 ;
        RECT 136.810 203.035 136.980 203.205 ;
        RECT 136.295 202.695 136.465 202.865 ;
        RECT 138.380 203.035 138.550 203.205 ;
        RECT 138.815 202.695 138.985 202.865 ;
        RECT 141.585 203.375 141.755 203.545 ;
        RECT 141.125 201.675 141.295 201.845 ;
        RECT 144.345 202.695 144.515 202.865 ;
        RECT 143.885 202.355 144.055 202.525 ;
        RECT 148.485 202.355 148.655 202.525 ;
        RECT 147.565 201.675 147.735 201.845 ;
        RECT 36.245 201.165 36.415 201.335 ;
        RECT 36.705 201.165 36.875 201.335 ;
        RECT 37.165 201.165 37.335 201.335 ;
        RECT 37.625 201.165 37.795 201.335 ;
        RECT 38.085 201.165 38.255 201.335 ;
        RECT 38.545 201.165 38.715 201.335 ;
        RECT 39.005 201.165 39.175 201.335 ;
        RECT 39.465 201.165 39.635 201.335 ;
        RECT 39.925 201.165 40.095 201.335 ;
        RECT 40.385 201.165 40.555 201.335 ;
        RECT 40.845 201.165 41.015 201.335 ;
        RECT 41.305 201.165 41.475 201.335 ;
        RECT 41.765 201.165 41.935 201.335 ;
        RECT 42.225 201.165 42.395 201.335 ;
        RECT 42.685 201.165 42.855 201.335 ;
        RECT 43.145 201.165 43.315 201.335 ;
        RECT 43.605 201.165 43.775 201.335 ;
        RECT 44.065 201.165 44.235 201.335 ;
        RECT 44.525 201.165 44.695 201.335 ;
        RECT 44.985 201.165 45.155 201.335 ;
        RECT 45.445 201.165 45.615 201.335 ;
        RECT 45.905 201.165 46.075 201.335 ;
        RECT 46.365 201.165 46.535 201.335 ;
        RECT 46.825 201.165 46.995 201.335 ;
        RECT 47.285 201.165 47.455 201.335 ;
        RECT 47.745 201.165 47.915 201.335 ;
        RECT 48.205 201.165 48.375 201.335 ;
        RECT 48.665 201.165 48.835 201.335 ;
        RECT 49.125 201.165 49.295 201.335 ;
        RECT 49.585 201.165 49.755 201.335 ;
        RECT 50.045 201.165 50.215 201.335 ;
        RECT 50.505 201.165 50.675 201.335 ;
        RECT 50.965 201.165 51.135 201.335 ;
        RECT 51.425 201.165 51.595 201.335 ;
        RECT 51.885 201.165 52.055 201.335 ;
        RECT 52.345 201.165 52.515 201.335 ;
        RECT 52.805 201.165 52.975 201.335 ;
        RECT 53.265 201.165 53.435 201.335 ;
        RECT 53.725 201.165 53.895 201.335 ;
        RECT 54.185 201.165 54.355 201.335 ;
        RECT 54.645 201.165 54.815 201.335 ;
        RECT 55.105 201.165 55.275 201.335 ;
        RECT 55.565 201.165 55.735 201.335 ;
        RECT 56.025 201.165 56.195 201.335 ;
        RECT 56.485 201.165 56.655 201.335 ;
        RECT 56.945 201.165 57.115 201.335 ;
        RECT 57.405 201.165 57.575 201.335 ;
        RECT 57.865 201.165 58.035 201.335 ;
        RECT 58.325 201.165 58.495 201.335 ;
        RECT 58.785 201.165 58.955 201.335 ;
        RECT 59.245 201.165 59.415 201.335 ;
        RECT 59.705 201.165 59.875 201.335 ;
        RECT 60.165 201.165 60.335 201.335 ;
        RECT 60.625 201.165 60.795 201.335 ;
        RECT 61.085 201.165 61.255 201.335 ;
        RECT 61.545 201.165 61.715 201.335 ;
        RECT 62.005 201.165 62.175 201.335 ;
        RECT 62.465 201.165 62.635 201.335 ;
        RECT 62.925 201.165 63.095 201.335 ;
        RECT 63.385 201.165 63.555 201.335 ;
        RECT 63.845 201.165 64.015 201.335 ;
        RECT 64.305 201.165 64.475 201.335 ;
        RECT 64.765 201.165 64.935 201.335 ;
        RECT 65.225 201.165 65.395 201.335 ;
        RECT 65.685 201.165 65.855 201.335 ;
        RECT 66.145 201.165 66.315 201.335 ;
        RECT 66.605 201.165 66.775 201.335 ;
        RECT 67.065 201.165 67.235 201.335 ;
        RECT 67.525 201.165 67.695 201.335 ;
        RECT 67.985 201.165 68.155 201.335 ;
        RECT 68.445 201.165 68.615 201.335 ;
        RECT 68.905 201.165 69.075 201.335 ;
        RECT 69.365 201.165 69.535 201.335 ;
        RECT 69.825 201.165 69.995 201.335 ;
        RECT 70.285 201.165 70.455 201.335 ;
        RECT 70.745 201.165 70.915 201.335 ;
        RECT 71.205 201.165 71.375 201.335 ;
        RECT 71.665 201.165 71.835 201.335 ;
        RECT 72.125 201.165 72.295 201.335 ;
        RECT 72.585 201.165 72.755 201.335 ;
        RECT 73.045 201.165 73.215 201.335 ;
        RECT 73.505 201.165 73.675 201.335 ;
        RECT 73.965 201.165 74.135 201.335 ;
        RECT 74.425 201.165 74.595 201.335 ;
        RECT 74.885 201.165 75.055 201.335 ;
        RECT 75.345 201.165 75.515 201.335 ;
        RECT 75.805 201.165 75.975 201.335 ;
        RECT 76.265 201.165 76.435 201.335 ;
        RECT 76.725 201.165 76.895 201.335 ;
        RECT 77.185 201.165 77.355 201.335 ;
        RECT 77.645 201.165 77.815 201.335 ;
        RECT 78.105 201.165 78.275 201.335 ;
        RECT 78.565 201.165 78.735 201.335 ;
        RECT 79.025 201.165 79.195 201.335 ;
        RECT 79.485 201.165 79.655 201.335 ;
        RECT 79.945 201.165 80.115 201.335 ;
        RECT 80.405 201.165 80.575 201.335 ;
        RECT 80.865 201.165 81.035 201.335 ;
        RECT 81.325 201.165 81.495 201.335 ;
        RECT 81.785 201.165 81.955 201.335 ;
        RECT 82.245 201.165 82.415 201.335 ;
        RECT 82.705 201.165 82.875 201.335 ;
        RECT 83.165 201.165 83.335 201.335 ;
        RECT 83.625 201.165 83.795 201.335 ;
        RECT 84.085 201.165 84.255 201.335 ;
        RECT 84.545 201.165 84.715 201.335 ;
        RECT 85.005 201.165 85.175 201.335 ;
        RECT 85.465 201.165 85.635 201.335 ;
        RECT 85.925 201.165 86.095 201.335 ;
        RECT 86.385 201.165 86.555 201.335 ;
        RECT 86.845 201.165 87.015 201.335 ;
        RECT 87.305 201.165 87.475 201.335 ;
        RECT 87.765 201.165 87.935 201.335 ;
        RECT 88.225 201.165 88.395 201.335 ;
        RECT 88.685 201.165 88.855 201.335 ;
        RECT 89.145 201.165 89.315 201.335 ;
        RECT 89.605 201.165 89.775 201.335 ;
        RECT 90.065 201.165 90.235 201.335 ;
        RECT 90.525 201.165 90.695 201.335 ;
        RECT 90.985 201.165 91.155 201.335 ;
        RECT 91.445 201.165 91.615 201.335 ;
        RECT 91.905 201.165 92.075 201.335 ;
        RECT 92.365 201.165 92.535 201.335 ;
        RECT 92.825 201.165 92.995 201.335 ;
        RECT 93.285 201.165 93.455 201.335 ;
        RECT 93.745 201.165 93.915 201.335 ;
        RECT 94.205 201.165 94.375 201.335 ;
        RECT 94.665 201.165 94.835 201.335 ;
        RECT 95.125 201.165 95.295 201.335 ;
        RECT 95.585 201.165 95.755 201.335 ;
        RECT 96.045 201.165 96.215 201.335 ;
        RECT 96.505 201.165 96.675 201.335 ;
        RECT 96.965 201.165 97.135 201.335 ;
        RECT 97.425 201.165 97.595 201.335 ;
        RECT 97.885 201.165 98.055 201.335 ;
        RECT 98.345 201.165 98.515 201.335 ;
        RECT 98.805 201.165 98.975 201.335 ;
        RECT 99.265 201.165 99.435 201.335 ;
        RECT 99.725 201.165 99.895 201.335 ;
        RECT 100.185 201.165 100.355 201.335 ;
        RECT 100.645 201.165 100.815 201.335 ;
        RECT 101.105 201.165 101.275 201.335 ;
        RECT 101.565 201.165 101.735 201.335 ;
        RECT 102.025 201.165 102.195 201.335 ;
        RECT 102.485 201.165 102.655 201.335 ;
        RECT 102.945 201.165 103.115 201.335 ;
        RECT 103.405 201.165 103.575 201.335 ;
        RECT 103.865 201.165 104.035 201.335 ;
        RECT 104.325 201.165 104.495 201.335 ;
        RECT 104.785 201.165 104.955 201.335 ;
        RECT 105.245 201.165 105.415 201.335 ;
        RECT 105.705 201.165 105.875 201.335 ;
        RECT 106.165 201.165 106.335 201.335 ;
        RECT 106.625 201.165 106.795 201.335 ;
        RECT 107.085 201.165 107.255 201.335 ;
        RECT 107.545 201.165 107.715 201.335 ;
        RECT 108.005 201.165 108.175 201.335 ;
        RECT 108.465 201.165 108.635 201.335 ;
        RECT 108.925 201.165 109.095 201.335 ;
        RECT 109.385 201.165 109.555 201.335 ;
        RECT 109.845 201.165 110.015 201.335 ;
        RECT 110.305 201.165 110.475 201.335 ;
        RECT 110.765 201.165 110.935 201.335 ;
        RECT 111.225 201.165 111.395 201.335 ;
        RECT 111.685 201.165 111.855 201.335 ;
        RECT 112.145 201.165 112.315 201.335 ;
        RECT 112.605 201.165 112.775 201.335 ;
        RECT 113.065 201.165 113.235 201.335 ;
        RECT 113.525 201.165 113.695 201.335 ;
        RECT 113.985 201.165 114.155 201.335 ;
        RECT 114.445 201.165 114.615 201.335 ;
        RECT 114.905 201.165 115.075 201.335 ;
        RECT 115.365 201.165 115.535 201.335 ;
        RECT 115.825 201.165 115.995 201.335 ;
        RECT 116.285 201.165 116.455 201.335 ;
        RECT 116.745 201.165 116.915 201.335 ;
        RECT 117.205 201.165 117.375 201.335 ;
        RECT 117.665 201.165 117.835 201.335 ;
        RECT 118.125 201.165 118.295 201.335 ;
        RECT 118.585 201.165 118.755 201.335 ;
        RECT 119.045 201.165 119.215 201.335 ;
        RECT 119.505 201.165 119.675 201.335 ;
        RECT 119.965 201.165 120.135 201.335 ;
        RECT 120.425 201.165 120.595 201.335 ;
        RECT 120.885 201.165 121.055 201.335 ;
        RECT 121.345 201.165 121.515 201.335 ;
        RECT 121.805 201.165 121.975 201.335 ;
        RECT 122.265 201.165 122.435 201.335 ;
        RECT 122.725 201.165 122.895 201.335 ;
        RECT 123.185 201.165 123.355 201.335 ;
        RECT 123.645 201.165 123.815 201.335 ;
        RECT 124.105 201.165 124.275 201.335 ;
        RECT 124.565 201.165 124.735 201.335 ;
        RECT 125.025 201.165 125.195 201.335 ;
        RECT 125.485 201.165 125.655 201.335 ;
        RECT 125.945 201.165 126.115 201.335 ;
        RECT 126.405 201.165 126.575 201.335 ;
        RECT 126.865 201.165 127.035 201.335 ;
        RECT 127.325 201.165 127.495 201.335 ;
        RECT 127.785 201.165 127.955 201.335 ;
        RECT 128.245 201.165 128.415 201.335 ;
        RECT 128.705 201.165 128.875 201.335 ;
        RECT 129.165 201.165 129.335 201.335 ;
        RECT 129.625 201.165 129.795 201.335 ;
        RECT 130.085 201.165 130.255 201.335 ;
        RECT 130.545 201.165 130.715 201.335 ;
        RECT 131.005 201.165 131.175 201.335 ;
        RECT 131.465 201.165 131.635 201.335 ;
        RECT 131.925 201.165 132.095 201.335 ;
        RECT 132.385 201.165 132.555 201.335 ;
        RECT 132.845 201.165 133.015 201.335 ;
        RECT 133.305 201.165 133.475 201.335 ;
        RECT 133.765 201.165 133.935 201.335 ;
        RECT 134.225 201.165 134.395 201.335 ;
        RECT 134.685 201.165 134.855 201.335 ;
        RECT 135.145 201.165 135.315 201.335 ;
        RECT 135.605 201.165 135.775 201.335 ;
        RECT 136.065 201.165 136.235 201.335 ;
        RECT 136.525 201.165 136.695 201.335 ;
        RECT 136.985 201.165 137.155 201.335 ;
        RECT 137.445 201.165 137.615 201.335 ;
        RECT 137.905 201.165 138.075 201.335 ;
        RECT 138.365 201.165 138.535 201.335 ;
        RECT 138.825 201.165 138.995 201.335 ;
        RECT 139.285 201.165 139.455 201.335 ;
        RECT 139.745 201.165 139.915 201.335 ;
        RECT 140.205 201.165 140.375 201.335 ;
        RECT 140.665 201.165 140.835 201.335 ;
        RECT 141.125 201.165 141.295 201.335 ;
        RECT 141.585 201.165 141.755 201.335 ;
        RECT 142.045 201.165 142.215 201.335 ;
        RECT 142.505 201.165 142.675 201.335 ;
        RECT 142.965 201.165 143.135 201.335 ;
        RECT 143.425 201.165 143.595 201.335 ;
        RECT 143.885 201.165 144.055 201.335 ;
        RECT 144.345 201.165 144.515 201.335 ;
        RECT 144.805 201.165 144.975 201.335 ;
        RECT 145.265 201.165 145.435 201.335 ;
        RECT 145.725 201.165 145.895 201.335 ;
        RECT 146.185 201.165 146.355 201.335 ;
        RECT 146.645 201.165 146.815 201.335 ;
        RECT 147.105 201.165 147.275 201.335 ;
        RECT 147.565 201.165 147.735 201.335 ;
        RECT 148.025 201.165 148.195 201.335 ;
        RECT 148.485 201.165 148.655 201.335 ;
        RECT 148.945 201.165 149.115 201.335 ;
        RECT 149.405 201.165 149.575 201.335 ;
        RECT 149.865 201.165 150.035 201.335 ;
        RECT 41.765 199.975 41.935 200.145 ;
        RECT 42.685 200.315 42.855 200.485 ;
        RECT 43.605 200.655 43.775 200.825 ;
        RECT 43.145 199.975 43.315 200.145 ;
        RECT 42.225 199.295 42.395 199.465 ;
        RECT 44.525 199.635 44.695 199.805 ;
        RECT 44.985 199.975 45.155 200.145 ;
        RECT 45.445 199.635 45.615 199.805 ;
        RECT 45.905 199.975 46.075 200.145 ;
        RECT 47.285 200.315 47.455 200.485 ;
        RECT 48.665 199.635 48.835 199.805 ;
        RECT 50.045 199.975 50.215 200.145 ;
        RECT 47.745 198.955 47.915 199.125 ;
        RECT 55.565 199.975 55.735 200.145 ;
        RECT 57.405 199.975 57.575 200.145 ;
        RECT 56.485 198.955 56.655 199.125 ;
        RECT 59.245 199.975 59.415 200.145 ;
        RECT 58.325 198.955 58.495 199.125 ;
        RECT 59.705 199.295 59.875 199.465 ;
        RECT 60.625 199.975 60.795 200.145 ;
        RECT 60.165 199.295 60.335 199.465 ;
        RECT 61.545 198.955 61.715 199.125 ;
        RECT 62.465 199.635 62.635 199.805 ;
        RECT 63.845 199.635 64.015 199.805 ;
        RECT 70.745 200.655 70.915 200.825 ;
        RECT 71.665 199.975 71.835 200.145 ;
        RECT 72.125 199.635 72.295 199.805 ;
        RECT 72.610 199.295 72.780 199.465 ;
        RECT 73.005 199.635 73.175 199.805 ;
        RECT 73.460 199.975 73.630 200.145 ;
        RECT 74.195 199.635 74.365 199.805 ;
        RECT 74.710 199.295 74.880 199.465 ;
        RECT 76.280 199.295 76.450 199.465 ;
        RECT 76.715 199.635 76.885 199.805 ;
        RECT 79.025 198.955 79.195 199.125 ;
        RECT 80.865 199.635 81.035 199.805 ;
        RECT 81.785 199.975 81.955 200.145 ;
        RECT 86.385 199.975 86.555 200.145 ;
        RECT 87.305 199.975 87.475 200.145 ;
        RECT 88.185 199.975 88.355 200.145 ;
        RECT 82.705 199.295 82.875 199.465 ;
        RECT 86.845 198.955 87.015 199.125 ;
        RECT 89.145 199.295 89.315 199.465 ;
        RECT 90.525 199.975 90.695 200.145 ;
        RECT 94.205 200.655 94.375 200.825 ;
        RECT 90.065 198.955 90.235 199.125 ;
        RECT 95.125 199.975 95.295 200.145 ;
        RECT 95.585 199.975 95.755 200.145 ;
        RECT 96.045 199.975 96.215 200.145 ;
        RECT 96.505 199.635 96.675 199.805 ;
        RECT 98.345 199.975 98.515 200.145 ;
        RECT 97.885 199.635 98.055 199.805 ;
        RECT 100.645 199.975 100.815 200.145 ;
        RECT 101.565 199.975 101.735 200.145 ;
        RECT 102.025 199.975 102.195 200.145 ;
        RECT 102.605 199.975 102.775 200.145 ;
        RECT 100.185 199.635 100.355 199.805 ;
        RECT 112.145 199.975 112.315 200.145 ;
        RECT 113.065 198.955 113.235 199.125 ;
        RECT 113.985 198.955 114.155 199.125 ;
        RECT 116.295 199.635 116.465 199.805 ;
        RECT 116.730 199.295 116.900 199.465 ;
        RECT 118.815 199.635 118.985 199.805 ;
        RECT 118.300 199.295 118.470 199.465 ;
        RECT 119.550 200.315 119.720 200.485 ;
        RECT 120.005 199.635 120.175 199.805 ;
        RECT 120.885 199.975 121.055 200.145 ;
        RECT 125.485 199.975 125.655 200.145 ;
        RECT 126.405 199.975 126.575 200.145 ;
        RECT 120.400 199.295 120.570 199.465 ;
        RECT 125.945 198.955 126.115 199.125 ;
        RECT 126.865 198.955 127.035 199.125 ;
        RECT 129.175 199.635 129.345 199.805 ;
        RECT 129.610 199.295 129.780 199.465 ;
        RECT 131.695 199.635 131.865 199.805 ;
        RECT 131.180 199.295 131.350 199.465 ;
        RECT 132.430 199.975 132.600 200.145 ;
        RECT 132.885 199.635 133.055 199.805 ;
        RECT 133.765 199.975 133.935 200.145 ;
        RECT 133.280 199.295 133.450 199.465 ;
        RECT 36.245 198.445 36.415 198.615 ;
        RECT 36.705 198.445 36.875 198.615 ;
        RECT 37.165 198.445 37.335 198.615 ;
        RECT 37.625 198.445 37.795 198.615 ;
        RECT 38.085 198.445 38.255 198.615 ;
        RECT 38.545 198.445 38.715 198.615 ;
        RECT 39.005 198.445 39.175 198.615 ;
        RECT 39.465 198.445 39.635 198.615 ;
        RECT 39.925 198.445 40.095 198.615 ;
        RECT 40.385 198.445 40.555 198.615 ;
        RECT 40.845 198.445 41.015 198.615 ;
        RECT 41.305 198.445 41.475 198.615 ;
        RECT 41.765 198.445 41.935 198.615 ;
        RECT 42.225 198.445 42.395 198.615 ;
        RECT 42.685 198.445 42.855 198.615 ;
        RECT 43.145 198.445 43.315 198.615 ;
        RECT 43.605 198.445 43.775 198.615 ;
        RECT 44.065 198.445 44.235 198.615 ;
        RECT 44.525 198.445 44.695 198.615 ;
        RECT 44.985 198.445 45.155 198.615 ;
        RECT 45.445 198.445 45.615 198.615 ;
        RECT 45.905 198.445 46.075 198.615 ;
        RECT 46.365 198.445 46.535 198.615 ;
        RECT 46.825 198.445 46.995 198.615 ;
        RECT 47.285 198.445 47.455 198.615 ;
        RECT 47.745 198.445 47.915 198.615 ;
        RECT 48.205 198.445 48.375 198.615 ;
        RECT 48.665 198.445 48.835 198.615 ;
        RECT 49.125 198.445 49.295 198.615 ;
        RECT 49.585 198.445 49.755 198.615 ;
        RECT 50.045 198.445 50.215 198.615 ;
        RECT 50.505 198.445 50.675 198.615 ;
        RECT 50.965 198.445 51.135 198.615 ;
        RECT 51.425 198.445 51.595 198.615 ;
        RECT 51.885 198.445 52.055 198.615 ;
        RECT 52.345 198.445 52.515 198.615 ;
        RECT 52.805 198.445 52.975 198.615 ;
        RECT 53.265 198.445 53.435 198.615 ;
        RECT 53.725 198.445 53.895 198.615 ;
        RECT 54.185 198.445 54.355 198.615 ;
        RECT 54.645 198.445 54.815 198.615 ;
        RECT 55.105 198.445 55.275 198.615 ;
        RECT 55.565 198.445 55.735 198.615 ;
        RECT 56.025 198.445 56.195 198.615 ;
        RECT 56.485 198.445 56.655 198.615 ;
        RECT 56.945 198.445 57.115 198.615 ;
        RECT 57.405 198.445 57.575 198.615 ;
        RECT 57.865 198.445 58.035 198.615 ;
        RECT 58.325 198.445 58.495 198.615 ;
        RECT 58.785 198.445 58.955 198.615 ;
        RECT 59.245 198.445 59.415 198.615 ;
        RECT 59.705 198.445 59.875 198.615 ;
        RECT 60.165 198.445 60.335 198.615 ;
        RECT 60.625 198.445 60.795 198.615 ;
        RECT 61.085 198.445 61.255 198.615 ;
        RECT 61.545 198.445 61.715 198.615 ;
        RECT 62.005 198.445 62.175 198.615 ;
        RECT 62.465 198.445 62.635 198.615 ;
        RECT 62.925 198.445 63.095 198.615 ;
        RECT 63.385 198.445 63.555 198.615 ;
        RECT 63.845 198.445 64.015 198.615 ;
        RECT 64.305 198.445 64.475 198.615 ;
        RECT 64.765 198.445 64.935 198.615 ;
        RECT 65.225 198.445 65.395 198.615 ;
        RECT 65.685 198.445 65.855 198.615 ;
        RECT 66.145 198.445 66.315 198.615 ;
        RECT 66.605 198.445 66.775 198.615 ;
        RECT 67.065 198.445 67.235 198.615 ;
        RECT 67.525 198.445 67.695 198.615 ;
        RECT 67.985 198.445 68.155 198.615 ;
        RECT 68.445 198.445 68.615 198.615 ;
        RECT 68.905 198.445 69.075 198.615 ;
        RECT 69.365 198.445 69.535 198.615 ;
        RECT 69.825 198.445 69.995 198.615 ;
        RECT 70.285 198.445 70.455 198.615 ;
        RECT 70.745 198.445 70.915 198.615 ;
        RECT 71.205 198.445 71.375 198.615 ;
        RECT 71.665 198.445 71.835 198.615 ;
        RECT 72.125 198.445 72.295 198.615 ;
        RECT 72.585 198.445 72.755 198.615 ;
        RECT 73.045 198.445 73.215 198.615 ;
        RECT 73.505 198.445 73.675 198.615 ;
        RECT 73.965 198.445 74.135 198.615 ;
        RECT 74.425 198.445 74.595 198.615 ;
        RECT 74.885 198.445 75.055 198.615 ;
        RECT 75.345 198.445 75.515 198.615 ;
        RECT 75.805 198.445 75.975 198.615 ;
        RECT 76.265 198.445 76.435 198.615 ;
        RECT 76.725 198.445 76.895 198.615 ;
        RECT 77.185 198.445 77.355 198.615 ;
        RECT 77.645 198.445 77.815 198.615 ;
        RECT 78.105 198.445 78.275 198.615 ;
        RECT 78.565 198.445 78.735 198.615 ;
        RECT 79.025 198.445 79.195 198.615 ;
        RECT 79.485 198.445 79.655 198.615 ;
        RECT 79.945 198.445 80.115 198.615 ;
        RECT 80.405 198.445 80.575 198.615 ;
        RECT 80.865 198.445 81.035 198.615 ;
        RECT 81.325 198.445 81.495 198.615 ;
        RECT 81.785 198.445 81.955 198.615 ;
        RECT 82.245 198.445 82.415 198.615 ;
        RECT 82.705 198.445 82.875 198.615 ;
        RECT 83.165 198.445 83.335 198.615 ;
        RECT 83.625 198.445 83.795 198.615 ;
        RECT 84.085 198.445 84.255 198.615 ;
        RECT 84.545 198.445 84.715 198.615 ;
        RECT 85.005 198.445 85.175 198.615 ;
        RECT 85.465 198.445 85.635 198.615 ;
        RECT 85.925 198.445 86.095 198.615 ;
        RECT 86.385 198.445 86.555 198.615 ;
        RECT 86.845 198.445 87.015 198.615 ;
        RECT 87.305 198.445 87.475 198.615 ;
        RECT 87.765 198.445 87.935 198.615 ;
        RECT 88.225 198.445 88.395 198.615 ;
        RECT 88.685 198.445 88.855 198.615 ;
        RECT 89.145 198.445 89.315 198.615 ;
        RECT 89.605 198.445 89.775 198.615 ;
        RECT 90.065 198.445 90.235 198.615 ;
        RECT 90.525 198.445 90.695 198.615 ;
        RECT 90.985 198.445 91.155 198.615 ;
        RECT 91.445 198.445 91.615 198.615 ;
        RECT 91.905 198.445 92.075 198.615 ;
        RECT 92.365 198.445 92.535 198.615 ;
        RECT 92.825 198.445 92.995 198.615 ;
        RECT 93.285 198.445 93.455 198.615 ;
        RECT 93.745 198.445 93.915 198.615 ;
        RECT 94.205 198.445 94.375 198.615 ;
        RECT 94.665 198.445 94.835 198.615 ;
        RECT 95.125 198.445 95.295 198.615 ;
        RECT 95.585 198.445 95.755 198.615 ;
        RECT 96.045 198.445 96.215 198.615 ;
        RECT 96.505 198.445 96.675 198.615 ;
        RECT 96.965 198.445 97.135 198.615 ;
        RECT 97.425 198.445 97.595 198.615 ;
        RECT 97.885 198.445 98.055 198.615 ;
        RECT 98.345 198.445 98.515 198.615 ;
        RECT 98.805 198.445 98.975 198.615 ;
        RECT 99.265 198.445 99.435 198.615 ;
        RECT 99.725 198.445 99.895 198.615 ;
        RECT 100.185 198.445 100.355 198.615 ;
        RECT 100.645 198.445 100.815 198.615 ;
        RECT 101.105 198.445 101.275 198.615 ;
        RECT 101.565 198.445 101.735 198.615 ;
        RECT 102.025 198.445 102.195 198.615 ;
        RECT 102.485 198.445 102.655 198.615 ;
        RECT 102.945 198.445 103.115 198.615 ;
        RECT 103.405 198.445 103.575 198.615 ;
        RECT 103.865 198.445 104.035 198.615 ;
        RECT 104.325 198.445 104.495 198.615 ;
        RECT 104.785 198.445 104.955 198.615 ;
        RECT 105.245 198.445 105.415 198.615 ;
        RECT 105.705 198.445 105.875 198.615 ;
        RECT 106.165 198.445 106.335 198.615 ;
        RECT 106.625 198.445 106.795 198.615 ;
        RECT 107.085 198.445 107.255 198.615 ;
        RECT 107.545 198.445 107.715 198.615 ;
        RECT 108.005 198.445 108.175 198.615 ;
        RECT 108.465 198.445 108.635 198.615 ;
        RECT 108.925 198.445 109.095 198.615 ;
        RECT 109.385 198.445 109.555 198.615 ;
        RECT 109.845 198.445 110.015 198.615 ;
        RECT 110.305 198.445 110.475 198.615 ;
        RECT 110.765 198.445 110.935 198.615 ;
        RECT 111.225 198.445 111.395 198.615 ;
        RECT 111.685 198.445 111.855 198.615 ;
        RECT 112.145 198.445 112.315 198.615 ;
        RECT 112.605 198.445 112.775 198.615 ;
        RECT 113.065 198.445 113.235 198.615 ;
        RECT 113.525 198.445 113.695 198.615 ;
        RECT 113.985 198.445 114.155 198.615 ;
        RECT 114.445 198.445 114.615 198.615 ;
        RECT 114.905 198.445 115.075 198.615 ;
        RECT 115.365 198.445 115.535 198.615 ;
        RECT 115.825 198.445 115.995 198.615 ;
        RECT 116.285 198.445 116.455 198.615 ;
        RECT 116.745 198.445 116.915 198.615 ;
        RECT 117.205 198.445 117.375 198.615 ;
        RECT 117.665 198.445 117.835 198.615 ;
        RECT 118.125 198.445 118.295 198.615 ;
        RECT 118.585 198.445 118.755 198.615 ;
        RECT 119.045 198.445 119.215 198.615 ;
        RECT 119.505 198.445 119.675 198.615 ;
        RECT 119.965 198.445 120.135 198.615 ;
        RECT 120.425 198.445 120.595 198.615 ;
        RECT 120.885 198.445 121.055 198.615 ;
        RECT 121.345 198.445 121.515 198.615 ;
        RECT 121.805 198.445 121.975 198.615 ;
        RECT 122.265 198.445 122.435 198.615 ;
        RECT 122.725 198.445 122.895 198.615 ;
        RECT 123.185 198.445 123.355 198.615 ;
        RECT 123.645 198.445 123.815 198.615 ;
        RECT 124.105 198.445 124.275 198.615 ;
        RECT 124.565 198.445 124.735 198.615 ;
        RECT 125.025 198.445 125.195 198.615 ;
        RECT 125.485 198.445 125.655 198.615 ;
        RECT 125.945 198.445 126.115 198.615 ;
        RECT 126.405 198.445 126.575 198.615 ;
        RECT 126.865 198.445 127.035 198.615 ;
        RECT 127.325 198.445 127.495 198.615 ;
        RECT 127.785 198.445 127.955 198.615 ;
        RECT 128.245 198.445 128.415 198.615 ;
        RECT 128.705 198.445 128.875 198.615 ;
        RECT 129.165 198.445 129.335 198.615 ;
        RECT 129.625 198.445 129.795 198.615 ;
        RECT 130.085 198.445 130.255 198.615 ;
        RECT 130.545 198.445 130.715 198.615 ;
        RECT 131.005 198.445 131.175 198.615 ;
        RECT 131.465 198.445 131.635 198.615 ;
        RECT 131.925 198.445 132.095 198.615 ;
        RECT 132.385 198.445 132.555 198.615 ;
        RECT 132.845 198.445 133.015 198.615 ;
        RECT 133.305 198.445 133.475 198.615 ;
        RECT 133.765 198.445 133.935 198.615 ;
        RECT 134.225 198.445 134.395 198.615 ;
        RECT 134.685 198.445 134.855 198.615 ;
        RECT 135.145 198.445 135.315 198.615 ;
        RECT 135.605 198.445 135.775 198.615 ;
        RECT 136.065 198.445 136.235 198.615 ;
        RECT 136.525 198.445 136.695 198.615 ;
        RECT 136.985 198.445 137.155 198.615 ;
        RECT 137.445 198.445 137.615 198.615 ;
        RECT 137.905 198.445 138.075 198.615 ;
        RECT 138.365 198.445 138.535 198.615 ;
        RECT 138.825 198.445 138.995 198.615 ;
        RECT 139.285 198.445 139.455 198.615 ;
        RECT 139.745 198.445 139.915 198.615 ;
        RECT 140.205 198.445 140.375 198.615 ;
        RECT 140.665 198.445 140.835 198.615 ;
        RECT 141.125 198.445 141.295 198.615 ;
        RECT 141.585 198.445 141.755 198.615 ;
        RECT 142.045 198.445 142.215 198.615 ;
        RECT 142.505 198.445 142.675 198.615 ;
        RECT 142.965 198.445 143.135 198.615 ;
        RECT 143.425 198.445 143.595 198.615 ;
        RECT 143.885 198.445 144.055 198.615 ;
        RECT 144.345 198.445 144.515 198.615 ;
        RECT 144.805 198.445 144.975 198.615 ;
        RECT 145.265 198.445 145.435 198.615 ;
        RECT 145.725 198.445 145.895 198.615 ;
        RECT 146.185 198.445 146.355 198.615 ;
        RECT 146.645 198.445 146.815 198.615 ;
        RECT 147.105 198.445 147.275 198.615 ;
        RECT 147.565 198.445 147.735 198.615 ;
        RECT 148.025 198.445 148.195 198.615 ;
        RECT 148.485 198.445 148.655 198.615 ;
        RECT 148.945 198.445 149.115 198.615 ;
        RECT 149.405 198.445 149.575 198.615 ;
        RECT 149.865 198.445 150.035 198.615 ;
        RECT 41.305 196.915 41.475 197.085 ;
        RECT 42.225 196.915 42.395 197.085 ;
        RECT 41.765 196.235 41.935 196.405 ;
        RECT 44.065 197.935 44.235 198.105 ;
        RECT 44.985 196.915 45.155 197.085 ;
        RECT 45.905 196.915 46.075 197.085 ;
        RECT 49.585 196.915 49.755 197.085 ;
        RECT 50.965 196.915 51.135 197.085 ;
        RECT 56.025 197.595 56.195 197.765 ;
        RECT 55.105 196.915 55.275 197.085 ;
        RECT 56.485 197.935 56.655 198.105 ;
        RECT 57.405 196.915 57.575 197.085 ;
        RECT 59.705 197.935 59.875 198.105 ;
        RECT 58.785 196.915 58.955 197.085 ;
        RECT 60.625 196.915 60.795 197.085 ;
        RECT 61.085 197.255 61.255 197.425 ;
        RECT 61.545 196.915 61.715 197.085 ;
        RECT 62.005 197.255 62.175 197.425 ;
        RECT 57.865 196.235 58.035 196.405 ;
        RECT 64.305 196.915 64.475 197.085 ;
        RECT 63.845 196.235 64.015 196.405 ;
        RECT 66.605 196.575 66.775 196.745 ;
        RECT 67.065 196.235 67.235 196.405 ;
        RECT 85.925 196.915 86.095 197.085 ;
        RECT 85.005 196.575 85.175 196.745 ;
        RECT 89.605 197.935 89.775 198.105 ;
        RECT 87.305 196.915 87.475 197.085 ;
        RECT 87.765 197.255 87.935 197.425 ;
        RECT 88.225 197.255 88.395 197.425 ;
        RECT 88.685 196.915 88.855 197.085 ;
        RECT 90.525 197.255 90.695 197.425 ;
        RECT 90.985 196.915 91.155 197.085 ;
        RECT 91.445 197.255 91.615 197.425 ;
        RECT 91.905 196.915 92.075 197.085 ;
        RECT 86.385 196.235 86.555 196.405 ;
        RECT 101.105 197.935 101.275 198.105 ;
        RECT 105.705 197.935 105.875 198.105 ;
        RECT 104.785 197.595 104.955 197.765 ;
        RECT 102.025 196.915 102.195 197.085 ;
        RECT 102.485 196.915 102.655 197.085 ;
        RECT 103.865 196.915 104.035 197.085 ;
        RECT 104.325 196.915 104.495 197.085 ;
        RECT 102.945 196.575 103.115 196.745 ;
        RECT 105.625 196.235 105.795 196.405 ;
        RECT 108.005 196.915 108.175 197.085 ;
        RECT 106.625 196.575 106.795 196.745 ;
        RECT 109.845 197.255 110.015 197.425 ;
        RECT 108.925 196.915 109.095 197.085 ;
        RECT 108.465 196.235 108.635 196.405 ;
        RECT 110.305 196.915 110.475 197.085 ;
        RECT 113.065 196.915 113.235 197.085 ;
        RECT 113.985 196.235 114.155 196.405 ;
        RECT 114.445 197.935 114.615 198.105 ;
        RECT 117.665 197.255 117.835 197.425 ;
        RECT 120.425 197.935 120.595 198.105 ;
        RECT 116.745 196.235 116.915 196.405 ;
        RECT 119.965 196.575 120.135 196.745 ;
        RECT 125.025 197.935 125.195 198.105 ;
        RECT 124.105 196.915 124.275 197.085 ;
        RECT 126.865 197.935 127.035 198.105 ;
        RECT 128.245 196.915 128.415 197.085 ;
        RECT 128.705 196.915 128.875 197.085 ;
        RECT 129.165 196.915 129.335 197.085 ;
        RECT 130.085 196.915 130.255 197.085 ;
        RECT 139.770 197.595 139.940 197.765 ;
        RECT 137.445 196.915 137.615 197.085 ;
        RECT 139.285 197.255 139.455 197.425 ;
        RECT 138.365 196.235 138.535 196.405 ;
        RECT 140.165 197.255 140.335 197.425 ;
        RECT 140.510 196.575 140.680 196.745 ;
        RECT 141.870 197.595 142.040 197.765 ;
        RECT 141.355 197.255 141.525 197.425 ;
        RECT 143.440 197.595 143.610 197.765 ;
        RECT 143.875 197.255 144.045 197.425 ;
        RECT 146.185 196.235 146.355 196.405 ;
        RECT 36.245 195.725 36.415 195.895 ;
        RECT 36.705 195.725 36.875 195.895 ;
        RECT 37.165 195.725 37.335 195.895 ;
        RECT 37.625 195.725 37.795 195.895 ;
        RECT 38.085 195.725 38.255 195.895 ;
        RECT 38.545 195.725 38.715 195.895 ;
        RECT 39.005 195.725 39.175 195.895 ;
        RECT 39.465 195.725 39.635 195.895 ;
        RECT 39.925 195.725 40.095 195.895 ;
        RECT 40.385 195.725 40.555 195.895 ;
        RECT 40.845 195.725 41.015 195.895 ;
        RECT 41.305 195.725 41.475 195.895 ;
        RECT 41.765 195.725 41.935 195.895 ;
        RECT 42.225 195.725 42.395 195.895 ;
        RECT 42.685 195.725 42.855 195.895 ;
        RECT 43.145 195.725 43.315 195.895 ;
        RECT 43.605 195.725 43.775 195.895 ;
        RECT 44.065 195.725 44.235 195.895 ;
        RECT 44.525 195.725 44.695 195.895 ;
        RECT 44.985 195.725 45.155 195.895 ;
        RECT 45.445 195.725 45.615 195.895 ;
        RECT 45.905 195.725 46.075 195.895 ;
        RECT 46.365 195.725 46.535 195.895 ;
        RECT 46.825 195.725 46.995 195.895 ;
        RECT 47.285 195.725 47.455 195.895 ;
        RECT 47.745 195.725 47.915 195.895 ;
        RECT 48.205 195.725 48.375 195.895 ;
        RECT 48.665 195.725 48.835 195.895 ;
        RECT 49.125 195.725 49.295 195.895 ;
        RECT 49.585 195.725 49.755 195.895 ;
        RECT 50.045 195.725 50.215 195.895 ;
        RECT 50.505 195.725 50.675 195.895 ;
        RECT 50.965 195.725 51.135 195.895 ;
        RECT 51.425 195.725 51.595 195.895 ;
        RECT 51.885 195.725 52.055 195.895 ;
        RECT 52.345 195.725 52.515 195.895 ;
        RECT 52.805 195.725 52.975 195.895 ;
        RECT 53.265 195.725 53.435 195.895 ;
        RECT 53.725 195.725 53.895 195.895 ;
        RECT 54.185 195.725 54.355 195.895 ;
        RECT 54.645 195.725 54.815 195.895 ;
        RECT 55.105 195.725 55.275 195.895 ;
        RECT 55.565 195.725 55.735 195.895 ;
        RECT 56.025 195.725 56.195 195.895 ;
        RECT 56.485 195.725 56.655 195.895 ;
        RECT 56.945 195.725 57.115 195.895 ;
        RECT 57.405 195.725 57.575 195.895 ;
        RECT 57.865 195.725 58.035 195.895 ;
        RECT 58.325 195.725 58.495 195.895 ;
        RECT 58.785 195.725 58.955 195.895 ;
        RECT 59.245 195.725 59.415 195.895 ;
        RECT 59.705 195.725 59.875 195.895 ;
        RECT 60.165 195.725 60.335 195.895 ;
        RECT 60.625 195.725 60.795 195.895 ;
        RECT 61.085 195.725 61.255 195.895 ;
        RECT 61.545 195.725 61.715 195.895 ;
        RECT 62.005 195.725 62.175 195.895 ;
        RECT 62.465 195.725 62.635 195.895 ;
        RECT 62.925 195.725 63.095 195.895 ;
        RECT 63.385 195.725 63.555 195.895 ;
        RECT 63.845 195.725 64.015 195.895 ;
        RECT 64.305 195.725 64.475 195.895 ;
        RECT 64.765 195.725 64.935 195.895 ;
        RECT 65.225 195.725 65.395 195.895 ;
        RECT 65.685 195.725 65.855 195.895 ;
        RECT 66.145 195.725 66.315 195.895 ;
        RECT 66.605 195.725 66.775 195.895 ;
        RECT 67.065 195.725 67.235 195.895 ;
        RECT 67.525 195.725 67.695 195.895 ;
        RECT 67.985 195.725 68.155 195.895 ;
        RECT 68.445 195.725 68.615 195.895 ;
        RECT 68.905 195.725 69.075 195.895 ;
        RECT 69.365 195.725 69.535 195.895 ;
        RECT 69.825 195.725 69.995 195.895 ;
        RECT 70.285 195.725 70.455 195.895 ;
        RECT 70.745 195.725 70.915 195.895 ;
        RECT 71.205 195.725 71.375 195.895 ;
        RECT 71.665 195.725 71.835 195.895 ;
        RECT 72.125 195.725 72.295 195.895 ;
        RECT 72.585 195.725 72.755 195.895 ;
        RECT 73.045 195.725 73.215 195.895 ;
        RECT 73.505 195.725 73.675 195.895 ;
        RECT 73.965 195.725 74.135 195.895 ;
        RECT 74.425 195.725 74.595 195.895 ;
        RECT 74.885 195.725 75.055 195.895 ;
        RECT 75.345 195.725 75.515 195.895 ;
        RECT 75.805 195.725 75.975 195.895 ;
        RECT 76.265 195.725 76.435 195.895 ;
        RECT 76.725 195.725 76.895 195.895 ;
        RECT 77.185 195.725 77.355 195.895 ;
        RECT 77.645 195.725 77.815 195.895 ;
        RECT 78.105 195.725 78.275 195.895 ;
        RECT 78.565 195.725 78.735 195.895 ;
        RECT 79.025 195.725 79.195 195.895 ;
        RECT 79.485 195.725 79.655 195.895 ;
        RECT 79.945 195.725 80.115 195.895 ;
        RECT 80.405 195.725 80.575 195.895 ;
        RECT 80.865 195.725 81.035 195.895 ;
        RECT 81.325 195.725 81.495 195.895 ;
        RECT 81.785 195.725 81.955 195.895 ;
        RECT 82.245 195.725 82.415 195.895 ;
        RECT 82.705 195.725 82.875 195.895 ;
        RECT 83.165 195.725 83.335 195.895 ;
        RECT 83.625 195.725 83.795 195.895 ;
        RECT 84.085 195.725 84.255 195.895 ;
        RECT 84.545 195.725 84.715 195.895 ;
        RECT 85.005 195.725 85.175 195.895 ;
        RECT 85.465 195.725 85.635 195.895 ;
        RECT 85.925 195.725 86.095 195.895 ;
        RECT 86.385 195.725 86.555 195.895 ;
        RECT 86.845 195.725 87.015 195.895 ;
        RECT 87.305 195.725 87.475 195.895 ;
        RECT 87.765 195.725 87.935 195.895 ;
        RECT 88.225 195.725 88.395 195.895 ;
        RECT 88.685 195.725 88.855 195.895 ;
        RECT 89.145 195.725 89.315 195.895 ;
        RECT 89.605 195.725 89.775 195.895 ;
        RECT 90.065 195.725 90.235 195.895 ;
        RECT 90.525 195.725 90.695 195.895 ;
        RECT 90.985 195.725 91.155 195.895 ;
        RECT 91.445 195.725 91.615 195.895 ;
        RECT 91.905 195.725 92.075 195.895 ;
        RECT 92.365 195.725 92.535 195.895 ;
        RECT 92.825 195.725 92.995 195.895 ;
        RECT 93.285 195.725 93.455 195.895 ;
        RECT 93.745 195.725 93.915 195.895 ;
        RECT 94.205 195.725 94.375 195.895 ;
        RECT 94.665 195.725 94.835 195.895 ;
        RECT 95.125 195.725 95.295 195.895 ;
        RECT 95.585 195.725 95.755 195.895 ;
        RECT 96.045 195.725 96.215 195.895 ;
        RECT 96.505 195.725 96.675 195.895 ;
        RECT 96.965 195.725 97.135 195.895 ;
        RECT 97.425 195.725 97.595 195.895 ;
        RECT 97.885 195.725 98.055 195.895 ;
        RECT 98.345 195.725 98.515 195.895 ;
        RECT 98.805 195.725 98.975 195.895 ;
        RECT 99.265 195.725 99.435 195.895 ;
        RECT 99.725 195.725 99.895 195.895 ;
        RECT 100.185 195.725 100.355 195.895 ;
        RECT 100.645 195.725 100.815 195.895 ;
        RECT 101.105 195.725 101.275 195.895 ;
        RECT 101.565 195.725 101.735 195.895 ;
        RECT 102.025 195.725 102.195 195.895 ;
        RECT 102.485 195.725 102.655 195.895 ;
        RECT 102.945 195.725 103.115 195.895 ;
        RECT 103.405 195.725 103.575 195.895 ;
        RECT 103.865 195.725 104.035 195.895 ;
        RECT 104.325 195.725 104.495 195.895 ;
        RECT 104.785 195.725 104.955 195.895 ;
        RECT 105.245 195.725 105.415 195.895 ;
        RECT 105.705 195.725 105.875 195.895 ;
        RECT 106.165 195.725 106.335 195.895 ;
        RECT 106.625 195.725 106.795 195.895 ;
        RECT 107.085 195.725 107.255 195.895 ;
        RECT 107.545 195.725 107.715 195.895 ;
        RECT 108.005 195.725 108.175 195.895 ;
        RECT 108.465 195.725 108.635 195.895 ;
        RECT 108.925 195.725 109.095 195.895 ;
        RECT 109.385 195.725 109.555 195.895 ;
        RECT 109.845 195.725 110.015 195.895 ;
        RECT 110.305 195.725 110.475 195.895 ;
        RECT 110.765 195.725 110.935 195.895 ;
        RECT 111.225 195.725 111.395 195.895 ;
        RECT 111.685 195.725 111.855 195.895 ;
        RECT 112.145 195.725 112.315 195.895 ;
        RECT 112.605 195.725 112.775 195.895 ;
        RECT 113.065 195.725 113.235 195.895 ;
        RECT 113.525 195.725 113.695 195.895 ;
        RECT 113.985 195.725 114.155 195.895 ;
        RECT 114.445 195.725 114.615 195.895 ;
        RECT 114.905 195.725 115.075 195.895 ;
        RECT 115.365 195.725 115.535 195.895 ;
        RECT 115.825 195.725 115.995 195.895 ;
        RECT 116.285 195.725 116.455 195.895 ;
        RECT 116.745 195.725 116.915 195.895 ;
        RECT 117.205 195.725 117.375 195.895 ;
        RECT 117.665 195.725 117.835 195.895 ;
        RECT 118.125 195.725 118.295 195.895 ;
        RECT 118.585 195.725 118.755 195.895 ;
        RECT 119.045 195.725 119.215 195.895 ;
        RECT 119.505 195.725 119.675 195.895 ;
        RECT 119.965 195.725 120.135 195.895 ;
        RECT 120.425 195.725 120.595 195.895 ;
        RECT 120.885 195.725 121.055 195.895 ;
        RECT 121.345 195.725 121.515 195.895 ;
        RECT 121.805 195.725 121.975 195.895 ;
        RECT 122.265 195.725 122.435 195.895 ;
        RECT 122.725 195.725 122.895 195.895 ;
        RECT 123.185 195.725 123.355 195.895 ;
        RECT 123.645 195.725 123.815 195.895 ;
        RECT 124.105 195.725 124.275 195.895 ;
        RECT 124.565 195.725 124.735 195.895 ;
        RECT 125.025 195.725 125.195 195.895 ;
        RECT 125.485 195.725 125.655 195.895 ;
        RECT 125.945 195.725 126.115 195.895 ;
        RECT 126.405 195.725 126.575 195.895 ;
        RECT 126.865 195.725 127.035 195.895 ;
        RECT 127.325 195.725 127.495 195.895 ;
        RECT 127.785 195.725 127.955 195.895 ;
        RECT 128.245 195.725 128.415 195.895 ;
        RECT 128.705 195.725 128.875 195.895 ;
        RECT 129.165 195.725 129.335 195.895 ;
        RECT 129.625 195.725 129.795 195.895 ;
        RECT 130.085 195.725 130.255 195.895 ;
        RECT 130.545 195.725 130.715 195.895 ;
        RECT 131.005 195.725 131.175 195.895 ;
        RECT 131.465 195.725 131.635 195.895 ;
        RECT 131.925 195.725 132.095 195.895 ;
        RECT 132.385 195.725 132.555 195.895 ;
        RECT 132.845 195.725 133.015 195.895 ;
        RECT 133.305 195.725 133.475 195.895 ;
        RECT 133.765 195.725 133.935 195.895 ;
        RECT 134.225 195.725 134.395 195.895 ;
        RECT 134.685 195.725 134.855 195.895 ;
        RECT 135.145 195.725 135.315 195.895 ;
        RECT 135.605 195.725 135.775 195.895 ;
        RECT 136.065 195.725 136.235 195.895 ;
        RECT 136.525 195.725 136.695 195.895 ;
        RECT 136.985 195.725 137.155 195.895 ;
        RECT 137.445 195.725 137.615 195.895 ;
        RECT 137.905 195.725 138.075 195.895 ;
        RECT 138.365 195.725 138.535 195.895 ;
        RECT 138.825 195.725 138.995 195.895 ;
        RECT 139.285 195.725 139.455 195.895 ;
        RECT 139.745 195.725 139.915 195.895 ;
        RECT 140.205 195.725 140.375 195.895 ;
        RECT 140.665 195.725 140.835 195.895 ;
        RECT 141.125 195.725 141.295 195.895 ;
        RECT 141.585 195.725 141.755 195.895 ;
        RECT 142.045 195.725 142.215 195.895 ;
        RECT 142.505 195.725 142.675 195.895 ;
        RECT 142.965 195.725 143.135 195.895 ;
        RECT 143.425 195.725 143.595 195.895 ;
        RECT 143.885 195.725 144.055 195.895 ;
        RECT 144.345 195.725 144.515 195.895 ;
        RECT 144.805 195.725 144.975 195.895 ;
        RECT 145.265 195.725 145.435 195.895 ;
        RECT 145.725 195.725 145.895 195.895 ;
        RECT 146.185 195.725 146.355 195.895 ;
        RECT 146.645 195.725 146.815 195.895 ;
        RECT 147.105 195.725 147.275 195.895 ;
        RECT 147.565 195.725 147.735 195.895 ;
        RECT 148.025 195.725 148.195 195.895 ;
        RECT 148.485 195.725 148.655 195.895 ;
        RECT 148.945 195.725 149.115 195.895 ;
        RECT 149.405 195.725 149.575 195.895 ;
        RECT 149.865 195.725 150.035 195.895 ;
        RECT 39.465 194.195 39.635 194.365 ;
        RECT 39.950 193.855 40.120 194.025 ;
        RECT 40.345 194.195 40.515 194.365 ;
        RECT 40.800 194.535 40.970 194.705 ;
        RECT 41.535 194.195 41.705 194.365 ;
        RECT 42.050 193.855 42.220 194.025 ;
        RECT 43.620 193.855 43.790 194.025 ;
        RECT 44.055 194.195 44.225 194.365 ;
        RECT 46.365 193.855 46.535 194.025 ;
        RECT 50.505 194.535 50.675 194.705 ;
        RECT 53.265 194.535 53.435 194.705 ;
        RECT 55.105 194.535 55.275 194.705 ;
        RECT 49.585 193.515 49.755 193.685 ;
        RECT 52.805 193.855 52.975 194.025 ;
        RECT 53.725 193.515 53.895 193.685 ;
        RECT 55.565 193.515 55.735 193.685 ;
        RECT 56.025 193.515 56.195 193.685 ;
        RECT 57.405 194.535 57.575 194.705 ;
        RECT 56.485 194.195 56.655 194.365 ;
        RECT 61.085 195.215 61.255 195.385 ;
        RECT 59.705 194.535 59.875 194.705 ;
        RECT 60.165 194.535 60.335 194.705 ;
        RECT 59.245 193.855 59.415 194.025 ;
        RECT 63.385 195.215 63.555 195.385 ;
        RECT 62.465 194.195 62.635 194.365 ;
        RECT 63.385 194.195 63.555 194.365 ;
        RECT 64.765 194.875 64.935 195.045 ;
        RECT 65.225 194.535 65.395 194.705 ;
        RECT 63.845 193.855 64.015 194.025 ;
        RECT 64.305 193.515 64.475 193.685 ;
        RECT 65.685 193.515 65.855 193.685 ;
        RECT 67.065 194.875 67.235 195.045 ;
        RECT 68.905 195.215 69.075 195.385 ;
        RECT 66.605 193.515 66.775 193.685 ;
        RECT 68.445 194.195 68.615 194.365 ;
        RECT 73.045 195.215 73.215 195.385 ;
        RECT 67.985 193.855 68.155 194.025 ;
        RECT 68.905 193.515 69.075 193.685 ;
        RECT 69.825 193.855 69.995 194.025 ;
        RECT 73.965 194.875 74.135 195.045 ;
        RECT 76.725 194.875 76.895 195.045 ;
        RECT 77.150 195.215 77.320 195.385 ;
        RECT 73.965 193.515 74.135 193.685 ;
        RECT 76.265 194.535 76.435 194.705 ;
        RECT 75.805 194.195 75.975 194.365 ;
        RECT 77.645 194.535 77.815 194.705 ;
        RECT 86.385 195.215 86.555 195.385 ;
        RECT 80.865 194.535 81.035 194.705 ;
        RECT 85.465 194.535 85.635 194.705 ;
        RECT 79.945 193.515 80.115 193.685 ;
        RECT 88.685 195.215 88.855 195.385 ;
        RECT 89.605 194.535 89.775 194.705 ;
        RECT 91.445 194.535 91.615 194.705 ;
        RECT 90.525 193.855 90.695 194.025 ;
        RECT 92.825 194.195 92.995 194.365 ;
        RECT 98.805 194.535 98.975 194.705 ;
        RECT 100.185 194.195 100.355 194.365 ;
        RECT 103.865 195.215 104.035 195.385 ;
        RECT 104.785 195.215 104.955 195.385 ;
        RECT 103.405 194.535 103.575 194.705 ;
        RECT 104.325 194.535 104.495 194.705 ;
        RECT 105.705 194.535 105.875 194.705 ;
        RECT 108.925 194.195 109.095 194.365 ;
        RECT 110.305 194.195 110.475 194.365 ;
        RECT 111.685 194.875 111.855 195.045 ;
        RECT 112.605 194.875 112.775 195.045 ;
        RECT 113.985 194.535 114.155 194.705 ;
        RECT 110.765 193.515 110.935 193.685 ;
        RECT 114.445 194.195 114.615 194.365 ;
        RECT 119.965 194.195 120.135 194.365 ;
        RECT 121.345 194.535 121.515 194.705 ;
        RECT 122.725 194.535 122.895 194.705 ;
        RECT 123.185 194.195 123.355 194.365 ;
        RECT 123.645 194.535 123.815 194.705 ;
        RECT 125.945 194.875 126.115 195.045 ;
        RECT 127.785 195.215 127.955 195.385 ;
        RECT 125.485 194.535 125.655 194.705 ;
        RECT 126.865 194.535 127.035 194.705 ;
        RECT 124.105 194.195 124.275 194.365 ;
        RECT 125.025 194.195 125.195 194.365 ;
        RECT 134.225 194.875 134.395 195.045 ;
        RECT 133.305 194.195 133.475 194.365 ;
        RECT 134.685 195.215 134.855 195.385 ;
        RECT 137.905 194.535 138.075 194.705 ;
        RECT 138.825 194.535 138.995 194.705 ;
        RECT 136.985 194.195 137.155 194.365 ;
        RECT 136.525 193.855 136.695 194.025 ;
        RECT 139.745 194.535 139.915 194.705 ;
        RECT 140.230 193.855 140.400 194.025 ;
        RECT 140.625 194.195 140.795 194.365 ;
        RECT 140.970 194.875 141.140 195.045 ;
        RECT 141.815 194.195 141.985 194.365 ;
        RECT 142.330 193.855 142.500 194.025 ;
        RECT 143.900 193.855 144.070 194.025 ;
        RECT 144.335 194.195 144.505 194.365 ;
        RECT 146.645 193.515 146.815 193.685 ;
        RECT 36.245 193.005 36.415 193.175 ;
        RECT 36.705 193.005 36.875 193.175 ;
        RECT 37.165 193.005 37.335 193.175 ;
        RECT 37.625 193.005 37.795 193.175 ;
        RECT 38.085 193.005 38.255 193.175 ;
        RECT 38.545 193.005 38.715 193.175 ;
        RECT 39.005 193.005 39.175 193.175 ;
        RECT 39.465 193.005 39.635 193.175 ;
        RECT 39.925 193.005 40.095 193.175 ;
        RECT 40.385 193.005 40.555 193.175 ;
        RECT 40.845 193.005 41.015 193.175 ;
        RECT 41.305 193.005 41.475 193.175 ;
        RECT 41.765 193.005 41.935 193.175 ;
        RECT 42.225 193.005 42.395 193.175 ;
        RECT 42.685 193.005 42.855 193.175 ;
        RECT 43.145 193.005 43.315 193.175 ;
        RECT 43.605 193.005 43.775 193.175 ;
        RECT 44.065 193.005 44.235 193.175 ;
        RECT 44.525 193.005 44.695 193.175 ;
        RECT 44.985 193.005 45.155 193.175 ;
        RECT 45.445 193.005 45.615 193.175 ;
        RECT 45.905 193.005 46.075 193.175 ;
        RECT 46.365 193.005 46.535 193.175 ;
        RECT 46.825 193.005 46.995 193.175 ;
        RECT 47.285 193.005 47.455 193.175 ;
        RECT 47.745 193.005 47.915 193.175 ;
        RECT 48.205 193.005 48.375 193.175 ;
        RECT 48.665 193.005 48.835 193.175 ;
        RECT 49.125 193.005 49.295 193.175 ;
        RECT 49.585 193.005 49.755 193.175 ;
        RECT 50.045 193.005 50.215 193.175 ;
        RECT 50.505 193.005 50.675 193.175 ;
        RECT 50.965 193.005 51.135 193.175 ;
        RECT 51.425 193.005 51.595 193.175 ;
        RECT 51.885 193.005 52.055 193.175 ;
        RECT 52.345 193.005 52.515 193.175 ;
        RECT 52.805 193.005 52.975 193.175 ;
        RECT 53.265 193.005 53.435 193.175 ;
        RECT 53.725 193.005 53.895 193.175 ;
        RECT 54.185 193.005 54.355 193.175 ;
        RECT 54.645 193.005 54.815 193.175 ;
        RECT 55.105 193.005 55.275 193.175 ;
        RECT 55.565 193.005 55.735 193.175 ;
        RECT 56.025 193.005 56.195 193.175 ;
        RECT 56.485 193.005 56.655 193.175 ;
        RECT 56.945 193.005 57.115 193.175 ;
        RECT 57.405 193.005 57.575 193.175 ;
        RECT 57.865 193.005 58.035 193.175 ;
        RECT 58.325 193.005 58.495 193.175 ;
        RECT 58.785 193.005 58.955 193.175 ;
        RECT 59.245 193.005 59.415 193.175 ;
        RECT 59.705 193.005 59.875 193.175 ;
        RECT 60.165 193.005 60.335 193.175 ;
        RECT 60.625 193.005 60.795 193.175 ;
        RECT 61.085 193.005 61.255 193.175 ;
        RECT 61.545 193.005 61.715 193.175 ;
        RECT 62.005 193.005 62.175 193.175 ;
        RECT 62.465 193.005 62.635 193.175 ;
        RECT 62.925 193.005 63.095 193.175 ;
        RECT 63.385 193.005 63.555 193.175 ;
        RECT 63.845 193.005 64.015 193.175 ;
        RECT 64.305 193.005 64.475 193.175 ;
        RECT 64.765 193.005 64.935 193.175 ;
        RECT 65.225 193.005 65.395 193.175 ;
        RECT 65.685 193.005 65.855 193.175 ;
        RECT 66.145 193.005 66.315 193.175 ;
        RECT 66.605 193.005 66.775 193.175 ;
        RECT 67.065 193.005 67.235 193.175 ;
        RECT 67.525 193.005 67.695 193.175 ;
        RECT 67.985 193.005 68.155 193.175 ;
        RECT 68.445 193.005 68.615 193.175 ;
        RECT 68.905 193.005 69.075 193.175 ;
        RECT 69.365 193.005 69.535 193.175 ;
        RECT 69.825 193.005 69.995 193.175 ;
        RECT 70.285 193.005 70.455 193.175 ;
        RECT 70.745 193.005 70.915 193.175 ;
        RECT 71.205 193.005 71.375 193.175 ;
        RECT 71.665 193.005 71.835 193.175 ;
        RECT 72.125 193.005 72.295 193.175 ;
        RECT 72.585 193.005 72.755 193.175 ;
        RECT 73.045 193.005 73.215 193.175 ;
        RECT 73.505 193.005 73.675 193.175 ;
        RECT 73.965 193.005 74.135 193.175 ;
        RECT 74.425 193.005 74.595 193.175 ;
        RECT 74.885 193.005 75.055 193.175 ;
        RECT 75.345 193.005 75.515 193.175 ;
        RECT 75.805 193.005 75.975 193.175 ;
        RECT 76.265 193.005 76.435 193.175 ;
        RECT 76.725 193.005 76.895 193.175 ;
        RECT 77.185 193.005 77.355 193.175 ;
        RECT 77.645 193.005 77.815 193.175 ;
        RECT 78.105 193.005 78.275 193.175 ;
        RECT 78.565 193.005 78.735 193.175 ;
        RECT 79.025 193.005 79.195 193.175 ;
        RECT 79.485 193.005 79.655 193.175 ;
        RECT 79.945 193.005 80.115 193.175 ;
        RECT 80.405 193.005 80.575 193.175 ;
        RECT 80.865 193.005 81.035 193.175 ;
        RECT 81.325 193.005 81.495 193.175 ;
        RECT 81.785 193.005 81.955 193.175 ;
        RECT 82.245 193.005 82.415 193.175 ;
        RECT 82.705 193.005 82.875 193.175 ;
        RECT 83.165 193.005 83.335 193.175 ;
        RECT 83.625 193.005 83.795 193.175 ;
        RECT 84.085 193.005 84.255 193.175 ;
        RECT 84.545 193.005 84.715 193.175 ;
        RECT 85.005 193.005 85.175 193.175 ;
        RECT 85.465 193.005 85.635 193.175 ;
        RECT 85.925 193.005 86.095 193.175 ;
        RECT 86.385 193.005 86.555 193.175 ;
        RECT 86.845 193.005 87.015 193.175 ;
        RECT 87.305 193.005 87.475 193.175 ;
        RECT 87.765 193.005 87.935 193.175 ;
        RECT 88.225 193.005 88.395 193.175 ;
        RECT 88.685 193.005 88.855 193.175 ;
        RECT 89.145 193.005 89.315 193.175 ;
        RECT 89.605 193.005 89.775 193.175 ;
        RECT 90.065 193.005 90.235 193.175 ;
        RECT 90.525 193.005 90.695 193.175 ;
        RECT 90.985 193.005 91.155 193.175 ;
        RECT 91.445 193.005 91.615 193.175 ;
        RECT 91.905 193.005 92.075 193.175 ;
        RECT 92.365 193.005 92.535 193.175 ;
        RECT 92.825 193.005 92.995 193.175 ;
        RECT 93.285 193.005 93.455 193.175 ;
        RECT 93.745 193.005 93.915 193.175 ;
        RECT 94.205 193.005 94.375 193.175 ;
        RECT 94.665 193.005 94.835 193.175 ;
        RECT 95.125 193.005 95.295 193.175 ;
        RECT 95.585 193.005 95.755 193.175 ;
        RECT 96.045 193.005 96.215 193.175 ;
        RECT 96.505 193.005 96.675 193.175 ;
        RECT 96.965 193.005 97.135 193.175 ;
        RECT 97.425 193.005 97.595 193.175 ;
        RECT 97.885 193.005 98.055 193.175 ;
        RECT 98.345 193.005 98.515 193.175 ;
        RECT 98.805 193.005 98.975 193.175 ;
        RECT 99.265 193.005 99.435 193.175 ;
        RECT 99.725 193.005 99.895 193.175 ;
        RECT 100.185 193.005 100.355 193.175 ;
        RECT 100.645 193.005 100.815 193.175 ;
        RECT 101.105 193.005 101.275 193.175 ;
        RECT 101.565 193.005 101.735 193.175 ;
        RECT 102.025 193.005 102.195 193.175 ;
        RECT 102.485 193.005 102.655 193.175 ;
        RECT 102.945 193.005 103.115 193.175 ;
        RECT 103.405 193.005 103.575 193.175 ;
        RECT 103.865 193.005 104.035 193.175 ;
        RECT 104.325 193.005 104.495 193.175 ;
        RECT 104.785 193.005 104.955 193.175 ;
        RECT 105.245 193.005 105.415 193.175 ;
        RECT 105.705 193.005 105.875 193.175 ;
        RECT 106.165 193.005 106.335 193.175 ;
        RECT 106.625 193.005 106.795 193.175 ;
        RECT 107.085 193.005 107.255 193.175 ;
        RECT 107.545 193.005 107.715 193.175 ;
        RECT 108.005 193.005 108.175 193.175 ;
        RECT 108.465 193.005 108.635 193.175 ;
        RECT 108.925 193.005 109.095 193.175 ;
        RECT 109.385 193.005 109.555 193.175 ;
        RECT 109.845 193.005 110.015 193.175 ;
        RECT 110.305 193.005 110.475 193.175 ;
        RECT 110.765 193.005 110.935 193.175 ;
        RECT 111.225 193.005 111.395 193.175 ;
        RECT 111.685 193.005 111.855 193.175 ;
        RECT 112.145 193.005 112.315 193.175 ;
        RECT 112.605 193.005 112.775 193.175 ;
        RECT 113.065 193.005 113.235 193.175 ;
        RECT 113.525 193.005 113.695 193.175 ;
        RECT 113.985 193.005 114.155 193.175 ;
        RECT 114.445 193.005 114.615 193.175 ;
        RECT 114.905 193.005 115.075 193.175 ;
        RECT 115.365 193.005 115.535 193.175 ;
        RECT 115.825 193.005 115.995 193.175 ;
        RECT 116.285 193.005 116.455 193.175 ;
        RECT 116.745 193.005 116.915 193.175 ;
        RECT 117.205 193.005 117.375 193.175 ;
        RECT 117.665 193.005 117.835 193.175 ;
        RECT 118.125 193.005 118.295 193.175 ;
        RECT 118.585 193.005 118.755 193.175 ;
        RECT 119.045 193.005 119.215 193.175 ;
        RECT 119.505 193.005 119.675 193.175 ;
        RECT 119.965 193.005 120.135 193.175 ;
        RECT 120.425 193.005 120.595 193.175 ;
        RECT 120.885 193.005 121.055 193.175 ;
        RECT 121.345 193.005 121.515 193.175 ;
        RECT 121.805 193.005 121.975 193.175 ;
        RECT 122.265 193.005 122.435 193.175 ;
        RECT 122.725 193.005 122.895 193.175 ;
        RECT 123.185 193.005 123.355 193.175 ;
        RECT 123.645 193.005 123.815 193.175 ;
        RECT 124.105 193.005 124.275 193.175 ;
        RECT 124.565 193.005 124.735 193.175 ;
        RECT 125.025 193.005 125.195 193.175 ;
        RECT 125.485 193.005 125.655 193.175 ;
        RECT 125.945 193.005 126.115 193.175 ;
        RECT 126.405 193.005 126.575 193.175 ;
        RECT 126.865 193.005 127.035 193.175 ;
        RECT 127.325 193.005 127.495 193.175 ;
        RECT 127.785 193.005 127.955 193.175 ;
        RECT 128.245 193.005 128.415 193.175 ;
        RECT 128.705 193.005 128.875 193.175 ;
        RECT 129.165 193.005 129.335 193.175 ;
        RECT 129.625 193.005 129.795 193.175 ;
        RECT 130.085 193.005 130.255 193.175 ;
        RECT 130.545 193.005 130.715 193.175 ;
        RECT 131.005 193.005 131.175 193.175 ;
        RECT 131.465 193.005 131.635 193.175 ;
        RECT 131.925 193.005 132.095 193.175 ;
        RECT 132.385 193.005 132.555 193.175 ;
        RECT 132.845 193.005 133.015 193.175 ;
        RECT 133.305 193.005 133.475 193.175 ;
        RECT 133.765 193.005 133.935 193.175 ;
        RECT 134.225 193.005 134.395 193.175 ;
        RECT 134.685 193.005 134.855 193.175 ;
        RECT 135.145 193.005 135.315 193.175 ;
        RECT 135.605 193.005 135.775 193.175 ;
        RECT 136.065 193.005 136.235 193.175 ;
        RECT 136.525 193.005 136.695 193.175 ;
        RECT 136.985 193.005 137.155 193.175 ;
        RECT 137.445 193.005 137.615 193.175 ;
        RECT 137.905 193.005 138.075 193.175 ;
        RECT 138.365 193.005 138.535 193.175 ;
        RECT 138.825 193.005 138.995 193.175 ;
        RECT 139.285 193.005 139.455 193.175 ;
        RECT 139.745 193.005 139.915 193.175 ;
        RECT 140.205 193.005 140.375 193.175 ;
        RECT 140.665 193.005 140.835 193.175 ;
        RECT 141.125 193.005 141.295 193.175 ;
        RECT 141.585 193.005 141.755 193.175 ;
        RECT 142.045 193.005 142.215 193.175 ;
        RECT 142.505 193.005 142.675 193.175 ;
        RECT 142.965 193.005 143.135 193.175 ;
        RECT 143.425 193.005 143.595 193.175 ;
        RECT 143.885 193.005 144.055 193.175 ;
        RECT 144.345 193.005 144.515 193.175 ;
        RECT 144.805 193.005 144.975 193.175 ;
        RECT 145.265 193.005 145.435 193.175 ;
        RECT 145.725 193.005 145.895 193.175 ;
        RECT 146.185 193.005 146.355 193.175 ;
        RECT 146.645 193.005 146.815 193.175 ;
        RECT 147.105 193.005 147.275 193.175 ;
        RECT 147.565 193.005 147.735 193.175 ;
        RECT 148.025 193.005 148.195 193.175 ;
        RECT 148.485 193.005 148.655 193.175 ;
        RECT 148.945 193.005 149.115 193.175 ;
        RECT 149.405 193.005 149.575 193.175 ;
        RECT 149.865 193.005 150.035 193.175 ;
        RECT 42.685 192.495 42.855 192.665 ;
        RECT 42.225 191.815 42.395 191.985 ;
        RECT 43.145 191.475 43.315 191.645 ;
        RECT 43.605 191.475 43.775 191.645 ;
        RECT 53.265 192.495 53.435 192.665 ;
        RECT 53.265 191.475 53.435 191.645 ;
        RECT 55.105 191.475 55.275 191.645 ;
        RECT 55.565 191.475 55.735 191.645 ;
        RECT 52.345 190.795 52.515 190.965 ;
        RECT 56.485 191.475 56.655 191.645 ;
        RECT 57.405 191.475 57.575 191.645 ;
        RECT 59.705 191.815 59.875 191.985 ;
        RECT 59.245 191.135 59.415 191.305 ;
        RECT 58.785 190.795 58.955 190.965 ;
        RECT 61.545 191.475 61.715 191.645 ;
        RECT 64.765 191.815 64.935 191.985 ;
        RECT 67.065 192.495 67.235 192.665 ;
        RECT 66.145 191.475 66.315 191.645 ;
        RECT 60.625 190.795 60.795 190.965 ;
        RECT 67.525 191.135 67.695 191.305 ;
        RECT 75.345 192.495 75.515 192.665 ;
        RECT 78.565 192.495 78.735 192.665 ;
        RECT 78.105 191.815 78.275 191.985 ;
        RECT 76.495 191.475 76.665 191.645 ;
        RECT 77.185 191.475 77.355 191.645 ;
        RECT 79.025 192.155 79.195 192.325 ;
        RECT 77.645 191.475 77.815 191.645 ;
        RECT 79.480 191.365 79.650 191.535 ;
        RECT 80.865 191.475 81.035 191.645 ;
        RECT 79.945 190.795 80.115 190.965 ;
        RECT 87.765 192.495 87.935 192.665 ;
        RECT 88.685 191.475 88.855 191.645 ;
        RECT 90.065 191.815 90.235 191.985 ;
        RECT 91.905 192.495 92.075 192.665 ;
        RECT 89.605 191.475 89.775 191.645 ;
        RECT 90.525 191.475 90.695 191.645 ;
        RECT 91.445 191.475 91.615 191.645 ;
        RECT 93.745 192.155 93.915 192.325 ;
        RECT 95.585 192.155 95.755 192.325 ;
        RECT 92.825 191.475 92.995 191.645 ;
        RECT 94.205 191.475 94.375 191.645 ;
        RECT 96.965 192.495 97.135 192.665 ;
        RECT 96.505 191.475 96.675 191.645 ;
        RECT 98.345 191.475 98.515 191.645 ;
        RECT 98.805 191.475 98.975 191.645 ;
        RECT 99.265 191.475 99.435 191.645 ;
        RECT 101.105 192.155 101.275 192.325 ;
        RECT 100.185 191.475 100.355 191.645 ;
        RECT 102.025 191.475 102.195 191.645 ;
        RECT 105.245 192.495 105.415 192.665 ;
        RECT 102.945 191.475 103.115 191.645 ;
        RECT 103.405 191.475 103.575 191.645 ;
        RECT 103.865 191.475 104.035 191.645 ;
        RECT 104.785 191.425 104.955 191.595 ;
        RECT 108.005 192.155 108.175 192.325 ;
        RECT 106.150 191.475 106.320 191.645 ;
        RECT 108.465 191.475 108.635 191.645 ;
        RECT 108.925 191.475 109.095 191.645 ;
        RECT 110.305 191.815 110.475 191.985 ;
        RECT 109.845 191.475 110.015 191.645 ;
        RECT 111.685 191.475 111.855 191.645 ;
        RECT 109.845 190.795 110.015 190.965 ;
        RECT 114.905 192.495 115.075 192.665 ;
        RECT 115.825 191.475 115.995 191.645 ;
        RECT 116.285 191.475 116.455 191.645 ;
        RECT 116.745 191.815 116.915 191.985 ;
        RECT 119.965 192.495 120.135 192.665 ;
        RECT 117.205 191.475 117.375 191.645 ;
        RECT 119.045 191.475 119.215 191.645 ;
        RECT 121.345 192.155 121.515 192.325 ;
        RECT 120.425 191.475 120.595 191.645 ;
        RECT 127.785 192.495 127.955 192.665 ;
        RECT 131.465 192.495 131.635 192.665 ;
        RECT 128.705 191.475 128.875 191.645 ;
        RECT 129.165 191.475 129.335 191.645 ;
        RECT 130.545 191.475 130.715 191.645 ;
        RECT 129.625 191.135 129.795 191.305 ;
        RECT 132.845 192.495 133.015 192.665 ;
        RECT 134.685 192.495 134.855 192.665 ;
        RECT 132.615 191.305 132.785 191.475 ;
        RECT 131.925 190.795 132.095 190.965 ;
        RECT 134.225 191.475 134.395 191.645 ;
        RECT 133.765 191.135 133.935 191.305 ;
        RECT 137.905 192.495 138.075 192.665 ;
        RECT 136.985 191.475 137.155 191.645 ;
        RECT 141.125 191.815 141.295 191.985 ;
        RECT 142.505 191.475 142.675 191.645 ;
        RECT 142.965 191.135 143.135 191.305 ;
        RECT 144.345 191.475 144.515 191.645 ;
        RECT 143.885 191.135 144.055 191.305 ;
        RECT 143.425 190.795 143.595 190.965 ;
        RECT 36.245 190.285 36.415 190.455 ;
        RECT 36.705 190.285 36.875 190.455 ;
        RECT 37.165 190.285 37.335 190.455 ;
        RECT 37.625 190.285 37.795 190.455 ;
        RECT 38.085 190.285 38.255 190.455 ;
        RECT 38.545 190.285 38.715 190.455 ;
        RECT 39.005 190.285 39.175 190.455 ;
        RECT 39.465 190.285 39.635 190.455 ;
        RECT 39.925 190.285 40.095 190.455 ;
        RECT 40.385 190.285 40.555 190.455 ;
        RECT 40.845 190.285 41.015 190.455 ;
        RECT 41.305 190.285 41.475 190.455 ;
        RECT 41.765 190.285 41.935 190.455 ;
        RECT 42.225 190.285 42.395 190.455 ;
        RECT 42.685 190.285 42.855 190.455 ;
        RECT 43.145 190.285 43.315 190.455 ;
        RECT 43.605 190.285 43.775 190.455 ;
        RECT 44.065 190.285 44.235 190.455 ;
        RECT 44.525 190.285 44.695 190.455 ;
        RECT 44.985 190.285 45.155 190.455 ;
        RECT 45.445 190.285 45.615 190.455 ;
        RECT 45.905 190.285 46.075 190.455 ;
        RECT 46.365 190.285 46.535 190.455 ;
        RECT 46.825 190.285 46.995 190.455 ;
        RECT 47.285 190.285 47.455 190.455 ;
        RECT 47.745 190.285 47.915 190.455 ;
        RECT 48.205 190.285 48.375 190.455 ;
        RECT 48.665 190.285 48.835 190.455 ;
        RECT 49.125 190.285 49.295 190.455 ;
        RECT 49.585 190.285 49.755 190.455 ;
        RECT 50.045 190.285 50.215 190.455 ;
        RECT 50.505 190.285 50.675 190.455 ;
        RECT 50.965 190.285 51.135 190.455 ;
        RECT 51.425 190.285 51.595 190.455 ;
        RECT 51.885 190.285 52.055 190.455 ;
        RECT 52.345 190.285 52.515 190.455 ;
        RECT 52.805 190.285 52.975 190.455 ;
        RECT 53.265 190.285 53.435 190.455 ;
        RECT 53.725 190.285 53.895 190.455 ;
        RECT 54.185 190.285 54.355 190.455 ;
        RECT 54.645 190.285 54.815 190.455 ;
        RECT 55.105 190.285 55.275 190.455 ;
        RECT 55.565 190.285 55.735 190.455 ;
        RECT 56.025 190.285 56.195 190.455 ;
        RECT 56.485 190.285 56.655 190.455 ;
        RECT 56.945 190.285 57.115 190.455 ;
        RECT 57.405 190.285 57.575 190.455 ;
        RECT 57.865 190.285 58.035 190.455 ;
        RECT 58.325 190.285 58.495 190.455 ;
        RECT 58.785 190.285 58.955 190.455 ;
        RECT 59.245 190.285 59.415 190.455 ;
        RECT 59.705 190.285 59.875 190.455 ;
        RECT 60.165 190.285 60.335 190.455 ;
        RECT 60.625 190.285 60.795 190.455 ;
        RECT 61.085 190.285 61.255 190.455 ;
        RECT 61.545 190.285 61.715 190.455 ;
        RECT 62.005 190.285 62.175 190.455 ;
        RECT 62.465 190.285 62.635 190.455 ;
        RECT 62.925 190.285 63.095 190.455 ;
        RECT 63.385 190.285 63.555 190.455 ;
        RECT 63.845 190.285 64.015 190.455 ;
        RECT 64.305 190.285 64.475 190.455 ;
        RECT 64.765 190.285 64.935 190.455 ;
        RECT 65.225 190.285 65.395 190.455 ;
        RECT 65.685 190.285 65.855 190.455 ;
        RECT 66.145 190.285 66.315 190.455 ;
        RECT 66.605 190.285 66.775 190.455 ;
        RECT 67.065 190.285 67.235 190.455 ;
        RECT 67.525 190.285 67.695 190.455 ;
        RECT 67.985 190.285 68.155 190.455 ;
        RECT 68.445 190.285 68.615 190.455 ;
        RECT 68.905 190.285 69.075 190.455 ;
        RECT 69.365 190.285 69.535 190.455 ;
        RECT 69.825 190.285 69.995 190.455 ;
        RECT 70.285 190.285 70.455 190.455 ;
        RECT 70.745 190.285 70.915 190.455 ;
        RECT 71.205 190.285 71.375 190.455 ;
        RECT 71.665 190.285 71.835 190.455 ;
        RECT 72.125 190.285 72.295 190.455 ;
        RECT 72.585 190.285 72.755 190.455 ;
        RECT 73.045 190.285 73.215 190.455 ;
        RECT 73.505 190.285 73.675 190.455 ;
        RECT 73.965 190.285 74.135 190.455 ;
        RECT 74.425 190.285 74.595 190.455 ;
        RECT 74.885 190.285 75.055 190.455 ;
        RECT 75.345 190.285 75.515 190.455 ;
        RECT 75.805 190.285 75.975 190.455 ;
        RECT 76.265 190.285 76.435 190.455 ;
        RECT 76.725 190.285 76.895 190.455 ;
        RECT 77.185 190.285 77.355 190.455 ;
        RECT 77.645 190.285 77.815 190.455 ;
        RECT 78.105 190.285 78.275 190.455 ;
        RECT 78.565 190.285 78.735 190.455 ;
        RECT 79.025 190.285 79.195 190.455 ;
        RECT 79.485 190.285 79.655 190.455 ;
        RECT 79.945 190.285 80.115 190.455 ;
        RECT 80.405 190.285 80.575 190.455 ;
        RECT 80.865 190.285 81.035 190.455 ;
        RECT 81.325 190.285 81.495 190.455 ;
        RECT 81.785 190.285 81.955 190.455 ;
        RECT 82.245 190.285 82.415 190.455 ;
        RECT 82.705 190.285 82.875 190.455 ;
        RECT 83.165 190.285 83.335 190.455 ;
        RECT 83.625 190.285 83.795 190.455 ;
        RECT 84.085 190.285 84.255 190.455 ;
        RECT 84.545 190.285 84.715 190.455 ;
        RECT 85.005 190.285 85.175 190.455 ;
        RECT 85.465 190.285 85.635 190.455 ;
        RECT 85.925 190.285 86.095 190.455 ;
        RECT 86.385 190.285 86.555 190.455 ;
        RECT 86.845 190.285 87.015 190.455 ;
        RECT 87.305 190.285 87.475 190.455 ;
        RECT 87.765 190.285 87.935 190.455 ;
        RECT 88.225 190.285 88.395 190.455 ;
        RECT 88.685 190.285 88.855 190.455 ;
        RECT 89.145 190.285 89.315 190.455 ;
        RECT 89.605 190.285 89.775 190.455 ;
        RECT 90.065 190.285 90.235 190.455 ;
        RECT 90.525 190.285 90.695 190.455 ;
        RECT 90.985 190.285 91.155 190.455 ;
        RECT 91.445 190.285 91.615 190.455 ;
        RECT 91.905 190.285 92.075 190.455 ;
        RECT 92.365 190.285 92.535 190.455 ;
        RECT 92.825 190.285 92.995 190.455 ;
        RECT 93.285 190.285 93.455 190.455 ;
        RECT 93.745 190.285 93.915 190.455 ;
        RECT 94.205 190.285 94.375 190.455 ;
        RECT 94.665 190.285 94.835 190.455 ;
        RECT 95.125 190.285 95.295 190.455 ;
        RECT 95.585 190.285 95.755 190.455 ;
        RECT 96.045 190.285 96.215 190.455 ;
        RECT 96.505 190.285 96.675 190.455 ;
        RECT 96.965 190.285 97.135 190.455 ;
        RECT 97.425 190.285 97.595 190.455 ;
        RECT 97.885 190.285 98.055 190.455 ;
        RECT 98.345 190.285 98.515 190.455 ;
        RECT 98.805 190.285 98.975 190.455 ;
        RECT 99.265 190.285 99.435 190.455 ;
        RECT 99.725 190.285 99.895 190.455 ;
        RECT 100.185 190.285 100.355 190.455 ;
        RECT 100.645 190.285 100.815 190.455 ;
        RECT 101.105 190.285 101.275 190.455 ;
        RECT 101.565 190.285 101.735 190.455 ;
        RECT 102.025 190.285 102.195 190.455 ;
        RECT 102.485 190.285 102.655 190.455 ;
        RECT 102.945 190.285 103.115 190.455 ;
        RECT 103.405 190.285 103.575 190.455 ;
        RECT 103.865 190.285 104.035 190.455 ;
        RECT 104.325 190.285 104.495 190.455 ;
        RECT 104.785 190.285 104.955 190.455 ;
        RECT 105.245 190.285 105.415 190.455 ;
        RECT 105.705 190.285 105.875 190.455 ;
        RECT 106.165 190.285 106.335 190.455 ;
        RECT 106.625 190.285 106.795 190.455 ;
        RECT 107.085 190.285 107.255 190.455 ;
        RECT 107.545 190.285 107.715 190.455 ;
        RECT 108.005 190.285 108.175 190.455 ;
        RECT 108.465 190.285 108.635 190.455 ;
        RECT 108.925 190.285 109.095 190.455 ;
        RECT 109.385 190.285 109.555 190.455 ;
        RECT 109.845 190.285 110.015 190.455 ;
        RECT 110.305 190.285 110.475 190.455 ;
        RECT 110.765 190.285 110.935 190.455 ;
        RECT 111.225 190.285 111.395 190.455 ;
        RECT 111.685 190.285 111.855 190.455 ;
        RECT 112.145 190.285 112.315 190.455 ;
        RECT 112.605 190.285 112.775 190.455 ;
        RECT 113.065 190.285 113.235 190.455 ;
        RECT 113.525 190.285 113.695 190.455 ;
        RECT 113.985 190.285 114.155 190.455 ;
        RECT 114.445 190.285 114.615 190.455 ;
        RECT 114.905 190.285 115.075 190.455 ;
        RECT 115.365 190.285 115.535 190.455 ;
        RECT 115.825 190.285 115.995 190.455 ;
        RECT 116.285 190.285 116.455 190.455 ;
        RECT 116.745 190.285 116.915 190.455 ;
        RECT 117.205 190.285 117.375 190.455 ;
        RECT 117.665 190.285 117.835 190.455 ;
        RECT 118.125 190.285 118.295 190.455 ;
        RECT 118.585 190.285 118.755 190.455 ;
        RECT 119.045 190.285 119.215 190.455 ;
        RECT 119.505 190.285 119.675 190.455 ;
        RECT 119.965 190.285 120.135 190.455 ;
        RECT 120.425 190.285 120.595 190.455 ;
        RECT 120.885 190.285 121.055 190.455 ;
        RECT 121.345 190.285 121.515 190.455 ;
        RECT 121.805 190.285 121.975 190.455 ;
        RECT 122.265 190.285 122.435 190.455 ;
        RECT 122.725 190.285 122.895 190.455 ;
        RECT 123.185 190.285 123.355 190.455 ;
        RECT 123.645 190.285 123.815 190.455 ;
        RECT 124.105 190.285 124.275 190.455 ;
        RECT 124.565 190.285 124.735 190.455 ;
        RECT 125.025 190.285 125.195 190.455 ;
        RECT 125.485 190.285 125.655 190.455 ;
        RECT 125.945 190.285 126.115 190.455 ;
        RECT 126.405 190.285 126.575 190.455 ;
        RECT 126.865 190.285 127.035 190.455 ;
        RECT 127.325 190.285 127.495 190.455 ;
        RECT 127.785 190.285 127.955 190.455 ;
        RECT 128.245 190.285 128.415 190.455 ;
        RECT 128.705 190.285 128.875 190.455 ;
        RECT 129.165 190.285 129.335 190.455 ;
        RECT 129.625 190.285 129.795 190.455 ;
        RECT 130.085 190.285 130.255 190.455 ;
        RECT 130.545 190.285 130.715 190.455 ;
        RECT 131.005 190.285 131.175 190.455 ;
        RECT 131.465 190.285 131.635 190.455 ;
        RECT 131.925 190.285 132.095 190.455 ;
        RECT 132.385 190.285 132.555 190.455 ;
        RECT 132.845 190.285 133.015 190.455 ;
        RECT 133.305 190.285 133.475 190.455 ;
        RECT 133.765 190.285 133.935 190.455 ;
        RECT 134.225 190.285 134.395 190.455 ;
        RECT 134.685 190.285 134.855 190.455 ;
        RECT 135.145 190.285 135.315 190.455 ;
        RECT 135.605 190.285 135.775 190.455 ;
        RECT 136.065 190.285 136.235 190.455 ;
        RECT 136.525 190.285 136.695 190.455 ;
        RECT 136.985 190.285 137.155 190.455 ;
        RECT 137.445 190.285 137.615 190.455 ;
        RECT 137.905 190.285 138.075 190.455 ;
        RECT 138.365 190.285 138.535 190.455 ;
        RECT 138.825 190.285 138.995 190.455 ;
        RECT 139.285 190.285 139.455 190.455 ;
        RECT 139.745 190.285 139.915 190.455 ;
        RECT 140.205 190.285 140.375 190.455 ;
        RECT 140.665 190.285 140.835 190.455 ;
        RECT 141.125 190.285 141.295 190.455 ;
        RECT 141.585 190.285 141.755 190.455 ;
        RECT 142.045 190.285 142.215 190.455 ;
        RECT 142.505 190.285 142.675 190.455 ;
        RECT 142.965 190.285 143.135 190.455 ;
        RECT 143.425 190.285 143.595 190.455 ;
        RECT 143.885 190.285 144.055 190.455 ;
        RECT 144.345 190.285 144.515 190.455 ;
        RECT 144.805 190.285 144.975 190.455 ;
        RECT 145.265 190.285 145.435 190.455 ;
        RECT 145.725 190.285 145.895 190.455 ;
        RECT 146.185 190.285 146.355 190.455 ;
        RECT 146.645 190.285 146.815 190.455 ;
        RECT 147.105 190.285 147.275 190.455 ;
        RECT 147.565 190.285 147.735 190.455 ;
        RECT 148.025 190.285 148.195 190.455 ;
        RECT 148.485 190.285 148.655 190.455 ;
        RECT 148.945 190.285 149.115 190.455 ;
        RECT 149.405 190.285 149.575 190.455 ;
        RECT 149.865 190.285 150.035 190.455 ;
        RECT 42.685 189.775 42.855 189.945 ;
        RECT 41.305 189.095 41.475 189.265 ;
        RECT 41.765 189.095 41.935 189.265 ;
        RECT 40.385 188.075 40.555 188.245 ;
        RECT 43.145 189.095 43.315 189.265 ;
        RECT 44.985 189.775 45.155 189.945 ;
        RECT 44.065 189.095 44.235 189.265 ;
        RECT 44.525 189.095 44.695 189.265 ;
        RECT 43.145 188.415 43.315 188.585 ;
        RECT 47.515 189.095 47.685 189.265 ;
        RECT 48.205 188.755 48.375 188.925 ;
        RECT 49.505 189.435 49.675 189.605 ;
        RECT 50.505 189.435 50.675 189.605 ;
        RECT 48.665 188.415 48.835 188.585 ;
        RECT 49.585 188.075 49.755 188.245 ;
        RECT 56.485 189.095 56.655 189.265 ;
        RECT 57.405 189.095 57.575 189.265 ;
        RECT 56.945 188.075 57.115 188.245 ;
        RECT 60.165 189.095 60.335 189.265 ;
        RECT 61.085 188.075 61.255 188.245 ;
        RECT 72.585 189.095 72.755 189.265 ;
        RECT 74.425 189.775 74.595 189.945 ;
        RECT 66.145 188.075 66.315 188.245 ;
        RECT 75.115 189.265 75.285 189.435 ;
        RECT 76.265 189.435 76.435 189.605 ;
        RECT 75.345 188.075 75.515 188.245 ;
        RECT 77.185 188.755 77.355 188.925 ;
        RECT 78.105 188.755 78.275 188.925 ;
        RECT 79.485 189.095 79.655 189.265 ;
        RECT 84.545 189.095 84.715 189.265 ;
        RECT 85.925 189.095 86.095 189.265 ;
        RECT 86.385 189.095 86.555 189.265 ;
        RECT 77.645 188.075 77.815 188.245 ;
        RECT 78.565 188.415 78.735 188.585 ;
        RECT 87.305 189.435 87.475 189.605 ;
        RECT 85.005 188.075 85.175 188.245 ;
        RECT 88.225 189.095 88.395 189.265 ;
        RECT 91.445 189.775 91.615 189.945 ;
        RECT 89.145 189.095 89.315 189.265 ;
        RECT 89.605 189.095 89.775 189.265 ;
        RECT 90.165 189.095 90.335 189.265 ;
        RECT 98.805 189.095 98.975 189.265 ;
        RECT 99.725 189.435 99.895 189.605 ;
        RECT 101.105 189.435 101.275 189.605 ;
        RECT 100.185 189.095 100.355 189.265 ;
        RECT 100.645 189.095 100.815 189.265 ;
        RECT 101.565 189.095 101.735 189.265 ;
        RECT 98.805 188.415 98.975 188.585 ;
        RECT 107.545 189.095 107.715 189.265 ;
        RECT 116.745 189.775 116.915 189.945 ;
        RECT 106.625 188.075 106.795 188.245 ;
        RECT 119.505 189.775 119.675 189.945 ;
        RECT 117.665 189.095 117.835 189.265 ;
        RECT 120.885 189.095 121.055 189.265 ;
        RECT 128.245 189.775 128.415 189.945 ;
        RECT 119.965 188.755 120.135 188.925 ;
        RECT 130.085 188.755 130.255 188.925 ;
        RECT 131.005 189.095 131.175 189.265 ;
        RECT 135.605 189.095 135.775 189.265 ;
        RECT 134.685 188.755 134.855 188.925 ;
        RECT 140.205 189.435 140.375 189.605 ;
        RECT 141.125 189.775 141.295 189.945 ;
        RECT 144.345 189.775 144.515 189.945 ;
        RECT 139.745 189.095 139.915 189.265 ;
        RECT 136.525 188.075 136.695 188.245 ;
        RECT 142.045 188.755 142.215 188.925 ;
        RECT 142.505 188.755 142.675 188.925 ;
        RECT 142.965 189.095 143.135 189.265 ;
        RECT 143.425 188.755 143.595 188.925 ;
        RECT 145.265 189.095 145.435 189.265 ;
        RECT 146.185 188.755 146.355 188.925 ;
        RECT 36.245 187.565 36.415 187.735 ;
        RECT 36.705 187.565 36.875 187.735 ;
        RECT 37.165 187.565 37.335 187.735 ;
        RECT 37.625 187.565 37.795 187.735 ;
        RECT 38.085 187.565 38.255 187.735 ;
        RECT 38.545 187.565 38.715 187.735 ;
        RECT 39.005 187.565 39.175 187.735 ;
        RECT 39.465 187.565 39.635 187.735 ;
        RECT 39.925 187.565 40.095 187.735 ;
        RECT 40.385 187.565 40.555 187.735 ;
        RECT 40.845 187.565 41.015 187.735 ;
        RECT 41.305 187.565 41.475 187.735 ;
        RECT 41.765 187.565 41.935 187.735 ;
        RECT 42.225 187.565 42.395 187.735 ;
        RECT 42.685 187.565 42.855 187.735 ;
        RECT 43.145 187.565 43.315 187.735 ;
        RECT 43.605 187.565 43.775 187.735 ;
        RECT 44.065 187.565 44.235 187.735 ;
        RECT 44.525 187.565 44.695 187.735 ;
        RECT 44.985 187.565 45.155 187.735 ;
        RECT 45.445 187.565 45.615 187.735 ;
        RECT 45.905 187.565 46.075 187.735 ;
        RECT 46.365 187.565 46.535 187.735 ;
        RECT 46.825 187.565 46.995 187.735 ;
        RECT 47.285 187.565 47.455 187.735 ;
        RECT 47.745 187.565 47.915 187.735 ;
        RECT 48.205 187.565 48.375 187.735 ;
        RECT 48.665 187.565 48.835 187.735 ;
        RECT 49.125 187.565 49.295 187.735 ;
        RECT 49.585 187.565 49.755 187.735 ;
        RECT 50.045 187.565 50.215 187.735 ;
        RECT 50.505 187.565 50.675 187.735 ;
        RECT 50.965 187.565 51.135 187.735 ;
        RECT 51.425 187.565 51.595 187.735 ;
        RECT 51.885 187.565 52.055 187.735 ;
        RECT 52.345 187.565 52.515 187.735 ;
        RECT 52.805 187.565 52.975 187.735 ;
        RECT 53.265 187.565 53.435 187.735 ;
        RECT 53.725 187.565 53.895 187.735 ;
        RECT 54.185 187.565 54.355 187.735 ;
        RECT 54.645 187.565 54.815 187.735 ;
        RECT 55.105 187.565 55.275 187.735 ;
        RECT 55.565 187.565 55.735 187.735 ;
        RECT 56.025 187.565 56.195 187.735 ;
        RECT 56.485 187.565 56.655 187.735 ;
        RECT 56.945 187.565 57.115 187.735 ;
        RECT 57.405 187.565 57.575 187.735 ;
        RECT 57.865 187.565 58.035 187.735 ;
        RECT 58.325 187.565 58.495 187.735 ;
        RECT 58.785 187.565 58.955 187.735 ;
        RECT 59.245 187.565 59.415 187.735 ;
        RECT 59.705 187.565 59.875 187.735 ;
        RECT 60.165 187.565 60.335 187.735 ;
        RECT 60.625 187.565 60.795 187.735 ;
        RECT 61.085 187.565 61.255 187.735 ;
        RECT 61.545 187.565 61.715 187.735 ;
        RECT 62.005 187.565 62.175 187.735 ;
        RECT 62.465 187.565 62.635 187.735 ;
        RECT 62.925 187.565 63.095 187.735 ;
        RECT 63.385 187.565 63.555 187.735 ;
        RECT 63.845 187.565 64.015 187.735 ;
        RECT 64.305 187.565 64.475 187.735 ;
        RECT 64.765 187.565 64.935 187.735 ;
        RECT 65.225 187.565 65.395 187.735 ;
        RECT 65.685 187.565 65.855 187.735 ;
        RECT 66.145 187.565 66.315 187.735 ;
        RECT 66.605 187.565 66.775 187.735 ;
        RECT 67.065 187.565 67.235 187.735 ;
        RECT 67.525 187.565 67.695 187.735 ;
        RECT 67.985 187.565 68.155 187.735 ;
        RECT 68.445 187.565 68.615 187.735 ;
        RECT 68.905 187.565 69.075 187.735 ;
        RECT 69.365 187.565 69.535 187.735 ;
        RECT 69.825 187.565 69.995 187.735 ;
        RECT 70.285 187.565 70.455 187.735 ;
        RECT 70.745 187.565 70.915 187.735 ;
        RECT 71.205 187.565 71.375 187.735 ;
        RECT 71.665 187.565 71.835 187.735 ;
        RECT 72.125 187.565 72.295 187.735 ;
        RECT 72.585 187.565 72.755 187.735 ;
        RECT 73.045 187.565 73.215 187.735 ;
        RECT 73.505 187.565 73.675 187.735 ;
        RECT 73.965 187.565 74.135 187.735 ;
        RECT 74.425 187.565 74.595 187.735 ;
        RECT 74.885 187.565 75.055 187.735 ;
        RECT 75.345 187.565 75.515 187.735 ;
        RECT 75.805 187.565 75.975 187.735 ;
        RECT 76.265 187.565 76.435 187.735 ;
        RECT 76.725 187.565 76.895 187.735 ;
        RECT 77.185 187.565 77.355 187.735 ;
        RECT 77.645 187.565 77.815 187.735 ;
        RECT 78.105 187.565 78.275 187.735 ;
        RECT 78.565 187.565 78.735 187.735 ;
        RECT 79.025 187.565 79.195 187.735 ;
        RECT 79.485 187.565 79.655 187.735 ;
        RECT 79.945 187.565 80.115 187.735 ;
        RECT 80.405 187.565 80.575 187.735 ;
        RECT 80.865 187.565 81.035 187.735 ;
        RECT 81.325 187.565 81.495 187.735 ;
        RECT 81.785 187.565 81.955 187.735 ;
        RECT 82.245 187.565 82.415 187.735 ;
        RECT 82.705 187.565 82.875 187.735 ;
        RECT 83.165 187.565 83.335 187.735 ;
        RECT 83.625 187.565 83.795 187.735 ;
        RECT 84.085 187.565 84.255 187.735 ;
        RECT 84.545 187.565 84.715 187.735 ;
        RECT 85.005 187.565 85.175 187.735 ;
        RECT 85.465 187.565 85.635 187.735 ;
        RECT 85.925 187.565 86.095 187.735 ;
        RECT 86.385 187.565 86.555 187.735 ;
        RECT 86.845 187.565 87.015 187.735 ;
        RECT 87.305 187.565 87.475 187.735 ;
        RECT 87.765 187.565 87.935 187.735 ;
        RECT 88.225 187.565 88.395 187.735 ;
        RECT 88.685 187.565 88.855 187.735 ;
        RECT 89.145 187.565 89.315 187.735 ;
        RECT 89.605 187.565 89.775 187.735 ;
        RECT 90.065 187.565 90.235 187.735 ;
        RECT 90.525 187.565 90.695 187.735 ;
        RECT 90.985 187.565 91.155 187.735 ;
        RECT 91.445 187.565 91.615 187.735 ;
        RECT 91.905 187.565 92.075 187.735 ;
        RECT 92.365 187.565 92.535 187.735 ;
        RECT 92.825 187.565 92.995 187.735 ;
        RECT 93.285 187.565 93.455 187.735 ;
        RECT 93.745 187.565 93.915 187.735 ;
        RECT 94.205 187.565 94.375 187.735 ;
        RECT 94.665 187.565 94.835 187.735 ;
        RECT 95.125 187.565 95.295 187.735 ;
        RECT 95.585 187.565 95.755 187.735 ;
        RECT 96.045 187.565 96.215 187.735 ;
        RECT 96.505 187.565 96.675 187.735 ;
        RECT 96.965 187.565 97.135 187.735 ;
        RECT 97.425 187.565 97.595 187.735 ;
        RECT 97.885 187.565 98.055 187.735 ;
        RECT 98.345 187.565 98.515 187.735 ;
        RECT 98.805 187.565 98.975 187.735 ;
        RECT 99.265 187.565 99.435 187.735 ;
        RECT 99.725 187.565 99.895 187.735 ;
        RECT 100.185 187.565 100.355 187.735 ;
        RECT 100.645 187.565 100.815 187.735 ;
        RECT 101.105 187.565 101.275 187.735 ;
        RECT 101.565 187.565 101.735 187.735 ;
        RECT 102.025 187.565 102.195 187.735 ;
        RECT 102.485 187.565 102.655 187.735 ;
        RECT 102.945 187.565 103.115 187.735 ;
        RECT 103.405 187.565 103.575 187.735 ;
        RECT 103.865 187.565 104.035 187.735 ;
        RECT 104.325 187.565 104.495 187.735 ;
        RECT 104.785 187.565 104.955 187.735 ;
        RECT 105.245 187.565 105.415 187.735 ;
        RECT 105.705 187.565 105.875 187.735 ;
        RECT 106.165 187.565 106.335 187.735 ;
        RECT 106.625 187.565 106.795 187.735 ;
        RECT 107.085 187.565 107.255 187.735 ;
        RECT 107.545 187.565 107.715 187.735 ;
        RECT 108.005 187.565 108.175 187.735 ;
        RECT 108.465 187.565 108.635 187.735 ;
        RECT 108.925 187.565 109.095 187.735 ;
        RECT 109.385 187.565 109.555 187.735 ;
        RECT 109.845 187.565 110.015 187.735 ;
        RECT 110.305 187.565 110.475 187.735 ;
        RECT 110.765 187.565 110.935 187.735 ;
        RECT 111.225 187.565 111.395 187.735 ;
        RECT 111.685 187.565 111.855 187.735 ;
        RECT 112.145 187.565 112.315 187.735 ;
        RECT 112.605 187.565 112.775 187.735 ;
        RECT 113.065 187.565 113.235 187.735 ;
        RECT 113.525 187.565 113.695 187.735 ;
        RECT 113.985 187.565 114.155 187.735 ;
        RECT 114.445 187.565 114.615 187.735 ;
        RECT 114.905 187.565 115.075 187.735 ;
        RECT 115.365 187.565 115.535 187.735 ;
        RECT 115.825 187.565 115.995 187.735 ;
        RECT 116.285 187.565 116.455 187.735 ;
        RECT 116.745 187.565 116.915 187.735 ;
        RECT 117.205 187.565 117.375 187.735 ;
        RECT 117.665 187.565 117.835 187.735 ;
        RECT 118.125 187.565 118.295 187.735 ;
        RECT 118.585 187.565 118.755 187.735 ;
        RECT 119.045 187.565 119.215 187.735 ;
        RECT 119.505 187.565 119.675 187.735 ;
        RECT 119.965 187.565 120.135 187.735 ;
        RECT 120.425 187.565 120.595 187.735 ;
        RECT 120.885 187.565 121.055 187.735 ;
        RECT 121.345 187.565 121.515 187.735 ;
        RECT 121.805 187.565 121.975 187.735 ;
        RECT 122.265 187.565 122.435 187.735 ;
        RECT 122.725 187.565 122.895 187.735 ;
        RECT 123.185 187.565 123.355 187.735 ;
        RECT 123.645 187.565 123.815 187.735 ;
        RECT 124.105 187.565 124.275 187.735 ;
        RECT 124.565 187.565 124.735 187.735 ;
        RECT 125.025 187.565 125.195 187.735 ;
        RECT 125.485 187.565 125.655 187.735 ;
        RECT 125.945 187.565 126.115 187.735 ;
        RECT 126.405 187.565 126.575 187.735 ;
        RECT 126.865 187.565 127.035 187.735 ;
        RECT 127.325 187.565 127.495 187.735 ;
        RECT 127.785 187.565 127.955 187.735 ;
        RECT 128.245 187.565 128.415 187.735 ;
        RECT 128.705 187.565 128.875 187.735 ;
        RECT 129.165 187.565 129.335 187.735 ;
        RECT 129.625 187.565 129.795 187.735 ;
        RECT 130.085 187.565 130.255 187.735 ;
        RECT 130.545 187.565 130.715 187.735 ;
        RECT 131.005 187.565 131.175 187.735 ;
        RECT 131.465 187.565 131.635 187.735 ;
        RECT 131.925 187.565 132.095 187.735 ;
        RECT 132.385 187.565 132.555 187.735 ;
        RECT 132.845 187.565 133.015 187.735 ;
        RECT 133.305 187.565 133.475 187.735 ;
        RECT 133.765 187.565 133.935 187.735 ;
        RECT 134.225 187.565 134.395 187.735 ;
        RECT 134.685 187.565 134.855 187.735 ;
        RECT 135.145 187.565 135.315 187.735 ;
        RECT 135.605 187.565 135.775 187.735 ;
        RECT 136.065 187.565 136.235 187.735 ;
        RECT 136.525 187.565 136.695 187.735 ;
        RECT 136.985 187.565 137.155 187.735 ;
        RECT 137.445 187.565 137.615 187.735 ;
        RECT 137.905 187.565 138.075 187.735 ;
        RECT 138.365 187.565 138.535 187.735 ;
        RECT 138.825 187.565 138.995 187.735 ;
        RECT 139.285 187.565 139.455 187.735 ;
        RECT 139.745 187.565 139.915 187.735 ;
        RECT 140.205 187.565 140.375 187.735 ;
        RECT 140.665 187.565 140.835 187.735 ;
        RECT 141.125 187.565 141.295 187.735 ;
        RECT 141.585 187.565 141.755 187.735 ;
        RECT 142.045 187.565 142.215 187.735 ;
        RECT 142.505 187.565 142.675 187.735 ;
        RECT 142.965 187.565 143.135 187.735 ;
        RECT 143.425 187.565 143.595 187.735 ;
        RECT 143.885 187.565 144.055 187.735 ;
        RECT 144.345 187.565 144.515 187.735 ;
        RECT 144.805 187.565 144.975 187.735 ;
        RECT 145.265 187.565 145.435 187.735 ;
        RECT 145.725 187.565 145.895 187.735 ;
        RECT 146.185 187.565 146.355 187.735 ;
        RECT 146.645 187.565 146.815 187.735 ;
        RECT 147.105 187.565 147.275 187.735 ;
        RECT 147.565 187.565 147.735 187.735 ;
        RECT 148.025 187.565 148.195 187.735 ;
        RECT 148.485 187.565 148.655 187.735 ;
        RECT 148.945 187.565 149.115 187.735 ;
        RECT 149.405 187.565 149.575 187.735 ;
        RECT 149.865 187.565 150.035 187.735 ;
        RECT 45.905 187.055 46.075 187.225 ;
        RECT 47.285 186.715 47.455 186.885 ;
        RECT 46.825 186.035 46.995 186.205 ;
        RECT 47.745 186.035 47.915 186.205 ;
        RECT 48.205 186.035 48.375 186.205 ;
        RECT 49.585 187.055 49.755 187.225 ;
        RECT 50.505 187.055 50.675 187.225 ;
        RECT 50.505 186.035 50.675 186.205 ;
        RECT 50.965 186.035 51.135 186.205 ;
        RECT 51.885 185.695 52.055 185.865 ;
        RECT 58.325 186.035 58.495 186.205 ;
        RECT 58.785 186.035 58.955 186.205 ;
        RECT 59.245 186.375 59.415 186.545 ;
        RECT 60.625 186.715 60.795 186.885 ;
        RECT 62.925 187.055 63.095 187.225 ;
        RECT 62.465 186.715 62.635 186.885 ;
        RECT 59.705 186.035 59.875 186.205 ;
        RECT 61.085 186.375 61.255 186.545 ;
        RECT 62.005 186.375 62.175 186.545 ;
        RECT 64.305 187.055 64.475 187.225 ;
        RECT 62.005 185.695 62.175 185.865 ;
        RECT 63.385 185.695 63.555 185.865 ;
        RECT 63.845 185.695 64.015 185.865 ;
        RECT 65.225 187.055 65.395 187.225 ;
        RECT 67.525 187.055 67.695 187.225 ;
        RECT 65.685 186.035 65.855 186.205 ;
        RECT 66.605 186.715 66.775 186.885 ;
        RECT 67.065 186.375 67.235 186.545 ;
        RECT 67.525 185.355 67.695 185.525 ;
        RECT 68.445 185.355 68.615 185.525 ;
        RECT 74.425 186.715 74.595 186.885 ;
        RECT 73.060 185.925 73.230 186.095 ;
        RECT 73.505 186.035 73.675 186.205 ;
        RECT 75.830 186.715 76.000 186.885 ;
        RECT 75.345 186.035 75.515 186.205 ;
        RECT 74.425 185.695 74.595 185.865 ;
        RECT 76.225 186.375 76.395 186.545 ;
        RECT 76.625 186.035 76.795 186.205 ;
        RECT 77.930 186.715 78.100 186.885 ;
        RECT 77.415 186.375 77.585 186.545 ;
        RECT 79.500 186.715 79.670 186.885 ;
        RECT 79.935 186.375 80.105 186.545 ;
        RECT 82.245 185.355 82.415 185.525 ;
        RECT 88.685 186.035 88.855 186.205 ;
        RECT 87.765 185.355 87.935 185.525 ;
        RECT 94.665 186.035 94.835 186.205 ;
        RECT 96.045 186.375 96.215 186.545 ;
        RECT 101.105 186.375 101.275 186.545 ;
        RECT 102.255 186.715 102.425 186.885 ;
        RECT 108.465 186.035 108.635 186.205 ;
        RECT 109.845 186.375 110.015 186.545 ;
        RECT 110.305 186.035 110.475 186.205 ;
        RECT 111.685 186.375 111.855 186.545 ;
        RECT 117.205 187.055 117.375 187.225 ;
        RECT 120.425 187.055 120.595 187.225 ;
        RECT 115.365 186.035 115.535 186.205 ;
        RECT 116.285 186.035 116.455 186.205 ;
        RECT 117.205 186.035 117.375 186.205 ;
        RECT 119.045 186.035 119.215 186.205 ;
        RECT 121.345 185.355 121.515 185.525 ;
        RECT 121.805 185.355 121.975 185.525 ;
        RECT 122.265 185.355 122.435 185.525 ;
        RECT 123.185 185.695 123.355 185.865 ;
        RECT 124.565 186.035 124.735 186.205 ;
        RECT 127.785 187.055 127.955 187.225 ;
        RECT 128.705 187.055 128.875 187.225 ;
        RECT 125.485 185.355 125.655 185.525 ;
        RECT 126.865 185.695 127.035 185.865 ;
        RECT 127.865 185.355 128.035 185.525 ;
        RECT 132.385 187.055 132.555 187.225 ;
        RECT 129.165 186.375 129.335 186.545 ;
        RECT 131.005 186.375 131.175 186.545 ;
        RECT 130.085 186.035 130.255 186.205 ;
        RECT 133.305 186.715 133.475 186.885 ;
        RECT 131.465 185.695 131.635 185.865 ;
        RECT 132.615 185.865 132.785 186.035 ;
        RECT 133.765 185.915 133.935 186.085 ;
        RECT 134.685 185.355 134.855 185.525 ;
        RECT 138.365 186.035 138.535 186.205 ;
        RECT 138.825 186.035 138.995 186.205 ;
        RECT 139.285 187.055 139.455 187.225 ;
        RECT 139.745 186.375 139.915 186.545 ;
        RECT 142.045 187.055 142.215 187.225 ;
        RECT 140.495 186.035 140.665 186.205 ;
        RECT 141.125 186.035 141.295 186.205 ;
        RECT 142.505 186.035 142.675 186.205 ;
        RECT 144.805 186.375 144.975 186.545 ;
        RECT 142.965 186.035 143.135 186.205 ;
        RECT 143.425 186.035 143.595 186.205 ;
        RECT 136.985 185.355 137.155 185.525 ;
        RECT 146.185 187.055 146.355 187.225 ;
        RECT 145.265 186.715 145.435 186.885 ;
        RECT 146.055 185.355 146.225 185.525 ;
        RECT 147.105 185.695 147.275 185.865 ;
        RECT 36.245 184.845 36.415 185.015 ;
        RECT 36.705 184.845 36.875 185.015 ;
        RECT 37.165 184.845 37.335 185.015 ;
        RECT 37.625 184.845 37.795 185.015 ;
        RECT 38.085 184.845 38.255 185.015 ;
        RECT 38.545 184.845 38.715 185.015 ;
        RECT 39.005 184.845 39.175 185.015 ;
        RECT 39.465 184.845 39.635 185.015 ;
        RECT 39.925 184.845 40.095 185.015 ;
        RECT 40.385 184.845 40.555 185.015 ;
        RECT 40.845 184.845 41.015 185.015 ;
        RECT 41.305 184.845 41.475 185.015 ;
        RECT 41.765 184.845 41.935 185.015 ;
        RECT 42.225 184.845 42.395 185.015 ;
        RECT 42.685 184.845 42.855 185.015 ;
        RECT 43.145 184.845 43.315 185.015 ;
        RECT 43.605 184.845 43.775 185.015 ;
        RECT 44.065 184.845 44.235 185.015 ;
        RECT 44.525 184.845 44.695 185.015 ;
        RECT 44.985 184.845 45.155 185.015 ;
        RECT 45.445 184.845 45.615 185.015 ;
        RECT 45.905 184.845 46.075 185.015 ;
        RECT 46.365 184.845 46.535 185.015 ;
        RECT 46.825 184.845 46.995 185.015 ;
        RECT 47.285 184.845 47.455 185.015 ;
        RECT 47.745 184.845 47.915 185.015 ;
        RECT 48.205 184.845 48.375 185.015 ;
        RECT 48.665 184.845 48.835 185.015 ;
        RECT 49.125 184.845 49.295 185.015 ;
        RECT 49.585 184.845 49.755 185.015 ;
        RECT 50.045 184.845 50.215 185.015 ;
        RECT 50.505 184.845 50.675 185.015 ;
        RECT 50.965 184.845 51.135 185.015 ;
        RECT 51.425 184.845 51.595 185.015 ;
        RECT 51.885 184.845 52.055 185.015 ;
        RECT 52.345 184.845 52.515 185.015 ;
        RECT 52.805 184.845 52.975 185.015 ;
        RECT 53.265 184.845 53.435 185.015 ;
        RECT 53.725 184.845 53.895 185.015 ;
        RECT 54.185 184.845 54.355 185.015 ;
        RECT 54.645 184.845 54.815 185.015 ;
        RECT 55.105 184.845 55.275 185.015 ;
        RECT 55.565 184.845 55.735 185.015 ;
        RECT 56.025 184.845 56.195 185.015 ;
        RECT 56.485 184.845 56.655 185.015 ;
        RECT 56.945 184.845 57.115 185.015 ;
        RECT 57.405 184.845 57.575 185.015 ;
        RECT 57.865 184.845 58.035 185.015 ;
        RECT 58.325 184.845 58.495 185.015 ;
        RECT 58.785 184.845 58.955 185.015 ;
        RECT 59.245 184.845 59.415 185.015 ;
        RECT 59.705 184.845 59.875 185.015 ;
        RECT 60.165 184.845 60.335 185.015 ;
        RECT 60.625 184.845 60.795 185.015 ;
        RECT 61.085 184.845 61.255 185.015 ;
        RECT 61.545 184.845 61.715 185.015 ;
        RECT 62.005 184.845 62.175 185.015 ;
        RECT 62.465 184.845 62.635 185.015 ;
        RECT 62.925 184.845 63.095 185.015 ;
        RECT 63.385 184.845 63.555 185.015 ;
        RECT 63.845 184.845 64.015 185.015 ;
        RECT 64.305 184.845 64.475 185.015 ;
        RECT 64.765 184.845 64.935 185.015 ;
        RECT 65.225 184.845 65.395 185.015 ;
        RECT 65.685 184.845 65.855 185.015 ;
        RECT 66.145 184.845 66.315 185.015 ;
        RECT 66.605 184.845 66.775 185.015 ;
        RECT 67.065 184.845 67.235 185.015 ;
        RECT 67.525 184.845 67.695 185.015 ;
        RECT 67.985 184.845 68.155 185.015 ;
        RECT 68.445 184.845 68.615 185.015 ;
        RECT 68.905 184.845 69.075 185.015 ;
        RECT 69.365 184.845 69.535 185.015 ;
        RECT 69.825 184.845 69.995 185.015 ;
        RECT 70.285 184.845 70.455 185.015 ;
        RECT 70.745 184.845 70.915 185.015 ;
        RECT 71.205 184.845 71.375 185.015 ;
        RECT 71.665 184.845 71.835 185.015 ;
        RECT 72.125 184.845 72.295 185.015 ;
        RECT 72.585 184.845 72.755 185.015 ;
        RECT 73.045 184.845 73.215 185.015 ;
        RECT 73.505 184.845 73.675 185.015 ;
        RECT 73.965 184.845 74.135 185.015 ;
        RECT 74.425 184.845 74.595 185.015 ;
        RECT 74.885 184.845 75.055 185.015 ;
        RECT 75.345 184.845 75.515 185.015 ;
        RECT 75.805 184.845 75.975 185.015 ;
        RECT 76.265 184.845 76.435 185.015 ;
        RECT 76.725 184.845 76.895 185.015 ;
        RECT 77.185 184.845 77.355 185.015 ;
        RECT 77.645 184.845 77.815 185.015 ;
        RECT 78.105 184.845 78.275 185.015 ;
        RECT 78.565 184.845 78.735 185.015 ;
        RECT 79.025 184.845 79.195 185.015 ;
        RECT 79.485 184.845 79.655 185.015 ;
        RECT 79.945 184.845 80.115 185.015 ;
        RECT 80.405 184.845 80.575 185.015 ;
        RECT 80.865 184.845 81.035 185.015 ;
        RECT 81.325 184.845 81.495 185.015 ;
        RECT 81.785 184.845 81.955 185.015 ;
        RECT 82.245 184.845 82.415 185.015 ;
        RECT 82.705 184.845 82.875 185.015 ;
        RECT 83.165 184.845 83.335 185.015 ;
        RECT 83.625 184.845 83.795 185.015 ;
        RECT 84.085 184.845 84.255 185.015 ;
        RECT 84.545 184.845 84.715 185.015 ;
        RECT 85.005 184.845 85.175 185.015 ;
        RECT 85.465 184.845 85.635 185.015 ;
        RECT 85.925 184.845 86.095 185.015 ;
        RECT 86.385 184.845 86.555 185.015 ;
        RECT 86.845 184.845 87.015 185.015 ;
        RECT 87.305 184.845 87.475 185.015 ;
        RECT 87.765 184.845 87.935 185.015 ;
        RECT 88.225 184.845 88.395 185.015 ;
        RECT 88.685 184.845 88.855 185.015 ;
        RECT 89.145 184.845 89.315 185.015 ;
        RECT 89.605 184.845 89.775 185.015 ;
        RECT 90.065 184.845 90.235 185.015 ;
        RECT 90.525 184.845 90.695 185.015 ;
        RECT 90.985 184.845 91.155 185.015 ;
        RECT 91.445 184.845 91.615 185.015 ;
        RECT 91.905 184.845 92.075 185.015 ;
        RECT 92.365 184.845 92.535 185.015 ;
        RECT 92.825 184.845 92.995 185.015 ;
        RECT 93.285 184.845 93.455 185.015 ;
        RECT 93.745 184.845 93.915 185.015 ;
        RECT 94.205 184.845 94.375 185.015 ;
        RECT 94.665 184.845 94.835 185.015 ;
        RECT 95.125 184.845 95.295 185.015 ;
        RECT 95.585 184.845 95.755 185.015 ;
        RECT 96.045 184.845 96.215 185.015 ;
        RECT 96.505 184.845 96.675 185.015 ;
        RECT 96.965 184.845 97.135 185.015 ;
        RECT 97.425 184.845 97.595 185.015 ;
        RECT 97.885 184.845 98.055 185.015 ;
        RECT 98.345 184.845 98.515 185.015 ;
        RECT 98.805 184.845 98.975 185.015 ;
        RECT 99.265 184.845 99.435 185.015 ;
        RECT 99.725 184.845 99.895 185.015 ;
        RECT 100.185 184.845 100.355 185.015 ;
        RECT 100.645 184.845 100.815 185.015 ;
        RECT 101.105 184.845 101.275 185.015 ;
        RECT 101.565 184.845 101.735 185.015 ;
        RECT 102.025 184.845 102.195 185.015 ;
        RECT 102.485 184.845 102.655 185.015 ;
        RECT 102.945 184.845 103.115 185.015 ;
        RECT 103.405 184.845 103.575 185.015 ;
        RECT 103.865 184.845 104.035 185.015 ;
        RECT 104.325 184.845 104.495 185.015 ;
        RECT 104.785 184.845 104.955 185.015 ;
        RECT 105.245 184.845 105.415 185.015 ;
        RECT 105.705 184.845 105.875 185.015 ;
        RECT 106.165 184.845 106.335 185.015 ;
        RECT 106.625 184.845 106.795 185.015 ;
        RECT 107.085 184.845 107.255 185.015 ;
        RECT 107.545 184.845 107.715 185.015 ;
        RECT 108.005 184.845 108.175 185.015 ;
        RECT 108.465 184.845 108.635 185.015 ;
        RECT 108.925 184.845 109.095 185.015 ;
        RECT 109.385 184.845 109.555 185.015 ;
        RECT 109.845 184.845 110.015 185.015 ;
        RECT 110.305 184.845 110.475 185.015 ;
        RECT 110.765 184.845 110.935 185.015 ;
        RECT 111.225 184.845 111.395 185.015 ;
        RECT 111.685 184.845 111.855 185.015 ;
        RECT 112.145 184.845 112.315 185.015 ;
        RECT 112.605 184.845 112.775 185.015 ;
        RECT 113.065 184.845 113.235 185.015 ;
        RECT 113.525 184.845 113.695 185.015 ;
        RECT 113.985 184.845 114.155 185.015 ;
        RECT 114.445 184.845 114.615 185.015 ;
        RECT 114.905 184.845 115.075 185.015 ;
        RECT 115.365 184.845 115.535 185.015 ;
        RECT 115.825 184.845 115.995 185.015 ;
        RECT 116.285 184.845 116.455 185.015 ;
        RECT 116.745 184.845 116.915 185.015 ;
        RECT 117.205 184.845 117.375 185.015 ;
        RECT 117.665 184.845 117.835 185.015 ;
        RECT 118.125 184.845 118.295 185.015 ;
        RECT 118.585 184.845 118.755 185.015 ;
        RECT 119.045 184.845 119.215 185.015 ;
        RECT 119.505 184.845 119.675 185.015 ;
        RECT 119.965 184.845 120.135 185.015 ;
        RECT 120.425 184.845 120.595 185.015 ;
        RECT 120.885 184.845 121.055 185.015 ;
        RECT 121.345 184.845 121.515 185.015 ;
        RECT 121.805 184.845 121.975 185.015 ;
        RECT 122.265 184.845 122.435 185.015 ;
        RECT 122.725 184.845 122.895 185.015 ;
        RECT 123.185 184.845 123.355 185.015 ;
        RECT 123.645 184.845 123.815 185.015 ;
        RECT 124.105 184.845 124.275 185.015 ;
        RECT 124.565 184.845 124.735 185.015 ;
        RECT 125.025 184.845 125.195 185.015 ;
        RECT 125.485 184.845 125.655 185.015 ;
        RECT 125.945 184.845 126.115 185.015 ;
        RECT 126.405 184.845 126.575 185.015 ;
        RECT 126.865 184.845 127.035 185.015 ;
        RECT 127.325 184.845 127.495 185.015 ;
        RECT 127.785 184.845 127.955 185.015 ;
        RECT 128.245 184.845 128.415 185.015 ;
        RECT 128.705 184.845 128.875 185.015 ;
        RECT 129.165 184.845 129.335 185.015 ;
        RECT 129.625 184.845 129.795 185.015 ;
        RECT 130.085 184.845 130.255 185.015 ;
        RECT 130.545 184.845 130.715 185.015 ;
        RECT 131.005 184.845 131.175 185.015 ;
        RECT 131.465 184.845 131.635 185.015 ;
        RECT 131.925 184.845 132.095 185.015 ;
        RECT 132.385 184.845 132.555 185.015 ;
        RECT 132.845 184.845 133.015 185.015 ;
        RECT 133.305 184.845 133.475 185.015 ;
        RECT 133.765 184.845 133.935 185.015 ;
        RECT 134.225 184.845 134.395 185.015 ;
        RECT 134.685 184.845 134.855 185.015 ;
        RECT 135.145 184.845 135.315 185.015 ;
        RECT 135.605 184.845 135.775 185.015 ;
        RECT 136.065 184.845 136.235 185.015 ;
        RECT 136.525 184.845 136.695 185.015 ;
        RECT 136.985 184.845 137.155 185.015 ;
        RECT 137.445 184.845 137.615 185.015 ;
        RECT 137.905 184.845 138.075 185.015 ;
        RECT 138.365 184.845 138.535 185.015 ;
        RECT 138.825 184.845 138.995 185.015 ;
        RECT 139.285 184.845 139.455 185.015 ;
        RECT 139.745 184.845 139.915 185.015 ;
        RECT 140.205 184.845 140.375 185.015 ;
        RECT 140.665 184.845 140.835 185.015 ;
        RECT 141.125 184.845 141.295 185.015 ;
        RECT 141.585 184.845 141.755 185.015 ;
        RECT 142.045 184.845 142.215 185.015 ;
        RECT 142.505 184.845 142.675 185.015 ;
        RECT 142.965 184.845 143.135 185.015 ;
        RECT 143.425 184.845 143.595 185.015 ;
        RECT 143.885 184.845 144.055 185.015 ;
        RECT 144.345 184.845 144.515 185.015 ;
        RECT 144.805 184.845 144.975 185.015 ;
        RECT 145.265 184.845 145.435 185.015 ;
        RECT 145.725 184.845 145.895 185.015 ;
        RECT 146.185 184.845 146.355 185.015 ;
        RECT 146.645 184.845 146.815 185.015 ;
        RECT 147.105 184.845 147.275 185.015 ;
        RECT 147.565 184.845 147.735 185.015 ;
        RECT 148.025 184.845 148.195 185.015 ;
        RECT 148.485 184.845 148.655 185.015 ;
        RECT 148.945 184.845 149.115 185.015 ;
        RECT 149.405 184.845 149.575 185.015 ;
        RECT 149.865 184.845 150.035 185.015 ;
        RECT 44.525 184.335 44.695 184.505 ;
        RECT 43.145 183.655 43.315 183.825 ;
        RECT 44.065 183.655 44.235 183.825 ;
        RECT 44.525 183.655 44.695 183.825 ;
        RECT 44.985 183.655 45.155 183.825 ;
        RECT 45.905 183.655 46.075 183.825 ;
        RECT 46.825 183.315 46.995 183.485 ;
        RECT 52.805 184.335 52.975 184.505 ;
        RECT 48.205 183.655 48.375 183.825 ;
        RECT 48.665 183.655 48.835 183.825 ;
        RECT 49.585 183.655 49.755 183.825 ;
        RECT 50.965 183.655 51.135 183.825 ;
        RECT 47.285 182.635 47.455 182.805 ;
        RECT 51.425 183.315 51.595 183.485 ;
        RECT 53.265 183.655 53.435 183.825 ;
        RECT 53.725 183.655 53.895 183.825 ;
        RECT 49.125 182.635 49.295 182.805 ;
        RECT 51.885 182.635 52.055 182.805 ;
        RECT 60.165 184.335 60.335 184.505 ;
        RECT 58.325 183.655 58.495 183.825 ;
        RECT 59.245 183.655 59.415 183.825 ;
        RECT 53.265 182.635 53.435 182.805 ;
        RECT 55.105 182.975 55.275 183.145 ;
        RECT 64.305 183.655 64.475 183.825 ;
        RECT 63.385 182.635 63.555 182.805 ;
        RECT 77.645 183.655 77.815 183.825 ;
        RECT 78.565 182.635 78.735 182.805 ;
        RECT 79.025 184.335 79.195 184.505 ;
        RECT 80.865 184.335 81.035 184.505 ;
        RECT 79.945 183.655 80.115 183.825 ;
        RECT 81.325 183.655 81.495 183.825 ;
        RECT 82.705 183.655 82.875 183.825 ;
        RECT 81.785 183.315 81.955 183.485 ;
        RECT 83.625 183.315 83.795 183.485 ;
        RECT 85.005 183.655 85.175 183.825 ;
        RECT 84.545 182.975 84.715 183.145 ;
        RECT 88.225 183.655 88.395 183.825 ;
        RECT 89.145 183.655 89.315 183.825 ;
        RECT 89.605 183.655 89.775 183.825 ;
        RECT 90.065 183.655 90.235 183.825 ;
        RECT 91.445 182.635 91.615 182.805 ;
        RECT 91.905 183.995 92.075 184.165 ;
        RECT 92.825 183.655 92.995 183.825 ;
        RECT 94.665 183.655 94.835 183.825 ;
        RECT 94.205 182.635 94.375 182.805 ;
        RECT 96.045 183.655 96.215 183.825 ;
        RECT 96.505 183.655 96.675 183.825 ;
        RECT 100.185 184.335 100.355 184.505 ;
        RECT 97.425 183.655 97.595 183.825 ;
        RECT 97.885 183.655 98.055 183.825 ;
        RECT 95.125 182.635 95.295 182.805 ;
        RECT 99.265 183.655 99.435 183.825 ;
        RECT 101.565 183.655 101.735 183.825 ;
        RECT 102.255 183.655 102.425 183.825 ;
        RECT 100.645 182.635 100.815 182.805 ;
        RECT 102.975 183.655 103.145 183.825 ;
        RECT 103.465 183.665 103.635 183.835 ;
        RECT 104.325 183.655 104.495 183.825 ;
        RECT 105.705 183.655 105.875 183.825 ;
        RECT 107.085 183.655 107.255 183.825 ;
        RECT 108.005 183.655 108.175 183.825 ;
        RECT 104.785 182.635 104.955 182.805 ;
        RECT 107.545 182.635 107.715 182.805 ;
        RECT 108.465 183.315 108.635 183.485 ;
        RECT 109.845 183.655 110.015 183.825 ;
        RECT 114.445 183.995 114.615 184.165 ;
        RECT 117.205 183.575 117.375 183.745 ;
        RECT 114.905 182.635 115.075 182.805 ;
        RECT 118.585 183.655 118.755 183.825 ;
        RECT 118.125 182.975 118.295 183.145 ;
        RECT 121.805 183.995 121.975 184.165 ;
        RECT 120.425 182.635 120.595 182.805 ;
        RECT 123.645 184.335 123.815 184.505 ;
        RECT 122.805 183.995 122.975 184.165 ;
        RECT 125.025 183.655 125.195 183.825 ;
        RECT 121.345 182.635 121.515 182.805 ;
        RECT 122.725 182.635 122.895 182.805 ;
        RECT 125.945 182.975 126.115 183.145 ;
        RECT 127.325 183.655 127.495 183.825 ;
        RECT 128.245 182.975 128.415 183.145 ;
        RECT 129.625 183.655 129.795 183.825 ;
        RECT 131.465 183.655 131.635 183.825 ;
        RECT 132.385 183.655 132.555 183.825 ;
        RECT 132.845 183.655 133.015 183.825 ;
        RECT 134.225 184.335 134.395 184.505 ;
        RECT 128.705 182.975 128.875 183.145 ;
        RECT 132.385 182.635 132.555 182.805 ;
        RECT 133.305 182.975 133.475 183.145 ;
        RECT 142.505 184.335 142.675 184.505 ;
        RECT 135.145 183.655 135.315 183.825 ;
        RECT 140.140 183.655 140.310 183.825 ;
        RECT 140.665 182.975 140.835 183.145 ;
        RECT 141.585 183.655 141.755 183.825 ;
        RECT 141.125 182.975 141.295 183.145 ;
        RECT 143.885 183.655 144.055 183.825 ;
        RECT 142.965 182.975 143.135 183.145 ;
        RECT 36.245 182.125 36.415 182.295 ;
        RECT 36.705 182.125 36.875 182.295 ;
        RECT 37.165 182.125 37.335 182.295 ;
        RECT 37.625 182.125 37.795 182.295 ;
        RECT 38.085 182.125 38.255 182.295 ;
        RECT 38.545 182.125 38.715 182.295 ;
        RECT 39.005 182.125 39.175 182.295 ;
        RECT 39.465 182.125 39.635 182.295 ;
        RECT 39.925 182.125 40.095 182.295 ;
        RECT 40.385 182.125 40.555 182.295 ;
        RECT 40.845 182.125 41.015 182.295 ;
        RECT 41.305 182.125 41.475 182.295 ;
        RECT 41.765 182.125 41.935 182.295 ;
        RECT 42.225 182.125 42.395 182.295 ;
        RECT 42.685 182.125 42.855 182.295 ;
        RECT 43.145 182.125 43.315 182.295 ;
        RECT 43.605 182.125 43.775 182.295 ;
        RECT 44.065 182.125 44.235 182.295 ;
        RECT 44.525 182.125 44.695 182.295 ;
        RECT 44.985 182.125 45.155 182.295 ;
        RECT 45.445 182.125 45.615 182.295 ;
        RECT 45.905 182.125 46.075 182.295 ;
        RECT 46.365 182.125 46.535 182.295 ;
        RECT 46.825 182.125 46.995 182.295 ;
        RECT 47.285 182.125 47.455 182.295 ;
        RECT 47.745 182.125 47.915 182.295 ;
        RECT 48.205 182.125 48.375 182.295 ;
        RECT 48.665 182.125 48.835 182.295 ;
        RECT 49.125 182.125 49.295 182.295 ;
        RECT 49.585 182.125 49.755 182.295 ;
        RECT 50.045 182.125 50.215 182.295 ;
        RECT 50.505 182.125 50.675 182.295 ;
        RECT 50.965 182.125 51.135 182.295 ;
        RECT 51.425 182.125 51.595 182.295 ;
        RECT 51.885 182.125 52.055 182.295 ;
        RECT 52.345 182.125 52.515 182.295 ;
        RECT 52.805 182.125 52.975 182.295 ;
        RECT 53.265 182.125 53.435 182.295 ;
        RECT 53.725 182.125 53.895 182.295 ;
        RECT 54.185 182.125 54.355 182.295 ;
        RECT 54.645 182.125 54.815 182.295 ;
        RECT 55.105 182.125 55.275 182.295 ;
        RECT 55.565 182.125 55.735 182.295 ;
        RECT 56.025 182.125 56.195 182.295 ;
        RECT 56.485 182.125 56.655 182.295 ;
        RECT 56.945 182.125 57.115 182.295 ;
        RECT 57.405 182.125 57.575 182.295 ;
        RECT 57.865 182.125 58.035 182.295 ;
        RECT 58.325 182.125 58.495 182.295 ;
        RECT 58.785 182.125 58.955 182.295 ;
        RECT 59.245 182.125 59.415 182.295 ;
        RECT 59.705 182.125 59.875 182.295 ;
        RECT 60.165 182.125 60.335 182.295 ;
        RECT 60.625 182.125 60.795 182.295 ;
        RECT 61.085 182.125 61.255 182.295 ;
        RECT 61.545 182.125 61.715 182.295 ;
        RECT 62.005 182.125 62.175 182.295 ;
        RECT 62.465 182.125 62.635 182.295 ;
        RECT 62.925 182.125 63.095 182.295 ;
        RECT 63.385 182.125 63.555 182.295 ;
        RECT 63.845 182.125 64.015 182.295 ;
        RECT 64.305 182.125 64.475 182.295 ;
        RECT 64.765 182.125 64.935 182.295 ;
        RECT 65.225 182.125 65.395 182.295 ;
        RECT 65.685 182.125 65.855 182.295 ;
        RECT 66.145 182.125 66.315 182.295 ;
        RECT 66.605 182.125 66.775 182.295 ;
        RECT 67.065 182.125 67.235 182.295 ;
        RECT 67.525 182.125 67.695 182.295 ;
        RECT 67.985 182.125 68.155 182.295 ;
        RECT 68.445 182.125 68.615 182.295 ;
        RECT 68.905 182.125 69.075 182.295 ;
        RECT 69.365 182.125 69.535 182.295 ;
        RECT 69.825 182.125 69.995 182.295 ;
        RECT 70.285 182.125 70.455 182.295 ;
        RECT 70.745 182.125 70.915 182.295 ;
        RECT 71.205 182.125 71.375 182.295 ;
        RECT 71.665 182.125 71.835 182.295 ;
        RECT 72.125 182.125 72.295 182.295 ;
        RECT 72.585 182.125 72.755 182.295 ;
        RECT 73.045 182.125 73.215 182.295 ;
        RECT 73.505 182.125 73.675 182.295 ;
        RECT 73.965 182.125 74.135 182.295 ;
        RECT 74.425 182.125 74.595 182.295 ;
        RECT 74.885 182.125 75.055 182.295 ;
        RECT 75.345 182.125 75.515 182.295 ;
        RECT 75.805 182.125 75.975 182.295 ;
        RECT 76.265 182.125 76.435 182.295 ;
        RECT 76.725 182.125 76.895 182.295 ;
        RECT 77.185 182.125 77.355 182.295 ;
        RECT 77.645 182.125 77.815 182.295 ;
        RECT 78.105 182.125 78.275 182.295 ;
        RECT 78.565 182.125 78.735 182.295 ;
        RECT 79.025 182.125 79.195 182.295 ;
        RECT 79.485 182.125 79.655 182.295 ;
        RECT 79.945 182.125 80.115 182.295 ;
        RECT 80.405 182.125 80.575 182.295 ;
        RECT 80.865 182.125 81.035 182.295 ;
        RECT 81.325 182.125 81.495 182.295 ;
        RECT 81.785 182.125 81.955 182.295 ;
        RECT 82.245 182.125 82.415 182.295 ;
        RECT 82.705 182.125 82.875 182.295 ;
        RECT 83.165 182.125 83.335 182.295 ;
        RECT 83.625 182.125 83.795 182.295 ;
        RECT 84.085 182.125 84.255 182.295 ;
        RECT 84.545 182.125 84.715 182.295 ;
        RECT 85.005 182.125 85.175 182.295 ;
        RECT 85.465 182.125 85.635 182.295 ;
        RECT 85.925 182.125 86.095 182.295 ;
        RECT 86.385 182.125 86.555 182.295 ;
        RECT 86.845 182.125 87.015 182.295 ;
        RECT 87.305 182.125 87.475 182.295 ;
        RECT 87.765 182.125 87.935 182.295 ;
        RECT 88.225 182.125 88.395 182.295 ;
        RECT 88.685 182.125 88.855 182.295 ;
        RECT 89.145 182.125 89.315 182.295 ;
        RECT 89.605 182.125 89.775 182.295 ;
        RECT 90.065 182.125 90.235 182.295 ;
        RECT 90.525 182.125 90.695 182.295 ;
        RECT 90.985 182.125 91.155 182.295 ;
        RECT 91.445 182.125 91.615 182.295 ;
        RECT 91.905 182.125 92.075 182.295 ;
        RECT 92.365 182.125 92.535 182.295 ;
        RECT 92.825 182.125 92.995 182.295 ;
        RECT 93.285 182.125 93.455 182.295 ;
        RECT 93.745 182.125 93.915 182.295 ;
        RECT 94.205 182.125 94.375 182.295 ;
        RECT 94.665 182.125 94.835 182.295 ;
        RECT 95.125 182.125 95.295 182.295 ;
        RECT 95.585 182.125 95.755 182.295 ;
        RECT 96.045 182.125 96.215 182.295 ;
        RECT 96.505 182.125 96.675 182.295 ;
        RECT 96.965 182.125 97.135 182.295 ;
        RECT 97.425 182.125 97.595 182.295 ;
        RECT 97.885 182.125 98.055 182.295 ;
        RECT 98.345 182.125 98.515 182.295 ;
        RECT 98.805 182.125 98.975 182.295 ;
        RECT 99.265 182.125 99.435 182.295 ;
        RECT 99.725 182.125 99.895 182.295 ;
        RECT 100.185 182.125 100.355 182.295 ;
        RECT 100.645 182.125 100.815 182.295 ;
        RECT 101.105 182.125 101.275 182.295 ;
        RECT 101.565 182.125 101.735 182.295 ;
        RECT 102.025 182.125 102.195 182.295 ;
        RECT 102.485 182.125 102.655 182.295 ;
        RECT 102.945 182.125 103.115 182.295 ;
        RECT 103.405 182.125 103.575 182.295 ;
        RECT 103.865 182.125 104.035 182.295 ;
        RECT 104.325 182.125 104.495 182.295 ;
        RECT 104.785 182.125 104.955 182.295 ;
        RECT 105.245 182.125 105.415 182.295 ;
        RECT 105.705 182.125 105.875 182.295 ;
        RECT 106.165 182.125 106.335 182.295 ;
        RECT 106.625 182.125 106.795 182.295 ;
        RECT 107.085 182.125 107.255 182.295 ;
        RECT 107.545 182.125 107.715 182.295 ;
        RECT 108.005 182.125 108.175 182.295 ;
        RECT 108.465 182.125 108.635 182.295 ;
        RECT 108.925 182.125 109.095 182.295 ;
        RECT 109.385 182.125 109.555 182.295 ;
        RECT 109.845 182.125 110.015 182.295 ;
        RECT 110.305 182.125 110.475 182.295 ;
        RECT 110.765 182.125 110.935 182.295 ;
        RECT 111.225 182.125 111.395 182.295 ;
        RECT 111.685 182.125 111.855 182.295 ;
        RECT 112.145 182.125 112.315 182.295 ;
        RECT 112.605 182.125 112.775 182.295 ;
        RECT 113.065 182.125 113.235 182.295 ;
        RECT 113.525 182.125 113.695 182.295 ;
        RECT 113.985 182.125 114.155 182.295 ;
        RECT 114.445 182.125 114.615 182.295 ;
        RECT 114.905 182.125 115.075 182.295 ;
        RECT 115.365 182.125 115.535 182.295 ;
        RECT 115.825 182.125 115.995 182.295 ;
        RECT 116.285 182.125 116.455 182.295 ;
        RECT 116.745 182.125 116.915 182.295 ;
        RECT 117.205 182.125 117.375 182.295 ;
        RECT 117.665 182.125 117.835 182.295 ;
        RECT 118.125 182.125 118.295 182.295 ;
        RECT 118.585 182.125 118.755 182.295 ;
        RECT 119.045 182.125 119.215 182.295 ;
        RECT 119.505 182.125 119.675 182.295 ;
        RECT 119.965 182.125 120.135 182.295 ;
        RECT 120.425 182.125 120.595 182.295 ;
        RECT 120.885 182.125 121.055 182.295 ;
        RECT 121.345 182.125 121.515 182.295 ;
        RECT 121.805 182.125 121.975 182.295 ;
        RECT 122.265 182.125 122.435 182.295 ;
        RECT 122.725 182.125 122.895 182.295 ;
        RECT 123.185 182.125 123.355 182.295 ;
        RECT 123.645 182.125 123.815 182.295 ;
        RECT 124.105 182.125 124.275 182.295 ;
        RECT 124.565 182.125 124.735 182.295 ;
        RECT 125.025 182.125 125.195 182.295 ;
        RECT 125.485 182.125 125.655 182.295 ;
        RECT 125.945 182.125 126.115 182.295 ;
        RECT 126.405 182.125 126.575 182.295 ;
        RECT 126.865 182.125 127.035 182.295 ;
        RECT 127.325 182.125 127.495 182.295 ;
        RECT 127.785 182.125 127.955 182.295 ;
        RECT 128.245 182.125 128.415 182.295 ;
        RECT 128.705 182.125 128.875 182.295 ;
        RECT 129.165 182.125 129.335 182.295 ;
        RECT 129.625 182.125 129.795 182.295 ;
        RECT 130.085 182.125 130.255 182.295 ;
        RECT 130.545 182.125 130.715 182.295 ;
        RECT 131.005 182.125 131.175 182.295 ;
        RECT 131.465 182.125 131.635 182.295 ;
        RECT 131.925 182.125 132.095 182.295 ;
        RECT 132.385 182.125 132.555 182.295 ;
        RECT 132.845 182.125 133.015 182.295 ;
        RECT 133.305 182.125 133.475 182.295 ;
        RECT 133.765 182.125 133.935 182.295 ;
        RECT 134.225 182.125 134.395 182.295 ;
        RECT 134.685 182.125 134.855 182.295 ;
        RECT 135.145 182.125 135.315 182.295 ;
        RECT 135.605 182.125 135.775 182.295 ;
        RECT 136.065 182.125 136.235 182.295 ;
        RECT 136.525 182.125 136.695 182.295 ;
        RECT 136.985 182.125 137.155 182.295 ;
        RECT 137.445 182.125 137.615 182.295 ;
        RECT 137.905 182.125 138.075 182.295 ;
        RECT 138.365 182.125 138.535 182.295 ;
        RECT 138.825 182.125 138.995 182.295 ;
        RECT 139.285 182.125 139.455 182.295 ;
        RECT 139.745 182.125 139.915 182.295 ;
        RECT 140.205 182.125 140.375 182.295 ;
        RECT 140.665 182.125 140.835 182.295 ;
        RECT 141.125 182.125 141.295 182.295 ;
        RECT 141.585 182.125 141.755 182.295 ;
        RECT 142.045 182.125 142.215 182.295 ;
        RECT 142.505 182.125 142.675 182.295 ;
        RECT 142.965 182.125 143.135 182.295 ;
        RECT 143.425 182.125 143.595 182.295 ;
        RECT 143.885 182.125 144.055 182.295 ;
        RECT 144.345 182.125 144.515 182.295 ;
        RECT 144.805 182.125 144.975 182.295 ;
        RECT 145.265 182.125 145.435 182.295 ;
        RECT 145.725 182.125 145.895 182.295 ;
        RECT 146.185 182.125 146.355 182.295 ;
        RECT 146.645 182.125 146.815 182.295 ;
        RECT 147.105 182.125 147.275 182.295 ;
        RECT 147.565 182.125 147.735 182.295 ;
        RECT 148.025 182.125 148.195 182.295 ;
        RECT 148.485 182.125 148.655 182.295 ;
        RECT 148.945 182.125 149.115 182.295 ;
        RECT 149.405 182.125 149.575 182.295 ;
        RECT 149.865 182.125 150.035 182.295 ;
        RECT 45.445 181.275 45.615 181.445 ;
        RECT 44.525 180.595 44.695 180.765 ;
        RECT 46.825 181.615 46.995 181.785 ;
        RECT 45.905 180.595 46.075 180.765 ;
        RECT 47.745 181.275 47.915 181.445 ;
        RECT 47.285 180.255 47.455 180.425 ;
        RECT 49.585 181.615 49.755 181.785 ;
        RECT 48.665 180.595 48.835 180.765 ;
        RECT 48.205 180.255 48.375 180.425 ;
        RECT 50.505 180.595 50.675 180.765 ;
        RECT 50.965 180.595 51.135 180.765 ;
        RECT 49.585 180.255 49.755 180.425 ;
        RECT 51.885 179.915 52.055 180.085 ;
        RECT 56.945 180.595 57.115 180.765 ;
        RECT 63.845 181.615 64.015 181.785 ;
        RECT 63.385 181.275 63.555 181.445 ;
        RECT 57.865 179.915 58.035 180.085 ;
        RECT 62.005 180.935 62.175 181.105 ;
        RECT 62.925 180.935 63.095 181.105 ;
        RECT 65.225 181.615 65.395 181.785 ;
        RECT 62.925 180.255 63.095 180.425 ;
        RECT 64.305 180.595 64.475 180.765 ;
        RECT 64.765 180.595 64.935 180.765 ;
        RECT 66.145 181.615 66.315 181.785 ;
        RECT 68.445 181.615 68.615 181.785 ;
        RECT 66.605 180.255 66.775 180.425 ;
        RECT 67.525 181.275 67.695 181.445 ;
        RECT 69.365 181.275 69.535 181.445 ;
        RECT 67.985 180.935 68.155 181.105 ;
        RECT 68.445 179.915 68.615 180.085 ;
        RECT 76.725 180.935 76.895 181.105 ;
        RECT 76.265 180.595 76.435 180.765 ;
        RECT 79.025 180.595 79.195 180.765 ;
        RECT 79.485 180.255 79.655 180.425 ;
        RECT 90.525 181.615 90.695 181.785 ;
        RECT 88.225 180.255 88.395 180.425 ;
        RECT 89.145 180.595 89.315 180.765 ;
        RECT 90.985 180.595 91.155 180.765 ;
        RECT 91.445 180.595 91.615 180.765 ;
        RECT 91.905 180.595 92.075 180.765 ;
        RECT 92.825 180.595 92.995 180.765 ;
        RECT 93.745 179.915 93.915 180.085 ;
        RECT 95.125 180.595 95.295 180.765 ;
        RECT 99.725 181.615 99.895 181.785 ;
        RECT 94.205 179.915 94.375 180.085 ;
        RECT 97.885 180.255 98.055 180.425 ;
        RECT 100.185 180.935 100.355 181.105 ;
        RECT 98.805 180.595 98.975 180.765 ;
        RECT 107.545 180.595 107.715 180.765 ;
        RECT 108.925 180.935 109.095 181.105 ;
        RECT 109.385 180.935 109.555 181.105 ;
        RECT 109.845 180.595 110.015 180.765 ;
        RECT 110.765 180.595 110.935 180.765 ;
        RECT 113.065 181.275 113.235 181.445 ;
        RECT 112.145 180.595 112.315 180.765 ;
        RECT 111.685 180.255 111.855 180.425 ;
        RECT 114.905 181.615 115.075 181.785 ;
        RECT 114.445 180.595 114.615 180.765 ;
        RECT 113.525 179.915 113.695 180.085 ;
        RECT 117.665 181.615 117.835 181.785 ;
        RECT 115.825 180.595 115.995 180.765 ;
        RECT 116.285 180.595 116.455 180.765 ;
        RECT 119.965 181.615 120.135 181.785 ;
        RECT 121.345 181.615 121.515 181.785 ;
        RECT 118.585 180.595 118.755 180.765 ;
        RECT 119.045 180.595 119.215 180.765 ;
        RECT 117.665 180.255 117.835 180.425 ;
        RECT 117.205 179.915 117.375 180.085 ;
        RECT 120.425 180.595 120.595 180.765 ;
        RECT 128.705 180.935 128.875 181.105 ;
        RECT 127.785 180.595 127.955 180.765 ;
        RECT 126.865 179.915 127.035 180.085 ;
        RECT 132.845 181.615 133.015 181.785 ;
        RECT 135.145 181.615 135.315 181.785 ;
        RECT 130.545 180.595 130.715 180.765 ;
        RECT 131.465 180.595 131.635 180.765 ;
        RECT 131.005 179.915 131.175 180.085 ;
        RECT 134.685 180.935 134.855 181.105 ;
        RECT 135.605 181.275 135.775 181.445 ;
        RECT 136.525 181.615 136.695 181.785 ;
        RECT 140.205 181.615 140.375 181.785 ;
        RECT 133.765 180.595 133.935 180.765 ;
        RECT 135.145 180.255 135.315 180.425 ;
        RECT 137.445 180.935 137.615 181.105 ;
        RECT 141.585 181.615 141.755 181.785 ;
        RECT 136.525 180.595 136.695 180.765 ;
        RECT 137.905 180.595 138.075 180.765 ;
        RECT 140.665 180.595 140.835 180.765 ;
        RECT 139.285 180.255 139.455 180.425 ;
        RECT 142.045 180.595 142.215 180.765 ;
        RECT 143.425 180.935 143.595 181.105 ;
        RECT 147.105 181.275 147.275 181.445 ;
        RECT 146.645 180.595 146.815 180.765 ;
        RECT 147.565 180.595 147.735 180.765 ;
        RECT 36.245 179.405 36.415 179.575 ;
        RECT 36.705 179.405 36.875 179.575 ;
        RECT 37.165 179.405 37.335 179.575 ;
        RECT 37.625 179.405 37.795 179.575 ;
        RECT 38.085 179.405 38.255 179.575 ;
        RECT 38.545 179.405 38.715 179.575 ;
        RECT 39.005 179.405 39.175 179.575 ;
        RECT 39.465 179.405 39.635 179.575 ;
        RECT 39.925 179.405 40.095 179.575 ;
        RECT 40.385 179.405 40.555 179.575 ;
        RECT 40.845 179.405 41.015 179.575 ;
        RECT 41.305 179.405 41.475 179.575 ;
        RECT 41.765 179.405 41.935 179.575 ;
        RECT 42.225 179.405 42.395 179.575 ;
        RECT 42.685 179.405 42.855 179.575 ;
        RECT 43.145 179.405 43.315 179.575 ;
        RECT 43.605 179.405 43.775 179.575 ;
        RECT 44.065 179.405 44.235 179.575 ;
        RECT 44.525 179.405 44.695 179.575 ;
        RECT 44.985 179.405 45.155 179.575 ;
        RECT 45.445 179.405 45.615 179.575 ;
        RECT 45.905 179.405 46.075 179.575 ;
        RECT 46.365 179.405 46.535 179.575 ;
        RECT 46.825 179.405 46.995 179.575 ;
        RECT 47.285 179.405 47.455 179.575 ;
        RECT 47.745 179.405 47.915 179.575 ;
        RECT 48.205 179.405 48.375 179.575 ;
        RECT 48.665 179.405 48.835 179.575 ;
        RECT 49.125 179.405 49.295 179.575 ;
        RECT 49.585 179.405 49.755 179.575 ;
        RECT 50.045 179.405 50.215 179.575 ;
        RECT 50.505 179.405 50.675 179.575 ;
        RECT 50.965 179.405 51.135 179.575 ;
        RECT 51.425 179.405 51.595 179.575 ;
        RECT 51.885 179.405 52.055 179.575 ;
        RECT 52.345 179.405 52.515 179.575 ;
        RECT 52.805 179.405 52.975 179.575 ;
        RECT 53.265 179.405 53.435 179.575 ;
        RECT 53.725 179.405 53.895 179.575 ;
        RECT 54.185 179.405 54.355 179.575 ;
        RECT 54.645 179.405 54.815 179.575 ;
        RECT 55.105 179.405 55.275 179.575 ;
        RECT 55.565 179.405 55.735 179.575 ;
        RECT 56.025 179.405 56.195 179.575 ;
        RECT 56.485 179.405 56.655 179.575 ;
        RECT 56.945 179.405 57.115 179.575 ;
        RECT 57.405 179.405 57.575 179.575 ;
        RECT 57.865 179.405 58.035 179.575 ;
        RECT 58.325 179.405 58.495 179.575 ;
        RECT 58.785 179.405 58.955 179.575 ;
        RECT 59.245 179.405 59.415 179.575 ;
        RECT 59.705 179.405 59.875 179.575 ;
        RECT 60.165 179.405 60.335 179.575 ;
        RECT 60.625 179.405 60.795 179.575 ;
        RECT 61.085 179.405 61.255 179.575 ;
        RECT 61.545 179.405 61.715 179.575 ;
        RECT 62.005 179.405 62.175 179.575 ;
        RECT 62.465 179.405 62.635 179.575 ;
        RECT 62.925 179.405 63.095 179.575 ;
        RECT 63.385 179.405 63.555 179.575 ;
        RECT 63.845 179.405 64.015 179.575 ;
        RECT 64.305 179.405 64.475 179.575 ;
        RECT 64.765 179.405 64.935 179.575 ;
        RECT 65.225 179.405 65.395 179.575 ;
        RECT 65.685 179.405 65.855 179.575 ;
        RECT 66.145 179.405 66.315 179.575 ;
        RECT 66.605 179.405 66.775 179.575 ;
        RECT 67.065 179.405 67.235 179.575 ;
        RECT 67.525 179.405 67.695 179.575 ;
        RECT 67.985 179.405 68.155 179.575 ;
        RECT 68.445 179.405 68.615 179.575 ;
        RECT 68.905 179.405 69.075 179.575 ;
        RECT 69.365 179.405 69.535 179.575 ;
        RECT 69.825 179.405 69.995 179.575 ;
        RECT 70.285 179.405 70.455 179.575 ;
        RECT 70.745 179.405 70.915 179.575 ;
        RECT 71.205 179.405 71.375 179.575 ;
        RECT 71.665 179.405 71.835 179.575 ;
        RECT 72.125 179.405 72.295 179.575 ;
        RECT 72.585 179.405 72.755 179.575 ;
        RECT 73.045 179.405 73.215 179.575 ;
        RECT 73.505 179.405 73.675 179.575 ;
        RECT 73.965 179.405 74.135 179.575 ;
        RECT 74.425 179.405 74.595 179.575 ;
        RECT 74.885 179.405 75.055 179.575 ;
        RECT 75.345 179.405 75.515 179.575 ;
        RECT 75.805 179.405 75.975 179.575 ;
        RECT 76.265 179.405 76.435 179.575 ;
        RECT 76.725 179.405 76.895 179.575 ;
        RECT 77.185 179.405 77.355 179.575 ;
        RECT 77.645 179.405 77.815 179.575 ;
        RECT 78.105 179.405 78.275 179.575 ;
        RECT 78.565 179.405 78.735 179.575 ;
        RECT 79.025 179.405 79.195 179.575 ;
        RECT 79.485 179.405 79.655 179.575 ;
        RECT 79.945 179.405 80.115 179.575 ;
        RECT 80.405 179.405 80.575 179.575 ;
        RECT 80.865 179.405 81.035 179.575 ;
        RECT 81.325 179.405 81.495 179.575 ;
        RECT 81.785 179.405 81.955 179.575 ;
        RECT 82.245 179.405 82.415 179.575 ;
        RECT 82.705 179.405 82.875 179.575 ;
        RECT 83.165 179.405 83.335 179.575 ;
        RECT 83.625 179.405 83.795 179.575 ;
        RECT 84.085 179.405 84.255 179.575 ;
        RECT 84.545 179.405 84.715 179.575 ;
        RECT 85.005 179.405 85.175 179.575 ;
        RECT 85.465 179.405 85.635 179.575 ;
        RECT 85.925 179.405 86.095 179.575 ;
        RECT 86.385 179.405 86.555 179.575 ;
        RECT 86.845 179.405 87.015 179.575 ;
        RECT 87.305 179.405 87.475 179.575 ;
        RECT 87.765 179.405 87.935 179.575 ;
        RECT 88.225 179.405 88.395 179.575 ;
        RECT 88.685 179.405 88.855 179.575 ;
        RECT 89.145 179.405 89.315 179.575 ;
        RECT 89.605 179.405 89.775 179.575 ;
        RECT 90.065 179.405 90.235 179.575 ;
        RECT 90.525 179.405 90.695 179.575 ;
        RECT 90.985 179.405 91.155 179.575 ;
        RECT 91.445 179.405 91.615 179.575 ;
        RECT 91.905 179.405 92.075 179.575 ;
        RECT 92.365 179.405 92.535 179.575 ;
        RECT 92.825 179.405 92.995 179.575 ;
        RECT 93.285 179.405 93.455 179.575 ;
        RECT 93.745 179.405 93.915 179.575 ;
        RECT 94.205 179.405 94.375 179.575 ;
        RECT 94.665 179.405 94.835 179.575 ;
        RECT 95.125 179.405 95.295 179.575 ;
        RECT 95.585 179.405 95.755 179.575 ;
        RECT 96.045 179.405 96.215 179.575 ;
        RECT 96.505 179.405 96.675 179.575 ;
        RECT 96.965 179.405 97.135 179.575 ;
        RECT 97.425 179.405 97.595 179.575 ;
        RECT 97.885 179.405 98.055 179.575 ;
        RECT 98.345 179.405 98.515 179.575 ;
        RECT 98.805 179.405 98.975 179.575 ;
        RECT 99.265 179.405 99.435 179.575 ;
        RECT 99.725 179.405 99.895 179.575 ;
        RECT 100.185 179.405 100.355 179.575 ;
        RECT 100.645 179.405 100.815 179.575 ;
        RECT 101.105 179.405 101.275 179.575 ;
        RECT 101.565 179.405 101.735 179.575 ;
        RECT 102.025 179.405 102.195 179.575 ;
        RECT 102.485 179.405 102.655 179.575 ;
        RECT 102.945 179.405 103.115 179.575 ;
        RECT 103.405 179.405 103.575 179.575 ;
        RECT 103.865 179.405 104.035 179.575 ;
        RECT 104.325 179.405 104.495 179.575 ;
        RECT 104.785 179.405 104.955 179.575 ;
        RECT 105.245 179.405 105.415 179.575 ;
        RECT 105.705 179.405 105.875 179.575 ;
        RECT 106.165 179.405 106.335 179.575 ;
        RECT 106.625 179.405 106.795 179.575 ;
        RECT 107.085 179.405 107.255 179.575 ;
        RECT 107.545 179.405 107.715 179.575 ;
        RECT 108.005 179.405 108.175 179.575 ;
        RECT 108.465 179.405 108.635 179.575 ;
        RECT 108.925 179.405 109.095 179.575 ;
        RECT 109.385 179.405 109.555 179.575 ;
        RECT 109.845 179.405 110.015 179.575 ;
        RECT 110.305 179.405 110.475 179.575 ;
        RECT 110.765 179.405 110.935 179.575 ;
        RECT 111.225 179.405 111.395 179.575 ;
        RECT 111.685 179.405 111.855 179.575 ;
        RECT 112.145 179.405 112.315 179.575 ;
        RECT 112.605 179.405 112.775 179.575 ;
        RECT 113.065 179.405 113.235 179.575 ;
        RECT 113.525 179.405 113.695 179.575 ;
        RECT 113.985 179.405 114.155 179.575 ;
        RECT 114.445 179.405 114.615 179.575 ;
        RECT 114.905 179.405 115.075 179.575 ;
        RECT 115.365 179.405 115.535 179.575 ;
        RECT 115.825 179.405 115.995 179.575 ;
        RECT 116.285 179.405 116.455 179.575 ;
        RECT 116.745 179.405 116.915 179.575 ;
        RECT 117.205 179.405 117.375 179.575 ;
        RECT 117.665 179.405 117.835 179.575 ;
        RECT 118.125 179.405 118.295 179.575 ;
        RECT 118.585 179.405 118.755 179.575 ;
        RECT 119.045 179.405 119.215 179.575 ;
        RECT 119.505 179.405 119.675 179.575 ;
        RECT 119.965 179.405 120.135 179.575 ;
        RECT 120.425 179.405 120.595 179.575 ;
        RECT 120.885 179.405 121.055 179.575 ;
        RECT 121.345 179.405 121.515 179.575 ;
        RECT 121.805 179.405 121.975 179.575 ;
        RECT 122.265 179.405 122.435 179.575 ;
        RECT 122.725 179.405 122.895 179.575 ;
        RECT 123.185 179.405 123.355 179.575 ;
        RECT 123.645 179.405 123.815 179.575 ;
        RECT 124.105 179.405 124.275 179.575 ;
        RECT 124.565 179.405 124.735 179.575 ;
        RECT 125.025 179.405 125.195 179.575 ;
        RECT 125.485 179.405 125.655 179.575 ;
        RECT 125.945 179.405 126.115 179.575 ;
        RECT 126.405 179.405 126.575 179.575 ;
        RECT 126.865 179.405 127.035 179.575 ;
        RECT 127.325 179.405 127.495 179.575 ;
        RECT 127.785 179.405 127.955 179.575 ;
        RECT 128.245 179.405 128.415 179.575 ;
        RECT 128.705 179.405 128.875 179.575 ;
        RECT 129.165 179.405 129.335 179.575 ;
        RECT 129.625 179.405 129.795 179.575 ;
        RECT 130.085 179.405 130.255 179.575 ;
        RECT 130.545 179.405 130.715 179.575 ;
        RECT 131.005 179.405 131.175 179.575 ;
        RECT 131.465 179.405 131.635 179.575 ;
        RECT 131.925 179.405 132.095 179.575 ;
        RECT 132.385 179.405 132.555 179.575 ;
        RECT 132.845 179.405 133.015 179.575 ;
        RECT 133.305 179.405 133.475 179.575 ;
        RECT 133.765 179.405 133.935 179.575 ;
        RECT 134.225 179.405 134.395 179.575 ;
        RECT 134.685 179.405 134.855 179.575 ;
        RECT 135.145 179.405 135.315 179.575 ;
        RECT 135.605 179.405 135.775 179.575 ;
        RECT 136.065 179.405 136.235 179.575 ;
        RECT 136.525 179.405 136.695 179.575 ;
        RECT 136.985 179.405 137.155 179.575 ;
        RECT 137.445 179.405 137.615 179.575 ;
        RECT 137.905 179.405 138.075 179.575 ;
        RECT 138.365 179.405 138.535 179.575 ;
        RECT 138.825 179.405 138.995 179.575 ;
        RECT 139.285 179.405 139.455 179.575 ;
        RECT 139.745 179.405 139.915 179.575 ;
        RECT 140.205 179.405 140.375 179.575 ;
        RECT 140.665 179.405 140.835 179.575 ;
        RECT 141.125 179.405 141.295 179.575 ;
        RECT 141.585 179.405 141.755 179.575 ;
        RECT 142.045 179.405 142.215 179.575 ;
        RECT 142.505 179.405 142.675 179.575 ;
        RECT 142.965 179.405 143.135 179.575 ;
        RECT 143.425 179.405 143.595 179.575 ;
        RECT 143.885 179.405 144.055 179.575 ;
        RECT 144.345 179.405 144.515 179.575 ;
        RECT 144.805 179.405 144.975 179.575 ;
        RECT 145.265 179.405 145.435 179.575 ;
        RECT 145.725 179.405 145.895 179.575 ;
        RECT 146.185 179.405 146.355 179.575 ;
        RECT 146.645 179.405 146.815 179.575 ;
        RECT 147.105 179.405 147.275 179.575 ;
        RECT 147.565 179.405 147.735 179.575 ;
        RECT 148.025 179.405 148.195 179.575 ;
        RECT 148.485 179.405 148.655 179.575 ;
        RECT 148.945 179.405 149.115 179.575 ;
        RECT 149.405 179.405 149.575 179.575 ;
        RECT 149.865 179.405 150.035 179.575 ;
        RECT 37.625 177.875 37.795 178.045 ;
        RECT 38.110 177.535 38.280 177.705 ;
        RECT 38.505 177.875 38.675 178.045 ;
        RECT 38.960 178.215 39.130 178.385 ;
        RECT 39.695 177.875 39.865 178.045 ;
        RECT 40.210 177.535 40.380 177.705 ;
        RECT 41.780 177.535 41.950 177.705 ;
        RECT 42.215 177.875 42.385 178.045 ;
        RECT 44.525 178.895 44.695 179.065 ;
        RECT 47.285 178.215 47.455 178.385 ;
        RECT 50.505 178.895 50.675 179.065 ;
        RECT 49.585 178.215 49.755 178.385 ;
        RECT 48.665 177.875 48.835 178.045 ;
        RECT 52.805 178.895 52.975 179.065 ;
        RECT 51.885 178.215 52.055 178.385 ;
        RECT 49.585 177.195 49.755 177.365 ;
        RECT 51.425 177.535 51.595 177.705 ;
        RECT 59.245 178.895 59.415 179.065 ;
        RECT 53.725 178.215 53.895 178.385 ;
        RECT 58.325 178.215 58.495 178.385 ;
        RECT 59.705 178.215 59.875 178.385 ;
        RECT 63.385 178.895 63.555 179.065 ;
        RECT 60.625 177.195 60.795 177.365 ;
        RECT 62.465 177.875 62.635 178.045 ;
        RECT 63.385 177.875 63.555 178.045 ;
        RECT 64.730 178.215 64.900 178.385 ;
        RECT 65.165 178.215 65.335 178.385 ;
        RECT 63.845 177.535 64.015 177.705 ;
        RECT 64.305 177.195 64.475 177.365 ;
        RECT 65.685 177.195 65.855 177.365 ;
        RECT 67.065 178.215 67.235 178.385 ;
        RECT 68.905 178.895 69.075 179.065 ;
        RECT 66.605 177.195 66.775 177.365 ;
        RECT 68.445 177.875 68.615 178.045 ;
        RECT 67.985 177.535 68.155 177.705 ;
        RECT 68.905 177.195 69.075 177.365 ;
        RECT 69.825 177.195 69.995 177.365 ;
        RECT 77.645 177.875 77.815 178.045 ;
        RECT 79.945 178.215 80.115 178.385 ;
        RECT 81.325 178.215 81.495 178.385 ;
        RECT 89.145 178.895 89.315 179.065 ;
        RECT 95.585 178.895 95.755 179.065 ;
        RECT 79.465 177.195 79.635 177.365 ;
        RECT 80.385 177.195 80.555 177.365 ;
        RECT 90.065 178.215 90.235 178.385 ;
        RECT 91.445 178.215 91.615 178.385 ;
        RECT 91.905 178.215 92.075 178.385 ;
        RECT 90.985 177.875 91.155 178.045 ;
        RECT 92.825 178.215 92.995 178.385 ;
        RECT 102.025 178.215 102.195 178.385 ;
        RECT 102.485 178.215 102.655 178.385 ;
        RECT 103.405 178.215 103.575 178.385 ;
        RECT 103.865 178.215 104.035 178.385 ;
        RECT 105.245 178.215 105.415 178.385 ;
        RECT 106.625 178.215 106.795 178.385 ;
        RECT 106.165 177.875 106.335 178.045 ;
        RECT 107.545 178.215 107.715 178.385 ;
        RECT 108.465 177.195 108.635 177.365 ;
        RECT 111.225 178.895 111.395 179.065 ;
        RECT 109.845 178.215 110.015 178.385 ;
        RECT 110.305 178.215 110.475 178.385 ;
        RECT 108.925 177.535 109.095 177.705 ;
        RECT 119.505 178.895 119.675 179.065 ;
        RECT 117.205 177.875 117.375 178.045 ;
        RECT 117.665 178.215 117.835 178.385 ;
        RECT 118.125 178.215 118.295 178.385 ;
        RECT 118.585 178.215 118.755 178.385 ;
        RECT 119.965 178.555 120.135 178.725 ;
        RECT 127.325 177.195 127.495 177.365 ;
        RECT 131.925 178.215 132.095 178.385 ;
        RECT 135.145 178.895 135.315 179.065 ;
        RECT 130.545 177.195 130.715 177.365 ;
        RECT 134.225 178.215 134.395 178.385 ;
        RECT 133.305 177.875 133.475 178.045 ;
        RECT 133.305 177.195 133.475 177.365 ;
        RECT 135.605 177.875 135.775 178.045 ;
        RECT 136.985 178.555 137.155 178.725 ;
        RECT 138.030 177.875 138.200 178.045 ;
        RECT 138.825 177.195 138.995 177.365 ;
        RECT 140.205 177.875 140.375 178.045 ;
        RECT 140.690 177.535 140.860 177.705 ;
        RECT 141.085 177.875 141.255 178.045 ;
        RECT 141.485 178.215 141.655 178.385 ;
        RECT 142.275 177.875 142.445 178.045 ;
        RECT 142.790 177.535 142.960 177.705 ;
        RECT 144.360 177.535 144.530 177.705 ;
        RECT 144.795 177.875 144.965 178.045 ;
        RECT 147.105 177.195 147.275 177.365 ;
        RECT 36.245 176.685 36.415 176.855 ;
        RECT 36.705 176.685 36.875 176.855 ;
        RECT 37.165 176.685 37.335 176.855 ;
        RECT 37.625 176.685 37.795 176.855 ;
        RECT 38.085 176.685 38.255 176.855 ;
        RECT 38.545 176.685 38.715 176.855 ;
        RECT 39.005 176.685 39.175 176.855 ;
        RECT 39.465 176.685 39.635 176.855 ;
        RECT 39.925 176.685 40.095 176.855 ;
        RECT 40.385 176.685 40.555 176.855 ;
        RECT 40.845 176.685 41.015 176.855 ;
        RECT 41.305 176.685 41.475 176.855 ;
        RECT 41.765 176.685 41.935 176.855 ;
        RECT 42.225 176.685 42.395 176.855 ;
        RECT 42.685 176.685 42.855 176.855 ;
        RECT 43.145 176.685 43.315 176.855 ;
        RECT 43.605 176.685 43.775 176.855 ;
        RECT 44.065 176.685 44.235 176.855 ;
        RECT 44.525 176.685 44.695 176.855 ;
        RECT 44.985 176.685 45.155 176.855 ;
        RECT 45.445 176.685 45.615 176.855 ;
        RECT 45.905 176.685 46.075 176.855 ;
        RECT 46.365 176.685 46.535 176.855 ;
        RECT 46.825 176.685 46.995 176.855 ;
        RECT 47.285 176.685 47.455 176.855 ;
        RECT 47.745 176.685 47.915 176.855 ;
        RECT 48.205 176.685 48.375 176.855 ;
        RECT 48.665 176.685 48.835 176.855 ;
        RECT 49.125 176.685 49.295 176.855 ;
        RECT 49.585 176.685 49.755 176.855 ;
        RECT 50.045 176.685 50.215 176.855 ;
        RECT 50.505 176.685 50.675 176.855 ;
        RECT 50.965 176.685 51.135 176.855 ;
        RECT 51.425 176.685 51.595 176.855 ;
        RECT 51.885 176.685 52.055 176.855 ;
        RECT 52.345 176.685 52.515 176.855 ;
        RECT 52.805 176.685 52.975 176.855 ;
        RECT 53.265 176.685 53.435 176.855 ;
        RECT 53.725 176.685 53.895 176.855 ;
        RECT 54.185 176.685 54.355 176.855 ;
        RECT 54.645 176.685 54.815 176.855 ;
        RECT 55.105 176.685 55.275 176.855 ;
        RECT 55.565 176.685 55.735 176.855 ;
        RECT 56.025 176.685 56.195 176.855 ;
        RECT 56.485 176.685 56.655 176.855 ;
        RECT 56.945 176.685 57.115 176.855 ;
        RECT 57.405 176.685 57.575 176.855 ;
        RECT 57.865 176.685 58.035 176.855 ;
        RECT 58.325 176.685 58.495 176.855 ;
        RECT 58.785 176.685 58.955 176.855 ;
        RECT 59.245 176.685 59.415 176.855 ;
        RECT 59.705 176.685 59.875 176.855 ;
        RECT 60.165 176.685 60.335 176.855 ;
        RECT 60.625 176.685 60.795 176.855 ;
        RECT 61.085 176.685 61.255 176.855 ;
        RECT 61.545 176.685 61.715 176.855 ;
        RECT 62.005 176.685 62.175 176.855 ;
        RECT 62.465 176.685 62.635 176.855 ;
        RECT 62.925 176.685 63.095 176.855 ;
        RECT 63.385 176.685 63.555 176.855 ;
        RECT 63.845 176.685 64.015 176.855 ;
        RECT 64.305 176.685 64.475 176.855 ;
        RECT 64.765 176.685 64.935 176.855 ;
        RECT 65.225 176.685 65.395 176.855 ;
        RECT 65.685 176.685 65.855 176.855 ;
        RECT 66.145 176.685 66.315 176.855 ;
        RECT 66.605 176.685 66.775 176.855 ;
        RECT 67.065 176.685 67.235 176.855 ;
        RECT 67.525 176.685 67.695 176.855 ;
        RECT 67.985 176.685 68.155 176.855 ;
        RECT 68.445 176.685 68.615 176.855 ;
        RECT 68.905 176.685 69.075 176.855 ;
        RECT 69.365 176.685 69.535 176.855 ;
        RECT 69.825 176.685 69.995 176.855 ;
        RECT 70.285 176.685 70.455 176.855 ;
        RECT 70.745 176.685 70.915 176.855 ;
        RECT 71.205 176.685 71.375 176.855 ;
        RECT 71.665 176.685 71.835 176.855 ;
        RECT 72.125 176.685 72.295 176.855 ;
        RECT 72.585 176.685 72.755 176.855 ;
        RECT 73.045 176.685 73.215 176.855 ;
        RECT 73.505 176.685 73.675 176.855 ;
        RECT 73.965 176.685 74.135 176.855 ;
        RECT 74.425 176.685 74.595 176.855 ;
        RECT 74.885 176.685 75.055 176.855 ;
        RECT 75.345 176.685 75.515 176.855 ;
        RECT 75.805 176.685 75.975 176.855 ;
        RECT 76.265 176.685 76.435 176.855 ;
        RECT 76.725 176.685 76.895 176.855 ;
        RECT 77.185 176.685 77.355 176.855 ;
        RECT 77.645 176.685 77.815 176.855 ;
        RECT 78.105 176.685 78.275 176.855 ;
        RECT 78.565 176.685 78.735 176.855 ;
        RECT 79.025 176.685 79.195 176.855 ;
        RECT 79.485 176.685 79.655 176.855 ;
        RECT 79.945 176.685 80.115 176.855 ;
        RECT 80.405 176.685 80.575 176.855 ;
        RECT 80.865 176.685 81.035 176.855 ;
        RECT 81.325 176.685 81.495 176.855 ;
        RECT 81.785 176.685 81.955 176.855 ;
        RECT 82.245 176.685 82.415 176.855 ;
        RECT 82.705 176.685 82.875 176.855 ;
        RECT 83.165 176.685 83.335 176.855 ;
        RECT 83.625 176.685 83.795 176.855 ;
        RECT 84.085 176.685 84.255 176.855 ;
        RECT 84.545 176.685 84.715 176.855 ;
        RECT 85.005 176.685 85.175 176.855 ;
        RECT 85.465 176.685 85.635 176.855 ;
        RECT 85.925 176.685 86.095 176.855 ;
        RECT 86.385 176.685 86.555 176.855 ;
        RECT 86.845 176.685 87.015 176.855 ;
        RECT 87.305 176.685 87.475 176.855 ;
        RECT 87.765 176.685 87.935 176.855 ;
        RECT 88.225 176.685 88.395 176.855 ;
        RECT 88.685 176.685 88.855 176.855 ;
        RECT 89.145 176.685 89.315 176.855 ;
        RECT 89.605 176.685 89.775 176.855 ;
        RECT 90.065 176.685 90.235 176.855 ;
        RECT 90.525 176.685 90.695 176.855 ;
        RECT 90.985 176.685 91.155 176.855 ;
        RECT 91.445 176.685 91.615 176.855 ;
        RECT 91.905 176.685 92.075 176.855 ;
        RECT 92.365 176.685 92.535 176.855 ;
        RECT 92.825 176.685 92.995 176.855 ;
        RECT 93.285 176.685 93.455 176.855 ;
        RECT 93.745 176.685 93.915 176.855 ;
        RECT 94.205 176.685 94.375 176.855 ;
        RECT 94.665 176.685 94.835 176.855 ;
        RECT 95.125 176.685 95.295 176.855 ;
        RECT 95.585 176.685 95.755 176.855 ;
        RECT 96.045 176.685 96.215 176.855 ;
        RECT 96.505 176.685 96.675 176.855 ;
        RECT 96.965 176.685 97.135 176.855 ;
        RECT 97.425 176.685 97.595 176.855 ;
        RECT 97.885 176.685 98.055 176.855 ;
        RECT 98.345 176.685 98.515 176.855 ;
        RECT 98.805 176.685 98.975 176.855 ;
        RECT 99.265 176.685 99.435 176.855 ;
        RECT 99.725 176.685 99.895 176.855 ;
        RECT 100.185 176.685 100.355 176.855 ;
        RECT 100.645 176.685 100.815 176.855 ;
        RECT 101.105 176.685 101.275 176.855 ;
        RECT 101.565 176.685 101.735 176.855 ;
        RECT 102.025 176.685 102.195 176.855 ;
        RECT 102.485 176.685 102.655 176.855 ;
        RECT 102.945 176.685 103.115 176.855 ;
        RECT 103.405 176.685 103.575 176.855 ;
        RECT 103.865 176.685 104.035 176.855 ;
        RECT 104.325 176.685 104.495 176.855 ;
        RECT 104.785 176.685 104.955 176.855 ;
        RECT 105.245 176.685 105.415 176.855 ;
        RECT 105.705 176.685 105.875 176.855 ;
        RECT 106.165 176.685 106.335 176.855 ;
        RECT 106.625 176.685 106.795 176.855 ;
        RECT 107.085 176.685 107.255 176.855 ;
        RECT 107.545 176.685 107.715 176.855 ;
        RECT 108.005 176.685 108.175 176.855 ;
        RECT 108.465 176.685 108.635 176.855 ;
        RECT 108.925 176.685 109.095 176.855 ;
        RECT 109.385 176.685 109.555 176.855 ;
        RECT 109.845 176.685 110.015 176.855 ;
        RECT 110.305 176.685 110.475 176.855 ;
        RECT 110.765 176.685 110.935 176.855 ;
        RECT 111.225 176.685 111.395 176.855 ;
        RECT 111.685 176.685 111.855 176.855 ;
        RECT 112.145 176.685 112.315 176.855 ;
        RECT 112.605 176.685 112.775 176.855 ;
        RECT 113.065 176.685 113.235 176.855 ;
        RECT 113.525 176.685 113.695 176.855 ;
        RECT 113.985 176.685 114.155 176.855 ;
        RECT 114.445 176.685 114.615 176.855 ;
        RECT 114.905 176.685 115.075 176.855 ;
        RECT 115.365 176.685 115.535 176.855 ;
        RECT 115.825 176.685 115.995 176.855 ;
        RECT 116.285 176.685 116.455 176.855 ;
        RECT 116.745 176.685 116.915 176.855 ;
        RECT 117.205 176.685 117.375 176.855 ;
        RECT 117.665 176.685 117.835 176.855 ;
        RECT 118.125 176.685 118.295 176.855 ;
        RECT 118.585 176.685 118.755 176.855 ;
        RECT 119.045 176.685 119.215 176.855 ;
        RECT 119.505 176.685 119.675 176.855 ;
        RECT 119.965 176.685 120.135 176.855 ;
        RECT 120.425 176.685 120.595 176.855 ;
        RECT 120.885 176.685 121.055 176.855 ;
        RECT 121.345 176.685 121.515 176.855 ;
        RECT 121.805 176.685 121.975 176.855 ;
        RECT 122.265 176.685 122.435 176.855 ;
        RECT 122.725 176.685 122.895 176.855 ;
        RECT 123.185 176.685 123.355 176.855 ;
        RECT 123.645 176.685 123.815 176.855 ;
        RECT 124.105 176.685 124.275 176.855 ;
        RECT 124.565 176.685 124.735 176.855 ;
        RECT 125.025 176.685 125.195 176.855 ;
        RECT 125.485 176.685 125.655 176.855 ;
        RECT 125.945 176.685 126.115 176.855 ;
        RECT 126.405 176.685 126.575 176.855 ;
        RECT 126.865 176.685 127.035 176.855 ;
        RECT 127.325 176.685 127.495 176.855 ;
        RECT 127.785 176.685 127.955 176.855 ;
        RECT 128.245 176.685 128.415 176.855 ;
        RECT 128.705 176.685 128.875 176.855 ;
        RECT 129.165 176.685 129.335 176.855 ;
        RECT 129.625 176.685 129.795 176.855 ;
        RECT 130.085 176.685 130.255 176.855 ;
        RECT 130.545 176.685 130.715 176.855 ;
        RECT 131.005 176.685 131.175 176.855 ;
        RECT 131.465 176.685 131.635 176.855 ;
        RECT 131.925 176.685 132.095 176.855 ;
        RECT 132.385 176.685 132.555 176.855 ;
        RECT 132.845 176.685 133.015 176.855 ;
        RECT 133.305 176.685 133.475 176.855 ;
        RECT 133.765 176.685 133.935 176.855 ;
        RECT 134.225 176.685 134.395 176.855 ;
        RECT 134.685 176.685 134.855 176.855 ;
        RECT 135.145 176.685 135.315 176.855 ;
        RECT 135.605 176.685 135.775 176.855 ;
        RECT 136.065 176.685 136.235 176.855 ;
        RECT 136.525 176.685 136.695 176.855 ;
        RECT 136.985 176.685 137.155 176.855 ;
        RECT 137.445 176.685 137.615 176.855 ;
        RECT 137.905 176.685 138.075 176.855 ;
        RECT 138.365 176.685 138.535 176.855 ;
        RECT 138.825 176.685 138.995 176.855 ;
        RECT 139.285 176.685 139.455 176.855 ;
        RECT 139.745 176.685 139.915 176.855 ;
        RECT 140.205 176.685 140.375 176.855 ;
        RECT 140.665 176.685 140.835 176.855 ;
        RECT 141.125 176.685 141.295 176.855 ;
        RECT 141.585 176.685 141.755 176.855 ;
        RECT 142.045 176.685 142.215 176.855 ;
        RECT 142.505 176.685 142.675 176.855 ;
        RECT 142.965 176.685 143.135 176.855 ;
        RECT 143.425 176.685 143.595 176.855 ;
        RECT 143.885 176.685 144.055 176.855 ;
        RECT 144.345 176.685 144.515 176.855 ;
        RECT 144.805 176.685 144.975 176.855 ;
        RECT 145.265 176.685 145.435 176.855 ;
        RECT 145.725 176.685 145.895 176.855 ;
        RECT 146.185 176.685 146.355 176.855 ;
        RECT 146.645 176.685 146.815 176.855 ;
        RECT 147.105 176.685 147.275 176.855 ;
        RECT 147.565 176.685 147.735 176.855 ;
        RECT 148.025 176.685 148.195 176.855 ;
        RECT 148.485 176.685 148.655 176.855 ;
        RECT 148.945 176.685 149.115 176.855 ;
        RECT 149.405 176.685 149.575 176.855 ;
        RECT 149.865 176.685 150.035 176.855 ;
        RECT 40.385 176.175 40.555 176.345 ;
        RECT 40.385 175.155 40.555 175.325 ;
        RECT 41.305 175.155 41.475 175.325 ;
        RECT 47.285 175.155 47.455 175.325 ;
        RECT 48.665 175.495 48.835 175.665 ;
        RECT 49.585 176.175 49.755 176.345 ;
        RECT 51.885 176.175 52.055 176.345 ;
        RECT 50.505 175.155 50.675 175.325 ;
        RECT 53.265 175.835 53.435 176.005 ;
        RECT 50.965 175.155 51.135 175.325 ;
        RECT 51.885 175.155 52.055 175.325 ;
        RECT 52.345 175.155 52.515 175.325 ;
        RECT 54.185 175.835 54.355 176.005 ;
        RECT 55.105 176.175 55.275 176.345 ;
        RECT 56.025 175.835 56.195 176.005 ;
        RECT 55.565 175.495 55.735 175.665 ;
        RECT 57.405 176.175 57.575 176.345 ;
        RECT 55.105 174.475 55.275 174.645 ;
        RECT 56.945 175.155 57.115 175.325 ;
        RECT 58.325 176.175 58.495 176.345 ;
        RECT 59.705 176.175 59.875 176.345 ;
        RECT 60.165 175.835 60.335 176.005 ;
        RECT 58.785 174.815 58.955 174.985 ;
        RECT 59.245 175.155 59.415 175.325 ;
        RECT 60.625 175.495 60.795 175.665 ;
        RECT 61.545 175.495 61.715 175.665 ;
        RECT 60.625 174.475 60.795 174.645 ;
        RECT 64.305 174.475 64.475 174.645 ;
        RECT 70.745 175.155 70.915 175.325 ;
        RECT 83.165 175.155 83.335 175.325 ;
        RECT 84.085 175.155 84.255 175.325 ;
        RECT 85.005 175.155 85.175 175.325 ;
        RECT 87.305 175.155 87.475 175.325 ;
        RECT 86.385 174.815 86.555 174.985 ;
        RECT 87.765 175.155 87.935 175.325 ;
        RECT 88.685 175.155 88.855 175.325 ;
        RECT 89.145 175.155 89.315 175.325 ;
        RECT 89.605 175.155 89.775 175.325 ;
        RECT 91.905 175.155 92.075 175.325 ;
        RECT 92.365 175.155 92.535 175.325 ;
        RECT 92.825 175.155 92.995 175.325 ;
        RECT 93.285 175.155 93.455 175.325 ;
        RECT 90.985 174.475 91.155 174.645 ;
        RECT 94.205 174.475 94.375 174.645 ;
        RECT 98.805 175.155 98.975 175.325 ;
        RECT 100.185 175.495 100.355 175.665 ;
        RECT 101.105 175.155 101.275 175.325 ;
        RECT 102.485 175.495 102.655 175.665 ;
        RECT 102.025 175.155 102.195 175.325 ;
        RECT 103.865 175.155 104.035 175.325 ;
        RECT 105.705 175.495 105.875 175.665 ;
        RECT 106.165 175.155 106.335 175.325 ;
        RECT 106.625 175.155 106.795 175.325 ;
        RECT 107.085 175.155 107.255 175.325 ;
        RECT 104.785 174.475 104.955 174.645 ;
        RECT 108.005 174.475 108.175 174.645 ;
        RECT 110.765 176.175 110.935 176.345 ;
        RECT 108.465 174.815 108.635 174.985 ;
        RECT 109.385 175.155 109.555 175.325 ;
        RECT 111.225 175.155 111.395 175.325 ;
        RECT 114.445 175.495 114.615 175.665 ;
        RECT 115.825 175.495 115.995 175.665 ;
        RECT 120.425 175.835 120.595 176.005 ;
        RECT 121.345 176.175 121.515 176.345 ;
        RECT 119.045 175.155 119.215 175.325 ;
        RECT 119.505 174.475 119.675 174.645 ;
        RECT 120.885 175.155 121.055 175.325 ;
        RECT 122.265 175.495 122.435 175.665 ;
        RECT 123.185 175.155 123.355 175.325 ;
        RECT 124.105 175.155 124.275 175.325 ;
        RECT 120.425 174.815 120.595 174.985 ;
        RECT 122.265 174.815 122.435 174.985 ;
        RECT 125.025 175.155 125.195 175.325 ;
        RECT 124.565 174.815 124.735 174.985 ;
        RECT 128.730 175.835 128.900 176.005 ;
        RECT 126.865 175.155 127.035 175.325 ;
        RECT 128.245 175.495 128.415 175.665 ;
        RECT 127.325 175.155 127.495 175.325 ;
        RECT 127.785 175.155 127.955 175.325 ;
        RECT 125.945 174.475 126.115 174.645 ;
        RECT 129.125 175.495 129.295 175.665 ;
        RECT 129.470 174.815 129.640 174.985 ;
        RECT 130.830 175.835 131.000 176.005 ;
        RECT 130.315 175.495 130.485 175.665 ;
        RECT 132.400 175.835 132.570 176.005 ;
        RECT 132.835 175.495 133.005 175.665 ;
        RECT 135.145 176.175 135.315 176.345 ;
        RECT 137.445 176.175 137.615 176.345 ;
        RECT 136.525 175.155 136.695 175.325 ;
        RECT 138.365 175.835 138.535 176.005 ;
        RECT 138.825 175.155 138.995 175.325 ;
        RECT 36.245 173.965 36.415 174.135 ;
        RECT 36.705 173.965 36.875 174.135 ;
        RECT 37.165 173.965 37.335 174.135 ;
        RECT 37.625 173.965 37.795 174.135 ;
        RECT 38.085 173.965 38.255 174.135 ;
        RECT 38.545 173.965 38.715 174.135 ;
        RECT 39.005 173.965 39.175 174.135 ;
        RECT 39.465 173.965 39.635 174.135 ;
        RECT 39.925 173.965 40.095 174.135 ;
        RECT 40.385 173.965 40.555 174.135 ;
        RECT 40.845 173.965 41.015 174.135 ;
        RECT 41.305 173.965 41.475 174.135 ;
        RECT 41.765 173.965 41.935 174.135 ;
        RECT 42.225 173.965 42.395 174.135 ;
        RECT 42.685 173.965 42.855 174.135 ;
        RECT 43.145 173.965 43.315 174.135 ;
        RECT 43.605 173.965 43.775 174.135 ;
        RECT 44.065 173.965 44.235 174.135 ;
        RECT 44.525 173.965 44.695 174.135 ;
        RECT 44.985 173.965 45.155 174.135 ;
        RECT 45.445 173.965 45.615 174.135 ;
        RECT 45.905 173.965 46.075 174.135 ;
        RECT 46.365 173.965 46.535 174.135 ;
        RECT 46.825 173.965 46.995 174.135 ;
        RECT 47.285 173.965 47.455 174.135 ;
        RECT 47.745 173.965 47.915 174.135 ;
        RECT 48.205 173.965 48.375 174.135 ;
        RECT 48.665 173.965 48.835 174.135 ;
        RECT 49.125 173.965 49.295 174.135 ;
        RECT 49.585 173.965 49.755 174.135 ;
        RECT 50.045 173.965 50.215 174.135 ;
        RECT 50.505 173.965 50.675 174.135 ;
        RECT 50.965 173.965 51.135 174.135 ;
        RECT 51.425 173.965 51.595 174.135 ;
        RECT 51.885 173.965 52.055 174.135 ;
        RECT 52.345 173.965 52.515 174.135 ;
        RECT 52.805 173.965 52.975 174.135 ;
        RECT 53.265 173.965 53.435 174.135 ;
        RECT 53.725 173.965 53.895 174.135 ;
        RECT 54.185 173.965 54.355 174.135 ;
        RECT 54.645 173.965 54.815 174.135 ;
        RECT 55.105 173.965 55.275 174.135 ;
        RECT 55.565 173.965 55.735 174.135 ;
        RECT 56.025 173.965 56.195 174.135 ;
        RECT 56.485 173.965 56.655 174.135 ;
        RECT 56.945 173.965 57.115 174.135 ;
        RECT 57.405 173.965 57.575 174.135 ;
        RECT 57.865 173.965 58.035 174.135 ;
        RECT 58.325 173.965 58.495 174.135 ;
        RECT 58.785 173.965 58.955 174.135 ;
        RECT 59.245 173.965 59.415 174.135 ;
        RECT 59.705 173.965 59.875 174.135 ;
        RECT 60.165 173.965 60.335 174.135 ;
        RECT 60.625 173.965 60.795 174.135 ;
        RECT 61.085 173.965 61.255 174.135 ;
        RECT 61.545 173.965 61.715 174.135 ;
        RECT 62.005 173.965 62.175 174.135 ;
        RECT 62.465 173.965 62.635 174.135 ;
        RECT 62.925 173.965 63.095 174.135 ;
        RECT 63.385 173.965 63.555 174.135 ;
        RECT 63.845 173.965 64.015 174.135 ;
        RECT 64.305 173.965 64.475 174.135 ;
        RECT 64.765 173.965 64.935 174.135 ;
        RECT 65.225 173.965 65.395 174.135 ;
        RECT 65.685 173.965 65.855 174.135 ;
        RECT 66.145 173.965 66.315 174.135 ;
        RECT 66.605 173.965 66.775 174.135 ;
        RECT 67.065 173.965 67.235 174.135 ;
        RECT 67.525 173.965 67.695 174.135 ;
        RECT 67.985 173.965 68.155 174.135 ;
        RECT 68.445 173.965 68.615 174.135 ;
        RECT 68.905 173.965 69.075 174.135 ;
        RECT 69.365 173.965 69.535 174.135 ;
        RECT 69.825 173.965 69.995 174.135 ;
        RECT 70.285 173.965 70.455 174.135 ;
        RECT 70.745 173.965 70.915 174.135 ;
        RECT 71.205 173.965 71.375 174.135 ;
        RECT 71.665 173.965 71.835 174.135 ;
        RECT 72.125 173.965 72.295 174.135 ;
        RECT 72.585 173.965 72.755 174.135 ;
        RECT 73.045 173.965 73.215 174.135 ;
        RECT 73.505 173.965 73.675 174.135 ;
        RECT 73.965 173.965 74.135 174.135 ;
        RECT 74.425 173.965 74.595 174.135 ;
        RECT 74.885 173.965 75.055 174.135 ;
        RECT 75.345 173.965 75.515 174.135 ;
        RECT 75.805 173.965 75.975 174.135 ;
        RECT 76.265 173.965 76.435 174.135 ;
        RECT 76.725 173.965 76.895 174.135 ;
        RECT 77.185 173.965 77.355 174.135 ;
        RECT 77.645 173.965 77.815 174.135 ;
        RECT 78.105 173.965 78.275 174.135 ;
        RECT 78.565 173.965 78.735 174.135 ;
        RECT 79.025 173.965 79.195 174.135 ;
        RECT 79.485 173.965 79.655 174.135 ;
        RECT 79.945 173.965 80.115 174.135 ;
        RECT 80.405 173.965 80.575 174.135 ;
        RECT 80.865 173.965 81.035 174.135 ;
        RECT 81.325 173.965 81.495 174.135 ;
        RECT 81.785 173.965 81.955 174.135 ;
        RECT 82.245 173.965 82.415 174.135 ;
        RECT 82.705 173.965 82.875 174.135 ;
        RECT 83.165 173.965 83.335 174.135 ;
        RECT 83.625 173.965 83.795 174.135 ;
        RECT 84.085 173.965 84.255 174.135 ;
        RECT 84.545 173.965 84.715 174.135 ;
        RECT 85.005 173.965 85.175 174.135 ;
        RECT 85.465 173.965 85.635 174.135 ;
        RECT 85.925 173.965 86.095 174.135 ;
        RECT 86.385 173.965 86.555 174.135 ;
        RECT 86.845 173.965 87.015 174.135 ;
        RECT 87.305 173.965 87.475 174.135 ;
        RECT 87.765 173.965 87.935 174.135 ;
        RECT 88.225 173.965 88.395 174.135 ;
        RECT 88.685 173.965 88.855 174.135 ;
        RECT 89.145 173.965 89.315 174.135 ;
        RECT 89.605 173.965 89.775 174.135 ;
        RECT 90.065 173.965 90.235 174.135 ;
        RECT 90.525 173.965 90.695 174.135 ;
        RECT 90.985 173.965 91.155 174.135 ;
        RECT 91.445 173.965 91.615 174.135 ;
        RECT 91.905 173.965 92.075 174.135 ;
        RECT 92.365 173.965 92.535 174.135 ;
        RECT 92.825 173.965 92.995 174.135 ;
        RECT 93.285 173.965 93.455 174.135 ;
        RECT 93.745 173.965 93.915 174.135 ;
        RECT 94.205 173.965 94.375 174.135 ;
        RECT 94.665 173.965 94.835 174.135 ;
        RECT 95.125 173.965 95.295 174.135 ;
        RECT 95.585 173.965 95.755 174.135 ;
        RECT 96.045 173.965 96.215 174.135 ;
        RECT 96.505 173.965 96.675 174.135 ;
        RECT 96.965 173.965 97.135 174.135 ;
        RECT 97.425 173.965 97.595 174.135 ;
        RECT 97.885 173.965 98.055 174.135 ;
        RECT 98.345 173.965 98.515 174.135 ;
        RECT 98.805 173.965 98.975 174.135 ;
        RECT 99.265 173.965 99.435 174.135 ;
        RECT 99.725 173.965 99.895 174.135 ;
        RECT 100.185 173.965 100.355 174.135 ;
        RECT 100.645 173.965 100.815 174.135 ;
        RECT 101.105 173.965 101.275 174.135 ;
        RECT 101.565 173.965 101.735 174.135 ;
        RECT 102.025 173.965 102.195 174.135 ;
        RECT 102.485 173.965 102.655 174.135 ;
        RECT 102.945 173.965 103.115 174.135 ;
        RECT 103.405 173.965 103.575 174.135 ;
        RECT 103.865 173.965 104.035 174.135 ;
        RECT 104.325 173.965 104.495 174.135 ;
        RECT 104.785 173.965 104.955 174.135 ;
        RECT 105.245 173.965 105.415 174.135 ;
        RECT 105.705 173.965 105.875 174.135 ;
        RECT 106.165 173.965 106.335 174.135 ;
        RECT 106.625 173.965 106.795 174.135 ;
        RECT 107.085 173.965 107.255 174.135 ;
        RECT 107.545 173.965 107.715 174.135 ;
        RECT 108.005 173.965 108.175 174.135 ;
        RECT 108.465 173.965 108.635 174.135 ;
        RECT 108.925 173.965 109.095 174.135 ;
        RECT 109.385 173.965 109.555 174.135 ;
        RECT 109.845 173.965 110.015 174.135 ;
        RECT 110.305 173.965 110.475 174.135 ;
        RECT 110.765 173.965 110.935 174.135 ;
        RECT 111.225 173.965 111.395 174.135 ;
        RECT 111.685 173.965 111.855 174.135 ;
        RECT 112.145 173.965 112.315 174.135 ;
        RECT 112.605 173.965 112.775 174.135 ;
        RECT 113.065 173.965 113.235 174.135 ;
        RECT 113.525 173.965 113.695 174.135 ;
        RECT 113.985 173.965 114.155 174.135 ;
        RECT 114.445 173.965 114.615 174.135 ;
        RECT 114.905 173.965 115.075 174.135 ;
        RECT 115.365 173.965 115.535 174.135 ;
        RECT 115.825 173.965 115.995 174.135 ;
        RECT 116.285 173.965 116.455 174.135 ;
        RECT 116.745 173.965 116.915 174.135 ;
        RECT 117.205 173.965 117.375 174.135 ;
        RECT 117.665 173.965 117.835 174.135 ;
        RECT 118.125 173.965 118.295 174.135 ;
        RECT 118.585 173.965 118.755 174.135 ;
        RECT 119.045 173.965 119.215 174.135 ;
        RECT 119.505 173.965 119.675 174.135 ;
        RECT 119.965 173.965 120.135 174.135 ;
        RECT 120.425 173.965 120.595 174.135 ;
        RECT 120.885 173.965 121.055 174.135 ;
        RECT 121.345 173.965 121.515 174.135 ;
        RECT 121.805 173.965 121.975 174.135 ;
        RECT 122.265 173.965 122.435 174.135 ;
        RECT 122.725 173.965 122.895 174.135 ;
        RECT 123.185 173.965 123.355 174.135 ;
        RECT 123.645 173.965 123.815 174.135 ;
        RECT 124.105 173.965 124.275 174.135 ;
        RECT 124.565 173.965 124.735 174.135 ;
        RECT 125.025 173.965 125.195 174.135 ;
        RECT 125.485 173.965 125.655 174.135 ;
        RECT 125.945 173.965 126.115 174.135 ;
        RECT 126.405 173.965 126.575 174.135 ;
        RECT 126.865 173.965 127.035 174.135 ;
        RECT 127.325 173.965 127.495 174.135 ;
        RECT 127.785 173.965 127.955 174.135 ;
        RECT 128.245 173.965 128.415 174.135 ;
        RECT 128.705 173.965 128.875 174.135 ;
        RECT 129.165 173.965 129.335 174.135 ;
        RECT 129.625 173.965 129.795 174.135 ;
        RECT 130.085 173.965 130.255 174.135 ;
        RECT 130.545 173.965 130.715 174.135 ;
        RECT 131.005 173.965 131.175 174.135 ;
        RECT 131.465 173.965 131.635 174.135 ;
        RECT 131.925 173.965 132.095 174.135 ;
        RECT 132.385 173.965 132.555 174.135 ;
        RECT 132.845 173.965 133.015 174.135 ;
        RECT 133.305 173.965 133.475 174.135 ;
        RECT 133.765 173.965 133.935 174.135 ;
        RECT 134.225 173.965 134.395 174.135 ;
        RECT 134.685 173.965 134.855 174.135 ;
        RECT 135.145 173.965 135.315 174.135 ;
        RECT 135.605 173.965 135.775 174.135 ;
        RECT 136.065 173.965 136.235 174.135 ;
        RECT 136.525 173.965 136.695 174.135 ;
        RECT 136.985 173.965 137.155 174.135 ;
        RECT 137.445 173.965 137.615 174.135 ;
        RECT 137.905 173.965 138.075 174.135 ;
        RECT 138.365 173.965 138.535 174.135 ;
        RECT 138.825 173.965 138.995 174.135 ;
        RECT 139.285 173.965 139.455 174.135 ;
        RECT 139.745 173.965 139.915 174.135 ;
        RECT 140.205 173.965 140.375 174.135 ;
        RECT 140.665 173.965 140.835 174.135 ;
        RECT 141.125 173.965 141.295 174.135 ;
        RECT 141.585 173.965 141.755 174.135 ;
        RECT 142.045 173.965 142.215 174.135 ;
        RECT 142.505 173.965 142.675 174.135 ;
        RECT 142.965 173.965 143.135 174.135 ;
        RECT 143.425 173.965 143.595 174.135 ;
        RECT 143.885 173.965 144.055 174.135 ;
        RECT 144.345 173.965 144.515 174.135 ;
        RECT 144.805 173.965 144.975 174.135 ;
        RECT 145.265 173.965 145.435 174.135 ;
        RECT 145.725 173.965 145.895 174.135 ;
        RECT 146.185 173.965 146.355 174.135 ;
        RECT 146.645 173.965 146.815 174.135 ;
        RECT 147.105 173.965 147.275 174.135 ;
        RECT 147.565 173.965 147.735 174.135 ;
        RECT 148.025 173.965 148.195 174.135 ;
        RECT 148.485 173.965 148.655 174.135 ;
        RECT 148.945 173.965 149.115 174.135 ;
        RECT 149.405 173.965 149.575 174.135 ;
        RECT 149.865 173.965 150.035 174.135 ;
        RECT 42.225 173.455 42.395 173.625 ;
        RECT 45.445 173.455 45.615 173.625 ;
        RECT 42.225 172.435 42.395 172.605 ;
        RECT 43.605 172.775 43.775 172.945 ;
        RECT 43.145 171.755 43.315 171.925 ;
        RECT 46.285 173.115 46.455 173.285 ;
        RECT 47.285 173.115 47.455 173.285 ;
        RECT 47.745 172.775 47.915 172.945 ;
        RECT 50.045 173.455 50.215 173.625 ;
        RECT 51.425 173.455 51.595 173.625 ;
        RECT 49.125 172.775 49.295 172.945 ;
        RECT 50.045 172.775 50.215 172.945 ;
        RECT 50.505 172.775 50.675 172.945 ;
        RECT 46.365 171.755 46.535 171.925 ;
        RECT 48.665 171.755 48.835 171.925 ;
        RECT 52.345 173.455 52.515 173.625 ;
        RECT 53.265 172.775 53.435 172.945 ;
        RECT 54.185 172.775 54.355 172.945 ;
        RECT 55.105 171.755 55.275 171.925 ;
        RECT 56.485 172.775 56.655 172.945 ;
        RECT 55.565 172.095 55.735 172.265 ;
        RECT 63.845 172.435 64.015 172.605 ;
        RECT 64.765 173.115 64.935 173.285 ;
        RECT 64.765 172.435 64.935 172.605 ;
        RECT 66.145 172.775 66.315 172.945 ;
        RECT 66.605 172.775 66.775 172.945 ;
        RECT 65.225 172.095 65.395 172.265 ;
        RECT 65.685 171.755 65.855 171.925 ;
        RECT 67.065 171.755 67.235 171.925 ;
        RECT 68.445 172.775 68.615 172.945 ;
        RECT 70.285 173.455 70.455 173.625 ;
        RECT 67.985 171.755 68.155 171.925 ;
        RECT 69.825 172.435 69.995 172.605 ;
        RECT 72.585 172.775 72.755 172.945 ;
        RECT 69.365 172.095 69.535 172.265 ;
        RECT 70.285 171.755 70.455 171.925 ;
        RECT 71.205 172.095 71.375 172.265 ;
        RECT 73.965 172.435 74.135 172.605 ;
        RECT 73.505 171.755 73.675 171.925 ;
        RECT 74.450 172.095 74.620 172.265 ;
        RECT 74.845 172.435 75.015 172.605 ;
        RECT 75.300 172.775 75.470 172.945 ;
        RECT 76.035 172.435 76.205 172.605 ;
        RECT 76.550 172.095 76.720 172.265 ;
        RECT 78.120 172.095 78.290 172.265 ;
        RECT 78.555 172.435 78.725 172.605 ;
        RECT 86.385 172.775 86.555 172.945 ;
        RECT 87.305 172.775 87.475 172.945 ;
        RECT 88.225 172.775 88.395 172.945 ;
        RECT 89.145 172.775 89.315 172.945 ;
        RECT 89.605 172.775 89.775 172.945 ;
        RECT 80.865 172.095 81.035 172.265 ;
        RECT 86.845 172.095 87.015 172.265 ;
        RECT 90.985 172.775 91.155 172.945 ;
        RECT 91.905 171.755 92.075 171.925 ;
        RECT 92.365 171.755 92.535 171.925 ;
        RECT 93.285 172.435 93.455 172.605 ;
        RECT 93.745 172.435 93.915 172.605 ;
        RECT 94.205 172.435 94.375 172.605 ;
        RECT 94.665 172.775 94.835 172.945 ;
        RECT 99.725 172.775 99.895 172.945 ;
        RECT 103.405 173.455 103.575 173.625 ;
        RECT 100.645 172.775 100.815 172.945 ;
        RECT 102.485 172.775 102.655 172.945 ;
        RECT 101.105 172.435 101.275 172.605 ;
        RECT 103.865 172.775 104.035 172.945 ;
        RECT 104.785 172.775 104.955 172.945 ;
        RECT 106.165 172.775 106.335 172.945 ;
        RECT 107.545 172.775 107.715 172.945 ;
        RECT 104.325 171.755 104.495 171.925 ;
        RECT 106.625 171.755 106.795 171.925 ;
        RECT 108.465 171.755 108.635 171.925 ;
        RECT 116.285 172.775 116.455 172.945 ;
        RECT 119.965 172.775 120.135 172.945 ;
        RECT 120.885 172.775 121.055 172.945 ;
        RECT 121.345 172.775 121.515 172.945 ;
        RECT 117.205 172.095 117.375 172.265 ;
        RECT 119.965 172.095 120.135 172.265 ;
        RECT 139.745 173.455 139.915 173.625 ;
        RECT 138.825 172.775 138.995 172.945 ;
        RECT 141.125 172.775 141.295 172.945 ;
        RECT 137.905 171.755 138.075 171.925 ;
        RECT 141.585 171.755 141.755 171.925 ;
        RECT 142.045 172.775 142.215 172.945 ;
        RECT 143.425 172.775 143.595 172.945 ;
        RECT 142.505 171.755 142.675 171.925 ;
        RECT 36.245 171.245 36.415 171.415 ;
        RECT 36.705 171.245 36.875 171.415 ;
        RECT 37.165 171.245 37.335 171.415 ;
        RECT 37.625 171.245 37.795 171.415 ;
        RECT 38.085 171.245 38.255 171.415 ;
        RECT 38.545 171.245 38.715 171.415 ;
        RECT 39.005 171.245 39.175 171.415 ;
        RECT 39.465 171.245 39.635 171.415 ;
        RECT 39.925 171.245 40.095 171.415 ;
        RECT 40.385 171.245 40.555 171.415 ;
        RECT 40.845 171.245 41.015 171.415 ;
        RECT 41.305 171.245 41.475 171.415 ;
        RECT 41.765 171.245 41.935 171.415 ;
        RECT 42.225 171.245 42.395 171.415 ;
        RECT 42.685 171.245 42.855 171.415 ;
        RECT 43.145 171.245 43.315 171.415 ;
        RECT 43.605 171.245 43.775 171.415 ;
        RECT 44.065 171.245 44.235 171.415 ;
        RECT 44.525 171.245 44.695 171.415 ;
        RECT 44.985 171.245 45.155 171.415 ;
        RECT 45.445 171.245 45.615 171.415 ;
        RECT 45.905 171.245 46.075 171.415 ;
        RECT 46.365 171.245 46.535 171.415 ;
        RECT 46.825 171.245 46.995 171.415 ;
        RECT 47.285 171.245 47.455 171.415 ;
        RECT 47.745 171.245 47.915 171.415 ;
        RECT 48.205 171.245 48.375 171.415 ;
        RECT 48.665 171.245 48.835 171.415 ;
        RECT 49.125 171.245 49.295 171.415 ;
        RECT 49.585 171.245 49.755 171.415 ;
        RECT 50.045 171.245 50.215 171.415 ;
        RECT 50.505 171.245 50.675 171.415 ;
        RECT 50.965 171.245 51.135 171.415 ;
        RECT 51.425 171.245 51.595 171.415 ;
        RECT 51.885 171.245 52.055 171.415 ;
        RECT 52.345 171.245 52.515 171.415 ;
        RECT 52.805 171.245 52.975 171.415 ;
        RECT 53.265 171.245 53.435 171.415 ;
        RECT 53.725 171.245 53.895 171.415 ;
        RECT 54.185 171.245 54.355 171.415 ;
        RECT 54.645 171.245 54.815 171.415 ;
        RECT 55.105 171.245 55.275 171.415 ;
        RECT 55.565 171.245 55.735 171.415 ;
        RECT 56.025 171.245 56.195 171.415 ;
        RECT 56.485 171.245 56.655 171.415 ;
        RECT 56.945 171.245 57.115 171.415 ;
        RECT 57.405 171.245 57.575 171.415 ;
        RECT 57.865 171.245 58.035 171.415 ;
        RECT 58.325 171.245 58.495 171.415 ;
        RECT 58.785 171.245 58.955 171.415 ;
        RECT 59.245 171.245 59.415 171.415 ;
        RECT 59.705 171.245 59.875 171.415 ;
        RECT 60.165 171.245 60.335 171.415 ;
        RECT 60.625 171.245 60.795 171.415 ;
        RECT 61.085 171.245 61.255 171.415 ;
        RECT 61.545 171.245 61.715 171.415 ;
        RECT 62.005 171.245 62.175 171.415 ;
        RECT 62.465 171.245 62.635 171.415 ;
        RECT 62.925 171.245 63.095 171.415 ;
        RECT 63.385 171.245 63.555 171.415 ;
        RECT 63.845 171.245 64.015 171.415 ;
        RECT 64.305 171.245 64.475 171.415 ;
        RECT 64.765 171.245 64.935 171.415 ;
        RECT 65.225 171.245 65.395 171.415 ;
        RECT 65.685 171.245 65.855 171.415 ;
        RECT 66.145 171.245 66.315 171.415 ;
        RECT 66.605 171.245 66.775 171.415 ;
        RECT 67.065 171.245 67.235 171.415 ;
        RECT 67.525 171.245 67.695 171.415 ;
        RECT 67.985 171.245 68.155 171.415 ;
        RECT 68.445 171.245 68.615 171.415 ;
        RECT 68.905 171.245 69.075 171.415 ;
        RECT 69.365 171.245 69.535 171.415 ;
        RECT 69.825 171.245 69.995 171.415 ;
        RECT 70.285 171.245 70.455 171.415 ;
        RECT 70.745 171.245 70.915 171.415 ;
        RECT 71.205 171.245 71.375 171.415 ;
        RECT 71.665 171.245 71.835 171.415 ;
        RECT 72.125 171.245 72.295 171.415 ;
        RECT 72.585 171.245 72.755 171.415 ;
        RECT 73.045 171.245 73.215 171.415 ;
        RECT 73.505 171.245 73.675 171.415 ;
        RECT 73.965 171.245 74.135 171.415 ;
        RECT 74.425 171.245 74.595 171.415 ;
        RECT 74.885 171.245 75.055 171.415 ;
        RECT 75.345 171.245 75.515 171.415 ;
        RECT 75.805 171.245 75.975 171.415 ;
        RECT 76.265 171.245 76.435 171.415 ;
        RECT 76.725 171.245 76.895 171.415 ;
        RECT 77.185 171.245 77.355 171.415 ;
        RECT 77.645 171.245 77.815 171.415 ;
        RECT 78.105 171.245 78.275 171.415 ;
        RECT 78.565 171.245 78.735 171.415 ;
        RECT 79.025 171.245 79.195 171.415 ;
        RECT 79.485 171.245 79.655 171.415 ;
        RECT 79.945 171.245 80.115 171.415 ;
        RECT 80.405 171.245 80.575 171.415 ;
        RECT 80.865 171.245 81.035 171.415 ;
        RECT 81.325 171.245 81.495 171.415 ;
        RECT 81.785 171.245 81.955 171.415 ;
        RECT 82.245 171.245 82.415 171.415 ;
        RECT 82.705 171.245 82.875 171.415 ;
        RECT 83.165 171.245 83.335 171.415 ;
        RECT 83.625 171.245 83.795 171.415 ;
        RECT 84.085 171.245 84.255 171.415 ;
        RECT 84.545 171.245 84.715 171.415 ;
        RECT 85.005 171.245 85.175 171.415 ;
        RECT 85.465 171.245 85.635 171.415 ;
        RECT 85.925 171.245 86.095 171.415 ;
        RECT 86.385 171.245 86.555 171.415 ;
        RECT 86.845 171.245 87.015 171.415 ;
        RECT 87.305 171.245 87.475 171.415 ;
        RECT 87.765 171.245 87.935 171.415 ;
        RECT 88.225 171.245 88.395 171.415 ;
        RECT 88.685 171.245 88.855 171.415 ;
        RECT 89.145 171.245 89.315 171.415 ;
        RECT 89.605 171.245 89.775 171.415 ;
        RECT 90.065 171.245 90.235 171.415 ;
        RECT 90.525 171.245 90.695 171.415 ;
        RECT 90.985 171.245 91.155 171.415 ;
        RECT 91.445 171.245 91.615 171.415 ;
        RECT 91.905 171.245 92.075 171.415 ;
        RECT 92.365 171.245 92.535 171.415 ;
        RECT 92.825 171.245 92.995 171.415 ;
        RECT 93.285 171.245 93.455 171.415 ;
        RECT 93.745 171.245 93.915 171.415 ;
        RECT 94.205 171.245 94.375 171.415 ;
        RECT 94.665 171.245 94.835 171.415 ;
        RECT 95.125 171.245 95.295 171.415 ;
        RECT 95.585 171.245 95.755 171.415 ;
        RECT 96.045 171.245 96.215 171.415 ;
        RECT 96.505 171.245 96.675 171.415 ;
        RECT 96.965 171.245 97.135 171.415 ;
        RECT 97.425 171.245 97.595 171.415 ;
        RECT 97.885 171.245 98.055 171.415 ;
        RECT 98.345 171.245 98.515 171.415 ;
        RECT 98.805 171.245 98.975 171.415 ;
        RECT 99.265 171.245 99.435 171.415 ;
        RECT 99.725 171.245 99.895 171.415 ;
        RECT 100.185 171.245 100.355 171.415 ;
        RECT 100.645 171.245 100.815 171.415 ;
        RECT 101.105 171.245 101.275 171.415 ;
        RECT 101.565 171.245 101.735 171.415 ;
        RECT 102.025 171.245 102.195 171.415 ;
        RECT 102.485 171.245 102.655 171.415 ;
        RECT 102.945 171.245 103.115 171.415 ;
        RECT 103.405 171.245 103.575 171.415 ;
        RECT 103.865 171.245 104.035 171.415 ;
        RECT 104.325 171.245 104.495 171.415 ;
        RECT 104.785 171.245 104.955 171.415 ;
        RECT 105.245 171.245 105.415 171.415 ;
        RECT 105.705 171.245 105.875 171.415 ;
        RECT 106.165 171.245 106.335 171.415 ;
        RECT 106.625 171.245 106.795 171.415 ;
        RECT 107.085 171.245 107.255 171.415 ;
        RECT 107.545 171.245 107.715 171.415 ;
        RECT 108.005 171.245 108.175 171.415 ;
        RECT 108.465 171.245 108.635 171.415 ;
        RECT 108.925 171.245 109.095 171.415 ;
        RECT 109.385 171.245 109.555 171.415 ;
        RECT 109.845 171.245 110.015 171.415 ;
        RECT 110.305 171.245 110.475 171.415 ;
        RECT 110.765 171.245 110.935 171.415 ;
        RECT 111.225 171.245 111.395 171.415 ;
        RECT 111.685 171.245 111.855 171.415 ;
        RECT 112.145 171.245 112.315 171.415 ;
        RECT 112.605 171.245 112.775 171.415 ;
        RECT 113.065 171.245 113.235 171.415 ;
        RECT 113.525 171.245 113.695 171.415 ;
        RECT 113.985 171.245 114.155 171.415 ;
        RECT 114.445 171.245 114.615 171.415 ;
        RECT 114.905 171.245 115.075 171.415 ;
        RECT 115.365 171.245 115.535 171.415 ;
        RECT 115.825 171.245 115.995 171.415 ;
        RECT 116.285 171.245 116.455 171.415 ;
        RECT 116.745 171.245 116.915 171.415 ;
        RECT 117.205 171.245 117.375 171.415 ;
        RECT 117.665 171.245 117.835 171.415 ;
        RECT 118.125 171.245 118.295 171.415 ;
        RECT 118.585 171.245 118.755 171.415 ;
        RECT 119.045 171.245 119.215 171.415 ;
        RECT 119.505 171.245 119.675 171.415 ;
        RECT 119.965 171.245 120.135 171.415 ;
        RECT 120.425 171.245 120.595 171.415 ;
        RECT 120.885 171.245 121.055 171.415 ;
        RECT 121.345 171.245 121.515 171.415 ;
        RECT 121.805 171.245 121.975 171.415 ;
        RECT 122.265 171.245 122.435 171.415 ;
        RECT 122.725 171.245 122.895 171.415 ;
        RECT 123.185 171.245 123.355 171.415 ;
        RECT 123.645 171.245 123.815 171.415 ;
        RECT 124.105 171.245 124.275 171.415 ;
        RECT 124.565 171.245 124.735 171.415 ;
        RECT 125.025 171.245 125.195 171.415 ;
        RECT 125.485 171.245 125.655 171.415 ;
        RECT 125.945 171.245 126.115 171.415 ;
        RECT 126.405 171.245 126.575 171.415 ;
        RECT 126.865 171.245 127.035 171.415 ;
        RECT 127.325 171.245 127.495 171.415 ;
        RECT 127.785 171.245 127.955 171.415 ;
        RECT 128.245 171.245 128.415 171.415 ;
        RECT 128.705 171.245 128.875 171.415 ;
        RECT 129.165 171.245 129.335 171.415 ;
        RECT 129.625 171.245 129.795 171.415 ;
        RECT 130.085 171.245 130.255 171.415 ;
        RECT 130.545 171.245 130.715 171.415 ;
        RECT 131.005 171.245 131.175 171.415 ;
        RECT 131.465 171.245 131.635 171.415 ;
        RECT 131.925 171.245 132.095 171.415 ;
        RECT 132.385 171.245 132.555 171.415 ;
        RECT 132.845 171.245 133.015 171.415 ;
        RECT 133.305 171.245 133.475 171.415 ;
        RECT 133.765 171.245 133.935 171.415 ;
        RECT 134.225 171.245 134.395 171.415 ;
        RECT 134.685 171.245 134.855 171.415 ;
        RECT 135.145 171.245 135.315 171.415 ;
        RECT 135.605 171.245 135.775 171.415 ;
        RECT 136.065 171.245 136.235 171.415 ;
        RECT 136.525 171.245 136.695 171.415 ;
        RECT 136.985 171.245 137.155 171.415 ;
        RECT 137.445 171.245 137.615 171.415 ;
        RECT 137.905 171.245 138.075 171.415 ;
        RECT 138.365 171.245 138.535 171.415 ;
        RECT 138.825 171.245 138.995 171.415 ;
        RECT 139.285 171.245 139.455 171.415 ;
        RECT 139.745 171.245 139.915 171.415 ;
        RECT 140.205 171.245 140.375 171.415 ;
        RECT 140.665 171.245 140.835 171.415 ;
        RECT 141.125 171.245 141.295 171.415 ;
        RECT 141.585 171.245 141.755 171.415 ;
        RECT 142.045 171.245 142.215 171.415 ;
        RECT 142.505 171.245 142.675 171.415 ;
        RECT 142.965 171.245 143.135 171.415 ;
        RECT 143.425 171.245 143.595 171.415 ;
        RECT 143.885 171.245 144.055 171.415 ;
        RECT 144.345 171.245 144.515 171.415 ;
        RECT 144.805 171.245 144.975 171.415 ;
        RECT 145.265 171.245 145.435 171.415 ;
        RECT 145.725 171.245 145.895 171.415 ;
        RECT 146.185 171.245 146.355 171.415 ;
        RECT 146.645 171.245 146.815 171.415 ;
        RECT 147.105 171.245 147.275 171.415 ;
        RECT 147.565 171.245 147.735 171.415 ;
        RECT 148.025 171.245 148.195 171.415 ;
        RECT 148.485 171.245 148.655 171.415 ;
        RECT 148.945 171.245 149.115 171.415 ;
        RECT 149.405 171.245 149.575 171.415 ;
        RECT 149.865 171.245 150.035 171.415 ;
        RECT 41.305 170.395 41.475 170.565 ;
        RECT 44.525 170.735 44.695 170.905 ;
        RECT 40.845 169.715 41.015 169.885 ;
        RECT 42.225 170.055 42.395 170.225 ;
        RECT 43.145 169.715 43.315 169.885 ;
        RECT 43.605 169.715 43.775 169.885 ;
        RECT 42.225 169.375 42.395 169.545 ;
        RECT 46.365 170.735 46.535 170.905 ;
        RECT 47.285 170.735 47.455 170.905 ;
        RECT 44.985 169.715 45.155 169.885 ;
        RECT 45.905 169.715 46.075 169.885 ;
        RECT 45.445 169.035 45.615 169.205 ;
        RECT 47.155 169.035 47.325 169.205 ;
        RECT 48.205 169.375 48.375 169.545 ;
        RECT 64.305 170.735 64.475 170.905 ;
        RECT 63.845 170.395 64.015 170.565 ;
        RECT 61.085 169.715 61.255 169.885 ;
        RECT 62.465 170.055 62.635 170.225 ;
        RECT 63.385 170.055 63.555 170.225 ;
        RECT 62.005 169.035 62.175 169.205 ;
        RECT 65.685 170.735 65.855 170.905 ;
        RECT 63.385 169.375 63.555 169.545 ;
        RECT 64.765 169.715 64.935 169.885 ;
        RECT 65.225 169.715 65.395 169.885 ;
        RECT 66.605 170.735 66.775 170.905 ;
        RECT 68.905 170.735 69.075 170.905 ;
        RECT 67.065 169.375 67.235 169.545 ;
        RECT 67.985 170.395 68.155 170.565 ;
        RECT 68.445 170.055 68.615 170.225 ;
        RECT 68.905 169.035 69.075 169.205 ;
        RECT 69.825 169.035 69.995 169.205 ;
        RECT 76.265 170.735 76.435 170.905 ;
        RECT 75.345 169.035 75.515 169.205 ;
        RECT 76.265 169.035 76.435 169.205 ;
        RECT 78.105 170.395 78.275 170.565 ;
        RECT 88.685 169.715 88.855 169.885 ;
        RECT 89.145 170.055 89.315 170.225 ;
        RECT 89.605 170.055 89.775 170.225 ;
        RECT 90.065 170.055 90.235 170.225 ;
        RECT 91.440 169.715 91.610 169.885 ;
        RECT 91.900 170.055 92.070 170.225 ;
        RECT 92.415 169.715 92.585 169.885 ;
        RECT 92.825 170.055 92.995 170.225 ;
        RECT 87.765 169.035 87.935 169.205 ;
        RECT 95.125 169.375 95.295 169.545 ;
        RECT 93.745 169.035 93.915 169.205 ;
        RECT 96.045 169.035 96.215 169.205 ;
        RECT 102.945 170.395 103.115 170.565 ;
        RECT 102.025 169.715 102.195 169.885 ;
        RECT 103.405 169.715 103.575 169.885 ;
        RECT 101.105 169.035 101.275 169.205 ;
        RECT 107.545 169.715 107.715 169.885 ;
        RECT 108.465 169.715 108.635 169.885 ;
        RECT 108.005 169.375 108.175 169.545 ;
        RECT 109.385 169.715 109.555 169.885 ;
        RECT 109.845 170.055 110.015 170.225 ;
        RECT 110.305 169.715 110.475 169.885 ;
        RECT 110.765 169.715 110.935 169.885 ;
        RECT 113.985 169.715 114.155 169.885 ;
        RECT 113.065 169.375 113.235 169.545 ;
        RECT 111.685 169.035 111.855 169.205 ;
        RECT 115.365 169.715 115.535 169.885 ;
        RECT 114.445 169.035 114.615 169.205 ;
        RECT 123.185 169.715 123.355 169.885 ;
        RECT 124.105 169.715 124.275 169.885 ;
        RECT 123.645 169.375 123.815 169.545 ;
        RECT 126.865 169.715 127.035 169.885 ;
        RECT 127.785 169.375 127.955 169.545 ;
        RECT 128.705 169.715 128.875 169.885 ;
        RECT 128.245 169.375 128.415 169.545 ;
        RECT 137.905 170.735 138.075 170.905 ;
        RECT 141.150 170.395 141.320 170.565 ;
        RECT 139.285 169.715 139.455 169.885 ;
        RECT 129.625 169.035 129.795 169.205 ;
        RECT 137.905 169.375 138.075 169.545 ;
        RECT 140.665 170.055 140.835 170.225 ;
        RECT 140.205 169.035 140.375 169.205 ;
        RECT 141.545 170.055 141.715 170.225 ;
        RECT 141.890 169.375 142.060 169.545 ;
        RECT 143.250 170.395 143.420 170.565 ;
        RECT 142.735 170.055 142.905 170.225 ;
        RECT 144.820 170.395 144.990 170.565 ;
        RECT 145.255 170.055 145.425 170.225 ;
        RECT 147.565 170.735 147.735 170.905 ;
        RECT 36.245 168.525 36.415 168.695 ;
        RECT 36.705 168.525 36.875 168.695 ;
        RECT 37.165 168.525 37.335 168.695 ;
        RECT 37.625 168.525 37.795 168.695 ;
        RECT 38.085 168.525 38.255 168.695 ;
        RECT 38.545 168.525 38.715 168.695 ;
        RECT 39.005 168.525 39.175 168.695 ;
        RECT 39.465 168.525 39.635 168.695 ;
        RECT 39.925 168.525 40.095 168.695 ;
        RECT 40.385 168.525 40.555 168.695 ;
        RECT 40.845 168.525 41.015 168.695 ;
        RECT 41.305 168.525 41.475 168.695 ;
        RECT 41.765 168.525 41.935 168.695 ;
        RECT 42.225 168.525 42.395 168.695 ;
        RECT 42.685 168.525 42.855 168.695 ;
        RECT 43.145 168.525 43.315 168.695 ;
        RECT 43.605 168.525 43.775 168.695 ;
        RECT 44.065 168.525 44.235 168.695 ;
        RECT 44.525 168.525 44.695 168.695 ;
        RECT 44.985 168.525 45.155 168.695 ;
        RECT 45.445 168.525 45.615 168.695 ;
        RECT 45.905 168.525 46.075 168.695 ;
        RECT 46.365 168.525 46.535 168.695 ;
        RECT 46.825 168.525 46.995 168.695 ;
        RECT 47.285 168.525 47.455 168.695 ;
        RECT 47.745 168.525 47.915 168.695 ;
        RECT 48.205 168.525 48.375 168.695 ;
        RECT 48.665 168.525 48.835 168.695 ;
        RECT 49.125 168.525 49.295 168.695 ;
        RECT 49.585 168.525 49.755 168.695 ;
        RECT 50.045 168.525 50.215 168.695 ;
        RECT 50.505 168.525 50.675 168.695 ;
        RECT 50.965 168.525 51.135 168.695 ;
        RECT 51.425 168.525 51.595 168.695 ;
        RECT 51.885 168.525 52.055 168.695 ;
        RECT 52.345 168.525 52.515 168.695 ;
        RECT 52.805 168.525 52.975 168.695 ;
        RECT 53.265 168.525 53.435 168.695 ;
        RECT 53.725 168.525 53.895 168.695 ;
        RECT 54.185 168.525 54.355 168.695 ;
        RECT 54.645 168.525 54.815 168.695 ;
        RECT 55.105 168.525 55.275 168.695 ;
        RECT 55.565 168.525 55.735 168.695 ;
        RECT 56.025 168.525 56.195 168.695 ;
        RECT 56.485 168.525 56.655 168.695 ;
        RECT 56.945 168.525 57.115 168.695 ;
        RECT 57.405 168.525 57.575 168.695 ;
        RECT 57.865 168.525 58.035 168.695 ;
        RECT 58.325 168.525 58.495 168.695 ;
        RECT 58.785 168.525 58.955 168.695 ;
        RECT 59.245 168.525 59.415 168.695 ;
        RECT 59.705 168.525 59.875 168.695 ;
        RECT 60.165 168.525 60.335 168.695 ;
        RECT 60.625 168.525 60.795 168.695 ;
        RECT 61.085 168.525 61.255 168.695 ;
        RECT 61.545 168.525 61.715 168.695 ;
        RECT 62.005 168.525 62.175 168.695 ;
        RECT 62.465 168.525 62.635 168.695 ;
        RECT 62.925 168.525 63.095 168.695 ;
        RECT 63.385 168.525 63.555 168.695 ;
        RECT 63.845 168.525 64.015 168.695 ;
        RECT 64.305 168.525 64.475 168.695 ;
        RECT 64.765 168.525 64.935 168.695 ;
        RECT 65.225 168.525 65.395 168.695 ;
        RECT 65.685 168.525 65.855 168.695 ;
        RECT 66.145 168.525 66.315 168.695 ;
        RECT 66.605 168.525 66.775 168.695 ;
        RECT 67.065 168.525 67.235 168.695 ;
        RECT 67.525 168.525 67.695 168.695 ;
        RECT 67.985 168.525 68.155 168.695 ;
        RECT 68.445 168.525 68.615 168.695 ;
        RECT 68.905 168.525 69.075 168.695 ;
        RECT 69.365 168.525 69.535 168.695 ;
        RECT 69.825 168.525 69.995 168.695 ;
        RECT 70.285 168.525 70.455 168.695 ;
        RECT 70.745 168.525 70.915 168.695 ;
        RECT 71.205 168.525 71.375 168.695 ;
        RECT 71.665 168.525 71.835 168.695 ;
        RECT 72.125 168.525 72.295 168.695 ;
        RECT 72.585 168.525 72.755 168.695 ;
        RECT 73.045 168.525 73.215 168.695 ;
        RECT 73.505 168.525 73.675 168.695 ;
        RECT 73.965 168.525 74.135 168.695 ;
        RECT 74.425 168.525 74.595 168.695 ;
        RECT 74.885 168.525 75.055 168.695 ;
        RECT 75.345 168.525 75.515 168.695 ;
        RECT 75.805 168.525 75.975 168.695 ;
        RECT 76.265 168.525 76.435 168.695 ;
        RECT 76.725 168.525 76.895 168.695 ;
        RECT 77.185 168.525 77.355 168.695 ;
        RECT 77.645 168.525 77.815 168.695 ;
        RECT 78.105 168.525 78.275 168.695 ;
        RECT 78.565 168.525 78.735 168.695 ;
        RECT 79.025 168.525 79.195 168.695 ;
        RECT 79.485 168.525 79.655 168.695 ;
        RECT 79.945 168.525 80.115 168.695 ;
        RECT 80.405 168.525 80.575 168.695 ;
        RECT 80.865 168.525 81.035 168.695 ;
        RECT 81.325 168.525 81.495 168.695 ;
        RECT 81.785 168.525 81.955 168.695 ;
        RECT 82.245 168.525 82.415 168.695 ;
        RECT 82.705 168.525 82.875 168.695 ;
        RECT 83.165 168.525 83.335 168.695 ;
        RECT 83.625 168.525 83.795 168.695 ;
        RECT 84.085 168.525 84.255 168.695 ;
        RECT 84.545 168.525 84.715 168.695 ;
        RECT 85.005 168.525 85.175 168.695 ;
        RECT 85.465 168.525 85.635 168.695 ;
        RECT 85.925 168.525 86.095 168.695 ;
        RECT 86.385 168.525 86.555 168.695 ;
        RECT 86.845 168.525 87.015 168.695 ;
        RECT 87.305 168.525 87.475 168.695 ;
        RECT 87.765 168.525 87.935 168.695 ;
        RECT 88.225 168.525 88.395 168.695 ;
        RECT 88.685 168.525 88.855 168.695 ;
        RECT 89.145 168.525 89.315 168.695 ;
        RECT 89.605 168.525 89.775 168.695 ;
        RECT 90.065 168.525 90.235 168.695 ;
        RECT 90.525 168.525 90.695 168.695 ;
        RECT 90.985 168.525 91.155 168.695 ;
        RECT 91.445 168.525 91.615 168.695 ;
        RECT 91.905 168.525 92.075 168.695 ;
        RECT 92.365 168.525 92.535 168.695 ;
        RECT 92.825 168.525 92.995 168.695 ;
        RECT 93.285 168.525 93.455 168.695 ;
        RECT 93.745 168.525 93.915 168.695 ;
        RECT 94.205 168.525 94.375 168.695 ;
        RECT 94.665 168.525 94.835 168.695 ;
        RECT 95.125 168.525 95.295 168.695 ;
        RECT 95.585 168.525 95.755 168.695 ;
        RECT 96.045 168.525 96.215 168.695 ;
        RECT 96.505 168.525 96.675 168.695 ;
        RECT 96.965 168.525 97.135 168.695 ;
        RECT 97.425 168.525 97.595 168.695 ;
        RECT 97.885 168.525 98.055 168.695 ;
        RECT 98.345 168.525 98.515 168.695 ;
        RECT 98.805 168.525 98.975 168.695 ;
        RECT 99.265 168.525 99.435 168.695 ;
        RECT 99.725 168.525 99.895 168.695 ;
        RECT 100.185 168.525 100.355 168.695 ;
        RECT 100.645 168.525 100.815 168.695 ;
        RECT 101.105 168.525 101.275 168.695 ;
        RECT 101.565 168.525 101.735 168.695 ;
        RECT 102.025 168.525 102.195 168.695 ;
        RECT 102.485 168.525 102.655 168.695 ;
        RECT 102.945 168.525 103.115 168.695 ;
        RECT 103.405 168.525 103.575 168.695 ;
        RECT 103.865 168.525 104.035 168.695 ;
        RECT 104.325 168.525 104.495 168.695 ;
        RECT 104.785 168.525 104.955 168.695 ;
        RECT 105.245 168.525 105.415 168.695 ;
        RECT 105.705 168.525 105.875 168.695 ;
        RECT 106.165 168.525 106.335 168.695 ;
        RECT 106.625 168.525 106.795 168.695 ;
        RECT 107.085 168.525 107.255 168.695 ;
        RECT 107.545 168.525 107.715 168.695 ;
        RECT 108.005 168.525 108.175 168.695 ;
        RECT 108.465 168.525 108.635 168.695 ;
        RECT 108.925 168.525 109.095 168.695 ;
        RECT 109.385 168.525 109.555 168.695 ;
        RECT 109.845 168.525 110.015 168.695 ;
        RECT 110.305 168.525 110.475 168.695 ;
        RECT 110.765 168.525 110.935 168.695 ;
        RECT 111.225 168.525 111.395 168.695 ;
        RECT 111.685 168.525 111.855 168.695 ;
        RECT 112.145 168.525 112.315 168.695 ;
        RECT 112.605 168.525 112.775 168.695 ;
        RECT 113.065 168.525 113.235 168.695 ;
        RECT 113.525 168.525 113.695 168.695 ;
        RECT 113.985 168.525 114.155 168.695 ;
        RECT 114.445 168.525 114.615 168.695 ;
        RECT 114.905 168.525 115.075 168.695 ;
        RECT 115.365 168.525 115.535 168.695 ;
        RECT 115.825 168.525 115.995 168.695 ;
        RECT 116.285 168.525 116.455 168.695 ;
        RECT 116.745 168.525 116.915 168.695 ;
        RECT 117.205 168.525 117.375 168.695 ;
        RECT 117.665 168.525 117.835 168.695 ;
        RECT 118.125 168.525 118.295 168.695 ;
        RECT 118.585 168.525 118.755 168.695 ;
        RECT 119.045 168.525 119.215 168.695 ;
        RECT 119.505 168.525 119.675 168.695 ;
        RECT 119.965 168.525 120.135 168.695 ;
        RECT 120.425 168.525 120.595 168.695 ;
        RECT 120.885 168.525 121.055 168.695 ;
        RECT 121.345 168.525 121.515 168.695 ;
        RECT 121.805 168.525 121.975 168.695 ;
        RECT 122.265 168.525 122.435 168.695 ;
        RECT 122.725 168.525 122.895 168.695 ;
        RECT 123.185 168.525 123.355 168.695 ;
        RECT 123.645 168.525 123.815 168.695 ;
        RECT 124.105 168.525 124.275 168.695 ;
        RECT 124.565 168.525 124.735 168.695 ;
        RECT 125.025 168.525 125.195 168.695 ;
        RECT 125.485 168.525 125.655 168.695 ;
        RECT 125.945 168.525 126.115 168.695 ;
        RECT 126.405 168.525 126.575 168.695 ;
        RECT 126.865 168.525 127.035 168.695 ;
        RECT 127.325 168.525 127.495 168.695 ;
        RECT 127.785 168.525 127.955 168.695 ;
        RECT 128.245 168.525 128.415 168.695 ;
        RECT 128.705 168.525 128.875 168.695 ;
        RECT 129.165 168.525 129.335 168.695 ;
        RECT 129.625 168.525 129.795 168.695 ;
        RECT 130.085 168.525 130.255 168.695 ;
        RECT 130.545 168.525 130.715 168.695 ;
        RECT 131.005 168.525 131.175 168.695 ;
        RECT 131.465 168.525 131.635 168.695 ;
        RECT 131.925 168.525 132.095 168.695 ;
        RECT 132.385 168.525 132.555 168.695 ;
        RECT 132.845 168.525 133.015 168.695 ;
        RECT 133.305 168.525 133.475 168.695 ;
        RECT 133.765 168.525 133.935 168.695 ;
        RECT 134.225 168.525 134.395 168.695 ;
        RECT 134.685 168.525 134.855 168.695 ;
        RECT 135.145 168.525 135.315 168.695 ;
        RECT 135.605 168.525 135.775 168.695 ;
        RECT 136.065 168.525 136.235 168.695 ;
        RECT 136.525 168.525 136.695 168.695 ;
        RECT 136.985 168.525 137.155 168.695 ;
        RECT 137.445 168.525 137.615 168.695 ;
        RECT 137.905 168.525 138.075 168.695 ;
        RECT 138.365 168.525 138.535 168.695 ;
        RECT 138.825 168.525 138.995 168.695 ;
        RECT 139.285 168.525 139.455 168.695 ;
        RECT 139.745 168.525 139.915 168.695 ;
        RECT 140.205 168.525 140.375 168.695 ;
        RECT 140.665 168.525 140.835 168.695 ;
        RECT 141.125 168.525 141.295 168.695 ;
        RECT 141.585 168.525 141.755 168.695 ;
        RECT 142.045 168.525 142.215 168.695 ;
        RECT 142.505 168.525 142.675 168.695 ;
        RECT 142.965 168.525 143.135 168.695 ;
        RECT 143.425 168.525 143.595 168.695 ;
        RECT 143.885 168.525 144.055 168.695 ;
        RECT 144.345 168.525 144.515 168.695 ;
        RECT 144.805 168.525 144.975 168.695 ;
        RECT 145.265 168.525 145.435 168.695 ;
        RECT 145.725 168.525 145.895 168.695 ;
        RECT 146.185 168.525 146.355 168.695 ;
        RECT 146.645 168.525 146.815 168.695 ;
        RECT 147.105 168.525 147.275 168.695 ;
        RECT 147.565 168.525 147.735 168.695 ;
        RECT 148.025 168.525 148.195 168.695 ;
        RECT 148.485 168.525 148.655 168.695 ;
        RECT 148.945 168.525 149.115 168.695 ;
        RECT 149.405 168.525 149.575 168.695 ;
        RECT 149.865 168.525 150.035 168.695 ;
        RECT 41.765 166.995 41.935 167.165 ;
        RECT 43.605 167.675 43.775 167.845 ;
        RECT 44.985 167.335 45.155 167.505 ;
        RECT 43.605 166.315 43.775 166.485 ;
        RECT 44.525 166.315 44.695 166.485 ;
        RECT 45.470 166.655 45.640 166.825 ;
        RECT 45.865 166.995 46.035 167.165 ;
        RECT 46.265 167.335 46.435 167.505 ;
        RECT 47.055 166.995 47.225 167.165 ;
        RECT 47.570 166.655 47.740 166.825 ;
        RECT 49.140 166.655 49.310 166.825 ;
        RECT 49.575 166.995 49.745 167.165 ;
        RECT 51.885 166.315 52.055 166.485 ;
        RECT 57.865 166.315 58.035 166.485 ;
        RECT 58.785 166.995 58.955 167.165 ;
        RECT 59.245 166.995 59.415 167.165 ;
        RECT 59.705 166.995 59.875 167.165 ;
        RECT 60.165 166.995 60.335 167.165 ;
        RECT 62.465 167.335 62.635 167.505 ;
        RECT 62.950 166.655 63.120 166.825 ;
        RECT 63.345 166.995 63.515 167.165 ;
        RECT 63.745 167.335 63.915 167.505 ;
        RECT 64.535 166.995 64.705 167.165 ;
        RECT 65.050 166.655 65.220 166.825 ;
        RECT 66.620 166.655 66.790 166.825 ;
        RECT 67.055 166.995 67.225 167.165 ;
        RECT 71.205 167.335 71.375 167.505 ;
        RECT 69.365 166.315 69.535 166.485 ;
        RECT 72.125 166.655 72.295 166.825 ;
        RECT 72.585 167.335 72.755 167.505 ;
        RECT 73.505 167.675 73.675 167.845 ;
        RECT 73.965 168.015 74.135 168.185 ;
        RECT 75.345 168.015 75.515 168.185 ;
        RECT 74.425 167.335 74.595 167.505 ;
        RECT 75.805 168.015 75.975 168.185 ;
        RECT 76.725 167.335 76.895 167.505 ;
        RECT 77.185 166.995 77.355 167.165 ;
        RECT 77.645 166.995 77.815 167.165 ;
        RECT 78.105 166.995 78.275 167.165 ;
        RECT 79.025 167.335 79.195 167.505 ;
        RECT 79.485 166.995 79.655 167.165 ;
        RECT 87.305 167.335 87.475 167.505 ;
        RECT 88.225 167.335 88.395 167.505 ;
        RECT 86.385 166.315 86.555 166.485 ;
        RECT 91.445 168.015 91.615 168.185 ;
        RECT 89.145 167.335 89.315 167.505 ;
        RECT 89.605 167.335 89.775 167.505 ;
        RECT 90.065 167.335 90.235 167.505 ;
        RECT 94.275 166.995 94.445 167.165 ;
        RECT 94.665 167.335 94.835 167.505 ;
        RECT 95.125 166.995 95.295 167.165 ;
        RECT 95.585 167.335 95.755 167.505 ;
        RECT 96.965 167.335 97.135 167.505 ;
        RECT 97.885 167.335 98.055 167.505 ;
        RECT 99.725 167.335 99.895 167.505 ;
        RECT 100.645 167.335 100.815 167.505 ;
        RECT 96.505 166.315 96.675 166.485 ;
        RECT 98.345 166.995 98.515 167.165 ;
        RECT 102.025 167.335 102.195 167.505 ;
        RECT 101.105 166.655 101.275 166.825 ;
        RECT 102.945 166.315 103.115 166.485 ;
        RECT 110.765 168.015 110.935 168.185 ;
        RECT 110.305 167.335 110.475 167.505 ;
        RECT 109.385 166.315 109.555 166.485 ;
        RECT 111.685 167.335 111.855 167.505 ;
        RECT 118.585 167.335 118.755 167.505 ;
        RECT 119.045 167.335 119.215 167.505 ;
        RECT 117.665 166.315 117.835 166.485 ;
        RECT 121.805 168.015 121.975 168.185 ;
        RECT 121.345 167.335 121.515 167.505 ;
        RECT 122.265 167.335 122.435 167.505 ;
        RECT 125.945 167.675 126.115 167.845 ;
        RECT 123.645 167.335 123.815 167.505 ;
        RECT 125.025 167.335 125.195 167.505 ;
        RECT 126.405 167.335 126.575 167.505 ;
        RECT 126.865 167.335 127.035 167.505 ;
        RECT 119.965 166.315 120.135 166.485 ;
        RECT 122.725 166.995 122.895 167.165 ;
        RECT 124.565 166.995 124.735 167.165 ;
        RECT 128.705 167.675 128.875 167.845 ;
        RECT 128.245 167.335 128.415 167.505 ;
        RECT 129.165 167.335 129.335 167.505 ;
        RECT 131.925 167.335 132.095 167.505 ;
        RECT 132.410 166.655 132.580 166.825 ;
        RECT 132.805 166.995 132.975 167.165 ;
        RECT 133.150 167.675 133.320 167.845 ;
        RECT 133.995 166.995 134.165 167.165 ;
        RECT 134.510 166.655 134.680 166.825 ;
        RECT 136.080 166.655 136.250 166.825 ;
        RECT 136.515 166.995 136.685 167.165 ;
        RECT 138.825 168.015 138.995 168.185 ;
        RECT 143.885 168.015 144.055 168.185 ;
        RECT 141.125 167.335 141.295 167.505 ;
        RECT 140.665 166.995 140.835 167.165 ;
        RECT 142.965 167.335 143.135 167.505 ;
        RECT 144.345 167.335 144.515 167.505 ;
        RECT 142.965 166.315 143.135 166.485 ;
        RECT 145.265 166.655 145.435 166.825 ;
        RECT 36.245 165.805 36.415 165.975 ;
        RECT 36.705 165.805 36.875 165.975 ;
        RECT 37.165 165.805 37.335 165.975 ;
        RECT 37.625 165.805 37.795 165.975 ;
        RECT 38.085 165.805 38.255 165.975 ;
        RECT 38.545 165.805 38.715 165.975 ;
        RECT 39.005 165.805 39.175 165.975 ;
        RECT 39.465 165.805 39.635 165.975 ;
        RECT 39.925 165.805 40.095 165.975 ;
        RECT 40.385 165.805 40.555 165.975 ;
        RECT 40.845 165.805 41.015 165.975 ;
        RECT 41.305 165.805 41.475 165.975 ;
        RECT 41.765 165.805 41.935 165.975 ;
        RECT 42.225 165.805 42.395 165.975 ;
        RECT 42.685 165.805 42.855 165.975 ;
        RECT 43.145 165.805 43.315 165.975 ;
        RECT 43.605 165.805 43.775 165.975 ;
        RECT 44.065 165.805 44.235 165.975 ;
        RECT 44.525 165.805 44.695 165.975 ;
        RECT 44.985 165.805 45.155 165.975 ;
        RECT 45.445 165.805 45.615 165.975 ;
        RECT 45.905 165.805 46.075 165.975 ;
        RECT 46.365 165.805 46.535 165.975 ;
        RECT 46.825 165.805 46.995 165.975 ;
        RECT 47.285 165.805 47.455 165.975 ;
        RECT 47.745 165.805 47.915 165.975 ;
        RECT 48.205 165.805 48.375 165.975 ;
        RECT 48.665 165.805 48.835 165.975 ;
        RECT 49.125 165.805 49.295 165.975 ;
        RECT 49.585 165.805 49.755 165.975 ;
        RECT 50.045 165.805 50.215 165.975 ;
        RECT 50.505 165.805 50.675 165.975 ;
        RECT 50.965 165.805 51.135 165.975 ;
        RECT 51.425 165.805 51.595 165.975 ;
        RECT 51.885 165.805 52.055 165.975 ;
        RECT 52.345 165.805 52.515 165.975 ;
        RECT 52.805 165.805 52.975 165.975 ;
        RECT 53.265 165.805 53.435 165.975 ;
        RECT 53.725 165.805 53.895 165.975 ;
        RECT 54.185 165.805 54.355 165.975 ;
        RECT 54.645 165.805 54.815 165.975 ;
        RECT 55.105 165.805 55.275 165.975 ;
        RECT 55.565 165.805 55.735 165.975 ;
        RECT 56.025 165.805 56.195 165.975 ;
        RECT 56.485 165.805 56.655 165.975 ;
        RECT 56.945 165.805 57.115 165.975 ;
        RECT 57.405 165.805 57.575 165.975 ;
        RECT 57.865 165.805 58.035 165.975 ;
        RECT 58.325 165.805 58.495 165.975 ;
        RECT 58.785 165.805 58.955 165.975 ;
        RECT 59.245 165.805 59.415 165.975 ;
        RECT 59.705 165.805 59.875 165.975 ;
        RECT 60.165 165.805 60.335 165.975 ;
        RECT 60.625 165.805 60.795 165.975 ;
        RECT 61.085 165.805 61.255 165.975 ;
        RECT 61.545 165.805 61.715 165.975 ;
        RECT 62.005 165.805 62.175 165.975 ;
        RECT 62.465 165.805 62.635 165.975 ;
        RECT 62.925 165.805 63.095 165.975 ;
        RECT 63.385 165.805 63.555 165.975 ;
        RECT 63.845 165.805 64.015 165.975 ;
        RECT 64.305 165.805 64.475 165.975 ;
        RECT 64.765 165.805 64.935 165.975 ;
        RECT 65.225 165.805 65.395 165.975 ;
        RECT 65.685 165.805 65.855 165.975 ;
        RECT 66.145 165.805 66.315 165.975 ;
        RECT 66.605 165.805 66.775 165.975 ;
        RECT 67.065 165.805 67.235 165.975 ;
        RECT 67.525 165.805 67.695 165.975 ;
        RECT 67.985 165.805 68.155 165.975 ;
        RECT 68.445 165.805 68.615 165.975 ;
        RECT 68.905 165.805 69.075 165.975 ;
        RECT 69.365 165.805 69.535 165.975 ;
        RECT 69.825 165.805 69.995 165.975 ;
        RECT 70.285 165.805 70.455 165.975 ;
        RECT 70.745 165.805 70.915 165.975 ;
        RECT 71.205 165.805 71.375 165.975 ;
        RECT 71.665 165.805 71.835 165.975 ;
        RECT 72.125 165.805 72.295 165.975 ;
        RECT 72.585 165.805 72.755 165.975 ;
        RECT 73.045 165.805 73.215 165.975 ;
        RECT 73.505 165.805 73.675 165.975 ;
        RECT 73.965 165.805 74.135 165.975 ;
        RECT 74.425 165.805 74.595 165.975 ;
        RECT 74.885 165.805 75.055 165.975 ;
        RECT 75.345 165.805 75.515 165.975 ;
        RECT 75.805 165.805 75.975 165.975 ;
        RECT 76.265 165.805 76.435 165.975 ;
        RECT 76.725 165.805 76.895 165.975 ;
        RECT 77.185 165.805 77.355 165.975 ;
        RECT 77.645 165.805 77.815 165.975 ;
        RECT 78.105 165.805 78.275 165.975 ;
        RECT 78.565 165.805 78.735 165.975 ;
        RECT 79.025 165.805 79.195 165.975 ;
        RECT 79.485 165.805 79.655 165.975 ;
        RECT 79.945 165.805 80.115 165.975 ;
        RECT 80.405 165.805 80.575 165.975 ;
        RECT 80.865 165.805 81.035 165.975 ;
        RECT 81.325 165.805 81.495 165.975 ;
        RECT 81.785 165.805 81.955 165.975 ;
        RECT 82.245 165.805 82.415 165.975 ;
        RECT 82.705 165.805 82.875 165.975 ;
        RECT 83.165 165.805 83.335 165.975 ;
        RECT 83.625 165.805 83.795 165.975 ;
        RECT 84.085 165.805 84.255 165.975 ;
        RECT 84.545 165.805 84.715 165.975 ;
        RECT 85.005 165.805 85.175 165.975 ;
        RECT 85.465 165.805 85.635 165.975 ;
        RECT 85.925 165.805 86.095 165.975 ;
        RECT 86.385 165.805 86.555 165.975 ;
        RECT 86.845 165.805 87.015 165.975 ;
        RECT 87.305 165.805 87.475 165.975 ;
        RECT 87.765 165.805 87.935 165.975 ;
        RECT 88.225 165.805 88.395 165.975 ;
        RECT 88.685 165.805 88.855 165.975 ;
        RECT 89.145 165.805 89.315 165.975 ;
        RECT 89.605 165.805 89.775 165.975 ;
        RECT 90.065 165.805 90.235 165.975 ;
        RECT 90.525 165.805 90.695 165.975 ;
        RECT 90.985 165.805 91.155 165.975 ;
        RECT 91.445 165.805 91.615 165.975 ;
        RECT 91.905 165.805 92.075 165.975 ;
        RECT 92.365 165.805 92.535 165.975 ;
        RECT 92.825 165.805 92.995 165.975 ;
        RECT 93.285 165.805 93.455 165.975 ;
        RECT 93.745 165.805 93.915 165.975 ;
        RECT 94.205 165.805 94.375 165.975 ;
        RECT 94.665 165.805 94.835 165.975 ;
        RECT 95.125 165.805 95.295 165.975 ;
        RECT 95.585 165.805 95.755 165.975 ;
        RECT 96.045 165.805 96.215 165.975 ;
        RECT 96.505 165.805 96.675 165.975 ;
        RECT 96.965 165.805 97.135 165.975 ;
        RECT 97.425 165.805 97.595 165.975 ;
        RECT 97.885 165.805 98.055 165.975 ;
        RECT 98.345 165.805 98.515 165.975 ;
        RECT 98.805 165.805 98.975 165.975 ;
        RECT 99.265 165.805 99.435 165.975 ;
        RECT 99.725 165.805 99.895 165.975 ;
        RECT 100.185 165.805 100.355 165.975 ;
        RECT 100.645 165.805 100.815 165.975 ;
        RECT 101.105 165.805 101.275 165.975 ;
        RECT 101.565 165.805 101.735 165.975 ;
        RECT 102.025 165.805 102.195 165.975 ;
        RECT 102.485 165.805 102.655 165.975 ;
        RECT 102.945 165.805 103.115 165.975 ;
        RECT 103.405 165.805 103.575 165.975 ;
        RECT 103.865 165.805 104.035 165.975 ;
        RECT 104.325 165.805 104.495 165.975 ;
        RECT 104.785 165.805 104.955 165.975 ;
        RECT 105.245 165.805 105.415 165.975 ;
        RECT 105.705 165.805 105.875 165.975 ;
        RECT 106.165 165.805 106.335 165.975 ;
        RECT 106.625 165.805 106.795 165.975 ;
        RECT 107.085 165.805 107.255 165.975 ;
        RECT 107.545 165.805 107.715 165.975 ;
        RECT 108.005 165.805 108.175 165.975 ;
        RECT 108.465 165.805 108.635 165.975 ;
        RECT 108.925 165.805 109.095 165.975 ;
        RECT 109.385 165.805 109.555 165.975 ;
        RECT 109.845 165.805 110.015 165.975 ;
        RECT 110.305 165.805 110.475 165.975 ;
        RECT 110.765 165.805 110.935 165.975 ;
        RECT 111.225 165.805 111.395 165.975 ;
        RECT 111.685 165.805 111.855 165.975 ;
        RECT 112.145 165.805 112.315 165.975 ;
        RECT 112.605 165.805 112.775 165.975 ;
        RECT 113.065 165.805 113.235 165.975 ;
        RECT 113.525 165.805 113.695 165.975 ;
        RECT 113.985 165.805 114.155 165.975 ;
        RECT 114.445 165.805 114.615 165.975 ;
        RECT 114.905 165.805 115.075 165.975 ;
        RECT 115.365 165.805 115.535 165.975 ;
        RECT 115.825 165.805 115.995 165.975 ;
        RECT 116.285 165.805 116.455 165.975 ;
        RECT 116.745 165.805 116.915 165.975 ;
        RECT 117.205 165.805 117.375 165.975 ;
        RECT 117.665 165.805 117.835 165.975 ;
        RECT 118.125 165.805 118.295 165.975 ;
        RECT 118.585 165.805 118.755 165.975 ;
        RECT 119.045 165.805 119.215 165.975 ;
        RECT 119.505 165.805 119.675 165.975 ;
        RECT 119.965 165.805 120.135 165.975 ;
        RECT 120.425 165.805 120.595 165.975 ;
        RECT 120.885 165.805 121.055 165.975 ;
        RECT 121.345 165.805 121.515 165.975 ;
        RECT 121.805 165.805 121.975 165.975 ;
        RECT 122.265 165.805 122.435 165.975 ;
        RECT 122.725 165.805 122.895 165.975 ;
        RECT 123.185 165.805 123.355 165.975 ;
        RECT 123.645 165.805 123.815 165.975 ;
        RECT 124.105 165.805 124.275 165.975 ;
        RECT 124.565 165.805 124.735 165.975 ;
        RECT 125.025 165.805 125.195 165.975 ;
        RECT 125.485 165.805 125.655 165.975 ;
        RECT 125.945 165.805 126.115 165.975 ;
        RECT 126.405 165.805 126.575 165.975 ;
        RECT 126.865 165.805 127.035 165.975 ;
        RECT 127.325 165.805 127.495 165.975 ;
        RECT 127.785 165.805 127.955 165.975 ;
        RECT 128.245 165.805 128.415 165.975 ;
        RECT 128.705 165.805 128.875 165.975 ;
        RECT 129.165 165.805 129.335 165.975 ;
        RECT 129.625 165.805 129.795 165.975 ;
        RECT 130.085 165.805 130.255 165.975 ;
        RECT 130.545 165.805 130.715 165.975 ;
        RECT 131.005 165.805 131.175 165.975 ;
        RECT 131.465 165.805 131.635 165.975 ;
        RECT 131.925 165.805 132.095 165.975 ;
        RECT 132.385 165.805 132.555 165.975 ;
        RECT 132.845 165.805 133.015 165.975 ;
        RECT 133.305 165.805 133.475 165.975 ;
        RECT 133.765 165.805 133.935 165.975 ;
        RECT 134.225 165.805 134.395 165.975 ;
        RECT 134.685 165.805 134.855 165.975 ;
        RECT 135.145 165.805 135.315 165.975 ;
        RECT 135.605 165.805 135.775 165.975 ;
        RECT 136.065 165.805 136.235 165.975 ;
        RECT 136.525 165.805 136.695 165.975 ;
        RECT 136.985 165.805 137.155 165.975 ;
        RECT 137.445 165.805 137.615 165.975 ;
        RECT 137.905 165.805 138.075 165.975 ;
        RECT 138.365 165.805 138.535 165.975 ;
        RECT 138.825 165.805 138.995 165.975 ;
        RECT 139.285 165.805 139.455 165.975 ;
        RECT 139.745 165.805 139.915 165.975 ;
        RECT 140.205 165.805 140.375 165.975 ;
        RECT 140.665 165.805 140.835 165.975 ;
        RECT 141.125 165.805 141.295 165.975 ;
        RECT 141.585 165.805 141.755 165.975 ;
        RECT 142.045 165.805 142.215 165.975 ;
        RECT 142.505 165.805 142.675 165.975 ;
        RECT 142.965 165.805 143.135 165.975 ;
        RECT 143.425 165.805 143.595 165.975 ;
        RECT 143.885 165.805 144.055 165.975 ;
        RECT 144.345 165.805 144.515 165.975 ;
        RECT 144.805 165.805 144.975 165.975 ;
        RECT 145.265 165.805 145.435 165.975 ;
        RECT 145.725 165.805 145.895 165.975 ;
        RECT 146.185 165.805 146.355 165.975 ;
        RECT 146.645 165.805 146.815 165.975 ;
        RECT 147.105 165.805 147.275 165.975 ;
        RECT 147.565 165.805 147.735 165.975 ;
        RECT 148.025 165.805 148.195 165.975 ;
        RECT 148.485 165.805 148.655 165.975 ;
        RECT 148.945 165.805 149.115 165.975 ;
        RECT 149.405 165.805 149.575 165.975 ;
        RECT 149.865 165.805 150.035 165.975 ;
        RECT 43.145 164.615 43.315 164.785 ;
        RECT 44.065 164.955 44.235 165.125 ;
        RECT 44.525 164.275 44.695 164.445 ;
        RECT 45.905 164.275 46.075 164.445 ;
        RECT 44.985 163.595 45.155 163.765 ;
        RECT 56.025 164.275 56.195 164.445 ;
        RECT 57.405 164.615 57.575 164.785 ;
        RECT 60.165 165.295 60.335 165.465 ;
        RECT 59.245 164.275 59.415 164.445 ;
        RECT 60.625 164.275 60.795 164.445 ;
        RECT 62.005 164.615 62.175 164.785 ;
        RECT 66.375 165.295 66.545 165.465 ;
        RECT 65.225 164.615 65.395 164.785 ;
        RECT 71.665 164.615 71.835 164.785 ;
        RECT 71.205 164.275 71.375 164.445 ;
        RECT 73.045 163.595 73.215 163.765 ;
        RECT 75.345 164.275 75.515 164.445 ;
        RECT 76.725 164.275 76.895 164.445 ;
        RECT 75.805 163.935 75.975 164.105 ;
        RECT 85.005 164.275 85.175 164.445 ;
        RECT 77.645 163.595 77.815 163.765 ;
        RECT 86.845 164.275 87.015 164.445 ;
        RECT 85.925 163.935 86.095 164.105 ;
        RECT 87.305 164.275 87.475 164.445 ;
        RECT 88.685 164.615 88.855 164.785 ;
        RECT 88.225 164.275 88.395 164.445 ;
        RECT 90.065 164.275 90.235 164.445 ;
        RECT 91.905 164.615 92.075 164.785 ;
        RECT 92.365 164.275 92.535 164.445 ;
        RECT 92.825 164.275 92.995 164.445 ;
        RECT 93.285 164.275 93.455 164.445 ;
        RECT 90.985 163.595 91.155 163.765 ;
        RECT 94.205 163.595 94.375 163.765 ;
        RECT 95.125 165.295 95.295 165.465 ;
        RECT 96.505 164.275 96.675 164.445 ;
        RECT 96.965 164.275 97.135 164.445 ;
        RECT 97.425 164.275 97.595 164.445 ;
        RECT 98.345 164.275 98.515 164.445 ;
        RECT 101.105 164.275 101.275 164.445 ;
        RECT 102.485 164.275 102.655 164.445 ;
        RECT 108.005 164.275 108.175 164.445 ;
        RECT 107.085 163.595 107.255 163.765 ;
        RECT 110.765 164.615 110.935 164.785 ;
        RECT 109.385 164.275 109.555 164.445 ;
        RECT 111.225 164.275 111.395 164.445 ;
        RECT 108.465 163.595 108.635 163.765 ;
        RECT 112.605 164.615 112.775 164.785 ;
        RECT 113.065 164.615 113.235 164.785 ;
        RECT 111.685 163.595 111.855 163.765 ;
        RECT 125.945 165.295 126.115 165.465 ;
        RECT 121.805 164.275 121.975 164.445 ;
        RECT 124.105 164.615 124.275 164.785 ;
        RECT 125.025 164.275 125.195 164.445 ;
        RECT 114.905 163.595 115.075 163.765 ;
        RECT 122.725 163.595 122.895 163.765 ;
        RECT 127.785 164.955 127.955 165.125 ;
        RECT 126.865 164.275 127.035 164.445 ;
        RECT 127.785 164.275 127.955 164.445 ;
        RECT 138.825 165.295 138.995 165.465 ;
        RECT 140.665 165.295 140.835 165.465 ;
        RECT 141.125 164.615 141.295 164.785 ;
        RECT 140.205 164.275 140.375 164.445 ;
        RECT 140.665 164.275 140.835 164.445 ;
        RECT 143.425 165.295 143.595 165.465 ;
        RECT 142.045 164.275 142.215 164.445 ;
        RECT 142.965 164.275 143.135 164.445 ;
        RECT 143.885 164.225 144.055 164.395 ;
        RECT 36.245 163.085 36.415 163.255 ;
        RECT 36.705 163.085 36.875 163.255 ;
        RECT 37.165 163.085 37.335 163.255 ;
        RECT 37.625 163.085 37.795 163.255 ;
        RECT 38.085 163.085 38.255 163.255 ;
        RECT 38.545 163.085 38.715 163.255 ;
        RECT 39.005 163.085 39.175 163.255 ;
        RECT 39.465 163.085 39.635 163.255 ;
        RECT 39.925 163.085 40.095 163.255 ;
        RECT 40.385 163.085 40.555 163.255 ;
        RECT 40.845 163.085 41.015 163.255 ;
        RECT 41.305 163.085 41.475 163.255 ;
        RECT 41.765 163.085 41.935 163.255 ;
        RECT 42.225 163.085 42.395 163.255 ;
        RECT 42.685 163.085 42.855 163.255 ;
        RECT 43.145 163.085 43.315 163.255 ;
        RECT 43.605 163.085 43.775 163.255 ;
        RECT 44.065 163.085 44.235 163.255 ;
        RECT 44.525 163.085 44.695 163.255 ;
        RECT 44.985 163.085 45.155 163.255 ;
        RECT 45.445 163.085 45.615 163.255 ;
        RECT 45.905 163.085 46.075 163.255 ;
        RECT 46.365 163.085 46.535 163.255 ;
        RECT 46.825 163.085 46.995 163.255 ;
        RECT 47.285 163.085 47.455 163.255 ;
        RECT 47.745 163.085 47.915 163.255 ;
        RECT 48.205 163.085 48.375 163.255 ;
        RECT 48.665 163.085 48.835 163.255 ;
        RECT 49.125 163.085 49.295 163.255 ;
        RECT 49.585 163.085 49.755 163.255 ;
        RECT 50.045 163.085 50.215 163.255 ;
        RECT 50.505 163.085 50.675 163.255 ;
        RECT 50.965 163.085 51.135 163.255 ;
        RECT 51.425 163.085 51.595 163.255 ;
        RECT 51.885 163.085 52.055 163.255 ;
        RECT 52.345 163.085 52.515 163.255 ;
        RECT 52.805 163.085 52.975 163.255 ;
        RECT 53.265 163.085 53.435 163.255 ;
        RECT 53.725 163.085 53.895 163.255 ;
        RECT 54.185 163.085 54.355 163.255 ;
        RECT 54.645 163.085 54.815 163.255 ;
        RECT 55.105 163.085 55.275 163.255 ;
        RECT 55.565 163.085 55.735 163.255 ;
        RECT 56.025 163.085 56.195 163.255 ;
        RECT 56.485 163.085 56.655 163.255 ;
        RECT 56.945 163.085 57.115 163.255 ;
        RECT 57.405 163.085 57.575 163.255 ;
        RECT 57.865 163.085 58.035 163.255 ;
        RECT 58.325 163.085 58.495 163.255 ;
        RECT 58.785 163.085 58.955 163.255 ;
        RECT 59.245 163.085 59.415 163.255 ;
        RECT 59.705 163.085 59.875 163.255 ;
        RECT 60.165 163.085 60.335 163.255 ;
        RECT 60.625 163.085 60.795 163.255 ;
        RECT 61.085 163.085 61.255 163.255 ;
        RECT 61.545 163.085 61.715 163.255 ;
        RECT 62.005 163.085 62.175 163.255 ;
        RECT 62.465 163.085 62.635 163.255 ;
        RECT 62.925 163.085 63.095 163.255 ;
        RECT 63.385 163.085 63.555 163.255 ;
        RECT 63.845 163.085 64.015 163.255 ;
        RECT 64.305 163.085 64.475 163.255 ;
        RECT 64.765 163.085 64.935 163.255 ;
        RECT 65.225 163.085 65.395 163.255 ;
        RECT 65.685 163.085 65.855 163.255 ;
        RECT 66.145 163.085 66.315 163.255 ;
        RECT 66.605 163.085 66.775 163.255 ;
        RECT 67.065 163.085 67.235 163.255 ;
        RECT 67.525 163.085 67.695 163.255 ;
        RECT 67.985 163.085 68.155 163.255 ;
        RECT 68.445 163.085 68.615 163.255 ;
        RECT 68.905 163.085 69.075 163.255 ;
        RECT 69.365 163.085 69.535 163.255 ;
        RECT 69.825 163.085 69.995 163.255 ;
        RECT 70.285 163.085 70.455 163.255 ;
        RECT 70.745 163.085 70.915 163.255 ;
        RECT 71.205 163.085 71.375 163.255 ;
        RECT 71.665 163.085 71.835 163.255 ;
        RECT 72.125 163.085 72.295 163.255 ;
        RECT 72.585 163.085 72.755 163.255 ;
        RECT 73.045 163.085 73.215 163.255 ;
        RECT 73.505 163.085 73.675 163.255 ;
        RECT 73.965 163.085 74.135 163.255 ;
        RECT 74.425 163.085 74.595 163.255 ;
        RECT 74.885 163.085 75.055 163.255 ;
        RECT 75.345 163.085 75.515 163.255 ;
        RECT 75.805 163.085 75.975 163.255 ;
        RECT 76.265 163.085 76.435 163.255 ;
        RECT 76.725 163.085 76.895 163.255 ;
        RECT 77.185 163.085 77.355 163.255 ;
        RECT 77.645 163.085 77.815 163.255 ;
        RECT 78.105 163.085 78.275 163.255 ;
        RECT 78.565 163.085 78.735 163.255 ;
        RECT 79.025 163.085 79.195 163.255 ;
        RECT 79.485 163.085 79.655 163.255 ;
        RECT 79.945 163.085 80.115 163.255 ;
        RECT 80.405 163.085 80.575 163.255 ;
        RECT 80.865 163.085 81.035 163.255 ;
        RECT 81.325 163.085 81.495 163.255 ;
        RECT 81.785 163.085 81.955 163.255 ;
        RECT 82.245 163.085 82.415 163.255 ;
        RECT 82.705 163.085 82.875 163.255 ;
        RECT 83.165 163.085 83.335 163.255 ;
        RECT 83.625 163.085 83.795 163.255 ;
        RECT 84.085 163.085 84.255 163.255 ;
        RECT 84.545 163.085 84.715 163.255 ;
        RECT 85.005 163.085 85.175 163.255 ;
        RECT 85.465 163.085 85.635 163.255 ;
        RECT 85.925 163.085 86.095 163.255 ;
        RECT 86.385 163.085 86.555 163.255 ;
        RECT 86.845 163.085 87.015 163.255 ;
        RECT 87.305 163.085 87.475 163.255 ;
        RECT 87.765 163.085 87.935 163.255 ;
        RECT 88.225 163.085 88.395 163.255 ;
        RECT 88.685 163.085 88.855 163.255 ;
        RECT 89.145 163.085 89.315 163.255 ;
        RECT 89.605 163.085 89.775 163.255 ;
        RECT 90.065 163.085 90.235 163.255 ;
        RECT 90.525 163.085 90.695 163.255 ;
        RECT 90.985 163.085 91.155 163.255 ;
        RECT 91.445 163.085 91.615 163.255 ;
        RECT 91.905 163.085 92.075 163.255 ;
        RECT 92.365 163.085 92.535 163.255 ;
        RECT 92.825 163.085 92.995 163.255 ;
        RECT 93.285 163.085 93.455 163.255 ;
        RECT 93.745 163.085 93.915 163.255 ;
        RECT 94.205 163.085 94.375 163.255 ;
        RECT 94.665 163.085 94.835 163.255 ;
        RECT 95.125 163.085 95.295 163.255 ;
        RECT 95.585 163.085 95.755 163.255 ;
        RECT 96.045 163.085 96.215 163.255 ;
        RECT 96.505 163.085 96.675 163.255 ;
        RECT 96.965 163.085 97.135 163.255 ;
        RECT 97.425 163.085 97.595 163.255 ;
        RECT 97.885 163.085 98.055 163.255 ;
        RECT 98.345 163.085 98.515 163.255 ;
        RECT 98.805 163.085 98.975 163.255 ;
        RECT 99.265 163.085 99.435 163.255 ;
        RECT 99.725 163.085 99.895 163.255 ;
        RECT 100.185 163.085 100.355 163.255 ;
        RECT 100.645 163.085 100.815 163.255 ;
        RECT 101.105 163.085 101.275 163.255 ;
        RECT 101.565 163.085 101.735 163.255 ;
        RECT 102.025 163.085 102.195 163.255 ;
        RECT 102.485 163.085 102.655 163.255 ;
        RECT 102.945 163.085 103.115 163.255 ;
        RECT 103.405 163.085 103.575 163.255 ;
        RECT 103.865 163.085 104.035 163.255 ;
        RECT 104.325 163.085 104.495 163.255 ;
        RECT 104.785 163.085 104.955 163.255 ;
        RECT 105.245 163.085 105.415 163.255 ;
        RECT 105.705 163.085 105.875 163.255 ;
        RECT 106.165 163.085 106.335 163.255 ;
        RECT 106.625 163.085 106.795 163.255 ;
        RECT 107.085 163.085 107.255 163.255 ;
        RECT 107.545 163.085 107.715 163.255 ;
        RECT 108.005 163.085 108.175 163.255 ;
        RECT 108.465 163.085 108.635 163.255 ;
        RECT 108.925 163.085 109.095 163.255 ;
        RECT 109.385 163.085 109.555 163.255 ;
        RECT 109.845 163.085 110.015 163.255 ;
        RECT 110.305 163.085 110.475 163.255 ;
        RECT 110.765 163.085 110.935 163.255 ;
        RECT 111.225 163.085 111.395 163.255 ;
        RECT 111.685 163.085 111.855 163.255 ;
        RECT 112.145 163.085 112.315 163.255 ;
        RECT 112.605 163.085 112.775 163.255 ;
        RECT 113.065 163.085 113.235 163.255 ;
        RECT 113.525 163.085 113.695 163.255 ;
        RECT 113.985 163.085 114.155 163.255 ;
        RECT 114.445 163.085 114.615 163.255 ;
        RECT 114.905 163.085 115.075 163.255 ;
        RECT 115.365 163.085 115.535 163.255 ;
        RECT 115.825 163.085 115.995 163.255 ;
        RECT 116.285 163.085 116.455 163.255 ;
        RECT 116.745 163.085 116.915 163.255 ;
        RECT 117.205 163.085 117.375 163.255 ;
        RECT 117.665 163.085 117.835 163.255 ;
        RECT 118.125 163.085 118.295 163.255 ;
        RECT 118.585 163.085 118.755 163.255 ;
        RECT 119.045 163.085 119.215 163.255 ;
        RECT 119.505 163.085 119.675 163.255 ;
        RECT 119.965 163.085 120.135 163.255 ;
        RECT 120.425 163.085 120.595 163.255 ;
        RECT 120.885 163.085 121.055 163.255 ;
        RECT 121.345 163.085 121.515 163.255 ;
        RECT 121.805 163.085 121.975 163.255 ;
        RECT 122.265 163.085 122.435 163.255 ;
        RECT 122.725 163.085 122.895 163.255 ;
        RECT 123.185 163.085 123.355 163.255 ;
        RECT 123.645 163.085 123.815 163.255 ;
        RECT 124.105 163.085 124.275 163.255 ;
        RECT 124.565 163.085 124.735 163.255 ;
        RECT 125.025 163.085 125.195 163.255 ;
        RECT 125.485 163.085 125.655 163.255 ;
        RECT 125.945 163.085 126.115 163.255 ;
        RECT 126.405 163.085 126.575 163.255 ;
        RECT 126.865 163.085 127.035 163.255 ;
        RECT 127.325 163.085 127.495 163.255 ;
        RECT 127.785 163.085 127.955 163.255 ;
        RECT 128.245 163.085 128.415 163.255 ;
        RECT 128.705 163.085 128.875 163.255 ;
        RECT 129.165 163.085 129.335 163.255 ;
        RECT 129.625 163.085 129.795 163.255 ;
        RECT 130.085 163.085 130.255 163.255 ;
        RECT 130.545 163.085 130.715 163.255 ;
        RECT 131.005 163.085 131.175 163.255 ;
        RECT 131.465 163.085 131.635 163.255 ;
        RECT 131.925 163.085 132.095 163.255 ;
        RECT 132.385 163.085 132.555 163.255 ;
        RECT 132.845 163.085 133.015 163.255 ;
        RECT 133.305 163.085 133.475 163.255 ;
        RECT 133.765 163.085 133.935 163.255 ;
        RECT 134.225 163.085 134.395 163.255 ;
        RECT 134.685 163.085 134.855 163.255 ;
        RECT 135.145 163.085 135.315 163.255 ;
        RECT 135.605 163.085 135.775 163.255 ;
        RECT 136.065 163.085 136.235 163.255 ;
        RECT 136.525 163.085 136.695 163.255 ;
        RECT 136.985 163.085 137.155 163.255 ;
        RECT 137.445 163.085 137.615 163.255 ;
        RECT 137.905 163.085 138.075 163.255 ;
        RECT 138.365 163.085 138.535 163.255 ;
        RECT 138.825 163.085 138.995 163.255 ;
        RECT 139.285 163.085 139.455 163.255 ;
        RECT 139.745 163.085 139.915 163.255 ;
        RECT 140.205 163.085 140.375 163.255 ;
        RECT 140.665 163.085 140.835 163.255 ;
        RECT 141.125 163.085 141.295 163.255 ;
        RECT 141.585 163.085 141.755 163.255 ;
        RECT 142.045 163.085 142.215 163.255 ;
        RECT 142.505 163.085 142.675 163.255 ;
        RECT 142.965 163.085 143.135 163.255 ;
        RECT 143.425 163.085 143.595 163.255 ;
        RECT 143.885 163.085 144.055 163.255 ;
        RECT 144.345 163.085 144.515 163.255 ;
        RECT 144.805 163.085 144.975 163.255 ;
        RECT 145.265 163.085 145.435 163.255 ;
        RECT 145.725 163.085 145.895 163.255 ;
        RECT 146.185 163.085 146.355 163.255 ;
        RECT 146.645 163.085 146.815 163.255 ;
        RECT 147.105 163.085 147.275 163.255 ;
        RECT 147.565 163.085 147.735 163.255 ;
        RECT 148.025 163.085 148.195 163.255 ;
        RECT 148.485 163.085 148.655 163.255 ;
        RECT 148.945 163.085 149.115 163.255 ;
        RECT 149.405 163.085 149.575 163.255 ;
        RECT 149.865 163.085 150.035 163.255 ;
        RECT 39.925 161.895 40.095 162.065 ;
        RECT 40.410 161.215 40.580 161.385 ;
        RECT 40.805 161.555 40.975 161.725 ;
        RECT 41.260 162.235 41.430 162.405 ;
        RECT 41.995 161.555 42.165 161.725 ;
        RECT 42.510 161.215 42.680 161.385 ;
        RECT 44.080 161.215 44.250 161.385 ;
        RECT 44.515 161.555 44.685 161.725 ;
        RECT 46.825 162.575 46.995 162.745 ;
        RECT 50.505 162.575 50.675 162.745 ;
        RECT 51.425 161.895 51.595 162.065 ;
        RECT 51.885 161.555 52.055 161.725 ;
        RECT 53.265 161.555 53.435 161.725 ;
        RECT 57.405 161.895 57.575 162.065 ;
        RECT 56.485 161.555 56.655 161.725 ;
        RECT 61.085 162.575 61.255 162.745 ;
        RECT 60.165 161.895 60.335 162.065 ;
        RECT 58.325 160.875 58.495 161.045 ;
        RECT 62.465 161.895 62.635 162.065 ;
        RECT 62.925 161.555 63.095 161.725 ;
        RECT 67.985 161.895 68.155 162.065 ;
        RECT 68.445 161.555 68.615 161.725 ;
        RECT 72.125 162.575 72.295 162.745 ;
        RECT 70.285 161.895 70.455 162.065 ;
        RECT 71.205 161.895 71.375 162.065 ;
        RECT 69.825 161.215 69.995 161.385 ;
        RECT 86.385 161.895 86.555 162.065 ;
        RECT 92.825 162.575 92.995 162.745 ;
        RECT 87.305 161.215 87.475 161.385 ;
        RECT 91.905 161.895 92.075 162.065 ;
        RECT 92.825 161.895 92.995 162.065 ;
        RECT 98.805 161.895 98.975 162.065 ;
        RECT 97.425 161.555 97.595 161.725 ;
        RECT 97.885 161.555 98.055 161.725 ;
        RECT 99.725 160.875 99.895 161.045 ;
        RECT 101.105 162.575 101.275 162.745 ;
        RECT 102.025 161.895 102.195 162.065 ;
        RECT 103.865 161.895 104.035 162.065 ;
        RECT 103.405 161.555 103.575 161.725 ;
        RECT 105.245 161.895 105.415 162.065 ;
        RECT 109.385 161.895 109.555 162.065 ;
        RECT 110.305 161.895 110.475 162.065 ;
        RECT 104.325 160.875 104.495 161.045 ;
        RECT 110.765 161.555 110.935 161.725 ;
        RECT 112.145 161.895 112.315 162.065 ;
        RECT 113.985 161.895 114.155 162.065 ;
        RECT 117.665 162.575 117.835 162.745 ;
        RECT 114.905 161.895 115.075 162.065 ;
        RECT 115.365 161.895 115.535 162.065 ;
        RECT 113.065 160.875 113.235 161.045 ;
        RECT 116.745 161.895 116.915 162.065 ;
        RECT 125.945 162.575 126.115 162.745 ;
        RECT 123.645 162.235 123.815 162.405 ;
        RECT 125.025 161.895 125.195 162.065 ;
        RECT 124.565 161.555 124.735 161.725 ;
        RECT 125.025 160.875 125.195 161.045 ;
        RECT 128.705 161.895 128.875 162.065 ;
        RECT 131.465 161.895 131.635 162.065 ;
        RECT 127.785 160.875 127.955 161.045 ;
        RECT 132.385 161.555 132.555 161.725 ;
        RECT 131.925 160.875 132.095 161.045 ;
        RECT 138.825 162.575 138.995 162.745 ;
        RECT 136.525 162.235 136.695 162.405 ;
        RECT 137.905 161.895 138.075 162.065 ;
        RECT 134.685 161.215 134.855 161.385 ;
        RECT 137.445 161.555 137.615 161.725 ;
        RECT 139.745 161.895 139.915 162.065 ;
        RECT 136.985 160.875 137.155 161.045 ;
        RECT 140.230 161.215 140.400 161.385 ;
        RECT 140.625 161.555 140.795 161.725 ;
        RECT 141.025 161.895 141.195 162.065 ;
        RECT 141.815 161.555 141.985 161.725 ;
        RECT 142.330 161.215 142.500 161.385 ;
        RECT 143.900 161.215 144.070 161.385 ;
        RECT 144.335 161.555 144.505 161.725 ;
        RECT 146.645 162.575 146.815 162.745 ;
        RECT 36.245 160.365 36.415 160.535 ;
        RECT 36.705 160.365 36.875 160.535 ;
        RECT 37.165 160.365 37.335 160.535 ;
        RECT 37.625 160.365 37.795 160.535 ;
        RECT 38.085 160.365 38.255 160.535 ;
        RECT 38.545 160.365 38.715 160.535 ;
        RECT 39.005 160.365 39.175 160.535 ;
        RECT 39.465 160.365 39.635 160.535 ;
        RECT 39.925 160.365 40.095 160.535 ;
        RECT 40.385 160.365 40.555 160.535 ;
        RECT 40.845 160.365 41.015 160.535 ;
        RECT 41.305 160.365 41.475 160.535 ;
        RECT 41.765 160.365 41.935 160.535 ;
        RECT 42.225 160.365 42.395 160.535 ;
        RECT 42.685 160.365 42.855 160.535 ;
        RECT 43.145 160.365 43.315 160.535 ;
        RECT 43.605 160.365 43.775 160.535 ;
        RECT 44.065 160.365 44.235 160.535 ;
        RECT 44.525 160.365 44.695 160.535 ;
        RECT 44.985 160.365 45.155 160.535 ;
        RECT 45.445 160.365 45.615 160.535 ;
        RECT 45.905 160.365 46.075 160.535 ;
        RECT 46.365 160.365 46.535 160.535 ;
        RECT 46.825 160.365 46.995 160.535 ;
        RECT 47.285 160.365 47.455 160.535 ;
        RECT 47.745 160.365 47.915 160.535 ;
        RECT 48.205 160.365 48.375 160.535 ;
        RECT 48.665 160.365 48.835 160.535 ;
        RECT 49.125 160.365 49.295 160.535 ;
        RECT 49.585 160.365 49.755 160.535 ;
        RECT 50.045 160.365 50.215 160.535 ;
        RECT 50.505 160.365 50.675 160.535 ;
        RECT 50.965 160.365 51.135 160.535 ;
        RECT 51.425 160.365 51.595 160.535 ;
        RECT 51.885 160.365 52.055 160.535 ;
        RECT 52.345 160.365 52.515 160.535 ;
        RECT 52.805 160.365 52.975 160.535 ;
        RECT 53.265 160.365 53.435 160.535 ;
        RECT 53.725 160.365 53.895 160.535 ;
        RECT 54.185 160.365 54.355 160.535 ;
        RECT 54.645 160.365 54.815 160.535 ;
        RECT 55.105 160.365 55.275 160.535 ;
        RECT 55.565 160.365 55.735 160.535 ;
        RECT 56.025 160.365 56.195 160.535 ;
        RECT 56.485 160.365 56.655 160.535 ;
        RECT 56.945 160.365 57.115 160.535 ;
        RECT 57.405 160.365 57.575 160.535 ;
        RECT 57.865 160.365 58.035 160.535 ;
        RECT 58.325 160.365 58.495 160.535 ;
        RECT 58.785 160.365 58.955 160.535 ;
        RECT 59.245 160.365 59.415 160.535 ;
        RECT 59.705 160.365 59.875 160.535 ;
        RECT 60.165 160.365 60.335 160.535 ;
        RECT 60.625 160.365 60.795 160.535 ;
        RECT 61.085 160.365 61.255 160.535 ;
        RECT 61.545 160.365 61.715 160.535 ;
        RECT 62.005 160.365 62.175 160.535 ;
        RECT 62.465 160.365 62.635 160.535 ;
        RECT 62.925 160.365 63.095 160.535 ;
        RECT 63.385 160.365 63.555 160.535 ;
        RECT 63.845 160.365 64.015 160.535 ;
        RECT 64.305 160.365 64.475 160.535 ;
        RECT 64.765 160.365 64.935 160.535 ;
        RECT 65.225 160.365 65.395 160.535 ;
        RECT 65.685 160.365 65.855 160.535 ;
        RECT 66.145 160.365 66.315 160.535 ;
        RECT 66.605 160.365 66.775 160.535 ;
        RECT 67.065 160.365 67.235 160.535 ;
        RECT 67.525 160.365 67.695 160.535 ;
        RECT 67.985 160.365 68.155 160.535 ;
        RECT 68.445 160.365 68.615 160.535 ;
        RECT 68.905 160.365 69.075 160.535 ;
        RECT 69.365 160.365 69.535 160.535 ;
        RECT 69.825 160.365 69.995 160.535 ;
        RECT 70.285 160.365 70.455 160.535 ;
        RECT 70.745 160.365 70.915 160.535 ;
        RECT 71.205 160.365 71.375 160.535 ;
        RECT 71.665 160.365 71.835 160.535 ;
        RECT 72.125 160.365 72.295 160.535 ;
        RECT 72.585 160.365 72.755 160.535 ;
        RECT 73.045 160.365 73.215 160.535 ;
        RECT 73.505 160.365 73.675 160.535 ;
        RECT 73.965 160.365 74.135 160.535 ;
        RECT 74.425 160.365 74.595 160.535 ;
        RECT 74.885 160.365 75.055 160.535 ;
        RECT 75.345 160.365 75.515 160.535 ;
        RECT 75.805 160.365 75.975 160.535 ;
        RECT 76.265 160.365 76.435 160.535 ;
        RECT 76.725 160.365 76.895 160.535 ;
        RECT 77.185 160.365 77.355 160.535 ;
        RECT 77.645 160.365 77.815 160.535 ;
        RECT 78.105 160.365 78.275 160.535 ;
        RECT 78.565 160.365 78.735 160.535 ;
        RECT 79.025 160.365 79.195 160.535 ;
        RECT 79.485 160.365 79.655 160.535 ;
        RECT 79.945 160.365 80.115 160.535 ;
        RECT 80.405 160.365 80.575 160.535 ;
        RECT 80.865 160.365 81.035 160.535 ;
        RECT 81.325 160.365 81.495 160.535 ;
        RECT 81.785 160.365 81.955 160.535 ;
        RECT 82.245 160.365 82.415 160.535 ;
        RECT 82.705 160.365 82.875 160.535 ;
        RECT 83.165 160.365 83.335 160.535 ;
        RECT 83.625 160.365 83.795 160.535 ;
        RECT 84.085 160.365 84.255 160.535 ;
        RECT 84.545 160.365 84.715 160.535 ;
        RECT 85.005 160.365 85.175 160.535 ;
        RECT 85.465 160.365 85.635 160.535 ;
        RECT 85.925 160.365 86.095 160.535 ;
        RECT 86.385 160.365 86.555 160.535 ;
        RECT 86.845 160.365 87.015 160.535 ;
        RECT 87.305 160.365 87.475 160.535 ;
        RECT 87.765 160.365 87.935 160.535 ;
        RECT 88.225 160.365 88.395 160.535 ;
        RECT 88.685 160.365 88.855 160.535 ;
        RECT 89.145 160.365 89.315 160.535 ;
        RECT 89.605 160.365 89.775 160.535 ;
        RECT 90.065 160.365 90.235 160.535 ;
        RECT 90.525 160.365 90.695 160.535 ;
        RECT 90.985 160.365 91.155 160.535 ;
        RECT 91.445 160.365 91.615 160.535 ;
        RECT 91.905 160.365 92.075 160.535 ;
        RECT 92.365 160.365 92.535 160.535 ;
        RECT 92.825 160.365 92.995 160.535 ;
        RECT 93.285 160.365 93.455 160.535 ;
        RECT 93.745 160.365 93.915 160.535 ;
        RECT 94.205 160.365 94.375 160.535 ;
        RECT 94.665 160.365 94.835 160.535 ;
        RECT 95.125 160.365 95.295 160.535 ;
        RECT 95.585 160.365 95.755 160.535 ;
        RECT 96.045 160.365 96.215 160.535 ;
        RECT 96.505 160.365 96.675 160.535 ;
        RECT 96.965 160.365 97.135 160.535 ;
        RECT 97.425 160.365 97.595 160.535 ;
        RECT 97.885 160.365 98.055 160.535 ;
        RECT 98.345 160.365 98.515 160.535 ;
        RECT 98.805 160.365 98.975 160.535 ;
        RECT 99.265 160.365 99.435 160.535 ;
        RECT 99.725 160.365 99.895 160.535 ;
        RECT 100.185 160.365 100.355 160.535 ;
        RECT 100.645 160.365 100.815 160.535 ;
        RECT 101.105 160.365 101.275 160.535 ;
        RECT 101.565 160.365 101.735 160.535 ;
        RECT 102.025 160.365 102.195 160.535 ;
        RECT 102.485 160.365 102.655 160.535 ;
        RECT 102.945 160.365 103.115 160.535 ;
        RECT 103.405 160.365 103.575 160.535 ;
        RECT 103.865 160.365 104.035 160.535 ;
        RECT 104.325 160.365 104.495 160.535 ;
        RECT 104.785 160.365 104.955 160.535 ;
        RECT 105.245 160.365 105.415 160.535 ;
        RECT 105.705 160.365 105.875 160.535 ;
        RECT 106.165 160.365 106.335 160.535 ;
        RECT 106.625 160.365 106.795 160.535 ;
        RECT 107.085 160.365 107.255 160.535 ;
        RECT 107.545 160.365 107.715 160.535 ;
        RECT 108.005 160.365 108.175 160.535 ;
        RECT 108.465 160.365 108.635 160.535 ;
        RECT 108.925 160.365 109.095 160.535 ;
        RECT 109.385 160.365 109.555 160.535 ;
        RECT 109.845 160.365 110.015 160.535 ;
        RECT 110.305 160.365 110.475 160.535 ;
        RECT 110.765 160.365 110.935 160.535 ;
        RECT 111.225 160.365 111.395 160.535 ;
        RECT 111.685 160.365 111.855 160.535 ;
        RECT 112.145 160.365 112.315 160.535 ;
        RECT 112.605 160.365 112.775 160.535 ;
        RECT 113.065 160.365 113.235 160.535 ;
        RECT 113.525 160.365 113.695 160.535 ;
        RECT 113.985 160.365 114.155 160.535 ;
        RECT 114.445 160.365 114.615 160.535 ;
        RECT 114.905 160.365 115.075 160.535 ;
        RECT 115.365 160.365 115.535 160.535 ;
        RECT 115.825 160.365 115.995 160.535 ;
        RECT 116.285 160.365 116.455 160.535 ;
        RECT 116.745 160.365 116.915 160.535 ;
        RECT 117.205 160.365 117.375 160.535 ;
        RECT 117.665 160.365 117.835 160.535 ;
        RECT 118.125 160.365 118.295 160.535 ;
        RECT 118.585 160.365 118.755 160.535 ;
        RECT 119.045 160.365 119.215 160.535 ;
        RECT 119.505 160.365 119.675 160.535 ;
        RECT 119.965 160.365 120.135 160.535 ;
        RECT 120.425 160.365 120.595 160.535 ;
        RECT 120.885 160.365 121.055 160.535 ;
        RECT 121.345 160.365 121.515 160.535 ;
        RECT 121.805 160.365 121.975 160.535 ;
        RECT 122.265 160.365 122.435 160.535 ;
        RECT 122.725 160.365 122.895 160.535 ;
        RECT 123.185 160.365 123.355 160.535 ;
        RECT 123.645 160.365 123.815 160.535 ;
        RECT 124.105 160.365 124.275 160.535 ;
        RECT 124.565 160.365 124.735 160.535 ;
        RECT 125.025 160.365 125.195 160.535 ;
        RECT 125.485 160.365 125.655 160.535 ;
        RECT 125.945 160.365 126.115 160.535 ;
        RECT 126.405 160.365 126.575 160.535 ;
        RECT 126.865 160.365 127.035 160.535 ;
        RECT 127.325 160.365 127.495 160.535 ;
        RECT 127.785 160.365 127.955 160.535 ;
        RECT 128.245 160.365 128.415 160.535 ;
        RECT 128.705 160.365 128.875 160.535 ;
        RECT 129.165 160.365 129.335 160.535 ;
        RECT 129.625 160.365 129.795 160.535 ;
        RECT 130.085 160.365 130.255 160.535 ;
        RECT 130.545 160.365 130.715 160.535 ;
        RECT 131.005 160.365 131.175 160.535 ;
        RECT 131.465 160.365 131.635 160.535 ;
        RECT 131.925 160.365 132.095 160.535 ;
        RECT 132.385 160.365 132.555 160.535 ;
        RECT 132.845 160.365 133.015 160.535 ;
        RECT 133.305 160.365 133.475 160.535 ;
        RECT 133.765 160.365 133.935 160.535 ;
        RECT 134.225 160.365 134.395 160.535 ;
        RECT 134.685 160.365 134.855 160.535 ;
        RECT 135.145 160.365 135.315 160.535 ;
        RECT 135.605 160.365 135.775 160.535 ;
        RECT 136.065 160.365 136.235 160.535 ;
        RECT 136.525 160.365 136.695 160.535 ;
        RECT 136.985 160.365 137.155 160.535 ;
        RECT 137.445 160.365 137.615 160.535 ;
        RECT 137.905 160.365 138.075 160.535 ;
        RECT 138.365 160.365 138.535 160.535 ;
        RECT 138.825 160.365 138.995 160.535 ;
        RECT 139.285 160.365 139.455 160.535 ;
        RECT 139.745 160.365 139.915 160.535 ;
        RECT 140.205 160.365 140.375 160.535 ;
        RECT 140.665 160.365 140.835 160.535 ;
        RECT 141.125 160.365 141.295 160.535 ;
        RECT 141.585 160.365 141.755 160.535 ;
        RECT 142.045 160.365 142.215 160.535 ;
        RECT 142.505 160.365 142.675 160.535 ;
        RECT 142.965 160.365 143.135 160.535 ;
        RECT 143.425 160.365 143.595 160.535 ;
        RECT 143.885 160.365 144.055 160.535 ;
        RECT 144.345 160.365 144.515 160.535 ;
        RECT 144.805 160.365 144.975 160.535 ;
        RECT 145.265 160.365 145.435 160.535 ;
        RECT 145.725 160.365 145.895 160.535 ;
        RECT 146.185 160.365 146.355 160.535 ;
        RECT 146.645 160.365 146.815 160.535 ;
        RECT 147.105 160.365 147.275 160.535 ;
        RECT 147.565 160.365 147.735 160.535 ;
        RECT 148.025 160.365 148.195 160.535 ;
        RECT 148.485 160.365 148.655 160.535 ;
        RECT 148.945 160.365 149.115 160.535 ;
        RECT 149.405 160.365 149.575 160.535 ;
        RECT 149.865 160.365 150.035 160.535 ;
        RECT 46.825 159.855 46.995 160.025 ;
        RECT 42.225 158.835 42.395 159.005 ;
        RECT 43.605 158.835 43.775 159.005 ;
        RECT 44.985 158.835 45.155 159.005 ;
        RECT 45.905 158.835 46.075 159.005 ;
        RECT 42.715 158.155 42.885 158.325 ;
        RECT 43.145 158.155 43.315 158.325 ;
        RECT 55.105 159.175 55.275 159.345 ;
        RECT 54.645 158.835 54.815 159.005 ;
        RECT 56.485 159.175 56.655 159.345 ;
        RECT 58.325 158.835 58.495 159.005 ;
        RECT 58.785 158.835 58.955 159.005 ;
        RECT 59.705 158.835 59.875 159.005 ;
        RECT 60.625 158.495 60.795 158.665 ;
        RECT 71.665 159.175 71.835 159.345 ;
        RECT 72.585 158.835 72.755 159.005 ;
        RECT 75.345 158.835 75.515 159.005 ;
        RECT 75.805 158.835 75.975 159.005 ;
        RECT 76.265 158.835 76.435 159.005 ;
        RECT 73.505 158.155 73.675 158.325 ;
        RECT 79.025 158.835 79.195 159.005 ;
        RECT 79.485 158.835 79.655 159.005 ;
        RECT 82.245 158.835 82.415 159.005 ;
        RECT 84.085 158.495 84.255 158.665 ;
        RECT 96.965 158.835 97.135 159.005 ;
        RECT 97.885 158.835 98.055 159.005 ;
        RECT 98.345 158.835 98.515 159.005 ;
        RECT 98.805 158.835 98.975 159.005 ;
        RECT 101.105 158.835 101.275 159.005 ;
        RECT 102.485 159.175 102.655 159.345 ;
        RECT 102.025 158.835 102.195 159.005 ;
        RECT 103.865 158.835 104.035 159.005 ;
        RECT 105.245 159.175 105.415 159.345 ;
        RECT 105.705 159.175 105.875 159.345 ;
        RECT 106.625 158.835 106.795 159.005 ;
        RECT 104.785 158.495 104.955 158.665 ;
        RECT 107.545 158.155 107.715 158.325 ;
        RECT 109.385 158.835 109.555 159.005 ;
        RECT 110.305 158.835 110.475 159.005 ;
        RECT 111.685 159.175 111.855 159.345 ;
        RECT 111.225 158.835 111.395 159.005 ;
        RECT 112.145 158.835 112.315 159.005 ;
        RECT 113.525 159.175 113.695 159.345 ;
        RECT 113.065 158.785 113.235 158.955 ;
        RECT 113.985 158.835 114.155 159.005 ;
        RECT 114.905 158.835 115.075 159.005 ;
        RECT 125.025 159.855 125.195 160.025 ;
        RECT 115.825 158.155 115.995 158.325 ;
        RECT 126.865 159.175 127.035 159.345 ;
        RECT 125.945 158.835 126.115 159.005 ;
        RECT 128.245 158.835 128.415 159.005 ;
        RECT 132.845 158.835 133.015 159.005 ;
        RECT 133.765 158.835 133.935 159.005 ;
        RECT 134.225 158.835 134.395 159.005 ;
        RECT 134.685 158.835 134.855 159.005 ;
        RECT 136.525 158.835 136.695 159.005 ;
        RECT 136.065 158.495 136.235 158.665 ;
        RECT 137.445 158.835 137.615 159.005 ;
        RECT 137.905 158.835 138.075 159.005 ;
        RECT 138.365 158.835 138.535 159.005 ;
        RECT 139.745 158.155 139.915 158.325 ;
        RECT 141.585 159.515 141.755 159.685 ;
        RECT 143.425 159.855 143.595 160.025 ;
        RECT 141.125 158.835 141.295 159.005 ;
        RECT 140.205 158.155 140.375 158.325 ;
        RECT 142.505 158.835 142.675 159.005 ;
        RECT 143.885 158.835 144.055 159.005 ;
        RECT 146.185 159.515 146.355 159.685 ;
        RECT 145.725 158.835 145.895 159.005 ;
        RECT 144.805 158.155 144.975 158.325 ;
        RECT 147.105 158.835 147.275 159.005 ;
        RECT 36.245 157.645 36.415 157.815 ;
        RECT 36.705 157.645 36.875 157.815 ;
        RECT 37.165 157.645 37.335 157.815 ;
        RECT 37.625 157.645 37.795 157.815 ;
        RECT 38.085 157.645 38.255 157.815 ;
        RECT 38.545 157.645 38.715 157.815 ;
        RECT 39.005 157.645 39.175 157.815 ;
        RECT 39.465 157.645 39.635 157.815 ;
        RECT 39.925 157.645 40.095 157.815 ;
        RECT 40.385 157.645 40.555 157.815 ;
        RECT 40.845 157.645 41.015 157.815 ;
        RECT 41.305 157.645 41.475 157.815 ;
        RECT 41.765 157.645 41.935 157.815 ;
        RECT 42.225 157.645 42.395 157.815 ;
        RECT 42.685 157.645 42.855 157.815 ;
        RECT 43.145 157.645 43.315 157.815 ;
        RECT 43.605 157.645 43.775 157.815 ;
        RECT 44.065 157.645 44.235 157.815 ;
        RECT 44.525 157.645 44.695 157.815 ;
        RECT 44.985 157.645 45.155 157.815 ;
        RECT 45.445 157.645 45.615 157.815 ;
        RECT 45.905 157.645 46.075 157.815 ;
        RECT 46.365 157.645 46.535 157.815 ;
        RECT 46.825 157.645 46.995 157.815 ;
        RECT 47.285 157.645 47.455 157.815 ;
        RECT 47.745 157.645 47.915 157.815 ;
        RECT 48.205 157.645 48.375 157.815 ;
        RECT 48.665 157.645 48.835 157.815 ;
        RECT 49.125 157.645 49.295 157.815 ;
        RECT 49.585 157.645 49.755 157.815 ;
        RECT 50.045 157.645 50.215 157.815 ;
        RECT 50.505 157.645 50.675 157.815 ;
        RECT 50.965 157.645 51.135 157.815 ;
        RECT 51.425 157.645 51.595 157.815 ;
        RECT 51.885 157.645 52.055 157.815 ;
        RECT 52.345 157.645 52.515 157.815 ;
        RECT 52.805 157.645 52.975 157.815 ;
        RECT 53.265 157.645 53.435 157.815 ;
        RECT 53.725 157.645 53.895 157.815 ;
        RECT 54.185 157.645 54.355 157.815 ;
        RECT 54.645 157.645 54.815 157.815 ;
        RECT 55.105 157.645 55.275 157.815 ;
        RECT 55.565 157.645 55.735 157.815 ;
        RECT 56.025 157.645 56.195 157.815 ;
        RECT 56.485 157.645 56.655 157.815 ;
        RECT 56.945 157.645 57.115 157.815 ;
        RECT 57.405 157.645 57.575 157.815 ;
        RECT 57.865 157.645 58.035 157.815 ;
        RECT 58.325 157.645 58.495 157.815 ;
        RECT 58.785 157.645 58.955 157.815 ;
        RECT 59.245 157.645 59.415 157.815 ;
        RECT 59.705 157.645 59.875 157.815 ;
        RECT 60.165 157.645 60.335 157.815 ;
        RECT 60.625 157.645 60.795 157.815 ;
        RECT 61.085 157.645 61.255 157.815 ;
        RECT 61.545 157.645 61.715 157.815 ;
        RECT 62.005 157.645 62.175 157.815 ;
        RECT 62.465 157.645 62.635 157.815 ;
        RECT 62.925 157.645 63.095 157.815 ;
        RECT 63.385 157.645 63.555 157.815 ;
        RECT 63.845 157.645 64.015 157.815 ;
        RECT 64.305 157.645 64.475 157.815 ;
        RECT 64.765 157.645 64.935 157.815 ;
        RECT 65.225 157.645 65.395 157.815 ;
        RECT 65.685 157.645 65.855 157.815 ;
        RECT 66.145 157.645 66.315 157.815 ;
        RECT 66.605 157.645 66.775 157.815 ;
        RECT 67.065 157.645 67.235 157.815 ;
        RECT 67.525 157.645 67.695 157.815 ;
        RECT 67.985 157.645 68.155 157.815 ;
        RECT 68.445 157.645 68.615 157.815 ;
        RECT 68.905 157.645 69.075 157.815 ;
        RECT 69.365 157.645 69.535 157.815 ;
        RECT 69.825 157.645 69.995 157.815 ;
        RECT 70.285 157.645 70.455 157.815 ;
        RECT 70.745 157.645 70.915 157.815 ;
        RECT 71.205 157.645 71.375 157.815 ;
        RECT 71.665 157.645 71.835 157.815 ;
        RECT 72.125 157.645 72.295 157.815 ;
        RECT 72.585 157.645 72.755 157.815 ;
        RECT 73.045 157.645 73.215 157.815 ;
        RECT 73.505 157.645 73.675 157.815 ;
        RECT 73.965 157.645 74.135 157.815 ;
        RECT 74.425 157.645 74.595 157.815 ;
        RECT 74.885 157.645 75.055 157.815 ;
        RECT 75.345 157.645 75.515 157.815 ;
        RECT 75.805 157.645 75.975 157.815 ;
        RECT 76.265 157.645 76.435 157.815 ;
        RECT 76.725 157.645 76.895 157.815 ;
        RECT 77.185 157.645 77.355 157.815 ;
        RECT 77.645 157.645 77.815 157.815 ;
        RECT 78.105 157.645 78.275 157.815 ;
        RECT 78.565 157.645 78.735 157.815 ;
        RECT 79.025 157.645 79.195 157.815 ;
        RECT 79.485 157.645 79.655 157.815 ;
        RECT 79.945 157.645 80.115 157.815 ;
        RECT 80.405 157.645 80.575 157.815 ;
        RECT 80.865 157.645 81.035 157.815 ;
        RECT 81.325 157.645 81.495 157.815 ;
        RECT 81.785 157.645 81.955 157.815 ;
        RECT 82.245 157.645 82.415 157.815 ;
        RECT 82.705 157.645 82.875 157.815 ;
        RECT 83.165 157.645 83.335 157.815 ;
        RECT 83.625 157.645 83.795 157.815 ;
        RECT 84.085 157.645 84.255 157.815 ;
        RECT 84.545 157.645 84.715 157.815 ;
        RECT 85.005 157.645 85.175 157.815 ;
        RECT 85.465 157.645 85.635 157.815 ;
        RECT 85.925 157.645 86.095 157.815 ;
        RECT 86.385 157.645 86.555 157.815 ;
        RECT 86.845 157.645 87.015 157.815 ;
        RECT 87.305 157.645 87.475 157.815 ;
        RECT 87.765 157.645 87.935 157.815 ;
        RECT 88.225 157.645 88.395 157.815 ;
        RECT 88.685 157.645 88.855 157.815 ;
        RECT 89.145 157.645 89.315 157.815 ;
        RECT 89.605 157.645 89.775 157.815 ;
        RECT 90.065 157.645 90.235 157.815 ;
        RECT 90.525 157.645 90.695 157.815 ;
        RECT 90.985 157.645 91.155 157.815 ;
        RECT 91.445 157.645 91.615 157.815 ;
        RECT 91.905 157.645 92.075 157.815 ;
        RECT 92.365 157.645 92.535 157.815 ;
        RECT 92.825 157.645 92.995 157.815 ;
        RECT 93.285 157.645 93.455 157.815 ;
        RECT 93.745 157.645 93.915 157.815 ;
        RECT 94.205 157.645 94.375 157.815 ;
        RECT 94.665 157.645 94.835 157.815 ;
        RECT 95.125 157.645 95.295 157.815 ;
        RECT 95.585 157.645 95.755 157.815 ;
        RECT 96.045 157.645 96.215 157.815 ;
        RECT 96.505 157.645 96.675 157.815 ;
        RECT 96.965 157.645 97.135 157.815 ;
        RECT 97.425 157.645 97.595 157.815 ;
        RECT 97.885 157.645 98.055 157.815 ;
        RECT 98.345 157.645 98.515 157.815 ;
        RECT 98.805 157.645 98.975 157.815 ;
        RECT 99.265 157.645 99.435 157.815 ;
        RECT 99.725 157.645 99.895 157.815 ;
        RECT 100.185 157.645 100.355 157.815 ;
        RECT 100.645 157.645 100.815 157.815 ;
        RECT 101.105 157.645 101.275 157.815 ;
        RECT 101.565 157.645 101.735 157.815 ;
        RECT 102.025 157.645 102.195 157.815 ;
        RECT 102.485 157.645 102.655 157.815 ;
        RECT 102.945 157.645 103.115 157.815 ;
        RECT 103.405 157.645 103.575 157.815 ;
        RECT 103.865 157.645 104.035 157.815 ;
        RECT 104.325 157.645 104.495 157.815 ;
        RECT 104.785 157.645 104.955 157.815 ;
        RECT 105.245 157.645 105.415 157.815 ;
        RECT 105.705 157.645 105.875 157.815 ;
        RECT 106.165 157.645 106.335 157.815 ;
        RECT 106.625 157.645 106.795 157.815 ;
        RECT 107.085 157.645 107.255 157.815 ;
        RECT 107.545 157.645 107.715 157.815 ;
        RECT 108.005 157.645 108.175 157.815 ;
        RECT 108.465 157.645 108.635 157.815 ;
        RECT 108.925 157.645 109.095 157.815 ;
        RECT 109.385 157.645 109.555 157.815 ;
        RECT 109.845 157.645 110.015 157.815 ;
        RECT 110.305 157.645 110.475 157.815 ;
        RECT 110.765 157.645 110.935 157.815 ;
        RECT 111.225 157.645 111.395 157.815 ;
        RECT 111.685 157.645 111.855 157.815 ;
        RECT 112.145 157.645 112.315 157.815 ;
        RECT 112.605 157.645 112.775 157.815 ;
        RECT 113.065 157.645 113.235 157.815 ;
        RECT 113.525 157.645 113.695 157.815 ;
        RECT 113.985 157.645 114.155 157.815 ;
        RECT 114.445 157.645 114.615 157.815 ;
        RECT 114.905 157.645 115.075 157.815 ;
        RECT 115.365 157.645 115.535 157.815 ;
        RECT 115.825 157.645 115.995 157.815 ;
        RECT 116.285 157.645 116.455 157.815 ;
        RECT 116.745 157.645 116.915 157.815 ;
        RECT 117.205 157.645 117.375 157.815 ;
        RECT 117.665 157.645 117.835 157.815 ;
        RECT 118.125 157.645 118.295 157.815 ;
        RECT 118.585 157.645 118.755 157.815 ;
        RECT 119.045 157.645 119.215 157.815 ;
        RECT 119.505 157.645 119.675 157.815 ;
        RECT 119.965 157.645 120.135 157.815 ;
        RECT 120.425 157.645 120.595 157.815 ;
        RECT 120.885 157.645 121.055 157.815 ;
        RECT 121.345 157.645 121.515 157.815 ;
        RECT 121.805 157.645 121.975 157.815 ;
        RECT 122.265 157.645 122.435 157.815 ;
        RECT 122.725 157.645 122.895 157.815 ;
        RECT 123.185 157.645 123.355 157.815 ;
        RECT 123.645 157.645 123.815 157.815 ;
        RECT 124.105 157.645 124.275 157.815 ;
        RECT 124.565 157.645 124.735 157.815 ;
        RECT 125.025 157.645 125.195 157.815 ;
        RECT 125.485 157.645 125.655 157.815 ;
        RECT 125.945 157.645 126.115 157.815 ;
        RECT 126.405 157.645 126.575 157.815 ;
        RECT 126.865 157.645 127.035 157.815 ;
        RECT 127.325 157.645 127.495 157.815 ;
        RECT 127.785 157.645 127.955 157.815 ;
        RECT 128.245 157.645 128.415 157.815 ;
        RECT 128.705 157.645 128.875 157.815 ;
        RECT 129.165 157.645 129.335 157.815 ;
        RECT 129.625 157.645 129.795 157.815 ;
        RECT 130.085 157.645 130.255 157.815 ;
        RECT 130.545 157.645 130.715 157.815 ;
        RECT 131.005 157.645 131.175 157.815 ;
        RECT 131.465 157.645 131.635 157.815 ;
        RECT 131.925 157.645 132.095 157.815 ;
        RECT 132.385 157.645 132.555 157.815 ;
        RECT 132.845 157.645 133.015 157.815 ;
        RECT 133.305 157.645 133.475 157.815 ;
        RECT 133.765 157.645 133.935 157.815 ;
        RECT 134.225 157.645 134.395 157.815 ;
        RECT 134.685 157.645 134.855 157.815 ;
        RECT 135.145 157.645 135.315 157.815 ;
        RECT 135.605 157.645 135.775 157.815 ;
        RECT 136.065 157.645 136.235 157.815 ;
        RECT 136.525 157.645 136.695 157.815 ;
        RECT 136.985 157.645 137.155 157.815 ;
        RECT 137.445 157.645 137.615 157.815 ;
        RECT 137.905 157.645 138.075 157.815 ;
        RECT 138.365 157.645 138.535 157.815 ;
        RECT 138.825 157.645 138.995 157.815 ;
        RECT 139.285 157.645 139.455 157.815 ;
        RECT 139.745 157.645 139.915 157.815 ;
        RECT 140.205 157.645 140.375 157.815 ;
        RECT 140.665 157.645 140.835 157.815 ;
        RECT 141.125 157.645 141.295 157.815 ;
        RECT 141.585 157.645 141.755 157.815 ;
        RECT 142.045 157.645 142.215 157.815 ;
        RECT 142.505 157.645 142.675 157.815 ;
        RECT 142.965 157.645 143.135 157.815 ;
        RECT 143.425 157.645 143.595 157.815 ;
        RECT 143.885 157.645 144.055 157.815 ;
        RECT 144.345 157.645 144.515 157.815 ;
        RECT 144.805 157.645 144.975 157.815 ;
        RECT 145.265 157.645 145.435 157.815 ;
        RECT 145.725 157.645 145.895 157.815 ;
        RECT 146.185 157.645 146.355 157.815 ;
        RECT 146.645 157.645 146.815 157.815 ;
        RECT 147.105 157.645 147.275 157.815 ;
        RECT 147.565 157.645 147.735 157.815 ;
        RECT 148.025 157.645 148.195 157.815 ;
        RECT 148.485 157.645 148.655 157.815 ;
        RECT 148.945 157.645 149.115 157.815 ;
        RECT 149.405 157.645 149.575 157.815 ;
        RECT 149.865 157.645 150.035 157.815 ;
        RECT 38.085 156.455 38.255 156.625 ;
        RECT 38.570 155.775 38.740 155.945 ;
        RECT 38.965 156.115 39.135 156.285 ;
        RECT 39.420 156.455 39.590 156.625 ;
        RECT 40.155 156.115 40.325 156.285 ;
        RECT 40.670 155.775 40.840 155.945 ;
        RECT 42.240 155.775 42.410 155.945 ;
        RECT 42.675 156.115 42.845 156.285 ;
        RECT 44.985 157.135 45.155 157.305 ;
        RECT 47.285 156.795 47.455 156.965 ;
        RECT 48.205 156.795 48.375 156.965 ;
        RECT 51.425 157.135 51.595 157.305 ;
        RECT 53.735 156.115 53.905 156.285 ;
        RECT 54.170 155.775 54.340 155.945 ;
        RECT 56.255 156.115 56.425 156.285 ;
        RECT 55.740 155.775 55.910 155.945 ;
        RECT 57.100 156.795 57.270 156.965 ;
        RECT 57.445 156.115 57.615 156.285 ;
        RECT 58.325 156.455 58.495 156.625 ;
        RECT 57.840 155.775 58.010 155.945 ;
        RECT 58.785 155.775 58.955 155.945 ;
        RECT 60.625 156.455 60.795 156.625 ;
        RECT 60.165 156.115 60.335 156.285 ;
        RECT 63.385 156.115 63.555 156.285 ;
        RECT 65.225 157.135 65.395 157.305 ;
        RECT 66.145 156.795 66.315 156.965 ;
        RECT 65.685 156.455 65.855 156.625 ;
        RECT 64.305 156.115 64.475 156.285 ;
        RECT 67.065 156.455 67.235 156.625 ;
        RECT 68.445 156.455 68.615 156.625 ;
        RECT 71.665 156.455 71.835 156.625 ;
        RECT 67.985 155.435 68.155 155.605 ;
        RECT 78.565 157.135 78.735 157.305 ;
        RECT 73.045 156.455 73.215 156.625 ;
        RECT 73.965 156.455 74.135 156.625 ;
        RECT 74.425 156.455 74.595 156.625 ;
        RECT 72.585 155.435 72.755 155.605 ;
        RECT 73.505 156.115 73.675 156.285 ;
        RECT 76.265 156.455 76.435 156.625 ;
        RECT 76.725 156.115 76.895 156.285 ;
        RECT 77.185 156.115 77.355 156.285 ;
        RECT 77.645 156.115 77.815 156.285 ;
        RECT 75.345 155.435 75.515 155.605 ;
        RECT 79.025 156.455 79.195 156.625 ;
        RECT 79.945 156.455 80.115 156.625 ;
        RECT 80.405 156.455 80.575 156.625 ;
        RECT 83.625 157.135 83.795 157.305 ;
        RECT 82.245 156.455 82.415 156.625 ;
        RECT 82.705 156.115 82.875 156.285 ;
        RECT 83.165 156.115 83.335 156.285 ;
        RECT 85.005 156.455 85.175 156.625 ;
        RECT 84.545 156.115 84.715 156.285 ;
        RECT 86.385 156.455 86.555 156.625 ;
        RECT 87.305 156.455 87.475 156.625 ;
        RECT 85.925 155.435 86.095 155.605 ;
        RECT 86.845 155.775 87.015 155.945 ;
        RECT 89.605 155.775 89.775 155.945 ;
        RECT 89.145 155.435 89.315 155.605 ;
        RECT 91.445 156.115 91.615 156.285 ;
        RECT 93.205 156.795 93.375 156.965 ;
        RECT 94.205 156.795 94.375 156.965 ;
        RECT 94.665 156.455 94.835 156.625 ;
        RECT 98.805 157.135 98.975 157.305 ;
        RECT 92.365 155.435 92.535 155.605 ;
        RECT 93.285 155.435 93.455 155.605 ;
        RECT 95.585 155.775 95.755 155.945 ;
        RECT 99.725 156.455 99.895 156.625 ;
        RECT 101.475 156.455 101.645 156.625 ;
        RECT 102.025 156.455 102.195 156.625 ;
        RECT 101.105 155.435 101.275 155.605 ;
        RECT 102.945 156.455 103.115 156.625 ;
        RECT 102.485 155.435 102.655 155.605 ;
        RECT 108.925 156.455 109.095 156.625 ;
        RECT 109.845 156.455 110.015 156.625 ;
        RECT 110.305 156.455 110.475 156.625 ;
        RECT 110.765 156.455 110.935 156.625 ;
        RECT 113.985 156.455 114.155 156.625 ;
        RECT 112.145 155.435 112.315 155.605 ;
        RECT 114.905 156.455 115.075 156.625 ;
        RECT 114.445 155.435 114.615 155.605 ;
        RECT 119.965 156.455 120.135 156.625 ;
        RECT 120.885 156.455 121.055 156.625 ;
        RECT 123.645 156.795 123.815 156.965 ;
        RECT 119.965 155.435 120.135 155.605 ;
        RECT 124.105 156.455 124.275 156.625 ;
        RECT 124.565 156.455 124.735 156.625 ;
        RECT 126.405 157.135 126.575 157.305 ;
        RECT 128.245 156.795 128.415 156.965 ;
        RECT 126.865 156.455 127.035 156.625 ;
        RECT 129.295 157.135 129.465 157.305 ;
        RECT 133.305 157.135 133.475 157.305 ;
        RECT 125.485 155.435 125.655 155.605 ;
        RECT 131.465 156.455 131.635 156.625 ;
        RECT 132.385 156.455 132.555 156.625 ;
        RECT 129.165 155.435 129.335 155.605 ;
        RECT 130.085 155.435 130.255 155.605 ;
        RECT 134.685 156.455 134.855 156.625 ;
        RECT 139.745 156.455 139.915 156.625 ;
        RECT 133.765 155.435 133.935 155.605 ;
        RECT 140.230 155.775 140.400 155.945 ;
        RECT 140.625 156.115 140.795 156.285 ;
        RECT 140.970 156.795 141.140 156.965 ;
        RECT 141.815 156.115 141.985 156.285 ;
        RECT 142.330 155.775 142.500 155.945 ;
        RECT 143.900 155.775 144.070 155.945 ;
        RECT 144.335 156.115 144.505 156.285 ;
        RECT 146.645 157.135 146.815 157.305 ;
        RECT 36.245 154.925 36.415 155.095 ;
        RECT 36.705 154.925 36.875 155.095 ;
        RECT 37.165 154.925 37.335 155.095 ;
        RECT 37.625 154.925 37.795 155.095 ;
        RECT 38.085 154.925 38.255 155.095 ;
        RECT 38.545 154.925 38.715 155.095 ;
        RECT 39.005 154.925 39.175 155.095 ;
        RECT 39.465 154.925 39.635 155.095 ;
        RECT 39.925 154.925 40.095 155.095 ;
        RECT 40.385 154.925 40.555 155.095 ;
        RECT 40.845 154.925 41.015 155.095 ;
        RECT 41.305 154.925 41.475 155.095 ;
        RECT 41.765 154.925 41.935 155.095 ;
        RECT 42.225 154.925 42.395 155.095 ;
        RECT 42.685 154.925 42.855 155.095 ;
        RECT 43.145 154.925 43.315 155.095 ;
        RECT 43.605 154.925 43.775 155.095 ;
        RECT 44.065 154.925 44.235 155.095 ;
        RECT 44.525 154.925 44.695 155.095 ;
        RECT 44.985 154.925 45.155 155.095 ;
        RECT 45.445 154.925 45.615 155.095 ;
        RECT 45.905 154.925 46.075 155.095 ;
        RECT 46.365 154.925 46.535 155.095 ;
        RECT 46.825 154.925 46.995 155.095 ;
        RECT 47.285 154.925 47.455 155.095 ;
        RECT 47.745 154.925 47.915 155.095 ;
        RECT 48.205 154.925 48.375 155.095 ;
        RECT 48.665 154.925 48.835 155.095 ;
        RECT 49.125 154.925 49.295 155.095 ;
        RECT 49.585 154.925 49.755 155.095 ;
        RECT 50.045 154.925 50.215 155.095 ;
        RECT 50.505 154.925 50.675 155.095 ;
        RECT 50.965 154.925 51.135 155.095 ;
        RECT 51.425 154.925 51.595 155.095 ;
        RECT 51.885 154.925 52.055 155.095 ;
        RECT 52.345 154.925 52.515 155.095 ;
        RECT 52.805 154.925 52.975 155.095 ;
        RECT 53.265 154.925 53.435 155.095 ;
        RECT 53.725 154.925 53.895 155.095 ;
        RECT 54.185 154.925 54.355 155.095 ;
        RECT 54.645 154.925 54.815 155.095 ;
        RECT 55.105 154.925 55.275 155.095 ;
        RECT 55.565 154.925 55.735 155.095 ;
        RECT 56.025 154.925 56.195 155.095 ;
        RECT 56.485 154.925 56.655 155.095 ;
        RECT 56.945 154.925 57.115 155.095 ;
        RECT 57.405 154.925 57.575 155.095 ;
        RECT 57.865 154.925 58.035 155.095 ;
        RECT 58.325 154.925 58.495 155.095 ;
        RECT 58.785 154.925 58.955 155.095 ;
        RECT 59.245 154.925 59.415 155.095 ;
        RECT 59.705 154.925 59.875 155.095 ;
        RECT 60.165 154.925 60.335 155.095 ;
        RECT 60.625 154.925 60.795 155.095 ;
        RECT 61.085 154.925 61.255 155.095 ;
        RECT 61.545 154.925 61.715 155.095 ;
        RECT 62.005 154.925 62.175 155.095 ;
        RECT 62.465 154.925 62.635 155.095 ;
        RECT 62.925 154.925 63.095 155.095 ;
        RECT 63.385 154.925 63.555 155.095 ;
        RECT 63.845 154.925 64.015 155.095 ;
        RECT 64.305 154.925 64.475 155.095 ;
        RECT 64.765 154.925 64.935 155.095 ;
        RECT 65.225 154.925 65.395 155.095 ;
        RECT 65.685 154.925 65.855 155.095 ;
        RECT 66.145 154.925 66.315 155.095 ;
        RECT 66.605 154.925 66.775 155.095 ;
        RECT 67.065 154.925 67.235 155.095 ;
        RECT 67.525 154.925 67.695 155.095 ;
        RECT 67.985 154.925 68.155 155.095 ;
        RECT 68.445 154.925 68.615 155.095 ;
        RECT 68.905 154.925 69.075 155.095 ;
        RECT 69.365 154.925 69.535 155.095 ;
        RECT 69.825 154.925 69.995 155.095 ;
        RECT 70.285 154.925 70.455 155.095 ;
        RECT 70.745 154.925 70.915 155.095 ;
        RECT 71.205 154.925 71.375 155.095 ;
        RECT 71.665 154.925 71.835 155.095 ;
        RECT 72.125 154.925 72.295 155.095 ;
        RECT 72.585 154.925 72.755 155.095 ;
        RECT 73.045 154.925 73.215 155.095 ;
        RECT 73.505 154.925 73.675 155.095 ;
        RECT 73.965 154.925 74.135 155.095 ;
        RECT 74.425 154.925 74.595 155.095 ;
        RECT 74.885 154.925 75.055 155.095 ;
        RECT 75.345 154.925 75.515 155.095 ;
        RECT 75.805 154.925 75.975 155.095 ;
        RECT 76.265 154.925 76.435 155.095 ;
        RECT 76.725 154.925 76.895 155.095 ;
        RECT 77.185 154.925 77.355 155.095 ;
        RECT 77.645 154.925 77.815 155.095 ;
        RECT 78.105 154.925 78.275 155.095 ;
        RECT 78.565 154.925 78.735 155.095 ;
        RECT 79.025 154.925 79.195 155.095 ;
        RECT 79.485 154.925 79.655 155.095 ;
        RECT 79.945 154.925 80.115 155.095 ;
        RECT 80.405 154.925 80.575 155.095 ;
        RECT 80.865 154.925 81.035 155.095 ;
        RECT 81.325 154.925 81.495 155.095 ;
        RECT 81.785 154.925 81.955 155.095 ;
        RECT 82.245 154.925 82.415 155.095 ;
        RECT 82.705 154.925 82.875 155.095 ;
        RECT 83.165 154.925 83.335 155.095 ;
        RECT 83.625 154.925 83.795 155.095 ;
        RECT 84.085 154.925 84.255 155.095 ;
        RECT 84.545 154.925 84.715 155.095 ;
        RECT 85.005 154.925 85.175 155.095 ;
        RECT 85.465 154.925 85.635 155.095 ;
        RECT 85.925 154.925 86.095 155.095 ;
        RECT 86.385 154.925 86.555 155.095 ;
        RECT 86.845 154.925 87.015 155.095 ;
        RECT 87.305 154.925 87.475 155.095 ;
        RECT 87.765 154.925 87.935 155.095 ;
        RECT 88.225 154.925 88.395 155.095 ;
        RECT 88.685 154.925 88.855 155.095 ;
        RECT 89.145 154.925 89.315 155.095 ;
        RECT 89.605 154.925 89.775 155.095 ;
        RECT 90.065 154.925 90.235 155.095 ;
        RECT 90.525 154.925 90.695 155.095 ;
        RECT 90.985 154.925 91.155 155.095 ;
        RECT 91.445 154.925 91.615 155.095 ;
        RECT 91.905 154.925 92.075 155.095 ;
        RECT 92.365 154.925 92.535 155.095 ;
        RECT 92.825 154.925 92.995 155.095 ;
        RECT 93.285 154.925 93.455 155.095 ;
        RECT 93.745 154.925 93.915 155.095 ;
        RECT 94.205 154.925 94.375 155.095 ;
        RECT 94.665 154.925 94.835 155.095 ;
        RECT 95.125 154.925 95.295 155.095 ;
        RECT 95.585 154.925 95.755 155.095 ;
        RECT 96.045 154.925 96.215 155.095 ;
        RECT 96.505 154.925 96.675 155.095 ;
        RECT 96.965 154.925 97.135 155.095 ;
        RECT 97.425 154.925 97.595 155.095 ;
        RECT 97.885 154.925 98.055 155.095 ;
        RECT 98.345 154.925 98.515 155.095 ;
        RECT 98.805 154.925 98.975 155.095 ;
        RECT 99.265 154.925 99.435 155.095 ;
        RECT 99.725 154.925 99.895 155.095 ;
        RECT 100.185 154.925 100.355 155.095 ;
        RECT 100.645 154.925 100.815 155.095 ;
        RECT 101.105 154.925 101.275 155.095 ;
        RECT 101.565 154.925 101.735 155.095 ;
        RECT 102.025 154.925 102.195 155.095 ;
        RECT 102.485 154.925 102.655 155.095 ;
        RECT 102.945 154.925 103.115 155.095 ;
        RECT 103.405 154.925 103.575 155.095 ;
        RECT 103.865 154.925 104.035 155.095 ;
        RECT 104.325 154.925 104.495 155.095 ;
        RECT 104.785 154.925 104.955 155.095 ;
        RECT 105.245 154.925 105.415 155.095 ;
        RECT 105.705 154.925 105.875 155.095 ;
        RECT 106.165 154.925 106.335 155.095 ;
        RECT 106.625 154.925 106.795 155.095 ;
        RECT 107.085 154.925 107.255 155.095 ;
        RECT 107.545 154.925 107.715 155.095 ;
        RECT 108.005 154.925 108.175 155.095 ;
        RECT 108.465 154.925 108.635 155.095 ;
        RECT 108.925 154.925 109.095 155.095 ;
        RECT 109.385 154.925 109.555 155.095 ;
        RECT 109.845 154.925 110.015 155.095 ;
        RECT 110.305 154.925 110.475 155.095 ;
        RECT 110.765 154.925 110.935 155.095 ;
        RECT 111.225 154.925 111.395 155.095 ;
        RECT 111.685 154.925 111.855 155.095 ;
        RECT 112.145 154.925 112.315 155.095 ;
        RECT 112.605 154.925 112.775 155.095 ;
        RECT 113.065 154.925 113.235 155.095 ;
        RECT 113.525 154.925 113.695 155.095 ;
        RECT 113.985 154.925 114.155 155.095 ;
        RECT 114.445 154.925 114.615 155.095 ;
        RECT 114.905 154.925 115.075 155.095 ;
        RECT 115.365 154.925 115.535 155.095 ;
        RECT 115.825 154.925 115.995 155.095 ;
        RECT 116.285 154.925 116.455 155.095 ;
        RECT 116.745 154.925 116.915 155.095 ;
        RECT 117.205 154.925 117.375 155.095 ;
        RECT 117.665 154.925 117.835 155.095 ;
        RECT 118.125 154.925 118.295 155.095 ;
        RECT 118.585 154.925 118.755 155.095 ;
        RECT 119.045 154.925 119.215 155.095 ;
        RECT 119.505 154.925 119.675 155.095 ;
        RECT 119.965 154.925 120.135 155.095 ;
        RECT 120.425 154.925 120.595 155.095 ;
        RECT 120.885 154.925 121.055 155.095 ;
        RECT 121.345 154.925 121.515 155.095 ;
        RECT 121.805 154.925 121.975 155.095 ;
        RECT 122.265 154.925 122.435 155.095 ;
        RECT 122.725 154.925 122.895 155.095 ;
        RECT 123.185 154.925 123.355 155.095 ;
        RECT 123.645 154.925 123.815 155.095 ;
        RECT 124.105 154.925 124.275 155.095 ;
        RECT 124.565 154.925 124.735 155.095 ;
        RECT 125.025 154.925 125.195 155.095 ;
        RECT 125.485 154.925 125.655 155.095 ;
        RECT 125.945 154.925 126.115 155.095 ;
        RECT 126.405 154.925 126.575 155.095 ;
        RECT 126.865 154.925 127.035 155.095 ;
        RECT 127.325 154.925 127.495 155.095 ;
        RECT 127.785 154.925 127.955 155.095 ;
        RECT 128.245 154.925 128.415 155.095 ;
        RECT 128.705 154.925 128.875 155.095 ;
        RECT 129.165 154.925 129.335 155.095 ;
        RECT 129.625 154.925 129.795 155.095 ;
        RECT 130.085 154.925 130.255 155.095 ;
        RECT 130.545 154.925 130.715 155.095 ;
        RECT 131.005 154.925 131.175 155.095 ;
        RECT 131.465 154.925 131.635 155.095 ;
        RECT 131.925 154.925 132.095 155.095 ;
        RECT 132.385 154.925 132.555 155.095 ;
        RECT 132.845 154.925 133.015 155.095 ;
        RECT 133.305 154.925 133.475 155.095 ;
        RECT 133.765 154.925 133.935 155.095 ;
        RECT 134.225 154.925 134.395 155.095 ;
        RECT 134.685 154.925 134.855 155.095 ;
        RECT 135.145 154.925 135.315 155.095 ;
        RECT 135.605 154.925 135.775 155.095 ;
        RECT 136.065 154.925 136.235 155.095 ;
        RECT 136.525 154.925 136.695 155.095 ;
        RECT 136.985 154.925 137.155 155.095 ;
        RECT 137.445 154.925 137.615 155.095 ;
        RECT 137.905 154.925 138.075 155.095 ;
        RECT 138.365 154.925 138.535 155.095 ;
        RECT 138.825 154.925 138.995 155.095 ;
        RECT 139.285 154.925 139.455 155.095 ;
        RECT 139.745 154.925 139.915 155.095 ;
        RECT 140.205 154.925 140.375 155.095 ;
        RECT 140.665 154.925 140.835 155.095 ;
        RECT 141.125 154.925 141.295 155.095 ;
        RECT 141.585 154.925 141.755 155.095 ;
        RECT 142.045 154.925 142.215 155.095 ;
        RECT 142.505 154.925 142.675 155.095 ;
        RECT 142.965 154.925 143.135 155.095 ;
        RECT 143.425 154.925 143.595 155.095 ;
        RECT 143.885 154.925 144.055 155.095 ;
        RECT 144.345 154.925 144.515 155.095 ;
        RECT 144.805 154.925 144.975 155.095 ;
        RECT 145.265 154.925 145.435 155.095 ;
        RECT 145.725 154.925 145.895 155.095 ;
        RECT 146.185 154.925 146.355 155.095 ;
        RECT 146.645 154.925 146.815 155.095 ;
        RECT 147.105 154.925 147.275 155.095 ;
        RECT 147.565 154.925 147.735 155.095 ;
        RECT 148.025 154.925 148.195 155.095 ;
        RECT 148.485 154.925 148.655 155.095 ;
        RECT 148.945 154.925 149.115 155.095 ;
        RECT 149.405 154.925 149.575 155.095 ;
        RECT 149.865 154.925 150.035 155.095 ;
        RECT 40.385 154.415 40.555 154.585 ;
        RECT 41.305 153.395 41.475 153.565 ;
        RECT 43.145 153.395 43.315 153.565 ;
        RECT 45.445 154.075 45.615 154.245 ;
        RECT 47.285 154.415 47.455 154.585 ;
        RECT 44.985 153.395 45.155 153.565 ;
        RECT 45.905 153.395 46.075 153.565 ;
        RECT 42.225 152.715 42.395 152.885 ;
        RECT 49.585 154.415 49.755 154.585 ;
        RECT 47.055 153.225 47.225 153.395 ;
        RECT 46.365 152.715 46.535 152.885 ;
        RECT 48.205 153.055 48.375 153.225 ;
        RECT 50.505 153.395 50.675 153.565 ;
        RECT 51.425 153.395 51.595 153.565 ;
        RECT 66.145 154.415 66.315 154.585 ;
        RECT 65.225 152.715 65.395 152.885 ;
        RECT 66.145 152.715 66.315 152.885 ;
        RECT 67.985 153.395 68.155 153.565 ;
        RECT 71.665 153.395 71.835 153.565 ;
        RECT 72.585 153.055 72.755 153.225 ;
        RECT 78.105 153.395 78.275 153.565 ;
        RECT 70.745 152.715 70.915 152.885 ;
        RECT 79.485 153.395 79.655 153.565 ;
        RECT 79.945 153.395 80.115 153.565 ;
        RECT 80.500 153.395 80.670 153.565 ;
        RECT 81.325 153.395 81.495 153.565 ;
        RECT 79.025 152.715 79.195 152.885 ;
        RECT 83.165 153.395 83.335 153.565 ;
        RECT 84.085 153.395 84.255 153.565 ;
        RECT 85.925 153.395 86.095 153.565 ;
        RECT 87.305 153.735 87.475 153.905 ;
        RECT 82.245 152.715 82.415 152.885 ;
        RECT 85.005 152.715 85.175 152.885 ;
        RECT 96.965 154.415 97.135 154.585 ;
        RECT 100.185 154.415 100.355 154.585 ;
        RECT 97.885 153.395 98.055 153.565 ;
        RECT 99.265 153.055 99.435 153.225 ;
        RECT 101.565 153.735 101.735 153.905 ;
        RECT 102.025 153.735 102.195 153.905 ;
        RECT 102.485 153.395 102.655 153.565 ;
        RECT 102.945 153.735 103.115 153.905 ;
        RECT 103.865 152.715 104.035 152.885 ;
        RECT 105.245 153.395 105.415 153.565 ;
        RECT 105.705 153.735 105.875 153.905 ;
        RECT 106.165 153.735 106.335 153.905 ;
        RECT 106.625 153.735 106.795 153.905 ;
        RECT 104.325 152.715 104.495 152.885 ;
        RECT 108.465 153.395 108.635 153.565 ;
        RECT 109.385 153.055 109.555 153.225 ;
        RECT 109.845 154.415 110.015 154.585 ;
        RECT 110.765 153.395 110.935 153.565 ;
        RECT 111.225 153.395 111.395 153.565 ;
        RECT 111.685 153.395 111.855 153.565 ;
        RECT 112.145 153.735 112.315 153.905 ;
        RECT 113.985 153.395 114.155 153.565 ;
        RECT 114.445 153.735 114.615 153.905 ;
        RECT 114.905 153.735 115.075 153.905 ;
        RECT 115.365 153.735 115.535 153.905 ;
        RECT 116.285 153.395 116.455 153.565 ;
        RECT 118.125 153.395 118.295 153.565 ;
        RECT 119.045 153.395 119.215 153.565 ;
        RECT 116.745 153.055 116.915 153.225 ;
        RECT 113.065 152.715 113.235 152.885 ;
        RECT 127.325 153.395 127.495 153.565 ;
        RECT 128.245 153.395 128.415 153.565 ;
        RECT 130.085 153.395 130.255 153.565 ;
        RECT 131.925 154.415 132.095 154.585 ;
        RECT 132.845 154.075 133.015 154.245 ;
        RECT 127.325 152.715 127.495 152.885 ;
        RECT 131.925 153.055 132.095 153.225 ;
        RECT 133.305 153.055 133.475 153.225 ;
        RECT 134.225 153.055 134.395 153.225 ;
        RECT 135.145 153.055 135.315 153.225 ;
        RECT 138.825 153.395 138.995 153.565 ;
        RECT 139.745 152.715 139.915 152.885 ;
        RECT 36.245 152.205 36.415 152.375 ;
        RECT 36.705 152.205 36.875 152.375 ;
        RECT 37.165 152.205 37.335 152.375 ;
        RECT 37.625 152.205 37.795 152.375 ;
        RECT 38.085 152.205 38.255 152.375 ;
        RECT 38.545 152.205 38.715 152.375 ;
        RECT 39.005 152.205 39.175 152.375 ;
        RECT 39.465 152.205 39.635 152.375 ;
        RECT 39.925 152.205 40.095 152.375 ;
        RECT 40.385 152.205 40.555 152.375 ;
        RECT 40.845 152.205 41.015 152.375 ;
        RECT 41.305 152.205 41.475 152.375 ;
        RECT 41.765 152.205 41.935 152.375 ;
        RECT 42.225 152.205 42.395 152.375 ;
        RECT 42.685 152.205 42.855 152.375 ;
        RECT 43.145 152.205 43.315 152.375 ;
        RECT 43.605 152.205 43.775 152.375 ;
        RECT 44.065 152.205 44.235 152.375 ;
        RECT 44.525 152.205 44.695 152.375 ;
        RECT 44.985 152.205 45.155 152.375 ;
        RECT 45.445 152.205 45.615 152.375 ;
        RECT 45.905 152.205 46.075 152.375 ;
        RECT 46.365 152.205 46.535 152.375 ;
        RECT 46.825 152.205 46.995 152.375 ;
        RECT 47.285 152.205 47.455 152.375 ;
        RECT 47.745 152.205 47.915 152.375 ;
        RECT 48.205 152.205 48.375 152.375 ;
        RECT 48.665 152.205 48.835 152.375 ;
        RECT 49.125 152.205 49.295 152.375 ;
        RECT 49.585 152.205 49.755 152.375 ;
        RECT 50.045 152.205 50.215 152.375 ;
        RECT 50.505 152.205 50.675 152.375 ;
        RECT 50.965 152.205 51.135 152.375 ;
        RECT 51.425 152.205 51.595 152.375 ;
        RECT 51.885 152.205 52.055 152.375 ;
        RECT 52.345 152.205 52.515 152.375 ;
        RECT 52.805 152.205 52.975 152.375 ;
        RECT 53.265 152.205 53.435 152.375 ;
        RECT 53.725 152.205 53.895 152.375 ;
        RECT 54.185 152.205 54.355 152.375 ;
        RECT 54.645 152.205 54.815 152.375 ;
        RECT 55.105 152.205 55.275 152.375 ;
        RECT 55.565 152.205 55.735 152.375 ;
        RECT 56.025 152.205 56.195 152.375 ;
        RECT 56.485 152.205 56.655 152.375 ;
        RECT 56.945 152.205 57.115 152.375 ;
        RECT 57.405 152.205 57.575 152.375 ;
        RECT 57.865 152.205 58.035 152.375 ;
        RECT 58.325 152.205 58.495 152.375 ;
        RECT 58.785 152.205 58.955 152.375 ;
        RECT 59.245 152.205 59.415 152.375 ;
        RECT 59.705 152.205 59.875 152.375 ;
        RECT 60.165 152.205 60.335 152.375 ;
        RECT 60.625 152.205 60.795 152.375 ;
        RECT 61.085 152.205 61.255 152.375 ;
        RECT 61.545 152.205 61.715 152.375 ;
        RECT 62.005 152.205 62.175 152.375 ;
        RECT 62.465 152.205 62.635 152.375 ;
        RECT 62.925 152.205 63.095 152.375 ;
        RECT 63.385 152.205 63.555 152.375 ;
        RECT 63.845 152.205 64.015 152.375 ;
        RECT 64.305 152.205 64.475 152.375 ;
        RECT 64.765 152.205 64.935 152.375 ;
        RECT 65.225 152.205 65.395 152.375 ;
        RECT 65.685 152.205 65.855 152.375 ;
        RECT 66.145 152.205 66.315 152.375 ;
        RECT 66.605 152.205 66.775 152.375 ;
        RECT 67.065 152.205 67.235 152.375 ;
        RECT 67.525 152.205 67.695 152.375 ;
        RECT 67.985 152.205 68.155 152.375 ;
        RECT 68.445 152.205 68.615 152.375 ;
        RECT 68.905 152.205 69.075 152.375 ;
        RECT 69.365 152.205 69.535 152.375 ;
        RECT 69.825 152.205 69.995 152.375 ;
        RECT 70.285 152.205 70.455 152.375 ;
        RECT 70.745 152.205 70.915 152.375 ;
        RECT 71.205 152.205 71.375 152.375 ;
        RECT 71.665 152.205 71.835 152.375 ;
        RECT 72.125 152.205 72.295 152.375 ;
        RECT 72.585 152.205 72.755 152.375 ;
        RECT 73.045 152.205 73.215 152.375 ;
        RECT 73.505 152.205 73.675 152.375 ;
        RECT 73.965 152.205 74.135 152.375 ;
        RECT 74.425 152.205 74.595 152.375 ;
        RECT 74.885 152.205 75.055 152.375 ;
        RECT 75.345 152.205 75.515 152.375 ;
        RECT 75.805 152.205 75.975 152.375 ;
        RECT 76.265 152.205 76.435 152.375 ;
        RECT 76.725 152.205 76.895 152.375 ;
        RECT 77.185 152.205 77.355 152.375 ;
        RECT 77.645 152.205 77.815 152.375 ;
        RECT 78.105 152.205 78.275 152.375 ;
        RECT 78.565 152.205 78.735 152.375 ;
        RECT 79.025 152.205 79.195 152.375 ;
        RECT 79.485 152.205 79.655 152.375 ;
        RECT 79.945 152.205 80.115 152.375 ;
        RECT 80.405 152.205 80.575 152.375 ;
        RECT 80.865 152.205 81.035 152.375 ;
        RECT 81.325 152.205 81.495 152.375 ;
        RECT 81.785 152.205 81.955 152.375 ;
        RECT 82.245 152.205 82.415 152.375 ;
        RECT 82.705 152.205 82.875 152.375 ;
        RECT 83.165 152.205 83.335 152.375 ;
        RECT 83.625 152.205 83.795 152.375 ;
        RECT 84.085 152.205 84.255 152.375 ;
        RECT 84.545 152.205 84.715 152.375 ;
        RECT 85.005 152.205 85.175 152.375 ;
        RECT 85.465 152.205 85.635 152.375 ;
        RECT 85.925 152.205 86.095 152.375 ;
        RECT 86.385 152.205 86.555 152.375 ;
        RECT 86.845 152.205 87.015 152.375 ;
        RECT 87.305 152.205 87.475 152.375 ;
        RECT 87.765 152.205 87.935 152.375 ;
        RECT 88.225 152.205 88.395 152.375 ;
        RECT 88.685 152.205 88.855 152.375 ;
        RECT 89.145 152.205 89.315 152.375 ;
        RECT 89.605 152.205 89.775 152.375 ;
        RECT 90.065 152.205 90.235 152.375 ;
        RECT 90.525 152.205 90.695 152.375 ;
        RECT 90.985 152.205 91.155 152.375 ;
        RECT 91.445 152.205 91.615 152.375 ;
        RECT 91.905 152.205 92.075 152.375 ;
        RECT 92.365 152.205 92.535 152.375 ;
        RECT 92.825 152.205 92.995 152.375 ;
        RECT 93.285 152.205 93.455 152.375 ;
        RECT 93.745 152.205 93.915 152.375 ;
        RECT 94.205 152.205 94.375 152.375 ;
        RECT 94.665 152.205 94.835 152.375 ;
        RECT 95.125 152.205 95.295 152.375 ;
        RECT 95.585 152.205 95.755 152.375 ;
        RECT 96.045 152.205 96.215 152.375 ;
        RECT 96.505 152.205 96.675 152.375 ;
        RECT 96.965 152.205 97.135 152.375 ;
        RECT 97.425 152.205 97.595 152.375 ;
        RECT 97.885 152.205 98.055 152.375 ;
        RECT 98.345 152.205 98.515 152.375 ;
        RECT 98.805 152.205 98.975 152.375 ;
        RECT 99.265 152.205 99.435 152.375 ;
        RECT 99.725 152.205 99.895 152.375 ;
        RECT 100.185 152.205 100.355 152.375 ;
        RECT 100.645 152.205 100.815 152.375 ;
        RECT 101.105 152.205 101.275 152.375 ;
        RECT 101.565 152.205 101.735 152.375 ;
        RECT 102.025 152.205 102.195 152.375 ;
        RECT 102.485 152.205 102.655 152.375 ;
        RECT 102.945 152.205 103.115 152.375 ;
        RECT 103.405 152.205 103.575 152.375 ;
        RECT 103.865 152.205 104.035 152.375 ;
        RECT 104.325 152.205 104.495 152.375 ;
        RECT 104.785 152.205 104.955 152.375 ;
        RECT 105.245 152.205 105.415 152.375 ;
        RECT 105.705 152.205 105.875 152.375 ;
        RECT 106.165 152.205 106.335 152.375 ;
        RECT 106.625 152.205 106.795 152.375 ;
        RECT 107.085 152.205 107.255 152.375 ;
        RECT 107.545 152.205 107.715 152.375 ;
        RECT 108.005 152.205 108.175 152.375 ;
        RECT 108.465 152.205 108.635 152.375 ;
        RECT 108.925 152.205 109.095 152.375 ;
        RECT 109.385 152.205 109.555 152.375 ;
        RECT 109.845 152.205 110.015 152.375 ;
        RECT 110.305 152.205 110.475 152.375 ;
        RECT 110.765 152.205 110.935 152.375 ;
        RECT 111.225 152.205 111.395 152.375 ;
        RECT 111.685 152.205 111.855 152.375 ;
        RECT 112.145 152.205 112.315 152.375 ;
        RECT 112.605 152.205 112.775 152.375 ;
        RECT 113.065 152.205 113.235 152.375 ;
        RECT 113.525 152.205 113.695 152.375 ;
        RECT 113.985 152.205 114.155 152.375 ;
        RECT 114.445 152.205 114.615 152.375 ;
        RECT 114.905 152.205 115.075 152.375 ;
        RECT 115.365 152.205 115.535 152.375 ;
        RECT 115.825 152.205 115.995 152.375 ;
        RECT 116.285 152.205 116.455 152.375 ;
        RECT 116.745 152.205 116.915 152.375 ;
        RECT 117.205 152.205 117.375 152.375 ;
        RECT 117.665 152.205 117.835 152.375 ;
        RECT 118.125 152.205 118.295 152.375 ;
        RECT 118.585 152.205 118.755 152.375 ;
        RECT 119.045 152.205 119.215 152.375 ;
        RECT 119.505 152.205 119.675 152.375 ;
        RECT 119.965 152.205 120.135 152.375 ;
        RECT 120.425 152.205 120.595 152.375 ;
        RECT 120.885 152.205 121.055 152.375 ;
        RECT 121.345 152.205 121.515 152.375 ;
        RECT 121.805 152.205 121.975 152.375 ;
        RECT 122.265 152.205 122.435 152.375 ;
        RECT 122.725 152.205 122.895 152.375 ;
        RECT 123.185 152.205 123.355 152.375 ;
        RECT 123.645 152.205 123.815 152.375 ;
        RECT 124.105 152.205 124.275 152.375 ;
        RECT 124.565 152.205 124.735 152.375 ;
        RECT 125.025 152.205 125.195 152.375 ;
        RECT 125.485 152.205 125.655 152.375 ;
        RECT 125.945 152.205 126.115 152.375 ;
        RECT 126.405 152.205 126.575 152.375 ;
        RECT 126.865 152.205 127.035 152.375 ;
        RECT 127.325 152.205 127.495 152.375 ;
        RECT 127.785 152.205 127.955 152.375 ;
        RECT 128.245 152.205 128.415 152.375 ;
        RECT 128.705 152.205 128.875 152.375 ;
        RECT 129.165 152.205 129.335 152.375 ;
        RECT 129.625 152.205 129.795 152.375 ;
        RECT 130.085 152.205 130.255 152.375 ;
        RECT 130.545 152.205 130.715 152.375 ;
        RECT 131.005 152.205 131.175 152.375 ;
        RECT 131.465 152.205 131.635 152.375 ;
        RECT 131.925 152.205 132.095 152.375 ;
        RECT 132.385 152.205 132.555 152.375 ;
        RECT 132.845 152.205 133.015 152.375 ;
        RECT 133.305 152.205 133.475 152.375 ;
        RECT 133.765 152.205 133.935 152.375 ;
        RECT 134.225 152.205 134.395 152.375 ;
        RECT 134.685 152.205 134.855 152.375 ;
        RECT 135.145 152.205 135.315 152.375 ;
        RECT 135.605 152.205 135.775 152.375 ;
        RECT 136.065 152.205 136.235 152.375 ;
        RECT 136.525 152.205 136.695 152.375 ;
        RECT 136.985 152.205 137.155 152.375 ;
        RECT 137.445 152.205 137.615 152.375 ;
        RECT 137.905 152.205 138.075 152.375 ;
        RECT 138.365 152.205 138.535 152.375 ;
        RECT 138.825 152.205 138.995 152.375 ;
        RECT 139.285 152.205 139.455 152.375 ;
        RECT 139.745 152.205 139.915 152.375 ;
        RECT 140.205 152.205 140.375 152.375 ;
        RECT 140.665 152.205 140.835 152.375 ;
        RECT 141.125 152.205 141.295 152.375 ;
        RECT 141.585 152.205 141.755 152.375 ;
        RECT 142.045 152.205 142.215 152.375 ;
        RECT 142.505 152.205 142.675 152.375 ;
        RECT 142.965 152.205 143.135 152.375 ;
        RECT 143.425 152.205 143.595 152.375 ;
        RECT 143.885 152.205 144.055 152.375 ;
        RECT 144.345 152.205 144.515 152.375 ;
        RECT 144.805 152.205 144.975 152.375 ;
        RECT 145.265 152.205 145.435 152.375 ;
        RECT 145.725 152.205 145.895 152.375 ;
        RECT 146.185 152.205 146.355 152.375 ;
        RECT 146.645 152.205 146.815 152.375 ;
        RECT 147.105 152.205 147.275 152.375 ;
        RECT 147.565 152.205 147.735 152.375 ;
        RECT 148.025 152.205 148.195 152.375 ;
        RECT 148.485 152.205 148.655 152.375 ;
        RECT 148.945 152.205 149.115 152.375 ;
        RECT 149.405 152.205 149.575 152.375 ;
        RECT 149.865 152.205 150.035 152.375 ;
        RECT 39.005 151.015 39.175 151.185 ;
        RECT 39.490 150.335 39.660 150.505 ;
        RECT 39.885 150.675 40.055 150.845 ;
        RECT 40.340 151.355 40.510 151.525 ;
        RECT 41.075 150.675 41.245 150.845 ;
        RECT 41.590 150.335 41.760 150.505 ;
        RECT 43.160 150.335 43.330 150.505 ;
        RECT 43.595 150.675 43.765 150.845 ;
        RECT 45.905 151.695 46.075 151.865 ;
        RECT 47.745 151.015 47.915 151.185 ;
        RECT 49.125 151.015 49.295 151.185 ;
        RECT 53.265 151.015 53.435 151.185 ;
        RECT 52.345 149.995 52.515 150.165 ;
        RECT 55.565 150.675 55.735 150.845 ;
        RECT 56.945 150.675 57.115 150.845 ;
        RECT 82.245 151.695 82.415 151.865 ;
        RECT 80.865 151.355 81.035 151.525 ;
        RECT 81.785 151.355 81.955 151.525 ;
        RECT 82.245 151.015 82.415 151.185 ;
        RECT 83.165 151.015 83.335 151.185 ;
        RECT 84.085 151.015 84.255 151.185 ;
        RECT 84.545 151.015 84.715 151.185 ;
        RECT 83.625 150.335 83.795 150.505 ;
        RECT 85.005 150.675 85.175 150.845 ;
        RECT 88.685 150.675 88.855 150.845 ;
        RECT 89.145 150.675 89.315 150.845 ;
        RECT 89.605 151.015 89.775 151.185 ;
        RECT 90.065 151.015 90.235 151.185 ;
        RECT 91.445 151.015 91.615 151.185 ;
        RECT 90.985 149.995 91.155 150.165 ;
        RECT 92.825 150.675 92.995 150.845 ;
        RECT 99.265 150.935 99.435 151.105 ;
        RECT 101.105 151.355 101.275 151.525 ;
        RECT 98.345 149.995 98.515 150.165 ;
        RECT 103.405 150.675 103.575 150.845 ;
        RECT 102.485 150.335 102.655 150.505 ;
        RECT 104.785 151.015 104.955 151.185 ;
        RECT 103.865 149.995 104.035 150.165 ;
        RECT 113.985 150.675 114.155 150.845 ;
        RECT 114.905 151.015 115.075 151.185 ;
        RECT 115.365 150.335 115.535 150.505 ;
        RECT 116.285 151.015 116.455 151.185 ;
        RECT 115.825 150.675 115.995 150.845 ;
        RECT 117.205 151.015 117.375 151.185 ;
        RECT 124.565 151.015 124.735 151.185 ;
        RECT 125.025 149.995 125.195 150.165 ;
        RECT 127.785 151.015 127.955 151.185 ;
        RECT 128.705 151.015 128.875 151.185 ;
        RECT 131.465 151.355 131.635 151.525 ;
        RECT 129.625 150.675 129.795 150.845 ;
        RECT 130.545 150.675 130.715 150.845 ;
        RECT 131.925 151.015 132.095 151.185 ;
        RECT 131.465 150.675 131.635 150.845 ;
        RECT 132.845 151.015 133.015 151.185 ;
        RECT 132.845 149.995 133.015 150.165 ;
        RECT 140.665 151.015 140.835 151.185 ;
        RECT 141.150 150.335 141.320 150.505 ;
        RECT 141.545 150.675 141.715 150.845 ;
        RECT 141.890 151.355 142.060 151.525 ;
        RECT 142.735 150.675 142.905 150.845 ;
        RECT 143.250 150.335 143.420 150.505 ;
        RECT 144.820 150.335 144.990 150.505 ;
        RECT 145.255 150.675 145.425 150.845 ;
        RECT 147.565 151.695 147.735 151.865 ;
        RECT 36.245 149.485 36.415 149.655 ;
        RECT 36.705 149.485 36.875 149.655 ;
        RECT 37.165 149.485 37.335 149.655 ;
        RECT 37.625 149.485 37.795 149.655 ;
        RECT 38.085 149.485 38.255 149.655 ;
        RECT 38.545 149.485 38.715 149.655 ;
        RECT 39.005 149.485 39.175 149.655 ;
        RECT 39.465 149.485 39.635 149.655 ;
        RECT 39.925 149.485 40.095 149.655 ;
        RECT 40.385 149.485 40.555 149.655 ;
        RECT 40.845 149.485 41.015 149.655 ;
        RECT 41.305 149.485 41.475 149.655 ;
        RECT 41.765 149.485 41.935 149.655 ;
        RECT 42.225 149.485 42.395 149.655 ;
        RECT 42.685 149.485 42.855 149.655 ;
        RECT 43.145 149.485 43.315 149.655 ;
        RECT 43.605 149.485 43.775 149.655 ;
        RECT 44.065 149.485 44.235 149.655 ;
        RECT 44.525 149.485 44.695 149.655 ;
        RECT 44.985 149.485 45.155 149.655 ;
        RECT 45.445 149.485 45.615 149.655 ;
        RECT 45.905 149.485 46.075 149.655 ;
        RECT 46.365 149.485 46.535 149.655 ;
        RECT 46.825 149.485 46.995 149.655 ;
        RECT 47.285 149.485 47.455 149.655 ;
        RECT 47.745 149.485 47.915 149.655 ;
        RECT 48.205 149.485 48.375 149.655 ;
        RECT 48.665 149.485 48.835 149.655 ;
        RECT 49.125 149.485 49.295 149.655 ;
        RECT 49.585 149.485 49.755 149.655 ;
        RECT 50.045 149.485 50.215 149.655 ;
        RECT 50.505 149.485 50.675 149.655 ;
        RECT 50.965 149.485 51.135 149.655 ;
        RECT 51.425 149.485 51.595 149.655 ;
        RECT 51.885 149.485 52.055 149.655 ;
        RECT 52.345 149.485 52.515 149.655 ;
        RECT 52.805 149.485 52.975 149.655 ;
        RECT 53.265 149.485 53.435 149.655 ;
        RECT 53.725 149.485 53.895 149.655 ;
        RECT 54.185 149.485 54.355 149.655 ;
        RECT 54.645 149.485 54.815 149.655 ;
        RECT 55.105 149.485 55.275 149.655 ;
        RECT 55.565 149.485 55.735 149.655 ;
        RECT 56.025 149.485 56.195 149.655 ;
        RECT 56.485 149.485 56.655 149.655 ;
        RECT 56.945 149.485 57.115 149.655 ;
        RECT 57.405 149.485 57.575 149.655 ;
        RECT 57.865 149.485 58.035 149.655 ;
        RECT 58.325 149.485 58.495 149.655 ;
        RECT 58.785 149.485 58.955 149.655 ;
        RECT 59.245 149.485 59.415 149.655 ;
        RECT 59.705 149.485 59.875 149.655 ;
        RECT 60.165 149.485 60.335 149.655 ;
        RECT 60.625 149.485 60.795 149.655 ;
        RECT 61.085 149.485 61.255 149.655 ;
        RECT 61.545 149.485 61.715 149.655 ;
        RECT 62.005 149.485 62.175 149.655 ;
        RECT 62.465 149.485 62.635 149.655 ;
        RECT 62.925 149.485 63.095 149.655 ;
        RECT 63.385 149.485 63.555 149.655 ;
        RECT 63.845 149.485 64.015 149.655 ;
        RECT 64.305 149.485 64.475 149.655 ;
        RECT 64.765 149.485 64.935 149.655 ;
        RECT 65.225 149.485 65.395 149.655 ;
        RECT 65.685 149.485 65.855 149.655 ;
        RECT 66.145 149.485 66.315 149.655 ;
        RECT 66.605 149.485 66.775 149.655 ;
        RECT 67.065 149.485 67.235 149.655 ;
        RECT 67.525 149.485 67.695 149.655 ;
        RECT 67.985 149.485 68.155 149.655 ;
        RECT 68.445 149.485 68.615 149.655 ;
        RECT 68.905 149.485 69.075 149.655 ;
        RECT 69.365 149.485 69.535 149.655 ;
        RECT 69.825 149.485 69.995 149.655 ;
        RECT 70.285 149.485 70.455 149.655 ;
        RECT 70.745 149.485 70.915 149.655 ;
        RECT 71.205 149.485 71.375 149.655 ;
        RECT 71.665 149.485 71.835 149.655 ;
        RECT 72.125 149.485 72.295 149.655 ;
        RECT 72.585 149.485 72.755 149.655 ;
        RECT 73.045 149.485 73.215 149.655 ;
        RECT 73.505 149.485 73.675 149.655 ;
        RECT 73.965 149.485 74.135 149.655 ;
        RECT 74.425 149.485 74.595 149.655 ;
        RECT 74.885 149.485 75.055 149.655 ;
        RECT 75.345 149.485 75.515 149.655 ;
        RECT 75.805 149.485 75.975 149.655 ;
        RECT 76.265 149.485 76.435 149.655 ;
        RECT 76.725 149.485 76.895 149.655 ;
        RECT 77.185 149.485 77.355 149.655 ;
        RECT 77.645 149.485 77.815 149.655 ;
        RECT 78.105 149.485 78.275 149.655 ;
        RECT 78.565 149.485 78.735 149.655 ;
        RECT 79.025 149.485 79.195 149.655 ;
        RECT 79.485 149.485 79.655 149.655 ;
        RECT 79.945 149.485 80.115 149.655 ;
        RECT 80.405 149.485 80.575 149.655 ;
        RECT 80.865 149.485 81.035 149.655 ;
        RECT 81.325 149.485 81.495 149.655 ;
        RECT 81.785 149.485 81.955 149.655 ;
        RECT 82.245 149.485 82.415 149.655 ;
        RECT 82.705 149.485 82.875 149.655 ;
        RECT 83.165 149.485 83.335 149.655 ;
        RECT 83.625 149.485 83.795 149.655 ;
        RECT 84.085 149.485 84.255 149.655 ;
        RECT 84.545 149.485 84.715 149.655 ;
        RECT 85.005 149.485 85.175 149.655 ;
        RECT 85.465 149.485 85.635 149.655 ;
        RECT 85.925 149.485 86.095 149.655 ;
        RECT 86.385 149.485 86.555 149.655 ;
        RECT 86.845 149.485 87.015 149.655 ;
        RECT 87.305 149.485 87.475 149.655 ;
        RECT 87.765 149.485 87.935 149.655 ;
        RECT 88.225 149.485 88.395 149.655 ;
        RECT 88.685 149.485 88.855 149.655 ;
        RECT 89.145 149.485 89.315 149.655 ;
        RECT 89.605 149.485 89.775 149.655 ;
        RECT 90.065 149.485 90.235 149.655 ;
        RECT 90.525 149.485 90.695 149.655 ;
        RECT 90.985 149.485 91.155 149.655 ;
        RECT 91.445 149.485 91.615 149.655 ;
        RECT 91.905 149.485 92.075 149.655 ;
        RECT 92.365 149.485 92.535 149.655 ;
        RECT 92.825 149.485 92.995 149.655 ;
        RECT 93.285 149.485 93.455 149.655 ;
        RECT 93.745 149.485 93.915 149.655 ;
        RECT 94.205 149.485 94.375 149.655 ;
        RECT 94.665 149.485 94.835 149.655 ;
        RECT 95.125 149.485 95.295 149.655 ;
        RECT 95.585 149.485 95.755 149.655 ;
        RECT 96.045 149.485 96.215 149.655 ;
        RECT 96.505 149.485 96.675 149.655 ;
        RECT 96.965 149.485 97.135 149.655 ;
        RECT 97.425 149.485 97.595 149.655 ;
        RECT 97.885 149.485 98.055 149.655 ;
        RECT 98.345 149.485 98.515 149.655 ;
        RECT 98.805 149.485 98.975 149.655 ;
        RECT 99.265 149.485 99.435 149.655 ;
        RECT 99.725 149.485 99.895 149.655 ;
        RECT 100.185 149.485 100.355 149.655 ;
        RECT 100.645 149.485 100.815 149.655 ;
        RECT 101.105 149.485 101.275 149.655 ;
        RECT 101.565 149.485 101.735 149.655 ;
        RECT 102.025 149.485 102.195 149.655 ;
        RECT 102.485 149.485 102.655 149.655 ;
        RECT 102.945 149.485 103.115 149.655 ;
        RECT 103.405 149.485 103.575 149.655 ;
        RECT 103.865 149.485 104.035 149.655 ;
        RECT 104.325 149.485 104.495 149.655 ;
        RECT 104.785 149.485 104.955 149.655 ;
        RECT 105.245 149.485 105.415 149.655 ;
        RECT 105.705 149.485 105.875 149.655 ;
        RECT 106.165 149.485 106.335 149.655 ;
        RECT 106.625 149.485 106.795 149.655 ;
        RECT 107.085 149.485 107.255 149.655 ;
        RECT 107.545 149.485 107.715 149.655 ;
        RECT 108.005 149.485 108.175 149.655 ;
        RECT 108.465 149.485 108.635 149.655 ;
        RECT 108.925 149.485 109.095 149.655 ;
        RECT 109.385 149.485 109.555 149.655 ;
        RECT 109.845 149.485 110.015 149.655 ;
        RECT 110.305 149.485 110.475 149.655 ;
        RECT 110.765 149.485 110.935 149.655 ;
        RECT 111.225 149.485 111.395 149.655 ;
        RECT 111.685 149.485 111.855 149.655 ;
        RECT 112.145 149.485 112.315 149.655 ;
        RECT 112.605 149.485 112.775 149.655 ;
        RECT 113.065 149.485 113.235 149.655 ;
        RECT 113.525 149.485 113.695 149.655 ;
        RECT 113.985 149.485 114.155 149.655 ;
        RECT 114.445 149.485 114.615 149.655 ;
        RECT 114.905 149.485 115.075 149.655 ;
        RECT 115.365 149.485 115.535 149.655 ;
        RECT 115.825 149.485 115.995 149.655 ;
        RECT 116.285 149.485 116.455 149.655 ;
        RECT 116.745 149.485 116.915 149.655 ;
        RECT 117.205 149.485 117.375 149.655 ;
        RECT 117.665 149.485 117.835 149.655 ;
        RECT 118.125 149.485 118.295 149.655 ;
        RECT 118.585 149.485 118.755 149.655 ;
        RECT 119.045 149.485 119.215 149.655 ;
        RECT 119.505 149.485 119.675 149.655 ;
        RECT 119.965 149.485 120.135 149.655 ;
        RECT 120.425 149.485 120.595 149.655 ;
        RECT 120.885 149.485 121.055 149.655 ;
        RECT 121.345 149.485 121.515 149.655 ;
        RECT 121.805 149.485 121.975 149.655 ;
        RECT 122.265 149.485 122.435 149.655 ;
        RECT 122.725 149.485 122.895 149.655 ;
        RECT 123.185 149.485 123.355 149.655 ;
        RECT 123.645 149.485 123.815 149.655 ;
        RECT 124.105 149.485 124.275 149.655 ;
        RECT 124.565 149.485 124.735 149.655 ;
        RECT 125.025 149.485 125.195 149.655 ;
        RECT 125.485 149.485 125.655 149.655 ;
        RECT 125.945 149.485 126.115 149.655 ;
        RECT 126.405 149.485 126.575 149.655 ;
        RECT 126.865 149.485 127.035 149.655 ;
        RECT 127.325 149.485 127.495 149.655 ;
        RECT 127.785 149.485 127.955 149.655 ;
        RECT 128.245 149.485 128.415 149.655 ;
        RECT 128.705 149.485 128.875 149.655 ;
        RECT 129.165 149.485 129.335 149.655 ;
        RECT 129.625 149.485 129.795 149.655 ;
        RECT 130.085 149.485 130.255 149.655 ;
        RECT 130.545 149.485 130.715 149.655 ;
        RECT 131.005 149.485 131.175 149.655 ;
        RECT 131.465 149.485 131.635 149.655 ;
        RECT 131.925 149.485 132.095 149.655 ;
        RECT 132.385 149.485 132.555 149.655 ;
        RECT 132.845 149.485 133.015 149.655 ;
        RECT 133.305 149.485 133.475 149.655 ;
        RECT 133.765 149.485 133.935 149.655 ;
        RECT 134.225 149.485 134.395 149.655 ;
        RECT 134.685 149.485 134.855 149.655 ;
        RECT 135.145 149.485 135.315 149.655 ;
        RECT 135.605 149.485 135.775 149.655 ;
        RECT 136.065 149.485 136.235 149.655 ;
        RECT 136.525 149.485 136.695 149.655 ;
        RECT 136.985 149.485 137.155 149.655 ;
        RECT 137.445 149.485 137.615 149.655 ;
        RECT 137.905 149.485 138.075 149.655 ;
        RECT 138.365 149.485 138.535 149.655 ;
        RECT 138.825 149.485 138.995 149.655 ;
        RECT 139.285 149.485 139.455 149.655 ;
        RECT 139.745 149.485 139.915 149.655 ;
        RECT 140.205 149.485 140.375 149.655 ;
        RECT 140.665 149.485 140.835 149.655 ;
        RECT 141.125 149.485 141.295 149.655 ;
        RECT 141.585 149.485 141.755 149.655 ;
        RECT 142.045 149.485 142.215 149.655 ;
        RECT 142.505 149.485 142.675 149.655 ;
        RECT 142.965 149.485 143.135 149.655 ;
        RECT 143.425 149.485 143.595 149.655 ;
        RECT 143.885 149.485 144.055 149.655 ;
        RECT 144.345 149.485 144.515 149.655 ;
        RECT 144.805 149.485 144.975 149.655 ;
        RECT 145.265 149.485 145.435 149.655 ;
        RECT 145.725 149.485 145.895 149.655 ;
        RECT 146.185 149.485 146.355 149.655 ;
        RECT 146.645 149.485 146.815 149.655 ;
        RECT 147.105 149.485 147.275 149.655 ;
        RECT 147.565 149.485 147.735 149.655 ;
        RECT 148.025 149.485 148.195 149.655 ;
        RECT 148.485 149.485 148.655 149.655 ;
        RECT 148.945 149.485 149.115 149.655 ;
        RECT 149.405 149.485 149.575 149.655 ;
        RECT 149.865 149.485 150.035 149.655 ;
        RECT 41.765 148.635 41.935 148.805 ;
        RECT 41.305 147.955 41.475 148.125 ;
        RECT 40.385 147.275 40.555 147.445 ;
        RECT 42.685 147.955 42.855 148.125 ;
        RECT 52.345 148.295 52.515 148.465 ;
        RECT 54.185 148.295 54.355 148.465 ;
        RECT 53.265 147.955 53.435 148.125 ;
        RECT 54.645 147.955 54.815 148.125 ;
        RECT 56.025 147.955 56.195 148.125 ;
        RECT 55.105 147.615 55.275 147.785 ;
        RECT 56.945 148.295 57.115 148.465 ;
        RECT 63.845 148.975 64.015 149.145 ;
        RECT 57.865 148.295 58.035 148.465 ;
        RECT 58.325 147.955 58.495 148.125 ;
        RECT 60.165 148.295 60.335 148.465 ;
        RECT 61.315 147.615 61.485 147.785 ;
        RECT 62.925 147.955 63.095 148.125 ;
        RECT 62.005 147.615 62.175 147.785 ;
        RECT 62.465 147.615 62.635 147.785 ;
        RECT 67.065 148.635 67.235 148.805 ;
        RECT 66.145 147.955 66.315 148.125 ;
        RECT 69.365 148.635 69.535 148.805 ;
        RECT 68.905 147.955 69.075 148.125 ;
        RECT 70.745 148.295 70.915 148.465 ;
        RECT 69.825 147.955 69.995 148.125 ;
        RECT 70.285 147.955 70.455 148.125 ;
        RECT 71.205 147.955 71.375 148.125 ;
        RECT 72.125 147.955 72.295 148.125 ;
        RECT 72.585 148.295 72.755 148.465 ;
        RECT 73.045 148.295 73.215 148.465 ;
        RECT 73.505 147.955 73.675 148.125 ;
        RECT 75.805 148.295 75.975 148.465 ;
        RECT 76.265 148.295 76.435 148.465 ;
        RECT 76.725 147.955 76.895 148.125 ;
        RECT 78.105 148.975 78.275 149.145 ;
        RECT 80.405 148.975 80.575 149.145 ;
        RECT 77.185 147.955 77.355 148.125 ;
        RECT 74.425 147.275 74.595 147.445 ;
        RECT 78.565 148.295 78.735 148.465 ;
        RECT 79.485 147.955 79.655 148.125 ;
        RECT 81.325 147.955 81.495 148.125 ;
        RECT 82.245 147.955 82.415 148.125 ;
        RECT 83.165 147.955 83.335 148.125 ;
        RECT 85.465 148.295 85.635 148.465 ;
        RECT 85.925 147.955 86.095 148.125 ;
        RECT 86.385 148.295 86.555 148.465 ;
        RECT 86.845 147.955 87.015 148.125 ;
        RECT 89.145 147.955 89.315 148.125 ;
        RECT 89.605 147.955 89.775 148.125 ;
        RECT 90.065 147.955 90.235 148.125 ;
        RECT 84.545 147.275 84.715 147.445 ;
        RECT 87.765 147.275 87.935 147.445 ;
        RECT 90.985 147.955 91.155 148.125 ;
        RECT 95.125 148.295 95.295 148.465 ;
        RECT 94.665 147.955 94.835 148.125 ;
        RECT 95.585 147.955 95.755 148.125 ;
        RECT 99.725 147.615 99.895 147.785 ;
        RECT 99.265 147.275 99.435 147.445 ;
        RECT 102.025 147.615 102.195 147.785 ;
        RECT 101.565 147.275 101.735 147.445 ;
        RECT 106.165 147.615 106.335 147.785 ;
        RECT 111.685 147.955 111.855 148.125 ;
        RECT 112.145 147.955 112.315 148.125 ;
        RECT 112.605 147.955 112.775 148.125 ;
        RECT 106.625 147.275 106.795 147.445 ;
        RECT 110.305 147.275 110.475 147.445 ;
        RECT 113.525 147.955 113.695 148.125 ;
        RECT 114.445 147.955 114.615 148.125 ;
        RECT 114.905 148.295 115.075 148.465 ;
        RECT 115.365 148.295 115.535 148.465 ;
        RECT 115.825 147.955 115.995 148.125 ;
        RECT 116.745 147.275 116.915 147.445 ;
        RECT 118.125 148.295 118.295 148.465 ;
        RECT 119.045 147.955 119.215 148.125 ;
        RECT 123.645 148.635 123.815 148.805 ;
        RECT 120.385 147.965 120.555 148.135 ;
        RECT 119.965 147.615 120.135 147.785 ;
        RECT 121.345 147.955 121.515 148.125 ;
        RECT 122.725 147.955 122.895 148.125 ;
        RECT 123.645 147.955 123.815 148.125 ;
        RECT 120.425 147.275 120.595 147.445 ;
        RECT 127.785 148.975 127.955 149.145 ;
        RECT 125.485 147.615 125.655 147.785 ;
        RECT 129.165 147.955 129.335 148.125 ;
        RECT 126.865 147.275 127.035 147.445 ;
        RECT 136.985 148.295 137.155 148.465 ;
        RECT 142.045 148.975 142.215 149.145 ;
        RECT 139.745 148.295 139.915 148.465 ;
        RECT 137.905 147.955 138.075 148.125 ;
        RECT 139.285 147.955 139.455 148.125 ;
        RECT 138.825 147.275 138.995 147.445 ;
        RECT 141.585 148.295 141.755 148.465 ;
        RECT 140.665 147.955 140.835 148.125 ;
        RECT 142.965 147.955 143.135 148.125 ;
        RECT 144.385 147.925 144.555 148.095 ;
        RECT 143.885 147.275 144.055 147.445 ;
        RECT 36.245 146.765 36.415 146.935 ;
        RECT 36.705 146.765 36.875 146.935 ;
        RECT 37.165 146.765 37.335 146.935 ;
        RECT 37.625 146.765 37.795 146.935 ;
        RECT 38.085 146.765 38.255 146.935 ;
        RECT 38.545 146.765 38.715 146.935 ;
        RECT 39.005 146.765 39.175 146.935 ;
        RECT 39.465 146.765 39.635 146.935 ;
        RECT 39.925 146.765 40.095 146.935 ;
        RECT 40.385 146.765 40.555 146.935 ;
        RECT 40.845 146.765 41.015 146.935 ;
        RECT 41.305 146.765 41.475 146.935 ;
        RECT 41.765 146.765 41.935 146.935 ;
        RECT 42.225 146.765 42.395 146.935 ;
        RECT 42.685 146.765 42.855 146.935 ;
        RECT 43.145 146.765 43.315 146.935 ;
        RECT 43.605 146.765 43.775 146.935 ;
        RECT 44.065 146.765 44.235 146.935 ;
        RECT 44.525 146.765 44.695 146.935 ;
        RECT 44.985 146.765 45.155 146.935 ;
        RECT 45.445 146.765 45.615 146.935 ;
        RECT 45.905 146.765 46.075 146.935 ;
        RECT 46.365 146.765 46.535 146.935 ;
        RECT 46.825 146.765 46.995 146.935 ;
        RECT 47.285 146.765 47.455 146.935 ;
        RECT 47.745 146.765 47.915 146.935 ;
        RECT 48.205 146.765 48.375 146.935 ;
        RECT 48.665 146.765 48.835 146.935 ;
        RECT 49.125 146.765 49.295 146.935 ;
        RECT 49.585 146.765 49.755 146.935 ;
        RECT 50.045 146.765 50.215 146.935 ;
        RECT 50.505 146.765 50.675 146.935 ;
        RECT 50.965 146.765 51.135 146.935 ;
        RECT 51.425 146.765 51.595 146.935 ;
        RECT 51.885 146.765 52.055 146.935 ;
        RECT 52.345 146.765 52.515 146.935 ;
        RECT 52.805 146.765 52.975 146.935 ;
        RECT 53.265 146.765 53.435 146.935 ;
        RECT 53.725 146.765 53.895 146.935 ;
        RECT 54.185 146.765 54.355 146.935 ;
        RECT 54.645 146.765 54.815 146.935 ;
        RECT 55.105 146.765 55.275 146.935 ;
        RECT 55.565 146.765 55.735 146.935 ;
        RECT 56.025 146.765 56.195 146.935 ;
        RECT 56.485 146.765 56.655 146.935 ;
        RECT 56.945 146.765 57.115 146.935 ;
        RECT 57.405 146.765 57.575 146.935 ;
        RECT 57.865 146.765 58.035 146.935 ;
        RECT 58.325 146.765 58.495 146.935 ;
        RECT 58.785 146.765 58.955 146.935 ;
        RECT 59.245 146.765 59.415 146.935 ;
        RECT 59.705 146.765 59.875 146.935 ;
        RECT 60.165 146.765 60.335 146.935 ;
        RECT 60.625 146.765 60.795 146.935 ;
        RECT 61.085 146.765 61.255 146.935 ;
        RECT 61.545 146.765 61.715 146.935 ;
        RECT 62.005 146.765 62.175 146.935 ;
        RECT 62.465 146.765 62.635 146.935 ;
        RECT 62.925 146.765 63.095 146.935 ;
        RECT 63.385 146.765 63.555 146.935 ;
        RECT 63.845 146.765 64.015 146.935 ;
        RECT 64.305 146.765 64.475 146.935 ;
        RECT 64.765 146.765 64.935 146.935 ;
        RECT 65.225 146.765 65.395 146.935 ;
        RECT 65.685 146.765 65.855 146.935 ;
        RECT 66.145 146.765 66.315 146.935 ;
        RECT 66.605 146.765 66.775 146.935 ;
        RECT 67.065 146.765 67.235 146.935 ;
        RECT 67.525 146.765 67.695 146.935 ;
        RECT 67.985 146.765 68.155 146.935 ;
        RECT 68.445 146.765 68.615 146.935 ;
        RECT 68.905 146.765 69.075 146.935 ;
        RECT 69.365 146.765 69.535 146.935 ;
        RECT 69.825 146.765 69.995 146.935 ;
        RECT 70.285 146.765 70.455 146.935 ;
        RECT 70.745 146.765 70.915 146.935 ;
        RECT 71.205 146.765 71.375 146.935 ;
        RECT 71.665 146.765 71.835 146.935 ;
        RECT 72.125 146.765 72.295 146.935 ;
        RECT 72.585 146.765 72.755 146.935 ;
        RECT 73.045 146.765 73.215 146.935 ;
        RECT 73.505 146.765 73.675 146.935 ;
        RECT 73.965 146.765 74.135 146.935 ;
        RECT 74.425 146.765 74.595 146.935 ;
        RECT 74.885 146.765 75.055 146.935 ;
        RECT 75.345 146.765 75.515 146.935 ;
        RECT 75.805 146.765 75.975 146.935 ;
        RECT 76.265 146.765 76.435 146.935 ;
        RECT 76.725 146.765 76.895 146.935 ;
        RECT 77.185 146.765 77.355 146.935 ;
        RECT 77.645 146.765 77.815 146.935 ;
        RECT 78.105 146.765 78.275 146.935 ;
        RECT 78.565 146.765 78.735 146.935 ;
        RECT 79.025 146.765 79.195 146.935 ;
        RECT 79.485 146.765 79.655 146.935 ;
        RECT 79.945 146.765 80.115 146.935 ;
        RECT 80.405 146.765 80.575 146.935 ;
        RECT 80.865 146.765 81.035 146.935 ;
        RECT 81.325 146.765 81.495 146.935 ;
        RECT 81.785 146.765 81.955 146.935 ;
        RECT 82.245 146.765 82.415 146.935 ;
        RECT 82.705 146.765 82.875 146.935 ;
        RECT 83.165 146.765 83.335 146.935 ;
        RECT 83.625 146.765 83.795 146.935 ;
        RECT 84.085 146.765 84.255 146.935 ;
        RECT 84.545 146.765 84.715 146.935 ;
        RECT 85.005 146.765 85.175 146.935 ;
        RECT 85.465 146.765 85.635 146.935 ;
        RECT 85.925 146.765 86.095 146.935 ;
        RECT 86.385 146.765 86.555 146.935 ;
        RECT 86.845 146.765 87.015 146.935 ;
        RECT 87.305 146.765 87.475 146.935 ;
        RECT 87.765 146.765 87.935 146.935 ;
        RECT 88.225 146.765 88.395 146.935 ;
        RECT 88.685 146.765 88.855 146.935 ;
        RECT 89.145 146.765 89.315 146.935 ;
        RECT 89.605 146.765 89.775 146.935 ;
        RECT 90.065 146.765 90.235 146.935 ;
        RECT 90.525 146.765 90.695 146.935 ;
        RECT 90.985 146.765 91.155 146.935 ;
        RECT 91.445 146.765 91.615 146.935 ;
        RECT 91.905 146.765 92.075 146.935 ;
        RECT 92.365 146.765 92.535 146.935 ;
        RECT 92.825 146.765 92.995 146.935 ;
        RECT 93.285 146.765 93.455 146.935 ;
        RECT 93.745 146.765 93.915 146.935 ;
        RECT 94.205 146.765 94.375 146.935 ;
        RECT 94.665 146.765 94.835 146.935 ;
        RECT 95.125 146.765 95.295 146.935 ;
        RECT 95.585 146.765 95.755 146.935 ;
        RECT 96.045 146.765 96.215 146.935 ;
        RECT 96.505 146.765 96.675 146.935 ;
        RECT 96.965 146.765 97.135 146.935 ;
        RECT 97.425 146.765 97.595 146.935 ;
        RECT 97.885 146.765 98.055 146.935 ;
        RECT 98.345 146.765 98.515 146.935 ;
        RECT 98.805 146.765 98.975 146.935 ;
        RECT 99.265 146.765 99.435 146.935 ;
        RECT 99.725 146.765 99.895 146.935 ;
        RECT 100.185 146.765 100.355 146.935 ;
        RECT 100.645 146.765 100.815 146.935 ;
        RECT 101.105 146.765 101.275 146.935 ;
        RECT 101.565 146.765 101.735 146.935 ;
        RECT 102.025 146.765 102.195 146.935 ;
        RECT 102.485 146.765 102.655 146.935 ;
        RECT 102.945 146.765 103.115 146.935 ;
        RECT 103.405 146.765 103.575 146.935 ;
        RECT 103.865 146.765 104.035 146.935 ;
        RECT 104.325 146.765 104.495 146.935 ;
        RECT 104.785 146.765 104.955 146.935 ;
        RECT 105.245 146.765 105.415 146.935 ;
        RECT 105.705 146.765 105.875 146.935 ;
        RECT 106.165 146.765 106.335 146.935 ;
        RECT 106.625 146.765 106.795 146.935 ;
        RECT 107.085 146.765 107.255 146.935 ;
        RECT 107.545 146.765 107.715 146.935 ;
        RECT 108.005 146.765 108.175 146.935 ;
        RECT 108.465 146.765 108.635 146.935 ;
        RECT 108.925 146.765 109.095 146.935 ;
        RECT 109.385 146.765 109.555 146.935 ;
        RECT 109.845 146.765 110.015 146.935 ;
        RECT 110.305 146.765 110.475 146.935 ;
        RECT 110.765 146.765 110.935 146.935 ;
        RECT 111.225 146.765 111.395 146.935 ;
        RECT 111.685 146.765 111.855 146.935 ;
        RECT 112.145 146.765 112.315 146.935 ;
        RECT 112.605 146.765 112.775 146.935 ;
        RECT 113.065 146.765 113.235 146.935 ;
        RECT 113.525 146.765 113.695 146.935 ;
        RECT 113.985 146.765 114.155 146.935 ;
        RECT 114.445 146.765 114.615 146.935 ;
        RECT 114.905 146.765 115.075 146.935 ;
        RECT 115.365 146.765 115.535 146.935 ;
        RECT 115.825 146.765 115.995 146.935 ;
        RECT 116.285 146.765 116.455 146.935 ;
        RECT 116.745 146.765 116.915 146.935 ;
        RECT 117.205 146.765 117.375 146.935 ;
        RECT 117.665 146.765 117.835 146.935 ;
        RECT 118.125 146.765 118.295 146.935 ;
        RECT 118.585 146.765 118.755 146.935 ;
        RECT 119.045 146.765 119.215 146.935 ;
        RECT 119.505 146.765 119.675 146.935 ;
        RECT 119.965 146.765 120.135 146.935 ;
        RECT 120.425 146.765 120.595 146.935 ;
        RECT 120.885 146.765 121.055 146.935 ;
        RECT 121.345 146.765 121.515 146.935 ;
        RECT 121.805 146.765 121.975 146.935 ;
        RECT 122.265 146.765 122.435 146.935 ;
        RECT 122.725 146.765 122.895 146.935 ;
        RECT 123.185 146.765 123.355 146.935 ;
        RECT 123.645 146.765 123.815 146.935 ;
        RECT 124.105 146.765 124.275 146.935 ;
        RECT 124.565 146.765 124.735 146.935 ;
        RECT 125.025 146.765 125.195 146.935 ;
        RECT 125.485 146.765 125.655 146.935 ;
        RECT 125.945 146.765 126.115 146.935 ;
        RECT 126.405 146.765 126.575 146.935 ;
        RECT 126.865 146.765 127.035 146.935 ;
        RECT 127.325 146.765 127.495 146.935 ;
        RECT 127.785 146.765 127.955 146.935 ;
        RECT 128.245 146.765 128.415 146.935 ;
        RECT 128.705 146.765 128.875 146.935 ;
        RECT 129.165 146.765 129.335 146.935 ;
        RECT 129.625 146.765 129.795 146.935 ;
        RECT 130.085 146.765 130.255 146.935 ;
        RECT 130.545 146.765 130.715 146.935 ;
        RECT 131.005 146.765 131.175 146.935 ;
        RECT 131.465 146.765 131.635 146.935 ;
        RECT 131.925 146.765 132.095 146.935 ;
        RECT 132.385 146.765 132.555 146.935 ;
        RECT 132.845 146.765 133.015 146.935 ;
        RECT 133.305 146.765 133.475 146.935 ;
        RECT 133.765 146.765 133.935 146.935 ;
        RECT 134.225 146.765 134.395 146.935 ;
        RECT 134.685 146.765 134.855 146.935 ;
        RECT 135.145 146.765 135.315 146.935 ;
        RECT 135.605 146.765 135.775 146.935 ;
        RECT 136.065 146.765 136.235 146.935 ;
        RECT 136.525 146.765 136.695 146.935 ;
        RECT 136.985 146.765 137.155 146.935 ;
        RECT 137.445 146.765 137.615 146.935 ;
        RECT 137.905 146.765 138.075 146.935 ;
        RECT 138.365 146.765 138.535 146.935 ;
        RECT 138.825 146.765 138.995 146.935 ;
        RECT 139.285 146.765 139.455 146.935 ;
        RECT 139.745 146.765 139.915 146.935 ;
        RECT 140.205 146.765 140.375 146.935 ;
        RECT 140.665 146.765 140.835 146.935 ;
        RECT 141.125 146.765 141.295 146.935 ;
        RECT 141.585 146.765 141.755 146.935 ;
        RECT 142.045 146.765 142.215 146.935 ;
        RECT 142.505 146.765 142.675 146.935 ;
        RECT 142.965 146.765 143.135 146.935 ;
        RECT 143.425 146.765 143.595 146.935 ;
        RECT 143.885 146.765 144.055 146.935 ;
        RECT 144.345 146.765 144.515 146.935 ;
        RECT 144.805 146.765 144.975 146.935 ;
        RECT 145.265 146.765 145.435 146.935 ;
        RECT 145.725 146.765 145.895 146.935 ;
        RECT 146.185 146.765 146.355 146.935 ;
        RECT 146.645 146.765 146.815 146.935 ;
        RECT 147.105 146.765 147.275 146.935 ;
        RECT 147.565 146.765 147.735 146.935 ;
        RECT 148.025 146.765 148.195 146.935 ;
        RECT 148.485 146.765 148.655 146.935 ;
        RECT 148.945 146.765 149.115 146.935 ;
        RECT 149.405 146.765 149.575 146.935 ;
        RECT 149.865 146.765 150.035 146.935 ;
        RECT 39.465 145.575 39.635 145.745 ;
        RECT 43.145 145.915 43.315 146.085 ;
        RECT 38.085 144.555 38.255 144.725 ;
        RECT 44.525 145.235 44.695 145.405 ;
        RECT 42.225 144.895 42.395 145.065 ;
        RECT 45.010 144.895 45.180 145.065 ;
        RECT 45.405 145.235 45.575 145.405 ;
        RECT 45.860 145.915 46.030 146.085 ;
        RECT 46.595 145.235 46.765 145.405 ;
        RECT 47.110 144.895 47.280 145.065 ;
        RECT 48.680 144.895 48.850 145.065 ;
        RECT 49.115 145.235 49.285 145.405 ;
        RECT 51.425 144.895 51.595 145.065 ;
        RECT 52.805 145.575 52.975 145.745 ;
        RECT 53.265 145.235 53.435 145.405 ;
        RECT 56.025 146.255 56.195 146.425 ;
        RECT 55.105 145.575 55.275 145.745 ;
        RECT 54.645 145.235 54.815 145.405 ;
        RECT 58.325 145.575 58.495 145.745 ;
        RECT 57.865 145.235 58.035 145.405 ;
        RECT 60.165 144.895 60.335 145.065 ;
        RECT 65.225 145.575 65.395 145.745 ;
        RECT 65.685 145.575 65.855 145.745 ;
        RECT 72.125 146.255 72.295 146.425 ;
        RECT 66.605 145.575 66.775 145.745 ;
        RECT 67.985 145.575 68.155 145.745 ;
        RECT 68.905 145.575 69.075 145.745 ;
        RECT 69.365 145.575 69.535 145.745 ;
        RECT 70.285 145.575 70.455 145.745 ;
        RECT 68.905 144.555 69.075 144.725 ;
        RECT 69.825 145.235 69.995 145.405 ;
        RECT 73.045 145.575 73.215 145.745 ;
        RECT 73.505 144.895 73.675 145.065 ;
        RECT 74.425 145.575 74.595 145.745 ;
        RECT 73.965 145.235 74.135 145.405 ;
        RECT 78.565 146.255 78.735 146.425 ;
        RECT 76.265 145.575 76.435 145.745 ;
        RECT 75.345 144.555 75.515 144.725 ;
        RECT 77.185 144.555 77.355 144.725 ;
        RECT 79.485 145.575 79.655 145.745 ;
        RECT 80.405 145.575 80.575 145.745 ;
        RECT 80.865 145.575 81.035 145.745 ;
        RECT 83.165 145.575 83.335 145.745 ;
        RECT 84.085 145.575 84.255 145.745 ;
        RECT 82.245 144.555 82.415 144.725 ;
        RECT 86.385 145.575 86.555 145.745 ;
        RECT 85.005 145.235 85.175 145.405 ;
        RECT 87.305 144.555 87.475 144.725 ;
        RECT 90.065 145.575 90.235 145.745 ;
        RECT 90.525 145.575 90.695 145.745 ;
        RECT 90.985 145.575 91.155 145.745 ;
        RECT 91.905 145.575 92.075 145.745 ;
        RECT 88.685 144.895 88.855 145.065 ;
        RECT 95.585 145.575 95.755 145.745 ;
        RECT 94.205 145.235 94.375 145.405 ;
        RECT 96.505 144.555 96.675 144.725 ;
        RECT 99.265 145.575 99.435 145.745 ;
        RECT 98.345 144.555 98.515 144.725 ;
        RECT 100.185 144.555 100.355 144.725 ;
        RECT 102.025 145.575 102.195 145.745 ;
        RECT 102.945 145.575 103.115 145.745 ;
        RECT 101.105 144.555 101.275 144.725 ;
        RECT 104.785 145.575 104.955 145.745 ;
        RECT 103.865 144.895 104.035 145.065 ;
        RECT 106.165 145.575 106.335 145.745 ;
        RECT 107.085 145.575 107.255 145.745 ;
        RECT 105.245 144.555 105.415 144.725 ;
        RECT 108.005 145.575 108.175 145.745 ;
        RECT 109.385 145.575 109.555 145.745 ;
        RECT 108.925 144.555 109.095 144.725 ;
        RECT 112.145 145.575 112.315 145.745 ;
        RECT 110.765 145.235 110.935 145.405 ;
        RECT 110.305 144.895 110.475 145.065 ;
        RECT 115.365 145.575 115.535 145.745 ;
        RECT 113.065 144.555 113.235 144.725 ;
        RECT 113.985 145.235 114.155 145.405 ;
        RECT 118.125 145.575 118.295 145.745 ;
        RECT 116.745 145.235 116.915 145.405 ;
        RECT 116.285 144.555 116.455 144.725 ;
        RECT 119.505 145.575 119.675 145.745 ;
        RECT 119.045 144.895 119.215 145.065 ;
        RECT 122.265 145.575 122.435 145.745 ;
        RECT 120.885 145.235 121.055 145.405 ;
        RECT 120.425 144.555 120.595 144.725 ;
        RECT 123.645 145.915 123.815 146.085 ;
        RECT 125.485 145.575 125.655 145.745 ;
        RECT 128.245 145.575 128.415 145.745 ;
        RECT 127.785 145.235 127.955 145.405 ;
        RECT 123.185 144.555 123.355 144.725 ;
        RECT 128.245 144.555 128.415 144.725 ;
        RECT 129.165 144.555 129.335 144.725 ;
        RECT 131.925 145.235 132.095 145.405 ;
        RECT 132.410 144.895 132.580 145.065 ;
        RECT 132.805 145.235 132.975 145.405 ;
        RECT 133.205 145.575 133.375 145.745 ;
        RECT 133.995 145.235 134.165 145.405 ;
        RECT 134.510 144.895 134.680 145.065 ;
        RECT 136.080 144.895 136.250 145.065 ;
        RECT 136.515 145.235 136.685 145.405 ;
        RECT 146.645 146.255 146.815 146.425 ;
        RECT 138.825 144.895 138.995 145.065 ;
        RECT 140.665 145.575 140.835 145.745 ;
        RECT 143.425 145.575 143.595 145.745 ;
        RECT 145.725 145.575 145.895 145.745 ;
        RECT 141.125 145.235 141.295 145.405 ;
        RECT 139.745 144.555 139.915 144.725 ;
        RECT 140.665 144.555 140.835 144.725 ;
        RECT 36.245 144.045 36.415 144.215 ;
        RECT 36.705 144.045 36.875 144.215 ;
        RECT 37.165 144.045 37.335 144.215 ;
        RECT 37.625 144.045 37.795 144.215 ;
        RECT 38.085 144.045 38.255 144.215 ;
        RECT 38.545 144.045 38.715 144.215 ;
        RECT 39.005 144.045 39.175 144.215 ;
        RECT 39.465 144.045 39.635 144.215 ;
        RECT 39.925 144.045 40.095 144.215 ;
        RECT 40.385 144.045 40.555 144.215 ;
        RECT 40.845 144.045 41.015 144.215 ;
        RECT 41.305 144.045 41.475 144.215 ;
        RECT 41.765 144.045 41.935 144.215 ;
        RECT 42.225 144.045 42.395 144.215 ;
        RECT 42.685 144.045 42.855 144.215 ;
        RECT 43.145 144.045 43.315 144.215 ;
        RECT 43.605 144.045 43.775 144.215 ;
        RECT 44.065 144.045 44.235 144.215 ;
        RECT 44.525 144.045 44.695 144.215 ;
        RECT 44.985 144.045 45.155 144.215 ;
        RECT 45.445 144.045 45.615 144.215 ;
        RECT 45.905 144.045 46.075 144.215 ;
        RECT 46.365 144.045 46.535 144.215 ;
        RECT 46.825 144.045 46.995 144.215 ;
        RECT 47.285 144.045 47.455 144.215 ;
        RECT 47.745 144.045 47.915 144.215 ;
        RECT 48.205 144.045 48.375 144.215 ;
        RECT 48.665 144.045 48.835 144.215 ;
        RECT 49.125 144.045 49.295 144.215 ;
        RECT 49.585 144.045 49.755 144.215 ;
        RECT 50.045 144.045 50.215 144.215 ;
        RECT 50.505 144.045 50.675 144.215 ;
        RECT 50.965 144.045 51.135 144.215 ;
        RECT 51.425 144.045 51.595 144.215 ;
        RECT 51.885 144.045 52.055 144.215 ;
        RECT 52.345 144.045 52.515 144.215 ;
        RECT 52.805 144.045 52.975 144.215 ;
        RECT 53.265 144.045 53.435 144.215 ;
        RECT 53.725 144.045 53.895 144.215 ;
        RECT 54.185 144.045 54.355 144.215 ;
        RECT 54.645 144.045 54.815 144.215 ;
        RECT 55.105 144.045 55.275 144.215 ;
        RECT 55.565 144.045 55.735 144.215 ;
        RECT 56.025 144.045 56.195 144.215 ;
        RECT 56.485 144.045 56.655 144.215 ;
        RECT 56.945 144.045 57.115 144.215 ;
        RECT 57.405 144.045 57.575 144.215 ;
        RECT 57.865 144.045 58.035 144.215 ;
        RECT 58.325 144.045 58.495 144.215 ;
        RECT 58.785 144.045 58.955 144.215 ;
        RECT 59.245 144.045 59.415 144.215 ;
        RECT 59.705 144.045 59.875 144.215 ;
        RECT 60.165 144.045 60.335 144.215 ;
        RECT 60.625 144.045 60.795 144.215 ;
        RECT 61.085 144.045 61.255 144.215 ;
        RECT 61.545 144.045 61.715 144.215 ;
        RECT 62.005 144.045 62.175 144.215 ;
        RECT 62.465 144.045 62.635 144.215 ;
        RECT 62.925 144.045 63.095 144.215 ;
        RECT 63.385 144.045 63.555 144.215 ;
        RECT 63.845 144.045 64.015 144.215 ;
        RECT 64.305 144.045 64.475 144.215 ;
        RECT 64.765 144.045 64.935 144.215 ;
        RECT 65.225 144.045 65.395 144.215 ;
        RECT 65.685 144.045 65.855 144.215 ;
        RECT 66.145 144.045 66.315 144.215 ;
        RECT 66.605 144.045 66.775 144.215 ;
        RECT 67.065 144.045 67.235 144.215 ;
        RECT 67.525 144.045 67.695 144.215 ;
        RECT 67.985 144.045 68.155 144.215 ;
        RECT 68.445 144.045 68.615 144.215 ;
        RECT 68.905 144.045 69.075 144.215 ;
        RECT 69.365 144.045 69.535 144.215 ;
        RECT 69.825 144.045 69.995 144.215 ;
        RECT 70.285 144.045 70.455 144.215 ;
        RECT 70.745 144.045 70.915 144.215 ;
        RECT 71.205 144.045 71.375 144.215 ;
        RECT 71.665 144.045 71.835 144.215 ;
        RECT 72.125 144.045 72.295 144.215 ;
        RECT 72.585 144.045 72.755 144.215 ;
        RECT 73.045 144.045 73.215 144.215 ;
        RECT 73.505 144.045 73.675 144.215 ;
        RECT 73.965 144.045 74.135 144.215 ;
        RECT 74.425 144.045 74.595 144.215 ;
        RECT 74.885 144.045 75.055 144.215 ;
        RECT 75.345 144.045 75.515 144.215 ;
        RECT 75.805 144.045 75.975 144.215 ;
        RECT 76.265 144.045 76.435 144.215 ;
        RECT 76.725 144.045 76.895 144.215 ;
        RECT 77.185 144.045 77.355 144.215 ;
        RECT 77.645 144.045 77.815 144.215 ;
        RECT 78.105 144.045 78.275 144.215 ;
        RECT 78.565 144.045 78.735 144.215 ;
        RECT 79.025 144.045 79.195 144.215 ;
        RECT 79.485 144.045 79.655 144.215 ;
        RECT 79.945 144.045 80.115 144.215 ;
        RECT 80.405 144.045 80.575 144.215 ;
        RECT 80.865 144.045 81.035 144.215 ;
        RECT 81.325 144.045 81.495 144.215 ;
        RECT 81.785 144.045 81.955 144.215 ;
        RECT 82.245 144.045 82.415 144.215 ;
        RECT 82.705 144.045 82.875 144.215 ;
        RECT 83.165 144.045 83.335 144.215 ;
        RECT 83.625 144.045 83.795 144.215 ;
        RECT 84.085 144.045 84.255 144.215 ;
        RECT 84.545 144.045 84.715 144.215 ;
        RECT 85.005 144.045 85.175 144.215 ;
        RECT 85.465 144.045 85.635 144.215 ;
        RECT 85.925 144.045 86.095 144.215 ;
        RECT 86.385 144.045 86.555 144.215 ;
        RECT 86.845 144.045 87.015 144.215 ;
        RECT 87.305 144.045 87.475 144.215 ;
        RECT 87.765 144.045 87.935 144.215 ;
        RECT 88.225 144.045 88.395 144.215 ;
        RECT 88.685 144.045 88.855 144.215 ;
        RECT 89.145 144.045 89.315 144.215 ;
        RECT 89.605 144.045 89.775 144.215 ;
        RECT 90.065 144.045 90.235 144.215 ;
        RECT 90.525 144.045 90.695 144.215 ;
        RECT 90.985 144.045 91.155 144.215 ;
        RECT 91.445 144.045 91.615 144.215 ;
        RECT 91.905 144.045 92.075 144.215 ;
        RECT 92.365 144.045 92.535 144.215 ;
        RECT 92.825 144.045 92.995 144.215 ;
        RECT 93.285 144.045 93.455 144.215 ;
        RECT 93.745 144.045 93.915 144.215 ;
        RECT 94.205 144.045 94.375 144.215 ;
        RECT 94.665 144.045 94.835 144.215 ;
        RECT 95.125 144.045 95.295 144.215 ;
        RECT 95.585 144.045 95.755 144.215 ;
        RECT 96.045 144.045 96.215 144.215 ;
        RECT 96.505 144.045 96.675 144.215 ;
        RECT 96.965 144.045 97.135 144.215 ;
        RECT 97.425 144.045 97.595 144.215 ;
        RECT 97.885 144.045 98.055 144.215 ;
        RECT 98.345 144.045 98.515 144.215 ;
        RECT 98.805 144.045 98.975 144.215 ;
        RECT 99.265 144.045 99.435 144.215 ;
        RECT 99.725 144.045 99.895 144.215 ;
        RECT 100.185 144.045 100.355 144.215 ;
        RECT 100.645 144.045 100.815 144.215 ;
        RECT 101.105 144.045 101.275 144.215 ;
        RECT 101.565 144.045 101.735 144.215 ;
        RECT 102.025 144.045 102.195 144.215 ;
        RECT 102.485 144.045 102.655 144.215 ;
        RECT 102.945 144.045 103.115 144.215 ;
        RECT 103.405 144.045 103.575 144.215 ;
        RECT 103.865 144.045 104.035 144.215 ;
        RECT 104.325 144.045 104.495 144.215 ;
        RECT 104.785 144.045 104.955 144.215 ;
        RECT 105.245 144.045 105.415 144.215 ;
        RECT 105.705 144.045 105.875 144.215 ;
        RECT 106.165 144.045 106.335 144.215 ;
        RECT 106.625 144.045 106.795 144.215 ;
        RECT 107.085 144.045 107.255 144.215 ;
        RECT 107.545 144.045 107.715 144.215 ;
        RECT 108.005 144.045 108.175 144.215 ;
        RECT 108.465 144.045 108.635 144.215 ;
        RECT 108.925 144.045 109.095 144.215 ;
        RECT 109.385 144.045 109.555 144.215 ;
        RECT 109.845 144.045 110.015 144.215 ;
        RECT 110.305 144.045 110.475 144.215 ;
        RECT 110.765 144.045 110.935 144.215 ;
        RECT 111.225 144.045 111.395 144.215 ;
        RECT 111.685 144.045 111.855 144.215 ;
        RECT 112.145 144.045 112.315 144.215 ;
        RECT 112.605 144.045 112.775 144.215 ;
        RECT 113.065 144.045 113.235 144.215 ;
        RECT 113.525 144.045 113.695 144.215 ;
        RECT 113.985 144.045 114.155 144.215 ;
        RECT 114.445 144.045 114.615 144.215 ;
        RECT 114.905 144.045 115.075 144.215 ;
        RECT 115.365 144.045 115.535 144.215 ;
        RECT 115.825 144.045 115.995 144.215 ;
        RECT 116.285 144.045 116.455 144.215 ;
        RECT 116.745 144.045 116.915 144.215 ;
        RECT 117.205 144.045 117.375 144.215 ;
        RECT 117.665 144.045 117.835 144.215 ;
        RECT 118.125 144.045 118.295 144.215 ;
        RECT 118.585 144.045 118.755 144.215 ;
        RECT 119.045 144.045 119.215 144.215 ;
        RECT 119.505 144.045 119.675 144.215 ;
        RECT 119.965 144.045 120.135 144.215 ;
        RECT 120.425 144.045 120.595 144.215 ;
        RECT 120.885 144.045 121.055 144.215 ;
        RECT 121.345 144.045 121.515 144.215 ;
        RECT 121.805 144.045 121.975 144.215 ;
        RECT 122.265 144.045 122.435 144.215 ;
        RECT 122.725 144.045 122.895 144.215 ;
        RECT 123.185 144.045 123.355 144.215 ;
        RECT 123.645 144.045 123.815 144.215 ;
        RECT 124.105 144.045 124.275 144.215 ;
        RECT 124.565 144.045 124.735 144.215 ;
        RECT 125.025 144.045 125.195 144.215 ;
        RECT 125.485 144.045 125.655 144.215 ;
        RECT 125.945 144.045 126.115 144.215 ;
        RECT 126.405 144.045 126.575 144.215 ;
        RECT 126.865 144.045 127.035 144.215 ;
        RECT 127.325 144.045 127.495 144.215 ;
        RECT 127.785 144.045 127.955 144.215 ;
        RECT 128.245 144.045 128.415 144.215 ;
        RECT 128.705 144.045 128.875 144.215 ;
        RECT 129.165 144.045 129.335 144.215 ;
        RECT 129.625 144.045 129.795 144.215 ;
        RECT 130.085 144.045 130.255 144.215 ;
        RECT 130.545 144.045 130.715 144.215 ;
        RECT 131.005 144.045 131.175 144.215 ;
        RECT 131.465 144.045 131.635 144.215 ;
        RECT 131.925 144.045 132.095 144.215 ;
        RECT 132.385 144.045 132.555 144.215 ;
        RECT 132.845 144.045 133.015 144.215 ;
        RECT 133.305 144.045 133.475 144.215 ;
        RECT 133.765 144.045 133.935 144.215 ;
        RECT 134.225 144.045 134.395 144.215 ;
        RECT 134.685 144.045 134.855 144.215 ;
        RECT 135.145 144.045 135.315 144.215 ;
        RECT 135.605 144.045 135.775 144.215 ;
        RECT 136.065 144.045 136.235 144.215 ;
        RECT 136.525 144.045 136.695 144.215 ;
        RECT 136.985 144.045 137.155 144.215 ;
        RECT 137.445 144.045 137.615 144.215 ;
        RECT 137.905 144.045 138.075 144.215 ;
        RECT 138.365 144.045 138.535 144.215 ;
        RECT 138.825 144.045 138.995 144.215 ;
        RECT 139.285 144.045 139.455 144.215 ;
        RECT 139.745 144.045 139.915 144.215 ;
        RECT 140.205 144.045 140.375 144.215 ;
        RECT 140.665 144.045 140.835 144.215 ;
        RECT 141.125 144.045 141.295 144.215 ;
        RECT 141.585 144.045 141.755 144.215 ;
        RECT 142.045 144.045 142.215 144.215 ;
        RECT 142.505 144.045 142.675 144.215 ;
        RECT 142.965 144.045 143.135 144.215 ;
        RECT 143.425 144.045 143.595 144.215 ;
        RECT 143.885 144.045 144.055 144.215 ;
        RECT 144.345 144.045 144.515 144.215 ;
        RECT 144.805 144.045 144.975 144.215 ;
        RECT 145.265 144.045 145.435 144.215 ;
        RECT 145.725 144.045 145.895 144.215 ;
        RECT 146.185 144.045 146.355 144.215 ;
        RECT 146.645 144.045 146.815 144.215 ;
        RECT 147.105 144.045 147.275 144.215 ;
        RECT 147.565 144.045 147.735 144.215 ;
        RECT 148.025 144.045 148.195 144.215 ;
        RECT 148.485 144.045 148.655 144.215 ;
        RECT 148.945 144.045 149.115 144.215 ;
        RECT 149.405 144.045 149.575 144.215 ;
        RECT 149.865 144.045 150.035 144.215 ;
        RECT 40.870 143.195 41.040 143.365 ;
        RECT 40.385 142.855 40.555 143.025 ;
        RECT 39.465 142.515 39.635 142.685 ;
        RECT 38.545 141.835 38.715 142.005 ;
        RECT 41.265 142.855 41.435 143.025 ;
        RECT 41.720 142.175 41.890 142.345 ;
        RECT 42.970 143.195 43.140 143.365 ;
        RECT 42.455 142.855 42.625 143.025 ;
        RECT 44.540 143.195 44.710 143.365 ;
        RECT 44.975 142.855 45.145 143.025 ;
        RECT 47.285 143.535 47.455 143.705 ;
        RECT 50.965 142.515 51.135 142.685 ;
        RECT 51.425 142.175 51.595 142.345 ;
        RECT 53.265 142.175 53.435 142.345 ;
        RECT 50.045 141.835 50.215 142.005 ;
        RECT 56.025 142.515 56.195 142.685 ;
        RECT 55.105 141.835 55.275 142.005 ;
        RECT 60.165 142.515 60.335 142.685 ;
        RECT 59.245 141.835 59.415 142.005 ;
        RECT 64.305 142.515 64.475 142.685 ;
        RECT 63.385 141.835 63.555 142.005 ;
        RECT 78.565 143.195 78.735 143.365 ;
        RECT 76.725 142.515 76.895 142.685 ;
        RECT 77.645 142.515 77.815 142.685 ;
        RECT 75.805 141.835 75.975 142.005 ;
        RECT 79.485 142.515 79.655 142.685 ;
        RECT 80.405 141.835 80.575 142.005 ;
        RECT 82.245 142.515 82.415 142.685 ;
        RECT 83.625 142.515 83.795 142.685 ;
        RECT 81.325 141.835 81.495 142.005 ;
        RECT 84.545 141.835 84.715 142.005 ;
        RECT 88.685 142.515 88.855 142.685 ;
        RECT 91.905 143.535 92.075 143.705 ;
        RECT 91.445 142.855 91.615 143.025 ;
        RECT 92.825 142.515 92.995 142.685 ;
        RECT 93.745 142.515 93.915 142.685 ;
        RECT 89.145 141.835 89.315 142.005 ;
        RECT 94.205 142.515 94.375 142.685 ;
        RECT 95.125 141.835 95.295 142.005 ;
        RECT 97.425 142.515 97.595 142.685 ;
        RECT 101.105 142.515 101.275 142.685 ;
        RECT 96.505 141.835 96.675 142.005 ;
        RECT 102.025 141.835 102.195 142.005 ;
        RECT 105.705 142.515 105.875 142.685 ;
        RECT 104.785 141.835 104.955 142.005 ;
        RECT 114.445 143.535 114.615 143.705 ;
        RECT 113.985 142.515 114.155 142.685 ;
        RECT 115.365 142.515 115.535 142.685 ;
        RECT 116.745 142.515 116.915 142.685 ;
        RECT 116.285 141.835 116.455 142.005 ;
        RECT 117.665 141.835 117.835 142.005 ;
        RECT 120.885 142.515 121.055 142.685 ;
        RECT 121.805 141.835 121.975 142.005 ;
        RECT 124.565 142.515 124.735 142.685 ;
        RECT 127.325 143.535 127.495 143.705 ;
        RECT 126.865 142.855 127.035 143.025 ;
        RECT 128.245 142.515 128.415 142.685 ;
        RECT 125.485 141.835 125.655 142.005 ;
        RECT 129.165 142.175 129.335 142.345 ;
        RECT 130.085 142.175 130.255 142.345 ;
        RECT 133.305 142.515 133.475 142.685 ;
        RECT 130.545 141.835 130.715 142.005 ;
        RECT 134.225 141.835 134.395 142.005 ;
        RECT 137.445 142.515 137.615 142.685 ;
        RECT 143.405 143.535 143.575 143.705 ;
        RECT 140.205 142.855 140.375 143.025 ;
        RECT 138.365 141.835 138.535 142.005 ;
        RECT 143.885 142.855 144.055 143.025 ;
        RECT 144.345 142.515 144.515 142.685 ;
        RECT 146.185 142.515 146.355 142.685 ;
        RECT 147.105 141.835 147.275 142.005 ;
        RECT 36.245 141.325 36.415 141.495 ;
        RECT 36.705 141.325 36.875 141.495 ;
        RECT 37.165 141.325 37.335 141.495 ;
        RECT 37.625 141.325 37.795 141.495 ;
        RECT 38.085 141.325 38.255 141.495 ;
        RECT 38.545 141.325 38.715 141.495 ;
        RECT 39.005 141.325 39.175 141.495 ;
        RECT 39.465 141.325 39.635 141.495 ;
        RECT 39.925 141.325 40.095 141.495 ;
        RECT 40.385 141.325 40.555 141.495 ;
        RECT 40.845 141.325 41.015 141.495 ;
        RECT 41.305 141.325 41.475 141.495 ;
        RECT 41.765 141.325 41.935 141.495 ;
        RECT 42.225 141.325 42.395 141.495 ;
        RECT 42.685 141.325 42.855 141.495 ;
        RECT 43.145 141.325 43.315 141.495 ;
        RECT 43.605 141.325 43.775 141.495 ;
        RECT 44.065 141.325 44.235 141.495 ;
        RECT 44.525 141.325 44.695 141.495 ;
        RECT 44.985 141.325 45.155 141.495 ;
        RECT 45.445 141.325 45.615 141.495 ;
        RECT 45.905 141.325 46.075 141.495 ;
        RECT 46.365 141.325 46.535 141.495 ;
        RECT 46.825 141.325 46.995 141.495 ;
        RECT 47.285 141.325 47.455 141.495 ;
        RECT 47.745 141.325 47.915 141.495 ;
        RECT 48.205 141.325 48.375 141.495 ;
        RECT 48.665 141.325 48.835 141.495 ;
        RECT 49.125 141.325 49.295 141.495 ;
        RECT 49.585 141.325 49.755 141.495 ;
        RECT 50.045 141.325 50.215 141.495 ;
        RECT 50.505 141.325 50.675 141.495 ;
        RECT 50.965 141.325 51.135 141.495 ;
        RECT 51.425 141.325 51.595 141.495 ;
        RECT 51.885 141.325 52.055 141.495 ;
        RECT 52.345 141.325 52.515 141.495 ;
        RECT 52.805 141.325 52.975 141.495 ;
        RECT 53.265 141.325 53.435 141.495 ;
        RECT 53.725 141.325 53.895 141.495 ;
        RECT 54.185 141.325 54.355 141.495 ;
        RECT 54.645 141.325 54.815 141.495 ;
        RECT 55.105 141.325 55.275 141.495 ;
        RECT 55.565 141.325 55.735 141.495 ;
        RECT 56.025 141.325 56.195 141.495 ;
        RECT 56.485 141.325 56.655 141.495 ;
        RECT 56.945 141.325 57.115 141.495 ;
        RECT 57.405 141.325 57.575 141.495 ;
        RECT 57.865 141.325 58.035 141.495 ;
        RECT 58.325 141.325 58.495 141.495 ;
        RECT 58.785 141.325 58.955 141.495 ;
        RECT 59.245 141.325 59.415 141.495 ;
        RECT 59.705 141.325 59.875 141.495 ;
        RECT 60.165 141.325 60.335 141.495 ;
        RECT 60.625 141.325 60.795 141.495 ;
        RECT 61.085 141.325 61.255 141.495 ;
        RECT 61.545 141.325 61.715 141.495 ;
        RECT 62.005 141.325 62.175 141.495 ;
        RECT 62.465 141.325 62.635 141.495 ;
        RECT 62.925 141.325 63.095 141.495 ;
        RECT 63.385 141.325 63.555 141.495 ;
        RECT 63.845 141.325 64.015 141.495 ;
        RECT 64.305 141.325 64.475 141.495 ;
        RECT 64.765 141.325 64.935 141.495 ;
        RECT 65.225 141.325 65.395 141.495 ;
        RECT 65.685 141.325 65.855 141.495 ;
        RECT 66.145 141.325 66.315 141.495 ;
        RECT 66.605 141.325 66.775 141.495 ;
        RECT 67.065 141.325 67.235 141.495 ;
        RECT 67.525 141.325 67.695 141.495 ;
        RECT 67.985 141.325 68.155 141.495 ;
        RECT 68.445 141.325 68.615 141.495 ;
        RECT 68.905 141.325 69.075 141.495 ;
        RECT 69.365 141.325 69.535 141.495 ;
        RECT 69.825 141.325 69.995 141.495 ;
        RECT 70.285 141.325 70.455 141.495 ;
        RECT 70.745 141.325 70.915 141.495 ;
        RECT 71.205 141.325 71.375 141.495 ;
        RECT 71.665 141.325 71.835 141.495 ;
        RECT 72.125 141.325 72.295 141.495 ;
        RECT 72.585 141.325 72.755 141.495 ;
        RECT 73.045 141.325 73.215 141.495 ;
        RECT 73.505 141.325 73.675 141.495 ;
        RECT 73.965 141.325 74.135 141.495 ;
        RECT 74.425 141.325 74.595 141.495 ;
        RECT 74.885 141.325 75.055 141.495 ;
        RECT 75.345 141.325 75.515 141.495 ;
        RECT 75.805 141.325 75.975 141.495 ;
        RECT 76.265 141.325 76.435 141.495 ;
        RECT 76.725 141.325 76.895 141.495 ;
        RECT 77.185 141.325 77.355 141.495 ;
        RECT 77.645 141.325 77.815 141.495 ;
        RECT 78.105 141.325 78.275 141.495 ;
        RECT 78.565 141.325 78.735 141.495 ;
        RECT 79.025 141.325 79.195 141.495 ;
        RECT 79.485 141.325 79.655 141.495 ;
        RECT 79.945 141.325 80.115 141.495 ;
        RECT 80.405 141.325 80.575 141.495 ;
        RECT 80.865 141.325 81.035 141.495 ;
        RECT 81.325 141.325 81.495 141.495 ;
        RECT 81.785 141.325 81.955 141.495 ;
        RECT 82.245 141.325 82.415 141.495 ;
        RECT 82.705 141.325 82.875 141.495 ;
        RECT 83.165 141.325 83.335 141.495 ;
        RECT 83.625 141.325 83.795 141.495 ;
        RECT 84.085 141.325 84.255 141.495 ;
        RECT 84.545 141.325 84.715 141.495 ;
        RECT 85.005 141.325 85.175 141.495 ;
        RECT 85.465 141.325 85.635 141.495 ;
        RECT 85.925 141.325 86.095 141.495 ;
        RECT 86.385 141.325 86.555 141.495 ;
        RECT 86.845 141.325 87.015 141.495 ;
        RECT 87.305 141.325 87.475 141.495 ;
        RECT 87.765 141.325 87.935 141.495 ;
        RECT 88.225 141.325 88.395 141.495 ;
        RECT 88.685 141.325 88.855 141.495 ;
        RECT 89.145 141.325 89.315 141.495 ;
        RECT 89.605 141.325 89.775 141.495 ;
        RECT 90.065 141.325 90.235 141.495 ;
        RECT 90.525 141.325 90.695 141.495 ;
        RECT 90.985 141.325 91.155 141.495 ;
        RECT 91.445 141.325 91.615 141.495 ;
        RECT 91.905 141.325 92.075 141.495 ;
        RECT 92.365 141.325 92.535 141.495 ;
        RECT 92.825 141.325 92.995 141.495 ;
        RECT 93.285 141.325 93.455 141.495 ;
        RECT 93.745 141.325 93.915 141.495 ;
        RECT 94.205 141.325 94.375 141.495 ;
        RECT 94.665 141.325 94.835 141.495 ;
        RECT 95.125 141.325 95.295 141.495 ;
        RECT 95.585 141.325 95.755 141.495 ;
        RECT 96.045 141.325 96.215 141.495 ;
        RECT 96.505 141.325 96.675 141.495 ;
        RECT 96.965 141.325 97.135 141.495 ;
        RECT 97.425 141.325 97.595 141.495 ;
        RECT 97.885 141.325 98.055 141.495 ;
        RECT 98.345 141.325 98.515 141.495 ;
        RECT 98.805 141.325 98.975 141.495 ;
        RECT 99.265 141.325 99.435 141.495 ;
        RECT 99.725 141.325 99.895 141.495 ;
        RECT 100.185 141.325 100.355 141.495 ;
        RECT 100.645 141.325 100.815 141.495 ;
        RECT 101.105 141.325 101.275 141.495 ;
        RECT 101.565 141.325 101.735 141.495 ;
        RECT 102.025 141.325 102.195 141.495 ;
        RECT 102.485 141.325 102.655 141.495 ;
        RECT 102.945 141.325 103.115 141.495 ;
        RECT 103.405 141.325 103.575 141.495 ;
        RECT 103.865 141.325 104.035 141.495 ;
        RECT 104.325 141.325 104.495 141.495 ;
        RECT 104.785 141.325 104.955 141.495 ;
        RECT 105.245 141.325 105.415 141.495 ;
        RECT 105.705 141.325 105.875 141.495 ;
        RECT 106.165 141.325 106.335 141.495 ;
        RECT 106.625 141.325 106.795 141.495 ;
        RECT 107.085 141.325 107.255 141.495 ;
        RECT 107.545 141.325 107.715 141.495 ;
        RECT 108.005 141.325 108.175 141.495 ;
        RECT 108.465 141.325 108.635 141.495 ;
        RECT 108.925 141.325 109.095 141.495 ;
        RECT 109.385 141.325 109.555 141.495 ;
        RECT 109.845 141.325 110.015 141.495 ;
        RECT 110.305 141.325 110.475 141.495 ;
        RECT 110.765 141.325 110.935 141.495 ;
        RECT 111.225 141.325 111.395 141.495 ;
        RECT 111.685 141.325 111.855 141.495 ;
        RECT 112.145 141.325 112.315 141.495 ;
        RECT 112.605 141.325 112.775 141.495 ;
        RECT 113.065 141.325 113.235 141.495 ;
        RECT 113.525 141.325 113.695 141.495 ;
        RECT 113.985 141.325 114.155 141.495 ;
        RECT 114.445 141.325 114.615 141.495 ;
        RECT 114.905 141.325 115.075 141.495 ;
        RECT 115.365 141.325 115.535 141.495 ;
        RECT 115.825 141.325 115.995 141.495 ;
        RECT 116.285 141.325 116.455 141.495 ;
        RECT 116.745 141.325 116.915 141.495 ;
        RECT 117.205 141.325 117.375 141.495 ;
        RECT 117.665 141.325 117.835 141.495 ;
        RECT 118.125 141.325 118.295 141.495 ;
        RECT 118.585 141.325 118.755 141.495 ;
        RECT 119.045 141.325 119.215 141.495 ;
        RECT 119.505 141.325 119.675 141.495 ;
        RECT 119.965 141.325 120.135 141.495 ;
        RECT 120.425 141.325 120.595 141.495 ;
        RECT 120.885 141.325 121.055 141.495 ;
        RECT 121.345 141.325 121.515 141.495 ;
        RECT 121.805 141.325 121.975 141.495 ;
        RECT 122.265 141.325 122.435 141.495 ;
        RECT 122.725 141.325 122.895 141.495 ;
        RECT 123.185 141.325 123.355 141.495 ;
        RECT 123.645 141.325 123.815 141.495 ;
        RECT 124.105 141.325 124.275 141.495 ;
        RECT 124.565 141.325 124.735 141.495 ;
        RECT 125.025 141.325 125.195 141.495 ;
        RECT 125.485 141.325 125.655 141.495 ;
        RECT 125.945 141.325 126.115 141.495 ;
        RECT 126.405 141.325 126.575 141.495 ;
        RECT 126.865 141.325 127.035 141.495 ;
        RECT 127.325 141.325 127.495 141.495 ;
        RECT 127.785 141.325 127.955 141.495 ;
        RECT 128.245 141.325 128.415 141.495 ;
        RECT 128.705 141.325 128.875 141.495 ;
        RECT 129.165 141.325 129.335 141.495 ;
        RECT 129.625 141.325 129.795 141.495 ;
        RECT 130.085 141.325 130.255 141.495 ;
        RECT 130.545 141.325 130.715 141.495 ;
        RECT 131.005 141.325 131.175 141.495 ;
        RECT 131.465 141.325 131.635 141.495 ;
        RECT 131.925 141.325 132.095 141.495 ;
        RECT 132.385 141.325 132.555 141.495 ;
        RECT 132.845 141.325 133.015 141.495 ;
        RECT 133.305 141.325 133.475 141.495 ;
        RECT 133.765 141.325 133.935 141.495 ;
        RECT 134.225 141.325 134.395 141.495 ;
        RECT 134.685 141.325 134.855 141.495 ;
        RECT 135.145 141.325 135.315 141.495 ;
        RECT 135.605 141.325 135.775 141.495 ;
        RECT 136.065 141.325 136.235 141.495 ;
        RECT 136.525 141.325 136.695 141.495 ;
        RECT 136.985 141.325 137.155 141.495 ;
        RECT 137.445 141.325 137.615 141.495 ;
        RECT 137.905 141.325 138.075 141.495 ;
        RECT 138.365 141.325 138.535 141.495 ;
        RECT 138.825 141.325 138.995 141.495 ;
        RECT 139.285 141.325 139.455 141.495 ;
        RECT 139.745 141.325 139.915 141.495 ;
        RECT 140.205 141.325 140.375 141.495 ;
        RECT 140.665 141.325 140.835 141.495 ;
        RECT 141.125 141.325 141.295 141.495 ;
        RECT 141.585 141.325 141.755 141.495 ;
        RECT 142.045 141.325 142.215 141.495 ;
        RECT 142.505 141.325 142.675 141.495 ;
        RECT 142.965 141.325 143.135 141.495 ;
        RECT 143.425 141.325 143.595 141.495 ;
        RECT 143.885 141.325 144.055 141.495 ;
        RECT 144.345 141.325 144.515 141.495 ;
        RECT 144.805 141.325 144.975 141.495 ;
        RECT 145.265 141.325 145.435 141.495 ;
        RECT 145.725 141.325 145.895 141.495 ;
        RECT 146.185 141.325 146.355 141.495 ;
        RECT 146.645 141.325 146.815 141.495 ;
        RECT 147.105 141.325 147.275 141.495 ;
        RECT 147.565 141.325 147.735 141.495 ;
        RECT 148.025 141.325 148.195 141.495 ;
        RECT 148.485 141.325 148.655 141.495 ;
        RECT 148.945 141.325 149.115 141.495 ;
        RECT 149.405 141.325 149.575 141.495 ;
        RECT 149.865 141.325 150.035 141.495 ;
        RECT 34.840 125.925 35.370 127.910 ;
        RECT 38.840 125.925 39.370 127.910 ;
        RECT 42.840 125.925 43.370 127.910 ;
        RECT 46.840 125.925 47.370 127.910 ;
        RECT 50.840 125.925 51.370 127.910 ;
        RECT 54.840 125.925 55.370 127.910 ;
        RECT 58.840 125.925 59.370 127.910 ;
        RECT 62.840 125.925 63.370 127.910 ;
        RECT 75.840 125.925 76.370 127.910 ;
        RECT 79.840 125.925 80.370 127.910 ;
        RECT 83.840 125.925 84.370 127.910 ;
        RECT 87.840 125.925 88.370 127.910 ;
        RECT 91.840 125.925 92.370 127.910 ;
        RECT 95.840 125.925 96.370 127.910 ;
        RECT 99.840 125.925 100.370 127.910 ;
        RECT 103.840 125.925 104.370 127.910 ;
        RECT 116.840 125.925 117.370 127.910 ;
        RECT 120.840 125.925 121.370 127.910 ;
        RECT 124.840 125.925 125.370 127.910 ;
        RECT 128.840 125.925 129.370 127.910 ;
        RECT 132.840 125.925 133.370 127.910 ;
        RECT 136.840 125.925 137.370 127.910 ;
        RECT 140.840 125.925 141.370 127.910 ;
        RECT 144.840 125.925 145.370 127.910 ;
        RECT 34.030 104.170 34.370 104.970 ;
        RECT 35.830 104.170 36.170 104.970 ;
        RECT 38.030 104.170 38.370 104.970 ;
        RECT 39.830 104.170 40.170 104.970 ;
        RECT 42.030 104.170 42.370 104.970 ;
        RECT 43.830 104.170 44.170 104.970 ;
        RECT 46.030 104.170 46.370 104.970 ;
        RECT 47.830 104.170 48.170 104.970 ;
        RECT 50.030 104.170 50.370 104.970 ;
        RECT 51.830 104.170 52.170 104.970 ;
        RECT 54.030 104.170 54.370 104.970 ;
        RECT 55.830 104.170 56.170 104.970 ;
        RECT 58.030 104.170 58.370 104.970 ;
        RECT 59.830 104.170 60.170 104.970 ;
        RECT 62.030 104.170 62.370 104.970 ;
        RECT 63.830 104.170 64.170 104.970 ;
        RECT 75.030 104.170 75.370 104.970 ;
        RECT 76.830 104.170 77.170 104.970 ;
        RECT 79.030 104.170 79.370 104.970 ;
        RECT 80.830 104.170 81.170 104.970 ;
        RECT 83.030 104.170 83.370 104.970 ;
        RECT 84.830 104.170 85.170 104.970 ;
        RECT 87.030 104.170 87.370 104.970 ;
        RECT 88.830 104.170 89.170 104.970 ;
        RECT 91.030 104.170 91.370 104.970 ;
        RECT 92.830 104.170 93.170 104.970 ;
        RECT 95.030 104.170 95.370 104.970 ;
        RECT 96.830 104.170 97.170 104.970 ;
        RECT 99.030 104.170 99.370 104.970 ;
        RECT 100.830 104.170 101.170 104.970 ;
        RECT 103.030 104.170 103.370 104.970 ;
        RECT 104.830 104.170 105.170 104.970 ;
        RECT 116.030 104.170 116.370 104.970 ;
        RECT 117.830 104.170 118.170 104.970 ;
        RECT 120.030 104.170 120.370 104.970 ;
        RECT 121.830 104.170 122.170 104.970 ;
        RECT 124.030 104.170 124.370 104.970 ;
        RECT 125.830 104.170 126.170 104.970 ;
        RECT 128.030 104.170 128.370 104.970 ;
        RECT 129.830 104.170 130.170 104.970 ;
        RECT 132.030 104.170 132.370 104.970 ;
        RECT 133.830 104.170 134.170 104.970 ;
        RECT 136.030 104.170 136.370 104.970 ;
        RECT 137.830 104.170 138.170 104.970 ;
        RECT 140.030 104.170 140.370 104.970 ;
        RECT 141.830 104.170 142.170 104.970 ;
        RECT 144.030 104.170 144.370 104.970 ;
        RECT 145.830 104.170 146.170 104.970 ;
        RECT 34.840 84.030 35.370 86.015 ;
        RECT 38.840 84.030 39.370 86.015 ;
        RECT 42.840 84.030 43.370 86.015 ;
        RECT 46.840 84.030 47.370 86.015 ;
        RECT 50.840 84.030 51.370 86.015 ;
        RECT 54.840 84.030 55.370 86.015 ;
        RECT 58.840 84.030 59.370 86.015 ;
        RECT 62.840 84.030 63.370 86.015 ;
        RECT 75.840 84.030 76.370 86.015 ;
        RECT 79.840 84.030 80.370 86.015 ;
        RECT 83.840 84.030 84.370 86.015 ;
        RECT 87.840 84.030 88.370 86.015 ;
        RECT 91.840 84.030 92.370 86.015 ;
        RECT 95.840 84.030 96.370 86.015 ;
        RECT 99.840 84.030 100.370 86.015 ;
        RECT 103.840 84.030 104.370 86.015 ;
        RECT 116.840 84.030 117.370 86.015 ;
        RECT 120.840 84.030 121.370 86.015 ;
        RECT 124.840 84.030 125.370 86.015 ;
        RECT 128.840 84.030 129.370 86.015 ;
        RECT 132.840 84.030 133.370 86.015 ;
        RECT 136.840 84.030 137.370 86.015 ;
        RECT 140.840 84.030 141.370 86.015 ;
        RECT 144.840 84.030 145.370 86.015 ;
        RECT 34.840 77.925 35.370 79.910 ;
        RECT 34.840 56.380 35.370 58.365 ;
        RECT 38.840 77.925 39.370 79.910 ;
        RECT 38.840 56.380 39.370 58.365 ;
        RECT 42.840 77.925 43.370 79.910 ;
        RECT 42.840 56.380 43.370 58.365 ;
        RECT 46.840 77.925 47.370 79.910 ;
        RECT 46.840 56.380 47.370 58.365 ;
        RECT 50.840 77.925 51.370 79.910 ;
        RECT 50.840 56.380 51.370 58.365 ;
        RECT 54.840 77.925 55.370 79.910 ;
        RECT 54.840 56.380 55.370 58.365 ;
        RECT 58.840 77.925 59.370 79.910 ;
        RECT 58.840 56.380 59.370 58.365 ;
        RECT 62.840 77.925 63.370 79.910 ;
        RECT 62.840 56.380 63.370 58.365 ;
        RECT 75.840 77.925 76.370 79.910 ;
        RECT 75.840 56.380 76.370 58.365 ;
        RECT 79.840 77.925 80.370 79.910 ;
        RECT 79.840 56.380 80.370 58.365 ;
        RECT 83.840 77.925 84.370 79.910 ;
        RECT 83.840 56.380 84.370 58.365 ;
        RECT 87.840 77.925 88.370 79.910 ;
        RECT 87.840 56.380 88.370 58.365 ;
        RECT 91.840 77.925 92.370 79.910 ;
        RECT 91.840 56.380 92.370 58.365 ;
        RECT 95.840 77.925 96.370 79.910 ;
        RECT 95.840 56.380 96.370 58.365 ;
        RECT 99.840 77.925 100.370 79.910 ;
        RECT 99.840 56.380 100.370 58.365 ;
        RECT 103.840 77.925 104.370 79.910 ;
        RECT 103.840 56.380 104.370 58.365 ;
        RECT 116.840 77.925 117.370 79.910 ;
        RECT 116.840 56.380 117.370 58.365 ;
        RECT 120.840 77.925 121.370 79.910 ;
        RECT 120.840 56.380 121.370 58.365 ;
        RECT 124.840 77.925 125.370 79.910 ;
        RECT 124.840 56.380 125.370 58.365 ;
        RECT 128.840 77.925 129.370 79.910 ;
        RECT 128.840 56.380 129.370 58.365 ;
        RECT 132.840 77.925 133.370 79.910 ;
        RECT 132.840 56.380 133.370 58.365 ;
        RECT 136.840 77.925 137.370 79.910 ;
        RECT 136.840 56.380 137.370 58.365 ;
        RECT 140.840 77.925 141.370 79.910 ;
        RECT 140.840 56.380 141.370 58.365 ;
        RECT 144.840 77.925 145.370 79.910 ;
        RECT 144.840 56.380 145.370 58.365 ;
        RECT 27.655 20.130 27.825 20.300 ;
        RECT 26.800 15.765 27.100 16.465 ;
        RECT 27.435 11.955 27.605 19.835 ;
        RECT 27.875 11.955 28.045 19.835 ;
        RECT 27.655 11.490 27.825 11.660 ;
        RECT 30.470 18.105 30.640 18.275 ;
        RECT 30.250 13.975 30.420 17.855 ;
        RECT 30.690 13.975 30.860 17.855 ;
        RECT 31.200 16.865 31.500 17.665 ;
        RECT 30.470 13.555 30.640 13.725 ;
      LAYER met1 ;
        RECT 114.370 215.770 114.690 215.830 ;
        RECT 66.160 215.630 114.690 215.770 ;
        RECT 66.160 215.490 66.300 215.630 ;
        RECT 114.370 215.570 114.690 215.630 ;
        RECT 119.430 215.770 119.750 215.830 ;
        RECT 119.430 215.630 144.960 215.770 ;
        RECT 119.430 215.570 119.750 215.630 ;
        RECT 144.820 215.490 144.960 215.630 ;
        RECT 66.070 215.230 66.390 215.490 ;
        RECT 66.990 215.430 67.310 215.490 ;
        RECT 105.630 215.430 105.950 215.490 ;
        RECT 66.990 215.290 105.950 215.430 ;
        RECT 66.990 215.230 67.310 215.290 ;
        RECT 105.630 215.230 105.950 215.290 ;
        RECT 107.010 215.430 107.330 215.490 ;
        RECT 123.570 215.430 123.890 215.490 ;
        RECT 107.010 215.290 123.890 215.430 ;
        RECT 107.010 215.230 107.330 215.290 ;
        RECT 123.570 215.230 123.890 215.290 ;
        RECT 144.730 215.230 145.050 215.490 ;
        RECT 36.100 214.610 150.180 215.090 ;
        RECT 56.410 214.210 56.730 214.470 ;
        RECT 59.170 214.210 59.490 214.470 ;
        RECT 64.230 214.210 64.550 214.470 ;
        RECT 66.530 214.210 66.850 214.470 ;
        RECT 69.750 214.410 70.070 214.470 ;
        RECT 71.145 214.410 71.435 214.455 ;
        RECT 69.750 214.270 71.435 214.410 ;
        RECT 69.750 214.210 70.070 214.270 ;
        RECT 71.145 214.225 71.435 214.270 ;
        RECT 73.890 214.410 74.210 214.470 ;
        RECT 75.745 214.410 76.035 214.455 ;
        RECT 73.890 214.270 76.035 214.410 ;
        RECT 73.890 214.210 74.210 214.270 ;
        RECT 75.745 214.225 76.035 214.270 ;
        RECT 78.950 214.210 79.270 214.470 ;
        RECT 81.250 214.210 81.570 214.470 ;
        RECT 84.930 214.410 85.250 214.470 ;
        RECT 85.865 214.410 86.155 214.455 ;
        RECT 84.930 214.270 86.155 214.410 ;
        RECT 84.930 214.210 85.250 214.270 ;
        RECT 85.865 214.225 86.155 214.270 ;
        RECT 88.610 214.210 88.930 214.470 ;
        RECT 105.630 214.410 105.950 214.470 ;
        RECT 126.330 214.410 126.650 214.470 ;
        RECT 140.605 214.410 140.895 214.455 ;
        RECT 105.630 214.270 114.600 214.410 ;
        RECT 105.630 214.210 105.950 214.270 ;
        RECT 113.925 214.070 114.215 214.115 ;
        RECT 68.920 213.930 114.215 214.070 ;
        RECT 32.470 149.430 33.130 213.760 ;
        RECT 44.450 213.390 44.770 213.450 ;
        RECT 44.925 213.390 45.215 213.435 ;
        RECT 44.450 213.250 45.215 213.390 ;
        RECT 44.450 213.190 44.770 213.250 ;
        RECT 44.925 213.205 45.215 213.250 ;
        RECT 57.345 213.205 57.635 213.435 ;
        RECT 57.790 213.390 58.110 213.450 ;
        RECT 63.325 213.390 63.615 213.435 ;
        RECT 57.790 213.250 63.615 213.390 ;
        RECT 57.420 213.050 57.560 213.205 ;
        RECT 57.790 213.190 58.110 213.250 ;
        RECT 63.325 213.205 63.615 213.250 ;
        RECT 60.565 213.050 60.855 213.095 ;
        RECT 66.990 213.050 67.310 213.110 ;
        RECT 57.420 212.910 59.400 213.050 ;
        RECT 59.260 212.770 59.400 212.910 ;
        RECT 60.565 212.910 67.310 213.050 ;
        RECT 60.565 212.865 60.855 212.910 ;
        RECT 66.990 212.850 67.310 212.910 ;
        RECT 67.910 212.850 68.230 213.110 ;
        RECT 68.920 212.770 69.060 213.930 ;
        RECT 113.925 213.885 114.215 213.930 ;
        RECT 71.590 213.730 71.910 213.790 ;
        RECT 114.460 213.730 114.600 214.270 ;
        RECT 126.330 214.270 150.020 214.410 ;
        RECT 126.330 214.210 126.650 214.270 ;
        RECT 140.605 214.225 140.895 214.270 ;
        RECT 118.510 214.070 118.830 214.130 ;
        RECT 116.760 213.930 118.830 214.070 ;
        RECT 116.760 213.775 116.900 213.930 ;
        RECT 118.510 213.870 118.830 213.930 ;
        RECT 119.890 214.070 120.210 214.130 ;
        RECT 139.685 214.070 139.975 214.115 ;
        RECT 119.890 213.930 139.975 214.070 ;
        RECT 119.890 213.870 120.210 213.930 ;
        RECT 139.685 213.885 139.975 213.930 ;
        RECT 144.285 213.885 144.575 214.115 ;
        RECT 144.730 214.070 145.050 214.130 ;
        RECT 147.505 214.070 147.795 214.115 ;
        RECT 144.730 213.930 147.795 214.070 ;
        RECT 116.225 213.730 116.515 213.775 ;
        RECT 71.590 213.590 113.680 213.730 ;
        RECT 114.460 213.590 116.515 213.730 ;
        RECT 71.590 213.530 71.910 213.590 ;
        RECT 72.065 213.205 72.355 213.435 ;
        RECT 72.140 213.050 72.280 213.205 ;
        RECT 72.510 213.190 72.830 213.450 ;
        RECT 73.445 213.390 73.735 213.435 ;
        RECT 76.190 213.390 76.510 213.450 ;
        RECT 73.445 213.250 76.510 213.390 ;
        RECT 73.445 213.205 73.735 213.250 ;
        RECT 76.190 213.190 76.510 213.250 ;
        RECT 78.030 213.190 78.350 213.450 ;
        RECT 84.010 213.390 84.330 213.450 ;
        RECT 86.785 213.390 87.075 213.435 ;
        RECT 84.010 213.250 87.075 213.390 ;
        RECT 84.010 213.190 84.330 213.250 ;
        RECT 86.785 213.205 87.075 213.250 ;
        RECT 99.205 213.205 99.495 213.435 ;
        RECT 99.650 213.390 99.970 213.450 ;
        RECT 101.045 213.390 101.335 213.435 ;
        RECT 99.650 213.250 101.335 213.390 ;
        RECT 76.650 213.050 76.970 213.110 ;
        RECT 72.140 212.910 76.970 213.050 ;
        RECT 76.650 212.850 76.970 212.910 ;
        RECT 77.125 213.050 77.415 213.095 ;
        RECT 80.790 213.050 81.110 213.110 ;
        RECT 77.125 212.910 81.110 213.050 ;
        RECT 77.125 212.865 77.415 212.910 ;
        RECT 80.790 212.850 81.110 212.910 ;
        RECT 81.710 213.050 82.030 213.110 ;
        RECT 82.645 213.050 82.935 213.095 ;
        RECT 81.710 212.910 82.935 213.050 ;
        RECT 81.710 212.850 82.030 212.910 ;
        RECT 82.645 212.865 82.935 212.910 ;
        RECT 90.005 213.050 90.295 213.095 ;
        RECT 93.210 213.050 93.530 213.110 ;
        RECT 90.005 212.910 93.530 213.050 ;
        RECT 99.280 213.050 99.420 213.205 ;
        RECT 99.650 213.190 99.970 213.250 ;
        RECT 101.045 213.205 101.335 213.250 ;
        RECT 102.425 213.205 102.715 213.435 ;
        RECT 113.540 213.390 113.680 213.590 ;
        RECT 116.225 213.545 116.515 213.590 ;
        RECT 116.685 213.545 116.975 213.775 ;
        RECT 117.130 213.730 117.450 213.790 ;
        RECT 144.360 213.730 144.500 213.885 ;
        RECT 144.730 213.870 145.050 213.930 ;
        RECT 147.505 213.885 147.795 213.930 ;
        RECT 117.130 213.590 144.500 213.730 ;
        RECT 117.130 213.530 117.450 213.590 ;
        RECT 117.590 213.390 117.910 213.450 ;
        RECT 113.540 213.250 117.910 213.390 ;
        RECT 102.500 213.050 102.640 213.205 ;
        RECT 117.590 213.190 117.910 213.250 ;
        RECT 121.730 213.390 122.050 213.450 ;
        RECT 122.205 213.390 122.495 213.435 ;
        RECT 121.730 213.250 122.495 213.390 ;
        RECT 121.730 213.190 122.050 213.250 ;
        RECT 122.205 213.205 122.495 213.250 ;
        RECT 125.410 213.390 125.730 213.450 ;
        RECT 126.805 213.390 127.095 213.435 ;
        RECT 125.410 213.250 127.095 213.390 ;
        RECT 125.410 213.190 125.730 213.250 ;
        RECT 126.805 213.205 127.095 213.250 ;
        RECT 129.090 213.390 129.410 213.450 ;
        RECT 130.485 213.390 130.775 213.435 ;
        RECT 129.090 213.250 130.775 213.390 ;
        RECT 129.090 213.190 129.410 213.250 ;
        RECT 130.485 213.205 130.775 213.250 ;
        RECT 133.690 213.190 134.010 213.450 ;
        RECT 134.150 213.390 134.470 213.450 ;
        RECT 135.085 213.390 135.375 213.435 ;
        RECT 134.150 213.250 135.375 213.390 ;
        RECT 134.150 213.190 134.470 213.250 ;
        RECT 135.085 213.205 135.375 213.250 ;
        RECT 136.450 213.390 136.770 213.450 ;
        RECT 137.845 213.390 138.135 213.435 ;
        RECT 136.450 213.250 138.135 213.390 ;
        RECT 136.450 213.190 136.770 213.250 ;
        RECT 137.845 213.205 138.135 213.250 ;
        RECT 140.130 213.190 140.450 213.450 ;
        RECT 140.590 213.390 140.910 213.450 ;
        RECT 141.985 213.390 142.275 213.435 ;
        RECT 140.590 213.250 142.275 213.390 ;
        RECT 140.590 213.190 140.910 213.250 ;
        RECT 141.985 213.205 142.275 213.250 ;
        RECT 143.365 213.205 143.655 213.435 ;
        RECT 143.810 213.390 144.130 213.450 ;
        RECT 145.205 213.390 145.495 213.435 ;
        RECT 143.810 213.250 145.495 213.390 ;
        RECT 99.280 212.910 102.640 213.050 ;
        RECT 90.005 212.865 90.295 212.910 ;
        RECT 93.210 212.850 93.530 212.910 ;
        RECT 102.500 212.770 102.640 212.910 ;
        RECT 115.765 213.050 116.055 213.095 ;
        RECT 124.490 213.050 124.810 213.110 ;
        RECT 140.220 213.050 140.360 213.190 ;
        RECT 143.440 213.050 143.580 213.205 ;
        RECT 143.810 213.190 144.130 213.250 ;
        RECT 145.205 213.205 145.495 213.250 ;
        RECT 147.490 213.390 147.810 213.450 ;
        RECT 148.425 213.390 148.715 213.435 ;
        RECT 147.490 213.250 148.715 213.390 ;
        RECT 147.490 213.190 147.810 213.250 ;
        RECT 148.425 213.205 148.715 213.250 ;
        RECT 115.765 212.910 137.140 213.050 ;
        RECT 140.220 212.910 143.580 213.050 ;
        RECT 115.765 212.865 116.055 212.910 ;
        RECT 124.490 212.850 124.810 212.910 ;
        RECT 45.830 212.710 46.150 212.770 ;
        RECT 48.145 212.710 48.435 212.755 ;
        RECT 45.830 212.570 48.435 212.710 ;
        RECT 45.830 212.510 46.150 212.570 ;
        RECT 48.145 212.525 48.435 212.570 ;
        RECT 59.170 212.510 59.490 212.770 ;
        RECT 68.830 212.510 69.150 212.770 ;
        RECT 72.970 212.510 73.290 212.770 ;
        RECT 92.750 212.710 93.070 212.770 ;
        RECT 98.745 212.710 99.035 212.755 ;
        RECT 92.750 212.570 99.035 212.710 ;
        RECT 92.750 212.510 93.070 212.570 ;
        RECT 98.745 212.525 99.035 212.570 ;
        RECT 102.410 212.510 102.730 212.770 ;
        RECT 123.125 212.710 123.415 212.755 ;
        RECT 125.870 212.710 126.190 212.770 ;
        RECT 123.125 212.570 126.190 212.710 ;
        RECT 123.125 212.525 123.415 212.570 ;
        RECT 125.870 212.510 126.190 212.570 ;
        RECT 127.710 212.510 128.030 212.770 ;
        RECT 129.550 212.510 129.870 212.770 ;
        RECT 132.785 212.710 133.075 212.755 ;
        RECT 133.230 212.710 133.550 212.770 ;
        RECT 132.785 212.570 133.550 212.710 ;
        RECT 132.785 212.525 133.075 212.570 ;
        RECT 133.230 212.510 133.550 212.570 ;
        RECT 134.150 212.510 134.470 212.770 ;
        RECT 137.000 212.755 137.140 212.910 ;
        RECT 136.925 212.525 137.215 212.755 ;
        RECT 141.050 212.710 141.370 212.770 ;
        RECT 142.445 212.710 142.735 212.755 ;
        RECT 141.050 212.570 142.735 212.710 ;
        RECT 149.880 212.710 150.020 214.270 ;
        RECT 149.880 212.570 150.480 212.710 ;
        RECT 141.050 212.510 141.370 212.570 ;
        RECT 142.445 212.525 142.735 212.570 ;
        RECT 36.100 211.890 150.180 212.370 ;
        RECT 44.450 211.490 44.770 211.750 ;
        RECT 45.370 211.690 45.690 211.750 ;
        RECT 57.790 211.690 58.110 211.750 ;
        RECT 45.370 211.550 58.110 211.690 ;
        RECT 45.370 211.490 45.690 211.550 ;
        RECT 57.790 211.490 58.110 211.550 ;
        RECT 61.485 211.505 61.775 211.735 ;
        RECT 64.245 211.690 64.535 211.735 ;
        RECT 66.530 211.690 66.850 211.750 ;
        RECT 64.245 211.550 66.850 211.690 ;
        RECT 64.245 211.505 64.535 211.550 ;
        RECT 61.560 211.350 61.700 211.505 ;
        RECT 66.530 211.490 66.850 211.550 ;
        RECT 67.005 211.690 67.295 211.735 ;
        RECT 71.590 211.690 71.910 211.750 ;
        RECT 67.005 211.550 71.910 211.690 ;
        RECT 67.005 211.505 67.295 211.550 ;
        RECT 71.590 211.490 71.910 211.550 ;
        RECT 72.970 211.490 73.290 211.750 ;
        RECT 78.030 211.490 78.350 211.750 ;
        RECT 84.485 211.690 84.775 211.735 ;
        RECT 85.405 211.690 85.695 211.735 ;
        RECT 86.770 211.690 87.090 211.750 ;
        RECT 88.625 211.690 88.915 211.735 ;
        RECT 107.010 211.690 107.330 211.750 ;
        RECT 84.485 211.550 85.160 211.690 ;
        RECT 84.485 211.505 84.775 211.550 ;
        RECT 63.770 211.350 64.090 211.410 ;
        RECT 46.380 211.210 54.800 211.350 ;
        RECT 61.560 211.210 64.090 211.350 ;
        RECT 73.060 211.350 73.200 211.490 ;
        RECT 73.060 211.210 74.120 211.350 ;
        RECT 38.900 211.010 39.190 211.055 ;
        RECT 38.900 210.870 42.840 211.010 ;
        RECT 38.900 210.825 39.190 210.870 ;
        RECT 37.565 210.485 37.855 210.715 ;
        RECT 38.445 210.670 38.735 210.715 ;
        RECT 39.635 210.670 39.925 210.715 ;
        RECT 42.155 210.670 42.445 210.715 ;
        RECT 38.445 210.530 42.445 210.670 ;
        RECT 38.445 210.485 38.735 210.530 ;
        RECT 39.635 210.485 39.925 210.530 ;
        RECT 42.155 210.485 42.445 210.530 ;
        RECT 37.640 209.990 37.780 210.485 ;
        RECT 38.050 210.330 38.340 210.375 ;
        RECT 40.150 210.330 40.440 210.375 ;
        RECT 41.720 210.330 42.010 210.375 ;
        RECT 38.050 210.190 42.010 210.330 ;
        RECT 38.050 210.145 38.340 210.190 ;
        RECT 40.150 210.145 40.440 210.190 ;
        RECT 41.720 210.145 42.010 210.190 ;
        RECT 42.700 210.050 42.840 210.870 ;
        RECT 45.830 210.810 46.150 211.070 ;
        RECT 46.380 211.055 46.520 211.210 ;
        RECT 47.670 211.055 47.990 211.070 ;
        RECT 54.660 211.055 54.800 211.210 ;
        RECT 63.770 211.150 64.090 211.210 ;
        RECT 46.305 210.825 46.595 211.055 ;
        RECT 47.640 210.825 47.990 211.055 ;
        RECT 54.585 211.010 54.875 211.055 ;
        RECT 55.030 211.010 55.350 211.070 ;
        RECT 54.585 210.870 55.350 211.010 ;
        RECT 54.585 210.825 54.875 210.870 ;
        RECT 47.670 210.810 47.990 210.825 ;
        RECT 55.030 210.810 55.350 210.870 ;
        RECT 55.920 211.010 56.210 211.055 ;
        RECT 55.920 210.870 59.860 211.010 ;
        RECT 55.920 210.825 56.210 210.870 ;
        RECT 47.185 210.670 47.475 210.715 ;
        RECT 48.375 210.670 48.665 210.715 ;
        RECT 50.895 210.670 51.185 210.715 ;
        RECT 47.185 210.530 51.185 210.670 ;
        RECT 47.185 210.485 47.475 210.530 ;
        RECT 48.375 210.485 48.665 210.530 ;
        RECT 50.895 210.485 51.185 210.530 ;
        RECT 55.465 210.670 55.755 210.715 ;
        RECT 56.655 210.670 56.945 210.715 ;
        RECT 59.175 210.670 59.465 210.715 ;
        RECT 55.465 210.530 59.465 210.670 ;
        RECT 55.465 210.485 55.755 210.530 ;
        RECT 56.655 210.485 56.945 210.530 ;
        RECT 59.175 210.485 59.465 210.530 ;
        RECT 46.790 210.330 47.080 210.375 ;
        RECT 48.890 210.330 49.180 210.375 ;
        RECT 50.460 210.330 50.750 210.375 ;
        RECT 46.790 210.190 50.750 210.330 ;
        RECT 46.790 210.145 47.080 210.190 ;
        RECT 48.890 210.145 49.180 210.190 ;
        RECT 50.460 210.145 50.750 210.190 ;
        RECT 55.070 210.330 55.360 210.375 ;
        RECT 57.170 210.330 57.460 210.375 ;
        RECT 58.740 210.330 59.030 210.375 ;
        RECT 55.070 210.190 59.030 210.330 ;
        RECT 59.720 210.330 59.860 210.870 ;
        RECT 60.090 210.810 60.410 211.070 ;
        RECT 66.070 210.810 66.390 211.070 ;
        RECT 66.545 210.825 66.835 211.055 ;
        RECT 66.990 211.010 67.310 211.070 ;
        RECT 67.465 211.010 67.755 211.055 ;
        RECT 66.990 210.870 67.755 211.010 ;
        RECT 60.180 210.670 60.320 210.810 ;
        RECT 66.620 210.670 66.760 210.825 ;
        RECT 66.990 210.810 67.310 210.870 ;
        RECT 67.465 210.825 67.755 210.870 ;
        RECT 68.830 210.810 69.150 211.070 ;
        RECT 71.145 211.010 71.435 211.055 ;
        RECT 73.430 211.010 73.750 211.070 ;
        RECT 71.145 210.870 73.750 211.010 ;
        RECT 71.145 210.825 71.435 210.870 ;
        RECT 73.430 210.810 73.750 210.870 ;
        RECT 73.980 210.715 74.120 211.210 ;
        RECT 74.365 211.010 74.655 211.055 ;
        RECT 77.110 211.010 77.430 211.070 ;
        RECT 74.365 210.870 77.430 211.010 ;
        RECT 74.365 210.825 74.655 210.870 ;
        RECT 77.110 210.810 77.430 210.870 ;
        RECT 60.180 210.530 66.760 210.670 ;
        RECT 71.605 210.485 71.895 210.715 ;
        RECT 73.905 210.485 74.195 210.715 ;
        RECT 78.120 210.670 78.260 211.490 ;
        RECT 85.020 211.350 85.160 211.550 ;
        RECT 85.405 211.550 88.915 211.690 ;
        RECT 85.405 211.505 85.695 211.550 ;
        RECT 86.770 211.490 87.090 211.550 ;
        RECT 88.625 211.505 88.915 211.550 ;
        RECT 93.760 211.550 107.330 211.690 ;
        RECT 88.165 211.350 88.455 211.395 ;
        RECT 85.020 211.210 88.455 211.350 ;
        RECT 80.805 211.010 81.095 211.055 ;
        RECT 79.040 210.870 81.095 211.010 ;
        RECT 79.040 210.730 79.180 210.870 ;
        RECT 80.805 210.825 81.095 210.870 ;
        RECT 84.470 211.010 84.790 211.070 ;
        RECT 85.020 211.055 85.160 211.210 ;
        RECT 88.165 211.165 88.455 211.210 ;
        RECT 93.760 211.055 93.900 211.550 ;
        RECT 107.010 211.490 107.330 211.550 ;
        RECT 112.070 211.690 112.390 211.750 ;
        RECT 116.225 211.690 116.515 211.735 ;
        RECT 112.070 211.550 116.515 211.690 ;
        RECT 112.070 211.490 112.390 211.550 ;
        RECT 116.225 211.505 116.515 211.550 ;
        RECT 118.050 211.490 118.370 211.750 ;
        RECT 123.570 211.490 123.890 211.750 ;
        RECT 125.410 211.690 125.730 211.750 ;
        RECT 129.550 211.690 129.870 211.750 ;
        RECT 125.410 211.550 129.870 211.690 ;
        RECT 125.410 211.490 125.730 211.550 ;
        RECT 129.550 211.490 129.870 211.550 ;
        RECT 138.765 211.690 139.055 211.735 ;
        RECT 140.590 211.690 140.910 211.750 ;
        RECT 138.765 211.550 140.910 211.690 ;
        RECT 138.765 211.505 139.055 211.550 ;
        RECT 140.590 211.490 140.910 211.550 ;
        RECT 141.065 211.690 141.355 211.735 ;
        RECT 148.425 211.690 148.715 211.735 ;
        RECT 150.340 211.690 150.480 212.570 ;
        RECT 141.065 211.550 142.200 211.690 ;
        RECT 141.065 211.505 141.355 211.550 ;
        RECT 120.350 211.350 120.670 211.410 ;
        RECT 142.060 211.350 142.200 211.550 ;
        RECT 148.425 211.550 150.480 211.690 ;
        RECT 148.425 211.505 148.715 211.550 ;
        RECT 142.750 211.350 143.040 211.395 ;
        RECT 95.140 211.210 102.640 211.350 ;
        RECT 95.140 211.055 95.280 211.210 ;
        RECT 102.500 211.055 102.640 211.210 ;
        RECT 107.560 211.210 141.740 211.350 ;
        RECT 142.060 211.210 143.040 211.350 ;
        RECT 84.945 211.010 85.235 211.055 ;
        RECT 84.470 210.870 85.235 211.010 ;
        RECT 84.470 210.810 84.790 210.870 ;
        RECT 84.945 210.825 85.235 210.870 ;
        RECT 86.325 210.825 86.615 211.055 ;
        RECT 93.685 210.825 93.975 211.055 ;
        RECT 95.065 210.825 95.355 211.055 ;
        RECT 96.345 211.010 96.635 211.055 ;
        RECT 95.600 210.870 96.635 211.010 ;
        RECT 75.360 210.530 78.260 210.670 ;
        RECT 67.925 210.330 68.215 210.375 ;
        RECT 59.720 210.190 68.215 210.330 ;
        RECT 55.070 210.145 55.360 210.190 ;
        RECT 57.170 210.145 57.460 210.190 ;
        RECT 58.740 210.145 59.030 210.190 ;
        RECT 67.925 210.145 68.215 210.190 ;
        RECT 38.470 209.990 38.790 210.050 ;
        RECT 37.640 209.850 38.790 209.990 ;
        RECT 38.470 209.790 38.790 209.850 ;
        RECT 42.610 209.790 42.930 210.050 ;
        RECT 53.205 209.990 53.495 210.035 ;
        RECT 54.570 209.990 54.890 210.050 ;
        RECT 53.205 209.850 54.890 209.990 ;
        RECT 53.205 209.805 53.495 209.850 ;
        RECT 54.570 209.790 54.890 209.850 ;
        RECT 64.230 209.990 64.550 210.050 ;
        RECT 65.165 209.990 65.455 210.035 ;
        RECT 64.230 209.850 65.455 209.990 ;
        RECT 71.680 209.990 71.820 210.485 ;
        RECT 72.985 210.330 73.275 210.375 ;
        RECT 75.360 210.330 75.500 210.530 ;
        RECT 78.950 210.470 79.270 210.730 ;
        RECT 79.870 210.470 80.190 210.730 ;
        RECT 81.725 210.670 82.015 210.715 ;
        RECT 82.185 210.670 82.475 210.715 ;
        RECT 86.400 210.670 86.540 210.825 ;
        RECT 90.005 210.670 90.295 210.715 ;
        RECT 95.600 210.670 95.740 210.870 ;
        RECT 96.345 210.825 96.635 210.870 ;
        RECT 102.425 210.825 102.715 211.055 ;
        RECT 103.760 211.010 104.050 211.055 ;
        RECT 106.090 211.010 106.410 211.070 ;
        RECT 103.760 210.870 106.410 211.010 ;
        RECT 103.760 210.825 104.050 210.870 ;
        RECT 81.725 210.530 90.295 210.670 ;
        RECT 81.725 210.485 82.015 210.530 ;
        RECT 82.185 210.485 82.475 210.530 ;
        RECT 90.005 210.485 90.295 210.530 ;
        RECT 94.680 210.530 95.740 210.670 ;
        RECT 95.945 210.670 96.235 210.715 ;
        RECT 97.135 210.670 97.425 210.715 ;
        RECT 99.655 210.670 99.945 210.715 ;
        RECT 95.945 210.530 99.945 210.670 ;
        RECT 72.985 210.190 75.500 210.330 ;
        RECT 72.985 210.145 73.275 210.190 ;
        RECT 83.550 210.130 83.870 210.390 ;
        RECT 94.680 210.375 94.820 210.530 ;
        RECT 95.945 210.485 96.235 210.530 ;
        RECT 97.135 210.485 97.425 210.530 ;
        RECT 99.655 210.485 99.945 210.530 ;
        RECT 94.605 210.145 94.895 210.375 ;
        RECT 95.550 210.330 95.840 210.375 ;
        RECT 97.650 210.330 97.940 210.375 ;
        RECT 99.220 210.330 99.510 210.375 ;
        RECT 95.550 210.190 99.510 210.330 ;
        RECT 95.550 210.145 95.840 210.190 ;
        RECT 97.650 210.145 97.940 210.190 ;
        RECT 99.220 210.145 99.510 210.190 ;
        RECT 73.890 209.990 74.210 210.050 ;
        RECT 71.680 209.850 74.210 209.990 ;
        RECT 64.230 209.790 64.550 209.850 ;
        RECT 65.165 209.805 65.455 209.850 ;
        RECT 73.890 209.790 74.210 209.850 ;
        RECT 75.745 209.990 76.035 210.035 ;
        RECT 79.870 209.990 80.190 210.050 ;
        RECT 75.745 209.850 80.190 209.990 ;
        RECT 75.745 209.805 76.035 209.850 ;
        RECT 79.870 209.790 80.190 209.850 ;
        RECT 87.230 209.790 87.550 210.050 ;
        RECT 87.690 209.990 88.010 210.050 ;
        RECT 89.545 209.990 89.835 210.035 ;
        RECT 87.690 209.850 89.835 209.990 ;
        RECT 87.690 209.790 88.010 209.850 ;
        RECT 89.545 209.805 89.835 209.850 ;
        RECT 89.990 209.790 90.310 210.050 ;
        RECT 99.650 209.990 99.970 210.050 ;
        RECT 101.965 209.990 102.255 210.035 ;
        RECT 99.650 209.850 102.255 209.990 ;
        RECT 102.500 209.990 102.640 210.825 ;
        RECT 106.090 210.810 106.410 210.870 ;
        RECT 103.305 210.670 103.595 210.715 ;
        RECT 104.495 210.670 104.785 210.715 ;
        RECT 107.015 210.670 107.305 210.715 ;
        RECT 103.305 210.530 107.305 210.670 ;
        RECT 103.305 210.485 103.595 210.530 ;
        RECT 104.495 210.485 104.785 210.530 ;
        RECT 107.015 210.485 107.305 210.530 ;
        RECT 102.910 210.330 103.200 210.375 ;
        RECT 105.010 210.330 105.300 210.375 ;
        RECT 106.580 210.330 106.870 210.375 ;
        RECT 102.910 210.190 106.870 210.330 ;
        RECT 102.910 210.145 103.200 210.190 ;
        RECT 105.010 210.145 105.300 210.190 ;
        RECT 106.580 210.145 106.870 210.190 ;
        RECT 107.560 209.990 107.700 211.210 ;
        RECT 120.350 211.150 120.670 211.210 ;
        RECT 111.625 211.010 111.915 211.055 ;
        RECT 111.625 210.870 115.520 211.010 ;
        RECT 111.625 210.825 111.915 210.870 ;
        RECT 109.310 210.670 109.630 210.730 ;
        RECT 110.705 210.670 110.995 210.715 ;
        RECT 109.310 210.530 110.995 210.670 ;
        RECT 109.310 210.470 109.630 210.530 ;
        RECT 110.705 210.485 110.995 210.530 ;
        RECT 113.005 210.670 113.295 210.715 ;
        RECT 114.830 210.670 115.150 210.730 ;
        RECT 113.005 210.530 115.150 210.670 ;
        RECT 115.380 210.670 115.520 210.870 ;
        RECT 115.750 210.810 116.070 211.070 ;
        RECT 118.985 211.010 119.275 211.055 ;
        RECT 121.270 211.010 121.590 211.070 ;
        RECT 121.745 211.010 122.035 211.055 ;
        RECT 124.490 211.010 124.810 211.070 ;
        RECT 116.300 210.870 122.035 211.010 ;
        RECT 116.300 210.670 116.440 210.870 ;
        RECT 118.985 210.825 119.275 210.870 ;
        RECT 121.270 210.810 121.590 210.870 ;
        RECT 121.745 210.825 122.035 210.870 ;
        RECT 122.740 210.870 124.810 211.010 ;
        RECT 115.380 210.530 116.440 210.670 ;
        RECT 117.145 210.670 117.435 210.715 ;
        RECT 118.510 210.670 118.830 210.730 ;
        RECT 117.145 210.530 118.830 210.670 ;
        RECT 113.005 210.485 113.295 210.530 ;
        RECT 114.830 210.470 115.150 210.530 ;
        RECT 117.145 210.485 117.435 210.530 ;
        RECT 118.510 210.470 118.830 210.530 ;
        RECT 120.365 210.670 120.655 210.715 ;
        RECT 122.740 210.670 122.880 210.870 ;
        RECT 124.490 210.810 124.810 210.870 ;
        RECT 126.330 211.010 126.650 211.070 ;
        RECT 131.940 211.055 132.080 211.210 ;
        RECT 133.230 211.055 133.550 211.070 ;
        RECT 141.600 211.055 141.740 211.210 ;
        RECT 142.750 211.165 143.040 211.210 ;
        RECT 129.105 211.010 129.395 211.055 ;
        RECT 126.330 210.870 129.395 211.010 ;
        RECT 126.330 210.810 126.650 210.870 ;
        RECT 129.105 210.825 129.395 210.870 ;
        RECT 129.565 210.825 129.855 211.055 ;
        RECT 131.865 210.825 132.155 211.055 ;
        RECT 133.200 211.010 133.550 211.055 ;
        RECT 140.145 211.010 140.435 211.055 ;
        RECT 133.035 210.870 133.550 211.010 ;
        RECT 133.200 210.825 133.550 210.870 ;
        RECT 120.365 210.530 122.880 210.670 ;
        RECT 120.365 210.485 120.655 210.530 ;
        RECT 123.110 210.470 123.430 210.730 ;
        RECT 125.885 210.670 126.175 210.715 ;
        RECT 125.500 210.530 126.175 210.670 ;
        RECT 112.530 210.130 112.850 210.390 ;
        RECT 118.970 210.130 119.290 210.390 ;
        RECT 120.810 210.130 121.130 210.390 ;
        RECT 102.500 209.850 107.700 209.990 ;
        RECT 109.325 209.990 109.615 210.035 ;
        RECT 110.230 209.990 110.550 210.050 ;
        RECT 109.325 209.850 110.550 209.990 ;
        RECT 99.650 209.790 99.970 209.850 ;
        RECT 101.965 209.805 102.255 209.850 ;
        RECT 109.325 209.805 109.615 209.850 ;
        RECT 110.230 209.790 110.550 209.850 ;
        RECT 113.910 209.790 114.230 210.050 ;
        RECT 119.060 209.990 119.200 210.130 ;
        RECT 119.905 209.990 120.195 210.035 ;
        RECT 122.650 209.990 122.970 210.050 ;
        RECT 119.060 209.850 122.970 209.990 ;
        RECT 125.500 209.990 125.640 210.530 ;
        RECT 125.885 210.485 126.175 210.530 ;
        RECT 126.805 210.670 127.095 210.715 ;
        RECT 127.250 210.670 127.570 210.730 ;
        RECT 128.185 210.670 128.475 210.715 ;
        RECT 129.640 210.670 129.780 210.825 ;
        RECT 133.230 210.810 133.550 210.825 ;
        RECT 137.000 210.870 140.435 211.010 ;
        RECT 126.805 210.530 128.475 210.670 ;
        RECT 126.805 210.485 127.095 210.530 ;
        RECT 127.250 210.470 127.570 210.530 ;
        RECT 128.185 210.485 128.475 210.530 ;
        RECT 129.180 210.530 129.780 210.670 ;
        RECT 132.745 210.670 133.035 210.715 ;
        RECT 133.935 210.670 134.225 210.715 ;
        RECT 136.455 210.670 136.745 210.715 ;
        RECT 132.745 210.530 136.745 210.670 ;
        RECT 127.710 210.330 128.030 210.390 ;
        RECT 129.180 210.330 129.320 210.530 ;
        RECT 132.745 210.485 133.035 210.530 ;
        RECT 133.935 210.485 134.225 210.530 ;
        RECT 136.455 210.485 136.745 210.530 ;
        RECT 127.710 210.190 129.320 210.330 ;
        RECT 132.350 210.330 132.640 210.375 ;
        RECT 134.450 210.330 134.740 210.375 ;
        RECT 136.020 210.330 136.310 210.375 ;
        RECT 132.350 210.190 136.310 210.330 ;
        RECT 127.710 210.130 128.030 210.190 ;
        RECT 132.350 210.145 132.640 210.190 ;
        RECT 134.450 210.145 134.740 210.190 ;
        RECT 136.020 210.145 136.310 210.190 ;
        RECT 126.330 209.990 126.650 210.050 ;
        RECT 125.500 209.850 126.650 209.990 ;
        RECT 119.905 209.805 120.195 209.850 ;
        RECT 122.650 209.790 122.970 209.850 ;
        RECT 126.330 209.790 126.650 209.850 ;
        RECT 131.405 209.990 131.695 210.035 ;
        RECT 137.000 209.990 137.140 210.870 ;
        RECT 140.145 210.825 140.435 210.870 ;
        RECT 141.525 210.825 141.815 211.055 ;
        RECT 142.405 210.670 142.695 210.715 ;
        RECT 143.595 210.670 143.885 210.715 ;
        RECT 146.115 210.670 146.405 210.715 ;
        RECT 142.405 210.530 146.405 210.670 ;
        RECT 142.405 210.485 142.695 210.530 ;
        RECT 143.595 210.485 143.885 210.530 ;
        RECT 146.115 210.485 146.405 210.530 ;
        RECT 142.010 210.330 142.300 210.375 ;
        RECT 144.110 210.330 144.400 210.375 ;
        RECT 145.680 210.330 145.970 210.375 ;
        RECT 142.010 210.190 145.970 210.330 ;
        RECT 142.010 210.145 142.300 210.190 ;
        RECT 144.110 210.145 144.400 210.190 ;
        RECT 145.680 210.145 145.970 210.190 ;
        RECT 131.405 209.850 137.140 209.990 ;
        RECT 131.405 209.805 131.695 209.850 ;
        RECT 36.100 209.170 150.180 209.650 ;
        RECT 42.610 208.770 42.930 209.030 ;
        RECT 45.370 208.770 45.690 209.030 ;
        RECT 47.670 208.770 47.990 209.030 ;
        RECT 72.510 208.970 72.830 209.030 ;
        RECT 75.745 208.970 76.035 209.015 ;
        RECT 72.510 208.830 76.035 208.970 ;
        RECT 72.510 208.770 72.830 208.830 ;
        RECT 75.745 208.785 76.035 208.830 ;
        RECT 76.190 208.970 76.510 209.030 ;
        RECT 78.505 208.970 78.795 209.015 ;
        RECT 76.190 208.830 78.795 208.970 ;
        RECT 76.190 208.770 76.510 208.830 ;
        RECT 78.505 208.785 78.795 208.830 ;
        RECT 82.185 208.970 82.475 209.015 ;
        RECT 83.550 208.970 83.870 209.030 ;
        RECT 82.185 208.830 83.870 208.970 ;
        RECT 82.185 208.785 82.475 208.830 ;
        RECT 83.550 208.770 83.870 208.830 ;
        RECT 87.690 208.770 88.010 209.030 ;
        RECT 88.165 208.970 88.455 209.015 ;
        RECT 89.990 208.970 90.310 209.030 ;
        RECT 88.165 208.830 90.310 208.970 ;
        RECT 88.165 208.785 88.455 208.830 ;
        RECT 89.990 208.770 90.310 208.830 ;
        RECT 91.000 208.830 98.960 208.970 ;
        RECT 45.460 208.290 45.600 208.770 ;
        RECT 60.550 208.630 60.840 208.675 ;
        RECT 62.120 208.630 62.410 208.675 ;
        RECT 64.220 208.630 64.510 208.675 ;
        RECT 60.550 208.490 64.510 208.630 ;
        RECT 60.550 208.445 60.840 208.490 ;
        RECT 62.120 208.445 62.410 208.490 ;
        RECT 64.220 208.445 64.510 208.490 ;
        RECT 64.690 208.630 65.010 208.690 ;
        RECT 65.165 208.630 65.455 208.675 ;
        RECT 85.850 208.630 86.170 208.690 ;
        RECT 64.690 208.490 86.170 208.630 ;
        RECT 64.690 208.430 65.010 208.490 ;
        RECT 65.165 208.445 65.455 208.490 ;
        RECT 85.850 208.430 86.170 208.490 ;
        RECT 86.325 208.630 86.615 208.675 ;
        RECT 87.780 208.630 87.920 208.770 ;
        RECT 86.325 208.490 87.920 208.630 ;
        RECT 89.070 208.630 89.390 208.690 ;
        RECT 90.465 208.630 90.755 208.675 ;
        RECT 89.070 208.490 90.755 208.630 ;
        RECT 86.325 208.445 86.615 208.490 ;
        RECT 43.620 208.150 45.600 208.290 ;
        RECT 60.115 208.290 60.405 208.335 ;
        RECT 62.635 208.290 62.925 208.335 ;
        RECT 63.825 208.290 64.115 208.335 ;
        RECT 60.115 208.150 64.115 208.290 ;
        RECT 39.390 207.950 39.710 208.010 ;
        RECT 43.620 207.995 43.760 208.150 ;
        RECT 60.115 208.105 60.405 208.150 ;
        RECT 62.635 208.105 62.925 208.150 ;
        RECT 63.825 208.105 64.115 208.150 ;
        RECT 77.585 208.290 77.875 208.335 ;
        RECT 84.945 208.290 85.235 208.335 ;
        RECT 77.585 208.150 81.480 208.290 ;
        RECT 77.585 208.105 77.875 208.150 ;
        RECT 42.625 207.950 42.915 207.995 ;
        RECT 39.390 207.810 42.915 207.950 ;
        RECT 39.390 207.750 39.710 207.810 ;
        RECT 42.625 207.765 42.915 207.810 ;
        RECT 43.545 207.765 43.835 207.995 ;
        RECT 43.990 207.750 44.310 208.010 ;
        RECT 44.925 207.765 45.215 207.995 ;
        RECT 42.150 207.610 42.470 207.670 ;
        RECT 45.000 207.610 45.140 207.765 ;
        RECT 46.750 207.750 47.070 208.010 ;
        RECT 52.730 207.950 53.050 208.010 ;
        RECT 55.030 207.950 55.350 208.010 ;
        RECT 64.705 207.950 64.995 207.995 ;
        RECT 67.450 207.950 67.770 208.010 ;
        RECT 52.730 207.810 67.770 207.950 ;
        RECT 52.730 207.750 53.050 207.810 ;
        RECT 55.030 207.750 55.350 207.810 ;
        RECT 64.705 207.765 64.995 207.810 ;
        RECT 67.450 207.750 67.770 207.810 ;
        RECT 72.050 207.950 72.370 208.010 ;
        RECT 72.525 207.950 72.815 207.995 ;
        RECT 72.050 207.810 72.815 207.950 ;
        RECT 72.050 207.750 72.370 207.810 ;
        RECT 72.525 207.765 72.815 207.810 ;
        RECT 73.445 207.950 73.735 207.995 ;
        RECT 74.350 207.950 74.670 208.010 ;
        RECT 73.445 207.810 74.670 207.950 ;
        RECT 73.445 207.765 73.735 207.810 ;
        RECT 74.350 207.750 74.670 207.810 ;
        RECT 75.285 207.765 75.575 207.995 ;
        RECT 76.190 207.950 76.510 208.010 ;
        RECT 76.665 207.950 76.955 207.995 ;
        RECT 78.045 207.950 78.335 207.995 ;
        RECT 76.190 207.810 78.335 207.950 ;
        RECT 42.150 207.470 45.140 207.610 ;
        RECT 63.480 207.610 63.770 207.655 ;
        RECT 64.230 207.610 64.550 207.670 ;
        RECT 66.085 207.610 66.375 207.655 ;
        RECT 63.480 207.470 64.550 207.610 ;
        RECT 42.150 207.410 42.470 207.470 ;
        RECT 63.480 207.425 63.770 207.470 ;
        RECT 64.230 207.410 64.550 207.470 ;
        RECT 65.240 207.470 66.375 207.610 ;
        RECT 45.845 207.270 46.135 207.315 ;
        RECT 46.290 207.270 46.610 207.330 ;
        RECT 45.845 207.130 46.610 207.270 ;
        RECT 45.845 207.085 46.135 207.130 ;
        RECT 46.290 207.070 46.610 207.130 ;
        RECT 57.805 207.270 58.095 207.315 ;
        RECT 61.010 207.270 61.330 207.330 ;
        RECT 65.240 207.270 65.380 207.470 ;
        RECT 66.085 207.425 66.375 207.470 ;
        RECT 57.805 207.130 65.380 207.270 ;
        RECT 75.360 207.270 75.500 207.765 ;
        RECT 76.190 207.750 76.510 207.810 ;
        RECT 76.665 207.765 76.955 207.810 ;
        RECT 78.045 207.765 78.335 207.810 ;
        RECT 78.950 207.950 79.270 208.010 ;
        RECT 79.870 207.950 80.190 208.010 ;
        RECT 81.340 207.950 81.480 208.150 ;
        RECT 84.945 208.150 86.540 208.290 ;
        RECT 84.945 208.105 85.235 208.150 ;
        RECT 84.485 207.950 84.775 207.995 ;
        RECT 78.950 207.810 79.640 207.950 ;
        RECT 78.950 207.750 79.270 207.810 ;
        RECT 79.500 207.610 79.640 207.810 ;
        RECT 79.870 207.810 81.020 207.950 ;
        RECT 81.340 207.810 84.775 207.950 ;
        RECT 79.870 207.750 80.190 207.810 ;
        RECT 80.345 207.610 80.635 207.655 ;
        RECT 79.500 207.470 80.635 207.610 ;
        RECT 80.880 207.610 81.020 207.810 ;
        RECT 84.485 207.765 84.775 207.810 ;
        RECT 81.265 207.610 81.555 207.655 ;
        RECT 80.880 207.470 81.555 207.610 ;
        RECT 86.400 207.610 86.540 208.150 ;
        RECT 86.860 207.995 87.000 208.490 ;
        RECT 89.070 208.430 89.390 208.490 ;
        RECT 90.465 208.445 90.755 208.490 ;
        RECT 88.625 208.290 88.915 208.335 ;
        RECT 91.000 208.290 91.140 208.830 ;
        RECT 92.750 208.430 93.070 208.690 ;
        RECT 92.840 208.290 92.980 208.430 ;
        RECT 88.625 208.150 91.140 208.290 ;
        RECT 88.625 208.105 88.915 208.150 ;
        RECT 91.000 208.030 91.140 208.150 ;
        RECT 91.920 208.150 92.980 208.290 ;
        RECT 86.785 207.765 87.075 207.995 ;
        RECT 87.230 207.950 87.550 208.010 ;
        RECT 87.705 207.950 87.995 207.995 ;
        RECT 87.230 207.810 87.995 207.950 ;
        RECT 87.230 207.750 87.550 207.810 ;
        RECT 87.705 207.765 87.995 207.810 ;
        RECT 89.085 207.950 89.375 207.995 ;
        RECT 90.450 207.950 90.770 208.010 ;
        RECT 91.000 207.995 91.170 208.030 ;
        RECT 89.085 207.810 90.770 207.950 ;
        RECT 89.085 207.765 89.375 207.810 ;
        RECT 90.450 207.750 90.770 207.810 ;
        RECT 90.925 207.765 91.215 207.995 ;
        RECT 91.370 207.950 91.690 208.010 ;
        RECT 91.920 207.995 92.060 208.150 ;
        RECT 91.845 207.950 92.135 207.995 ;
        RECT 98.270 207.950 98.590 208.010 ;
        RECT 98.820 207.995 98.960 208.830 ;
        RECT 106.090 208.770 106.410 209.030 ;
        RECT 114.370 208.970 114.690 209.030 ;
        RECT 114.845 208.970 115.135 209.015 ;
        RECT 114.370 208.830 115.135 208.970 ;
        RECT 114.370 208.770 114.690 208.830 ;
        RECT 114.845 208.785 115.135 208.830 ;
        RECT 117.590 208.770 117.910 209.030 ;
        RECT 121.270 208.770 121.590 209.030 ;
        RECT 122.650 208.970 122.970 209.030 ;
        RECT 124.505 208.970 124.795 209.015 ;
        RECT 122.650 208.830 124.795 208.970 ;
        RECT 122.650 208.770 122.970 208.830 ;
        RECT 124.505 208.785 124.795 208.830 ;
        RECT 125.410 208.770 125.730 209.030 ;
        RECT 126.330 208.970 126.650 209.030 ;
        RECT 127.725 208.970 128.015 209.015 ;
        RECT 126.330 208.830 128.015 208.970 ;
        RECT 126.330 208.770 126.650 208.830 ;
        RECT 127.725 208.785 128.015 208.830 ;
        RECT 133.690 208.770 134.010 209.030 ;
        RECT 140.590 208.770 140.910 209.030 ;
        RECT 101.965 208.630 102.255 208.675 ;
        RECT 104.250 208.630 104.570 208.690 ;
        RECT 101.965 208.490 104.570 208.630 ;
        RECT 101.965 208.445 102.255 208.490 ;
        RECT 104.250 208.430 104.570 208.490 ;
        RECT 110.230 208.090 110.550 208.350 ;
        RECT 111.625 208.290 111.915 208.335 ;
        RECT 112.070 208.290 112.390 208.350 ;
        RECT 111.625 208.150 112.390 208.290 ;
        RECT 111.625 208.105 111.915 208.150 ;
        RECT 112.070 208.090 112.390 208.150 ;
        RECT 112.530 208.290 112.850 208.350 ;
        RECT 117.145 208.290 117.435 208.335 ;
        RECT 112.530 208.150 117.435 208.290 ;
        RECT 112.530 208.090 112.850 208.150 ;
        RECT 117.145 208.105 117.435 208.150 ;
        RECT 91.370 207.810 92.135 207.950 ;
        RECT 91.370 207.750 91.690 207.810 ;
        RECT 91.845 207.765 92.135 207.810 ;
        RECT 92.380 207.810 98.590 207.950 ;
        RECT 92.380 207.610 92.520 207.810 ;
        RECT 98.270 207.750 98.590 207.810 ;
        RECT 98.745 207.765 99.035 207.995 ;
        RECT 86.400 207.470 92.520 207.610 ;
        RECT 98.820 207.610 98.960 207.765 ;
        RECT 99.190 207.750 99.510 208.010 ;
        RECT 99.650 207.750 99.970 208.010 ;
        RECT 102.410 207.750 102.730 208.010 ;
        RECT 103.345 207.950 103.635 207.995 ;
        RECT 106.550 207.950 106.870 208.010 ;
        RECT 103.345 207.810 106.870 207.950 ;
        RECT 103.345 207.765 103.635 207.810 ;
        RECT 106.550 207.750 106.870 207.810 ;
        RECT 107.025 207.950 107.315 207.995 ;
        RECT 113.910 207.950 114.230 208.010 ;
        RECT 107.025 207.810 114.230 207.950 ;
        RECT 117.680 207.950 117.820 208.770 ;
        RECT 118.065 208.290 118.355 208.335 ;
        RECT 118.510 208.290 118.830 208.350 ;
        RECT 121.360 208.290 121.500 208.770 ;
        RECT 124.965 208.290 125.255 208.335 ;
        RECT 125.500 208.290 125.640 208.770 ;
        RECT 118.065 208.150 121.040 208.290 ;
        RECT 121.360 208.150 123.800 208.290 ;
        RECT 118.065 208.105 118.355 208.150 ;
        RECT 118.510 208.090 118.830 208.150 ;
        RECT 119.905 207.950 120.195 207.995 ;
        RECT 120.365 207.950 120.655 207.995 ;
        RECT 117.680 207.810 120.655 207.950 ;
        RECT 120.900 207.950 121.040 208.150 ;
        RECT 120.900 207.810 121.960 207.950 ;
        RECT 107.025 207.765 107.315 207.810 ;
        RECT 113.910 207.750 114.230 207.810 ;
        RECT 119.905 207.765 120.195 207.810 ;
        RECT 120.365 207.765 120.655 207.810 ;
        RECT 121.820 207.610 121.960 207.810 ;
        RECT 122.650 207.750 122.970 208.010 ;
        RECT 123.660 207.995 123.800 208.150 ;
        RECT 124.965 208.150 125.640 208.290 ;
        RECT 128.720 208.490 131.620 208.630 ;
        RECT 124.965 208.105 125.255 208.150 ;
        RECT 123.585 207.765 123.875 207.995 ;
        RECT 126.790 207.950 127.110 208.010 ;
        RECT 127.725 207.950 128.015 207.995 ;
        RECT 126.790 207.810 128.015 207.950 ;
        RECT 126.790 207.750 127.110 207.810 ;
        RECT 127.725 207.765 128.015 207.810 ;
        RECT 128.170 207.950 128.490 208.010 ;
        RECT 128.720 207.995 128.860 208.490 ;
        RECT 129.090 208.290 129.410 208.350 ;
        RECT 131.480 208.335 131.620 208.490 ;
        RECT 130.485 208.290 130.775 208.335 ;
        RECT 129.090 208.150 130.775 208.290 ;
        RECT 129.090 208.090 129.410 208.150 ;
        RECT 130.485 208.105 130.775 208.150 ;
        RECT 131.405 208.290 131.695 208.335 ;
        RECT 136.465 208.290 136.755 208.335 ;
        RECT 131.405 208.150 136.755 208.290 ;
        RECT 131.405 208.105 131.695 208.150 ;
        RECT 136.465 208.105 136.755 208.150 ;
        RECT 128.645 207.950 128.935 207.995 ;
        RECT 128.170 207.810 128.935 207.950 ;
        RECT 128.170 207.750 128.490 207.810 ;
        RECT 128.645 207.765 128.935 207.810 ;
        RECT 129.180 207.610 129.320 208.090 ;
        RECT 131.865 207.950 132.155 207.995 ;
        RECT 134.150 207.950 134.470 208.010 ;
        RECT 131.865 207.810 134.470 207.950 ;
        RECT 131.865 207.765 132.155 207.810 ;
        RECT 134.150 207.750 134.470 207.810 ;
        RECT 137.385 207.950 137.675 207.995 ;
        RECT 140.680 207.950 140.820 208.770 ;
        RECT 137.385 207.810 140.820 207.950 ;
        RECT 137.385 207.765 137.675 207.810 ;
        RECT 98.820 207.470 103.560 207.610 ;
        RECT 80.345 207.425 80.635 207.470 ;
        RECT 81.265 207.425 81.555 207.470 ;
        RECT 83.090 207.270 83.410 207.330 ;
        RECT 75.360 207.130 83.410 207.270 ;
        RECT 57.805 207.085 58.095 207.130 ;
        RECT 61.010 207.070 61.330 207.130 ;
        RECT 83.090 207.070 83.410 207.130 ;
        RECT 88.150 207.270 88.470 207.330 ;
        RECT 91.385 207.270 91.675 207.315 ;
        RECT 88.150 207.130 91.675 207.270 ;
        RECT 103.420 207.270 103.560 207.470 ;
        RECT 115.840 207.470 120.120 207.610 ;
        RECT 121.820 207.470 129.320 207.610 ;
        RECT 115.840 207.270 115.980 207.470 ;
        RECT 119.980 207.330 120.120 207.470 ;
        RECT 103.420 207.130 115.980 207.270 ;
        RECT 116.685 207.270 116.975 207.315 ;
        RECT 117.130 207.270 117.450 207.330 ;
        RECT 116.685 207.130 117.450 207.270 ;
        RECT 88.150 207.070 88.470 207.130 ;
        RECT 91.385 207.085 91.675 207.130 ;
        RECT 116.685 207.085 116.975 207.130 ;
        RECT 117.130 207.070 117.450 207.130 ;
        RECT 117.590 207.270 117.910 207.330 ;
        RECT 118.985 207.270 119.275 207.315 ;
        RECT 117.590 207.130 119.275 207.270 ;
        RECT 117.590 207.070 117.910 207.130 ;
        RECT 118.985 207.085 119.275 207.130 ;
        RECT 119.890 207.070 120.210 207.330 ;
        RECT 126.790 207.070 127.110 207.330 ;
        RECT 36.100 206.450 150.180 206.930 ;
        RECT 52.730 206.250 53.050 206.310 ;
        RECT 45.000 206.110 53.050 206.250 ;
        RECT 38.930 205.910 39.250 205.970 ;
        RECT 42.625 205.910 42.915 205.955 ;
        RECT 38.930 205.770 42.915 205.910 ;
        RECT 38.930 205.710 39.250 205.770 ;
        RECT 42.625 205.725 42.915 205.770 ;
        RECT 43.705 205.910 43.995 205.955 ;
        RECT 44.450 205.910 44.770 205.970 ;
        RECT 43.705 205.770 44.770 205.910 ;
        RECT 43.705 205.725 43.995 205.770 ;
        RECT 44.450 205.710 44.770 205.770 ;
        RECT 38.470 205.570 38.790 205.630 ;
        RECT 45.000 205.615 45.140 206.110 ;
        RECT 52.730 206.050 53.050 206.110 ;
        RECT 72.525 206.250 72.815 206.295 ;
        RECT 76.190 206.250 76.510 206.310 ;
        RECT 98.730 206.250 99.050 206.310 ;
        RECT 120.810 206.250 121.130 206.310 ;
        RECT 72.525 206.110 76.510 206.250 ;
        RECT 72.525 206.065 72.815 206.110 ;
        RECT 76.190 206.050 76.510 206.110 ;
        RECT 76.740 206.110 95.510 206.250 ;
        RECT 46.290 205.955 46.610 205.970 ;
        RECT 46.260 205.910 46.610 205.955 ;
        RECT 67.910 205.910 68.230 205.970 ;
        RECT 72.050 205.910 72.370 205.970 ;
        RECT 46.260 205.770 46.760 205.910 ;
        RECT 50.520 205.770 68.230 205.910 ;
        RECT 46.260 205.725 46.610 205.770 ;
        RECT 46.290 205.710 46.610 205.725 ;
        RECT 44.925 205.570 45.215 205.615 ;
        RECT 38.470 205.430 45.215 205.570 ;
        RECT 38.470 205.370 38.790 205.430 ;
        RECT 44.925 205.385 45.215 205.430 ;
        RECT 45.805 205.230 46.095 205.275 ;
        RECT 46.995 205.230 47.285 205.275 ;
        RECT 49.515 205.230 49.805 205.275 ;
        RECT 45.805 205.090 49.805 205.230 ;
        RECT 45.805 205.045 46.095 205.090 ;
        RECT 46.995 205.045 47.285 205.090 ;
        RECT 49.515 205.045 49.805 205.090 ;
        RECT 45.410 204.890 45.700 204.935 ;
        RECT 47.510 204.890 47.800 204.935 ;
        RECT 49.080 204.890 49.370 204.935 ;
        RECT 45.410 204.750 49.370 204.890 ;
        RECT 45.410 204.705 45.700 204.750 ;
        RECT 47.510 204.705 47.800 204.750 ;
        RECT 49.080 204.705 49.370 204.750 ;
        RECT 50.520 204.610 50.660 205.770 ;
        RECT 67.910 205.710 68.230 205.770 ;
        RECT 71.680 205.770 72.370 205.910 ;
        RECT 63.770 205.570 64.090 205.630 ;
        RECT 71.680 205.615 71.820 205.770 ;
        RECT 72.050 205.710 72.370 205.770 ;
        RECT 73.890 205.910 74.210 205.970 ;
        RECT 76.740 205.910 76.880 206.110 ;
        RECT 73.890 205.770 76.880 205.910 ;
        RECT 84.470 205.910 84.790 205.970 ;
        RECT 85.405 205.910 85.695 205.955 ;
        RECT 93.670 205.910 93.990 205.970 ;
        RECT 84.470 205.770 85.695 205.910 ;
        RECT 73.890 205.710 74.210 205.770 ;
        RECT 84.470 205.710 84.790 205.770 ;
        RECT 64.705 205.570 64.995 205.615 ;
        RECT 65.165 205.570 65.455 205.615 ;
        RECT 63.770 205.430 65.455 205.570 ;
        RECT 63.770 205.370 64.090 205.430 ;
        RECT 64.705 205.385 64.995 205.430 ;
        RECT 65.165 205.385 65.455 205.430 ;
        RECT 71.605 205.385 71.895 205.615 ;
        RECT 72.525 205.385 72.815 205.615 ;
        RECT 54.110 205.230 54.430 205.290 ;
        RECT 62.390 205.230 62.710 205.290 ;
        RECT 71.680 205.230 71.820 205.385 ;
        RECT 54.110 205.090 71.820 205.230 ;
        RECT 72.600 205.230 72.740 205.385 ;
        RECT 77.110 205.370 77.430 205.630 ;
        RECT 85.020 205.615 85.160 205.770 ;
        RECT 85.405 205.725 85.695 205.770 ;
        RECT 88.240 205.770 93.990 205.910 ;
        RECT 95.370 205.910 95.510 206.110 ;
        RECT 98.730 206.110 121.130 206.250 ;
        RECT 98.730 206.050 99.050 206.110 ;
        RECT 120.810 206.050 121.130 206.110 ;
        RECT 122.190 206.250 122.510 206.310 ;
        RECT 122.665 206.250 122.955 206.295 ;
        RECT 122.190 206.110 122.955 206.250 ;
        RECT 122.190 206.050 122.510 206.110 ;
        RECT 122.665 206.065 122.955 206.110 ;
        RECT 123.570 206.250 123.890 206.310 ;
        RECT 125.410 206.250 125.730 206.310 ;
        RECT 123.570 206.110 125.730 206.250 ;
        RECT 123.570 206.050 123.890 206.110 ;
        RECT 125.410 206.050 125.730 206.110 ;
        RECT 125.870 206.050 126.190 206.310 ;
        RECT 126.790 206.050 127.110 206.310 ;
        RECT 127.725 206.065 128.015 206.295 ;
        RECT 113.925 205.910 114.215 205.955 ;
        RECT 123.110 205.910 123.430 205.970 ;
        RECT 126.880 205.910 127.020 206.050 ;
        RECT 95.370 205.770 113.680 205.910 ;
        RECT 84.025 205.385 84.315 205.615 ;
        RECT 84.945 205.570 85.235 205.615 ;
        RECT 86.325 205.570 86.615 205.615 ;
        RECT 87.230 205.570 87.550 205.630 ;
        RECT 84.945 205.430 85.345 205.570 ;
        RECT 86.325 205.430 87.550 205.570 ;
        RECT 84.945 205.385 85.235 205.430 ;
        RECT 86.325 205.385 86.615 205.430 ;
        RECT 74.350 205.230 74.670 205.290 ;
        RECT 72.600 205.090 74.670 205.230 ;
        RECT 77.200 205.230 77.340 205.370 ;
        RECT 79.870 205.230 80.190 205.290 ;
        RECT 77.200 205.090 80.190 205.230 ;
        RECT 54.110 205.030 54.430 205.090 ;
        RECT 62.390 205.030 62.710 205.090 ;
        RECT 74.350 205.030 74.670 205.090 ;
        RECT 79.870 205.030 80.190 205.090 ;
        RECT 81.250 205.230 81.570 205.290 ;
        RECT 84.100 205.230 84.240 205.385 ;
        RECT 86.400 205.230 86.540 205.385 ;
        RECT 87.230 205.370 87.550 205.430 ;
        RECT 81.250 205.090 86.540 205.230 ;
        RECT 81.250 205.030 81.570 205.090 ;
        RECT 62.850 204.890 63.170 204.950 ;
        RECT 88.240 204.890 88.380 205.770 ;
        RECT 93.670 205.710 93.990 205.770 ;
        RECT 89.070 205.370 89.390 205.630 ;
        RECT 88.625 205.045 88.915 205.275 ;
        RECT 91.845 205.045 92.135 205.275 ;
        RECT 92.290 205.230 92.610 205.290 ;
        RECT 112.990 205.230 113.310 205.290 ;
        RECT 92.290 205.090 113.310 205.230 ;
        RECT 113.540 205.230 113.680 205.770 ;
        RECT 113.925 205.770 123.430 205.910 ;
        RECT 113.925 205.725 114.215 205.770 ;
        RECT 123.110 205.710 123.430 205.770 ;
        RECT 123.660 205.770 127.020 205.910 ;
        RECT 127.800 205.910 127.940 206.065 ;
        RECT 129.090 206.050 129.410 206.310 ;
        RECT 141.065 206.065 141.355 206.295 ;
        RECT 140.590 205.910 140.910 205.970 ;
        RECT 127.800 205.770 133.460 205.910 ;
        RECT 114.845 205.570 115.135 205.615 ;
        RECT 117.590 205.570 117.910 205.630 ;
        RECT 123.660 205.615 123.800 205.770 ;
        RECT 114.845 205.430 117.910 205.570 ;
        RECT 114.845 205.385 115.135 205.430 ;
        RECT 117.590 205.370 117.910 205.430 ;
        RECT 118.985 205.570 119.275 205.615 ;
        RECT 122.205 205.570 122.495 205.615 ;
        RECT 123.585 205.570 123.875 205.615 ;
        RECT 125.870 205.570 126.190 205.630 ;
        RECT 118.985 205.430 121.960 205.570 ;
        RECT 118.985 205.385 119.275 205.430 ;
        RECT 116.225 205.230 116.515 205.275 ;
        RECT 117.130 205.230 117.450 205.290 ;
        RECT 121.820 205.230 121.960 205.430 ;
        RECT 122.205 205.430 123.875 205.570 ;
        RECT 122.205 205.385 122.495 205.430 ;
        RECT 123.585 205.385 123.875 205.430 ;
        RECT 124.120 205.430 126.190 205.570 ;
        RECT 124.120 205.230 124.260 205.430 ;
        RECT 125.870 205.370 126.190 205.430 ;
        RECT 129.565 205.570 129.855 205.615 ;
        RECT 132.310 205.570 132.630 205.630 ;
        RECT 133.320 205.615 133.460 205.770 ;
        RECT 134.240 205.770 140.910 205.910 ;
        RECT 141.140 205.910 141.280 206.065 ;
        RECT 142.750 205.910 143.040 205.955 ;
        RECT 141.140 205.770 143.040 205.910 ;
        RECT 129.565 205.430 132.630 205.570 ;
        RECT 129.565 205.385 129.855 205.430 ;
        RECT 132.310 205.370 132.630 205.430 ;
        RECT 133.245 205.385 133.535 205.615 ;
        RECT 113.540 205.090 115.520 205.230 ;
        RECT 62.850 204.750 88.380 204.890 ;
        RECT 62.850 204.690 63.170 204.750 ;
        RECT 43.530 204.350 43.850 204.610 ;
        RECT 44.465 204.550 44.755 204.595 ;
        RECT 46.750 204.550 47.070 204.610 ;
        RECT 44.465 204.410 47.070 204.550 ;
        RECT 44.465 204.365 44.755 204.410 ;
        RECT 46.750 204.350 47.070 204.410 ;
        RECT 50.430 204.350 50.750 204.610 ;
        RECT 51.825 204.550 52.115 204.595 ;
        RECT 60.090 204.550 60.410 204.610 ;
        RECT 51.825 204.410 60.410 204.550 ;
        RECT 51.825 204.365 52.115 204.410 ;
        RECT 60.090 204.350 60.410 204.410 ;
        RECT 63.770 204.350 64.090 204.610 ;
        RECT 65.610 204.350 65.930 204.610 ;
        RECT 67.910 204.550 68.230 204.610 ;
        RECT 73.430 204.550 73.750 204.610 ;
        RECT 67.910 204.410 73.750 204.550 ;
        RECT 67.910 204.350 68.230 204.410 ;
        RECT 73.430 204.350 73.750 204.410 ;
        RECT 78.045 204.550 78.335 204.595 ;
        RECT 83.090 204.550 83.410 204.610 ;
        RECT 78.045 204.410 83.410 204.550 ;
        RECT 78.045 204.365 78.335 204.410 ;
        RECT 83.090 204.350 83.410 204.410 ;
        RECT 84.485 204.550 84.775 204.595 ;
        RECT 86.770 204.550 87.090 204.610 ;
        RECT 84.485 204.410 87.090 204.550 ;
        RECT 84.485 204.365 84.775 204.410 ;
        RECT 86.770 204.350 87.090 204.410 ;
        RECT 87.245 204.550 87.535 204.595 ;
        RECT 87.690 204.550 88.010 204.610 ;
        RECT 87.245 204.410 88.010 204.550 ;
        RECT 88.700 204.550 88.840 205.045 ;
        RECT 89.070 204.890 89.390 204.950 ;
        RECT 90.465 204.890 90.755 204.935 ;
        RECT 89.070 204.750 90.755 204.890 ;
        RECT 89.070 204.690 89.390 204.750 ;
        RECT 90.465 204.705 90.755 204.750 ;
        RECT 90.910 204.890 91.230 204.950 ;
        RECT 91.920 204.890 92.060 205.045 ;
        RECT 92.290 205.030 92.610 205.090 ;
        RECT 112.990 205.030 113.310 205.090 ;
        RECT 115.380 204.950 115.520 205.090 ;
        RECT 116.225 205.090 119.200 205.230 ;
        RECT 121.820 205.090 124.260 205.230 ;
        RECT 116.225 205.045 116.515 205.090 ;
        RECT 117.130 205.030 117.450 205.090 ;
        RECT 90.910 204.750 105.860 204.890 ;
        RECT 90.910 204.690 91.230 204.750 ;
        RECT 105.720 204.610 105.860 204.750 ;
        RECT 115.290 204.690 115.610 204.950 ;
        RECT 115.765 204.890 116.055 204.935 ;
        RECT 119.060 204.890 119.200 205.090 ;
        RECT 124.950 205.030 125.270 205.290 ;
        RECT 125.410 205.230 125.730 205.290 ;
        RECT 134.240 205.230 134.380 205.770 ;
        RECT 140.590 205.710 140.910 205.770 ;
        RECT 142.750 205.725 143.040 205.770 ;
        RECT 140.130 205.370 140.450 205.630 ;
        RECT 125.410 205.090 134.380 205.230 ;
        RECT 134.610 205.230 134.930 205.290 ;
        RECT 141.525 205.230 141.815 205.275 ;
        RECT 134.610 205.090 141.815 205.230 ;
        RECT 125.410 205.030 125.730 205.090 ;
        RECT 134.610 205.030 134.930 205.090 ;
        RECT 141.525 205.045 141.815 205.090 ;
        RECT 142.405 205.230 142.695 205.275 ;
        RECT 143.595 205.230 143.885 205.275 ;
        RECT 146.115 205.230 146.405 205.275 ;
        RECT 142.405 205.090 146.405 205.230 ;
        RECT 142.405 205.045 142.695 205.090 ;
        RECT 143.595 205.045 143.885 205.090 ;
        RECT 146.115 205.045 146.405 205.090 ;
        RECT 141.050 204.890 141.370 204.950 ;
        RECT 115.765 204.750 118.740 204.890 ;
        RECT 119.060 204.750 141.370 204.890 ;
        RECT 115.765 204.705 116.055 204.750 ;
        RECT 96.890 204.550 97.210 204.610 ;
        RECT 88.700 204.410 97.210 204.550 ;
        RECT 87.245 204.365 87.535 204.410 ;
        RECT 87.690 204.350 88.010 204.410 ;
        RECT 96.890 204.350 97.210 204.410 ;
        RECT 105.630 204.550 105.950 204.610 ;
        RECT 118.600 204.595 118.740 204.750 ;
        RECT 141.050 204.690 141.370 204.750 ;
        RECT 142.010 204.890 142.300 204.935 ;
        RECT 144.110 204.890 144.400 204.935 ;
        RECT 145.680 204.890 145.970 204.935 ;
        RECT 142.010 204.750 145.970 204.890 ;
        RECT 142.010 204.705 142.300 204.750 ;
        RECT 144.110 204.705 144.400 204.750 ;
        RECT 145.680 204.705 145.970 204.750 ;
        RECT 116.685 204.550 116.975 204.595 ;
        RECT 105.630 204.410 116.975 204.550 ;
        RECT 105.630 204.350 105.950 204.410 ;
        RECT 116.685 204.365 116.975 204.410 ;
        RECT 118.525 204.550 118.815 204.595 ;
        RECT 121.270 204.550 121.590 204.610 ;
        RECT 118.525 204.410 121.590 204.550 ;
        RECT 118.525 204.365 118.815 204.410 ;
        RECT 121.270 204.350 121.590 204.410 ;
        RECT 134.165 204.550 134.455 204.595 ;
        RECT 135.530 204.550 135.850 204.610 ;
        RECT 134.165 204.410 135.850 204.550 ;
        RECT 134.165 204.365 134.455 204.410 ;
        RECT 135.530 204.350 135.850 204.410 ;
        RECT 148.425 204.550 148.715 204.595 ;
        RECT 148.425 204.410 150.480 204.550 ;
        RECT 148.425 204.365 148.715 204.410 ;
        RECT 36.100 203.730 150.180 204.210 ;
        RECT 41.690 203.330 42.010 203.590 ;
        RECT 42.150 203.530 42.470 203.590 ;
        RECT 42.625 203.530 42.915 203.575 ;
        RECT 42.150 203.390 42.915 203.530 ;
        RECT 42.150 203.330 42.470 203.390 ;
        RECT 42.625 203.345 42.915 203.390 ;
        RECT 43.530 203.330 43.850 203.590 ;
        RECT 44.450 203.530 44.770 203.590 ;
        RECT 44.925 203.530 45.215 203.575 ;
        RECT 49.985 203.530 50.275 203.575 ;
        RECT 52.730 203.530 53.050 203.590 ;
        RECT 61.010 203.530 61.330 203.590 ;
        RECT 44.450 203.390 45.215 203.530 ;
        RECT 44.450 203.330 44.770 203.390 ;
        RECT 44.925 203.345 45.215 203.390 ;
        RECT 45.920 203.390 50.275 203.530 ;
        RECT 39.865 203.190 40.155 203.235 ;
        RECT 43.620 203.190 43.760 203.330 ;
        RECT 45.370 203.190 45.690 203.250 ;
        RECT 39.865 203.050 43.760 203.190 ;
        RECT 44.080 203.050 45.690 203.190 ;
        RECT 39.865 203.005 40.155 203.050 ;
        RECT 41.230 202.850 41.550 202.910 ;
        RECT 39.480 202.710 43.300 202.850 ;
        RECT 39.480 202.555 39.620 202.710 ;
        RECT 41.230 202.650 41.550 202.710 ;
        RECT 43.160 202.555 43.300 202.710 ;
        RECT 44.080 202.555 44.220 203.050 ;
        RECT 45.370 202.990 45.690 203.050 ;
        RECT 39.405 202.325 39.695 202.555 ;
        RECT 40.325 202.510 40.615 202.555 ;
        RECT 40.325 202.370 42.840 202.510 ;
        RECT 40.325 202.325 40.615 202.370 ;
        RECT 38.930 202.170 39.250 202.230 ;
        RECT 40.785 202.170 41.075 202.215 ;
        RECT 38.930 202.030 41.075 202.170 ;
        RECT 42.700 202.170 42.840 202.370 ;
        RECT 43.085 202.325 43.375 202.555 ;
        RECT 44.005 202.325 44.295 202.555 ;
        RECT 45.385 202.510 45.675 202.555 ;
        RECT 45.000 202.370 45.675 202.510 ;
        RECT 45.920 202.510 46.060 203.390 ;
        RECT 49.985 203.345 50.275 203.390 ;
        RECT 50.980 203.390 53.050 203.530 ;
        RECT 48.130 203.190 48.450 203.250 ;
        RECT 46.435 203.050 48.450 203.190 ;
        RECT 46.435 202.850 46.575 203.050 ;
        RECT 48.130 202.990 48.450 203.050 ;
        RECT 50.980 202.895 51.120 203.390 ;
        RECT 52.730 203.330 53.050 203.390 ;
        RECT 59.260 203.390 61.330 203.530 ;
        RECT 51.390 203.190 51.680 203.235 ;
        RECT 53.490 203.190 53.780 203.235 ;
        RECT 55.060 203.190 55.350 203.235 ;
        RECT 51.390 203.050 55.350 203.190 ;
        RECT 51.390 203.005 51.680 203.050 ;
        RECT 53.490 203.005 53.780 203.050 ;
        RECT 55.060 203.005 55.350 203.050 ;
        RECT 59.260 202.895 59.400 203.390 ;
        RECT 61.010 203.330 61.330 203.390 ;
        RECT 62.850 203.330 63.170 203.590 ;
        RECT 65.610 203.330 65.930 203.590 ;
        RECT 68.370 203.530 68.690 203.590 ;
        RECT 79.425 203.530 79.715 203.575 ;
        RECT 68.370 203.390 79.715 203.530 ;
        RECT 68.370 203.330 68.690 203.390 ;
        RECT 79.425 203.345 79.715 203.390 ;
        RECT 83.550 203.530 83.870 203.590 ;
        RECT 98.270 203.530 98.590 203.590 ;
        RECT 101.505 203.530 101.795 203.575 ;
        RECT 83.550 203.390 87.000 203.530 ;
        RECT 83.550 203.330 83.870 203.390 ;
        RECT 64.705 203.190 64.995 203.235 ;
        RECT 65.700 203.190 65.840 203.330 ;
        RECT 64.705 203.050 65.840 203.190 ;
        RECT 64.705 203.005 64.995 203.050 ;
        RECT 46.435 202.710 46.995 202.850 ;
        RECT 46.855 202.555 46.995 202.710 ;
        RECT 50.905 202.665 51.195 202.895 ;
        RECT 51.785 202.850 52.075 202.895 ;
        RECT 52.975 202.850 53.265 202.895 ;
        RECT 55.495 202.850 55.785 202.895 ;
        RECT 51.785 202.710 55.785 202.850 ;
        RECT 51.785 202.665 52.075 202.710 ;
        RECT 52.975 202.665 53.265 202.710 ;
        RECT 55.495 202.665 55.785 202.710 ;
        RECT 59.185 202.665 59.475 202.895 ;
        RECT 60.090 202.650 60.410 202.910 ;
        RECT 46.305 202.510 46.595 202.555 ;
        RECT 45.920 202.370 46.595 202.510 ;
        RECT 42.700 202.030 43.300 202.170 ;
        RECT 38.930 201.970 39.250 202.030 ;
        RECT 40.785 201.985 41.075 202.030 ;
        RECT 43.160 201.890 43.300 202.030 ;
        RECT 41.690 201.875 42.010 201.890 ;
        RECT 41.690 201.645 42.075 201.875 ;
        RECT 41.690 201.630 42.010 201.645 ;
        RECT 43.070 201.630 43.390 201.890 ;
        RECT 45.000 201.830 45.140 202.370 ;
        RECT 45.385 202.325 45.675 202.370 ;
        RECT 46.305 202.325 46.595 202.370 ;
        RECT 46.765 202.325 47.055 202.555 ;
        RECT 47.455 202.510 47.745 202.555 ;
        RECT 48.130 202.510 48.450 202.570 ;
        RECT 49.525 202.510 49.815 202.555 ;
        RECT 47.455 202.325 47.855 202.510 ;
        RECT 47.715 202.170 47.855 202.325 ;
        RECT 48.130 202.370 49.815 202.510 ;
        RECT 48.130 202.310 48.450 202.370 ;
        RECT 49.525 202.325 49.815 202.370 ;
        RECT 50.445 202.510 50.735 202.555 ;
        RECT 57.330 202.510 57.650 202.570 ;
        RECT 60.565 202.510 60.855 202.555 ;
        RECT 63.785 202.510 64.075 202.555 ;
        RECT 50.445 202.370 53.420 202.510 ;
        RECT 50.445 202.325 50.735 202.370 ;
        RECT 50.520 202.170 50.660 202.325 ;
        RECT 47.715 202.030 50.660 202.170 ;
        RECT 52.185 201.985 52.475 202.215 ;
        RECT 53.280 202.170 53.420 202.370 ;
        RECT 57.330 202.370 60.855 202.510 ;
        RECT 57.330 202.310 57.650 202.370 ;
        RECT 60.565 202.325 60.855 202.370 ;
        RECT 61.100 202.370 64.075 202.510 ;
        RECT 61.100 202.170 61.240 202.370 ;
        RECT 63.785 202.325 64.075 202.370 ;
        RECT 64.245 202.510 64.535 202.555 ;
        RECT 64.690 202.510 65.010 202.570 ;
        RECT 64.245 202.370 65.010 202.510 ;
        RECT 64.245 202.325 64.535 202.370 ;
        RECT 64.690 202.310 65.010 202.370 ;
        RECT 65.165 202.325 65.455 202.555 ;
        RECT 65.700 202.510 65.840 203.050 ;
        RECT 66.990 202.990 67.310 203.250 ;
        RECT 67.950 203.190 68.240 203.235 ;
        RECT 70.050 203.190 70.340 203.235 ;
        RECT 71.620 203.190 71.910 203.235 ;
        RECT 84.010 203.190 84.330 203.250 ;
        RECT 67.950 203.050 71.910 203.190 ;
        RECT 67.950 203.005 68.240 203.050 ;
        RECT 70.050 203.005 70.340 203.050 ;
        RECT 71.620 203.005 71.910 203.050 ;
        RECT 72.600 203.050 84.330 203.190 ;
        RECT 86.860 203.190 87.000 203.390 ;
        RECT 98.270 203.390 101.795 203.530 ;
        RECT 98.270 203.330 98.590 203.390 ;
        RECT 101.505 203.345 101.795 203.390 ;
        RECT 112.990 203.330 113.310 203.590 ;
        RECT 116.225 203.530 116.515 203.575 ;
        RECT 121.270 203.530 121.590 203.590 ;
        RECT 125.425 203.530 125.715 203.575 ;
        RECT 140.130 203.530 140.450 203.590 ;
        RECT 141.525 203.530 141.815 203.575 ;
        RECT 150.340 203.530 150.480 204.410 ;
        RECT 116.225 203.390 125.715 203.530 ;
        RECT 116.225 203.345 116.515 203.390 ;
        RECT 121.270 203.330 121.590 203.390 ;
        RECT 125.425 203.345 125.715 203.390 ;
        RECT 125.960 203.390 139.440 203.530 ;
        RECT 86.860 203.050 89.760 203.190 ;
        RECT 67.080 202.850 67.220 202.990 ;
        RECT 68.345 202.850 68.635 202.895 ;
        RECT 69.535 202.850 69.825 202.895 ;
        RECT 72.055 202.850 72.345 202.895 ;
        RECT 67.080 202.710 68.140 202.850 ;
        RECT 66.085 202.510 66.375 202.555 ;
        RECT 65.700 202.370 66.375 202.510 ;
        RECT 66.085 202.325 66.375 202.370 ;
        RECT 67.005 202.325 67.295 202.555 ;
        RECT 65.240 202.170 65.380 202.325 ;
        RECT 66.545 202.170 66.835 202.215 ;
        RECT 53.280 202.030 61.240 202.170 ;
        RECT 62.480 202.030 64.920 202.170 ;
        RECT 65.240 202.030 66.835 202.170 ;
        RECT 48.130 201.830 48.450 201.890 ;
        RECT 45.000 201.690 48.450 201.830 ;
        RECT 48.130 201.630 48.450 201.690 ;
        RECT 48.605 201.830 48.895 201.875 ;
        RECT 52.260 201.830 52.400 201.985 ;
        RECT 53.280 201.890 53.420 202.030 ;
        RECT 48.605 201.690 52.400 201.830 ;
        RECT 48.605 201.645 48.895 201.690 ;
        RECT 53.190 201.630 53.510 201.890 ;
        RECT 57.790 201.630 58.110 201.890 ;
        RECT 62.480 201.875 62.620 202.030 ;
        RECT 62.405 201.645 62.695 201.875 ;
        RECT 64.780 201.830 64.920 202.030 ;
        RECT 66.545 201.985 66.835 202.030 ;
        RECT 67.080 201.830 67.220 202.325 ;
        RECT 67.450 202.310 67.770 202.570 ;
        RECT 68.000 202.510 68.140 202.710 ;
        RECT 68.345 202.710 72.345 202.850 ;
        RECT 68.345 202.665 68.635 202.710 ;
        RECT 69.535 202.665 69.825 202.710 ;
        RECT 72.055 202.665 72.345 202.710 ;
        RECT 72.600 202.510 72.740 203.050 ;
        RECT 84.010 202.990 84.330 203.050 ;
        RECT 81.265 202.850 81.555 202.895 ;
        RECT 86.325 202.850 86.615 202.895 ;
        RECT 81.265 202.710 86.615 202.850 ;
        RECT 81.265 202.665 81.555 202.710 ;
        RECT 86.325 202.665 86.615 202.710 ;
        RECT 86.770 202.650 87.090 202.910 ;
        RECT 87.690 202.650 88.010 202.910 ;
        RECT 89.620 202.895 89.760 203.050 ;
        RECT 97.810 202.990 98.130 203.250 ;
        RECT 100.200 203.050 104.480 203.190 ;
        RECT 88.625 202.850 88.915 202.895 ;
        RECT 88.625 202.710 89.300 202.850 ;
        RECT 88.625 202.665 88.915 202.710 ;
        RECT 68.000 202.370 72.740 202.510 ;
        RECT 80.345 202.325 80.635 202.555 ;
        RECT 81.725 202.510 82.015 202.555 ;
        RECT 82.630 202.510 82.950 202.570 ;
        RECT 81.725 202.370 82.950 202.510 ;
        RECT 86.860 202.510 87.000 202.650 ;
        RECT 87.245 202.510 87.535 202.555 ;
        RECT 86.860 202.370 87.535 202.510 ;
        RECT 81.725 202.325 82.015 202.370 ;
        RECT 64.780 201.690 67.220 201.830 ;
        RECT 67.540 201.830 67.680 202.310 ;
        RECT 68.800 202.170 69.090 202.215 ;
        RECT 70.670 202.170 70.990 202.230 ;
        RECT 68.800 202.030 70.990 202.170 ;
        RECT 80.420 202.170 80.560 202.325 ;
        RECT 82.630 202.310 82.950 202.370 ;
        RECT 87.245 202.325 87.535 202.370 ;
        RECT 88.165 202.325 88.455 202.555 ;
        RECT 89.160 202.510 89.300 202.710 ;
        RECT 89.545 202.665 89.835 202.895 ;
        RECT 92.750 202.850 93.070 202.910 ;
        RECT 100.200 202.895 100.340 203.050 ;
        RECT 99.665 202.850 99.955 202.895 ;
        RECT 92.750 202.710 99.955 202.850 ;
        RECT 92.750 202.650 93.070 202.710 ;
        RECT 99.665 202.665 99.955 202.710 ;
        RECT 100.125 202.665 100.415 202.895 ;
        RECT 102.410 202.650 102.730 202.910 ;
        RECT 104.340 202.895 104.480 203.050 ;
        RECT 104.265 202.850 104.555 202.895 ;
        RECT 113.080 202.850 113.220 203.330 ;
        RECT 115.290 203.190 115.610 203.250 ;
        RECT 125.960 203.190 126.100 203.390 ;
        RECT 131.405 203.190 131.695 203.235 ;
        RECT 115.290 203.050 126.100 203.190 ;
        RECT 131.020 203.050 131.695 203.190 ;
        RECT 115.290 202.990 115.610 203.050 ;
        RECT 123.570 202.850 123.890 202.910 ;
        RECT 104.265 202.710 105.400 202.850 ;
        RECT 113.080 202.710 123.890 202.850 ;
        RECT 104.265 202.665 104.555 202.710 ;
        RECT 105.260 202.570 105.400 202.710 ;
        RECT 123.570 202.650 123.890 202.710 ;
        RECT 124.950 202.850 125.270 202.910 ;
        RECT 127.250 202.850 127.570 202.910 ;
        RECT 131.020 202.895 131.160 203.050 ;
        RECT 131.405 203.005 131.695 203.050 ;
        RECT 134.650 203.190 134.940 203.235 ;
        RECT 136.750 203.190 137.040 203.235 ;
        RECT 138.320 203.190 138.610 203.235 ;
        RECT 134.650 203.050 138.610 203.190 ;
        RECT 134.650 203.005 134.940 203.050 ;
        RECT 136.750 203.005 137.040 203.050 ;
        RECT 138.320 203.005 138.610 203.050 ;
        RECT 130.945 202.850 131.235 202.895 ;
        RECT 124.950 202.710 131.235 202.850 ;
        RECT 124.950 202.650 125.270 202.710 ;
        RECT 127.250 202.650 127.570 202.710 ;
        RECT 130.945 202.665 131.235 202.710 ;
        RECT 135.045 202.850 135.335 202.895 ;
        RECT 136.235 202.850 136.525 202.895 ;
        RECT 138.755 202.850 139.045 202.895 ;
        RECT 135.045 202.710 139.045 202.850 ;
        RECT 135.045 202.665 135.335 202.710 ;
        RECT 136.235 202.665 136.525 202.710 ;
        RECT 138.755 202.665 139.045 202.710 ;
        RECT 89.990 202.510 90.310 202.570 ;
        RECT 89.160 202.370 90.310 202.510 ;
        RECT 88.240 202.170 88.380 202.325 ;
        RECT 89.990 202.310 90.310 202.370 ;
        RECT 90.465 202.510 90.755 202.555 ;
        RECT 90.910 202.510 91.230 202.570 ;
        RECT 90.465 202.370 91.230 202.510 ;
        RECT 90.465 202.325 90.755 202.370 ;
        RECT 90.910 202.310 91.230 202.370 ;
        RECT 91.370 202.310 91.690 202.570 ;
        RECT 91.830 202.310 92.150 202.570 ;
        RECT 98.730 202.510 99.050 202.570 ;
        RECT 95.600 202.370 99.050 202.510 ;
        RECT 89.530 202.170 89.850 202.230 ;
        RECT 95.600 202.170 95.740 202.370 ;
        RECT 98.730 202.310 99.050 202.370 ;
        RECT 102.870 202.310 103.190 202.570 ;
        RECT 104.710 202.310 105.030 202.570 ;
        RECT 105.170 202.310 105.490 202.570 ;
        RECT 105.630 202.310 105.950 202.570 ;
        RECT 115.305 202.325 115.595 202.555 ;
        RECT 116.685 202.510 116.975 202.555 ;
        RECT 119.430 202.510 119.750 202.570 ;
        RECT 116.685 202.370 119.750 202.510 ;
        RECT 116.685 202.325 116.975 202.370 ;
        RECT 115.380 202.170 115.520 202.325 ;
        RECT 119.430 202.310 119.750 202.370 ;
        RECT 124.505 202.325 124.795 202.555 ;
        RECT 125.885 202.510 126.175 202.555 ;
        RECT 125.885 202.370 129.320 202.510 ;
        RECT 125.885 202.325 126.175 202.370 ;
        RECT 117.590 202.170 117.910 202.230 ;
        RECT 124.580 202.170 124.720 202.325 ;
        RECT 80.420 202.030 81.710 202.170 ;
        RECT 88.240 202.030 89.850 202.170 ;
        RECT 68.800 201.985 69.090 202.030 ;
        RECT 70.670 201.970 70.990 202.030 ;
        RECT 69.750 201.830 70.070 201.890 ;
        RECT 67.540 201.690 70.070 201.830 ;
        RECT 69.750 201.630 70.070 201.690 ;
        RECT 74.350 201.830 74.670 201.890 ;
        RECT 80.790 201.830 81.110 201.890 ;
        RECT 74.350 201.690 81.110 201.830 ;
        RECT 81.570 201.830 81.710 202.030 ;
        RECT 89.530 201.970 89.850 202.030 ;
        RECT 90.080 202.030 95.740 202.170 ;
        RECT 97.440 202.030 106.780 202.170 ;
        RECT 115.380 202.030 124.720 202.170 ;
        RECT 84.470 201.830 84.790 201.890 ;
        RECT 90.080 201.830 90.220 202.030 ;
        RECT 81.570 201.690 90.220 201.830 ;
        RECT 93.210 201.830 93.530 201.890 ;
        RECT 97.440 201.830 97.580 202.030 ;
        RECT 106.640 201.890 106.780 202.030 ;
        RECT 117.590 201.970 117.910 202.030 ;
        RECT 93.210 201.690 97.580 201.830 ;
        RECT 74.350 201.630 74.670 201.690 ;
        RECT 80.790 201.630 81.110 201.690 ;
        RECT 84.470 201.630 84.790 201.690 ;
        RECT 93.210 201.630 93.530 201.690 ;
        RECT 106.550 201.630 106.870 201.890 ;
        RECT 114.385 201.830 114.675 201.875 ;
        RECT 119.890 201.830 120.210 201.890 ;
        RECT 114.385 201.690 120.210 201.830 ;
        RECT 114.385 201.645 114.675 201.690 ;
        RECT 119.890 201.630 120.210 201.690 ;
        RECT 123.585 201.830 123.875 201.875 ;
        RECT 127.250 201.830 127.570 201.890 ;
        RECT 123.585 201.690 127.570 201.830 ;
        RECT 129.180 201.830 129.320 202.370 ;
        RECT 129.565 202.325 129.855 202.555 ;
        RECT 132.310 202.510 132.630 202.570 ;
        RECT 134.165 202.510 134.455 202.555 ;
        RECT 134.610 202.510 134.930 202.570 ;
        RECT 135.530 202.555 135.850 202.570 ;
        RECT 135.500 202.510 135.850 202.555 ;
        RECT 132.310 202.370 133.460 202.510 ;
        RECT 129.640 202.170 129.780 202.325 ;
        RECT 132.310 202.310 132.630 202.370 ;
        RECT 133.320 202.230 133.460 202.370 ;
        RECT 134.165 202.370 134.930 202.510 ;
        RECT 135.335 202.370 135.850 202.510 ;
        RECT 139.300 202.510 139.440 203.390 ;
        RECT 140.130 203.390 141.815 203.530 ;
        RECT 140.130 203.330 140.450 203.390 ;
        RECT 141.525 203.345 141.815 203.390 ;
        RECT 148.040 203.390 150.480 203.530 ;
        RECT 141.050 202.850 141.370 202.910 ;
        RECT 144.285 202.850 144.575 202.895 ;
        RECT 141.050 202.710 144.575 202.850 ;
        RECT 141.050 202.650 141.370 202.710 ;
        RECT 144.285 202.665 144.575 202.710 ;
        RECT 143.825 202.510 144.115 202.555 ;
        RECT 148.040 202.510 148.180 203.390 ;
        RECT 149.790 202.850 150.110 202.910 ;
        RECT 148.500 202.710 150.110 202.850 ;
        RECT 148.500 202.555 148.640 202.710 ;
        RECT 149.790 202.650 150.110 202.710 ;
        RECT 139.300 202.370 148.180 202.510 ;
        RECT 134.165 202.325 134.455 202.370 ;
        RECT 134.610 202.310 134.930 202.370 ;
        RECT 135.500 202.325 135.850 202.370 ;
        RECT 143.825 202.325 144.115 202.370 ;
        RECT 148.425 202.325 148.715 202.555 ;
        RECT 135.530 202.310 135.850 202.325 ;
        RECT 132.770 202.170 133.090 202.230 ;
        RECT 129.640 202.030 133.090 202.170 ;
        RECT 132.770 201.970 133.090 202.030 ;
        RECT 133.230 201.970 133.550 202.230 ;
        RECT 143.365 202.170 143.655 202.215 ;
        RECT 144.270 202.170 144.590 202.230 ;
        RECT 143.365 202.030 144.590 202.170 ;
        RECT 143.365 201.985 143.655 202.030 ;
        RECT 144.270 201.970 144.590 202.030 ;
        RECT 134.150 201.830 134.470 201.890 ;
        RECT 129.180 201.690 134.470 201.830 ;
        RECT 123.585 201.645 123.875 201.690 ;
        RECT 127.250 201.630 127.570 201.690 ;
        RECT 134.150 201.630 134.470 201.690 ;
        RECT 136.910 201.830 137.230 201.890 ;
        RECT 141.065 201.830 141.355 201.875 ;
        RECT 136.910 201.690 141.355 201.830 ;
        RECT 136.910 201.630 137.230 201.690 ;
        RECT 141.065 201.645 141.355 201.690 ;
        RECT 147.490 201.630 147.810 201.890 ;
        RECT 36.100 201.010 150.180 201.490 ;
        RECT 41.690 200.810 42.010 200.870 ;
        RECT 43.545 200.810 43.835 200.855 ;
        RECT 57.330 200.810 57.650 200.870 ;
        RECT 60.090 200.810 60.410 200.870 ;
        RECT 41.690 200.670 43.835 200.810 ;
        RECT 41.690 200.610 42.010 200.670 ;
        RECT 43.545 200.625 43.835 200.670 ;
        RECT 45.000 200.670 50.200 200.810 ;
        RECT 41.230 200.270 41.550 200.530 ;
        RECT 42.610 200.270 42.930 200.530 ;
        RECT 41.320 200.130 41.460 200.270 ;
        RECT 41.705 200.130 41.995 200.175 ;
        RECT 41.320 199.990 41.995 200.130 ;
        RECT 41.705 199.945 41.995 199.990 ;
        RECT 43.070 200.130 43.390 200.190 ;
        RECT 45.000 200.175 45.140 200.670 ;
        RECT 45.370 200.470 45.690 200.530 ;
        RECT 47.225 200.470 47.515 200.515 ;
        RECT 45.370 200.330 47.515 200.470 ;
        RECT 45.370 200.270 45.690 200.330 ;
        RECT 47.225 200.285 47.515 200.330 ;
        RECT 50.060 200.470 50.200 200.670 ;
        RECT 57.330 200.670 60.410 200.810 ;
        RECT 57.330 200.610 57.650 200.670 ;
        RECT 60.090 200.610 60.410 200.670 ;
        RECT 70.670 200.610 70.990 200.870 ;
        RECT 91.370 200.810 91.690 200.870 ;
        RECT 94.145 200.810 94.435 200.855 ;
        RECT 71.220 200.670 88.840 200.810 ;
        RECT 71.220 200.470 71.360 200.670 ;
        RECT 87.690 200.470 88.010 200.530 ;
        RECT 50.060 200.330 71.360 200.470 ;
        RECT 85.940 200.330 88.010 200.470 ;
        RECT 88.700 200.470 88.840 200.670 ;
        RECT 91.370 200.670 94.435 200.810 ;
        RECT 91.370 200.610 91.690 200.670 ;
        RECT 94.145 200.625 94.435 200.670 ;
        RECT 102.410 200.610 102.730 200.870 ;
        RECT 103.345 200.810 103.635 200.855 ;
        RECT 104.710 200.810 105.030 200.870 ;
        RECT 103.345 200.670 105.030 200.810 ;
        RECT 103.345 200.625 103.635 200.670 ;
        RECT 104.710 200.610 105.030 200.670 ;
        RECT 112.070 200.610 112.390 200.870 ;
        RECT 120.350 200.610 120.670 200.870 ;
        RECT 102.500 200.470 102.640 200.610 ;
        RECT 88.700 200.330 95.740 200.470 ;
        RECT 44.925 200.130 45.215 200.175 ;
        RECT 43.070 199.990 45.215 200.130 ;
        RECT 41.780 199.790 41.920 199.945 ;
        RECT 43.070 199.930 43.390 199.990 ;
        RECT 44.925 199.945 45.215 199.990 ;
        RECT 45.830 199.930 46.150 200.190 ;
        RECT 50.060 200.175 50.200 200.330 ;
        RECT 49.985 199.945 50.275 200.175 ;
        RECT 54.570 200.130 54.890 200.190 ;
        RECT 55.505 200.130 55.795 200.175 ;
        RECT 54.570 199.990 55.795 200.130 ;
        RECT 54.570 199.930 54.890 199.990 ;
        RECT 55.505 199.945 55.795 199.990 ;
        RECT 56.410 200.130 56.730 200.190 ;
        RECT 57.345 200.130 57.635 200.175 ;
        RECT 56.410 199.990 57.635 200.130 ;
        RECT 43.530 199.790 43.850 199.850 ;
        RECT 41.780 199.650 43.850 199.790 ;
        RECT 43.530 199.590 43.850 199.650 ;
        RECT 44.465 199.605 44.755 199.835 ;
        RECT 45.385 199.605 45.675 199.835 ;
        RECT 46.290 199.790 46.610 199.850 ;
        RECT 48.605 199.790 48.895 199.835 ;
        RECT 55.580 199.790 55.720 199.945 ;
        RECT 56.410 199.930 56.730 199.990 ;
        RECT 57.345 199.945 57.635 199.990 ;
        RECT 57.790 200.130 58.110 200.190 ;
        RECT 59.185 200.130 59.475 200.175 ;
        RECT 57.790 199.990 59.475 200.130 ;
        RECT 57.790 199.930 58.110 199.990 ;
        RECT 59.185 199.945 59.475 199.990 ;
        RECT 60.090 199.930 60.410 200.190 ;
        RECT 60.565 200.130 60.855 200.175 ;
        RECT 62.850 200.130 63.170 200.190 ;
        RECT 60.565 199.990 63.170 200.130 ;
        RECT 60.565 199.945 60.855 199.990 ;
        RECT 62.850 199.930 63.170 199.990 ;
        RECT 71.605 200.130 71.895 200.175 ;
        RECT 72.510 200.130 72.830 200.190 ;
        RECT 71.605 199.990 72.830 200.130 ;
        RECT 71.605 199.945 71.895 199.990 ;
        RECT 72.510 199.930 72.830 199.990 ;
        RECT 73.400 200.130 73.690 200.175 ;
        RECT 75.730 200.130 76.050 200.190 ;
        RECT 73.400 199.990 76.050 200.130 ;
        RECT 73.400 199.945 73.690 199.990 ;
        RECT 75.730 199.930 76.050 199.990 ;
        RECT 81.725 200.130 82.015 200.175 ;
        RECT 84.470 200.130 84.790 200.190 ;
        RECT 81.725 199.990 84.790 200.130 ;
        RECT 81.725 199.945 82.015 199.990 ;
        RECT 84.470 199.930 84.790 199.990 ;
        RECT 56.870 199.790 57.190 199.850 ;
        RECT 46.290 199.650 52.400 199.790 ;
        RECT 55.580 199.650 57.190 199.790 ;
        RECT 60.180 199.790 60.320 199.930 ;
        RECT 62.405 199.790 62.695 199.835 ;
        RECT 60.180 199.650 62.695 199.790 ;
        RECT 38.930 199.250 39.250 199.510 ;
        RECT 42.150 199.250 42.470 199.510 ;
        RECT 44.540 199.450 44.680 199.605 ;
        RECT 44.910 199.450 45.230 199.510 ;
        RECT 44.540 199.310 45.230 199.450 ;
        RECT 45.460 199.450 45.600 199.605 ;
        RECT 46.290 199.590 46.610 199.650 ;
        RECT 48.605 199.605 48.895 199.650 ;
        RECT 52.260 199.450 52.400 199.650 ;
        RECT 56.870 199.590 57.190 199.650 ;
        RECT 62.405 199.605 62.695 199.650 ;
        RECT 63.785 199.605 64.075 199.835 ;
        RECT 69.750 199.790 70.070 199.850 ;
        RECT 72.065 199.790 72.355 199.835 ;
        RECT 69.750 199.650 72.355 199.790 ;
        RECT 58.710 199.450 59.030 199.510 ;
        RECT 59.645 199.450 59.935 199.495 ;
        RECT 45.460 199.310 51.120 199.450 ;
        RECT 52.260 199.310 58.020 199.450 ;
        RECT 44.910 199.250 45.230 199.310 ;
        RECT 39.020 199.110 39.160 199.250 ;
        RECT 50.980 199.170 51.120 199.310 ;
        RECT 45.370 199.110 45.690 199.170 ;
        RECT 39.020 198.970 45.690 199.110 ;
        RECT 45.370 198.910 45.690 198.970 ;
        RECT 47.685 199.110 47.975 199.155 ;
        RECT 48.130 199.110 48.450 199.170 ;
        RECT 47.685 198.970 48.450 199.110 ;
        RECT 47.685 198.925 47.975 198.970 ;
        RECT 48.130 198.910 48.450 198.970 ;
        RECT 50.890 198.910 51.210 199.170 ;
        RECT 54.110 199.110 54.430 199.170 ;
        RECT 56.410 199.110 56.730 199.170 ;
        RECT 54.110 198.970 56.730 199.110 ;
        RECT 57.880 199.110 58.020 199.310 ;
        RECT 58.710 199.310 59.935 199.450 ;
        RECT 58.710 199.250 59.030 199.310 ;
        RECT 59.645 199.265 59.935 199.310 ;
        RECT 60.105 199.450 60.395 199.495 ;
        RECT 63.310 199.450 63.630 199.510 ;
        RECT 63.860 199.450 64.000 199.605 ;
        RECT 69.750 199.590 70.070 199.650 ;
        RECT 72.065 199.605 72.355 199.650 ;
        RECT 72.945 199.790 73.235 199.835 ;
        RECT 74.135 199.790 74.425 199.835 ;
        RECT 76.655 199.790 76.945 199.835 ;
        RECT 72.945 199.650 76.945 199.790 ;
        RECT 72.945 199.605 73.235 199.650 ;
        RECT 74.135 199.605 74.425 199.650 ;
        RECT 76.655 199.605 76.945 199.650 ;
        RECT 77.110 199.790 77.430 199.850 ;
        RECT 80.805 199.790 81.095 199.835 ;
        RECT 77.110 199.650 81.095 199.790 ;
        RECT 77.110 199.590 77.430 199.650 ;
        RECT 80.805 199.605 81.095 199.650 ;
        RECT 82.170 199.790 82.490 199.850 ;
        RECT 83.105 199.790 83.395 199.835 ;
        RECT 82.170 199.650 83.395 199.790 ;
        RECT 82.170 199.590 82.490 199.650 ;
        RECT 83.105 199.605 83.395 199.650 ;
        RECT 84.010 199.790 84.330 199.850 ;
        RECT 85.940 199.790 86.080 200.330 ;
        RECT 87.690 200.270 88.010 200.330 ;
        RECT 86.325 200.130 86.615 200.175 ;
        RECT 86.325 199.990 87.000 200.130 ;
        RECT 86.325 199.945 86.615 199.990 ;
        RECT 86.860 199.850 87.000 199.990 ;
        RECT 87.245 199.945 87.535 200.175 ;
        RECT 87.780 200.130 87.920 200.270 ;
        RECT 95.600 200.175 95.740 200.330 ;
        RECT 100.200 200.330 102.640 200.470 ;
        RECT 88.125 200.130 88.415 200.175 ;
        RECT 87.780 199.990 88.415 200.130 ;
        RECT 88.125 199.945 88.415 199.990 ;
        RECT 90.465 200.130 90.755 200.175 ;
        RECT 95.065 200.130 95.355 200.175 ;
        RECT 90.465 199.990 95.355 200.130 ;
        RECT 90.465 199.945 90.755 199.990 ;
        RECT 84.010 199.650 86.080 199.790 ;
        RECT 84.010 199.590 84.330 199.650 ;
        RECT 86.770 199.590 87.090 199.850 ;
        RECT 87.320 199.790 87.460 199.945 ;
        RECT 90.910 199.790 91.230 199.850 ;
        RECT 87.320 199.650 91.230 199.790 ;
        RECT 90.910 199.590 91.230 199.650 ;
        RECT 60.105 199.310 64.000 199.450 ;
        RECT 60.105 199.265 60.395 199.310 ;
        RECT 63.310 199.250 63.630 199.310 ;
        RECT 58.265 199.110 58.555 199.155 ;
        RECT 60.550 199.110 60.870 199.170 ;
        RECT 57.880 198.970 60.870 199.110 ;
        RECT 54.110 198.910 54.430 198.970 ;
        RECT 56.410 198.910 56.730 198.970 ;
        RECT 58.265 198.925 58.555 198.970 ;
        RECT 60.550 198.910 60.870 198.970 ;
        RECT 61.470 198.910 61.790 199.170 ;
        RECT 63.860 199.110 64.000 199.310 ;
        RECT 72.550 199.450 72.840 199.495 ;
        RECT 74.650 199.450 74.940 199.495 ;
        RECT 76.220 199.450 76.510 199.495 ;
        RECT 72.550 199.310 76.510 199.450 ;
        RECT 72.550 199.265 72.840 199.310 ;
        RECT 74.650 199.265 74.940 199.310 ;
        RECT 76.220 199.265 76.510 199.310 ;
        RECT 79.870 199.450 80.190 199.510 ;
        RECT 82.645 199.450 82.935 199.495 ;
        RECT 87.690 199.450 88.010 199.510 ;
        RECT 79.870 199.310 81.020 199.450 ;
        RECT 79.870 199.250 80.190 199.310 ;
        RECT 66.530 199.110 66.850 199.170 ;
        RECT 72.970 199.110 73.290 199.170 ;
        RECT 63.860 198.970 73.290 199.110 ;
        RECT 66.530 198.910 66.850 198.970 ;
        RECT 72.970 198.910 73.290 198.970 ;
        RECT 78.965 199.110 79.255 199.155 ;
        RECT 80.330 199.110 80.650 199.170 ;
        RECT 78.965 198.970 80.650 199.110 ;
        RECT 80.880 199.110 81.020 199.310 ;
        RECT 82.645 199.310 88.010 199.450 ;
        RECT 82.645 199.265 82.935 199.310 ;
        RECT 87.690 199.250 88.010 199.310 ;
        RECT 89.085 199.450 89.375 199.495 ;
        RECT 90.450 199.450 90.770 199.510 ;
        RECT 91.460 199.450 91.600 199.990 ;
        RECT 95.065 199.945 95.355 199.990 ;
        RECT 95.525 199.945 95.815 200.175 ;
        RECT 95.985 200.130 96.275 200.175 ;
        RECT 95.985 199.990 97.580 200.130 ;
        RECT 95.985 199.945 96.275 199.990 ;
        RECT 97.440 199.850 97.580 199.990 ;
        RECT 98.270 199.930 98.590 200.190 ;
        RECT 96.430 199.590 96.750 199.850 ;
        RECT 97.350 199.590 97.670 199.850 ;
        RECT 100.200 199.835 100.340 200.330 ;
        RECT 100.585 199.945 100.875 200.175 ;
        RECT 101.505 199.945 101.795 200.175 ;
        RECT 97.825 199.605 98.115 199.835 ;
        RECT 100.125 199.605 100.415 199.835 ;
        RECT 89.085 199.310 91.600 199.450 ;
        RECT 94.130 199.450 94.450 199.510 ;
        RECT 97.900 199.450 98.040 199.605 ;
        RECT 94.130 199.310 98.040 199.450 ;
        RECT 98.730 199.450 99.050 199.510 ;
        RECT 100.660 199.450 100.800 199.945 ;
        RECT 98.730 199.310 100.800 199.450 ;
        RECT 89.085 199.265 89.375 199.310 ;
        RECT 90.450 199.250 90.770 199.310 ;
        RECT 94.130 199.250 94.450 199.310 ;
        RECT 98.730 199.250 99.050 199.310 ;
        RECT 86.310 199.110 86.630 199.170 ;
        RECT 80.880 198.970 86.630 199.110 ;
        RECT 78.965 198.925 79.255 198.970 ;
        RECT 80.330 198.910 80.650 198.970 ;
        RECT 86.310 198.910 86.630 198.970 ;
        RECT 86.785 199.110 87.075 199.155 ;
        RECT 87.230 199.110 87.550 199.170 ;
        RECT 86.785 198.970 87.550 199.110 ;
        RECT 86.785 198.925 87.075 198.970 ;
        RECT 87.230 198.910 87.550 198.970 ;
        RECT 89.530 199.110 89.850 199.170 ;
        RECT 90.005 199.110 90.295 199.155 ;
        RECT 94.590 199.110 94.910 199.170 ;
        RECT 89.530 198.970 94.910 199.110 ;
        RECT 89.530 198.910 89.850 198.970 ;
        RECT 90.005 198.925 90.295 198.970 ;
        RECT 94.590 198.910 94.910 198.970 ;
        RECT 99.650 199.110 99.970 199.170 ;
        RECT 101.580 199.110 101.720 199.945 ;
        RECT 101.950 199.930 102.270 200.190 ;
        RECT 102.500 200.175 102.640 200.330 ;
        RECT 103.790 200.470 104.110 200.530 ;
        RECT 107.010 200.470 107.330 200.530 ;
        RECT 112.160 200.470 112.300 200.610 ;
        RECT 103.790 200.330 112.300 200.470 ;
        RECT 112.990 200.470 113.310 200.530 ;
        RECT 119.490 200.470 119.780 200.515 ;
        RECT 112.990 200.330 119.780 200.470 ;
        RECT 103.790 200.270 104.110 200.330 ;
        RECT 107.010 200.270 107.330 200.330 ;
        RECT 112.990 200.270 113.310 200.330 ;
        RECT 119.490 200.285 119.780 200.330 ;
        RECT 120.440 200.470 120.580 200.610 ;
        RECT 128.630 200.470 128.950 200.530 ;
        RECT 134.610 200.470 134.930 200.530 ;
        RECT 120.440 200.330 134.930 200.470 ;
        RECT 102.500 199.990 102.835 200.175 ;
        RECT 102.545 199.945 102.835 199.990 ;
        RECT 112.085 200.130 112.375 200.175 ;
        RECT 114.370 200.130 114.690 200.190 ;
        RECT 112.085 199.990 114.690 200.130 ;
        RECT 120.440 200.130 120.580 200.330 ;
        RECT 128.630 200.270 128.950 200.330 ;
        RECT 120.825 200.130 121.115 200.175 ;
        RECT 120.440 199.990 121.115 200.130 ;
        RECT 112.085 199.945 112.375 199.990 ;
        RECT 114.370 199.930 114.690 199.990 ;
        RECT 120.825 199.945 121.115 199.990 ;
        RECT 124.950 199.930 125.270 200.190 ;
        RECT 125.410 199.930 125.730 200.190 ;
        RECT 126.345 199.945 126.635 200.175 ;
        RECT 126.790 200.130 127.110 200.190 ;
        RECT 133.780 200.175 133.920 200.330 ;
        RECT 134.610 200.270 134.930 200.330 ;
        RECT 132.370 200.130 132.660 200.175 ;
        RECT 126.790 199.990 132.660 200.130 ;
        RECT 116.235 199.790 116.525 199.835 ;
        RECT 118.755 199.790 119.045 199.835 ;
        RECT 119.945 199.790 120.235 199.835 ;
        RECT 116.235 199.650 120.235 199.790 ;
        RECT 125.040 199.790 125.180 199.930 ;
        RECT 126.420 199.790 126.560 199.945 ;
        RECT 126.790 199.930 127.110 199.990 ;
        RECT 132.370 199.945 132.660 199.990 ;
        RECT 133.705 199.945 133.995 200.175 ;
        RECT 127.250 199.790 127.570 199.850 ;
        RECT 125.040 199.650 127.570 199.790 ;
        RECT 116.235 199.605 116.525 199.650 ;
        RECT 118.755 199.605 119.045 199.650 ;
        RECT 119.945 199.605 120.235 199.650 ;
        RECT 127.250 199.590 127.570 199.650 ;
        RECT 129.115 199.790 129.405 199.835 ;
        RECT 131.635 199.790 131.925 199.835 ;
        RECT 132.825 199.790 133.115 199.835 ;
        RECT 129.115 199.650 133.115 199.790 ;
        RECT 129.115 199.605 129.405 199.650 ;
        RECT 131.635 199.605 131.925 199.650 ;
        RECT 132.825 199.605 133.115 199.650 ;
        RECT 116.670 199.450 116.960 199.495 ;
        RECT 118.240 199.450 118.530 199.495 ;
        RECT 120.340 199.450 120.630 199.495 ;
        RECT 116.670 199.310 120.630 199.450 ;
        RECT 116.670 199.265 116.960 199.310 ;
        RECT 118.240 199.265 118.530 199.310 ;
        RECT 120.340 199.265 120.630 199.310 ;
        RECT 121.270 199.450 121.590 199.510 ;
        RECT 129.550 199.450 129.840 199.495 ;
        RECT 131.120 199.450 131.410 199.495 ;
        RECT 133.220 199.450 133.510 199.495 ;
        RECT 121.270 199.310 127.480 199.450 ;
        RECT 121.270 199.250 121.590 199.310 ;
        RECT 99.650 198.970 101.720 199.110 ;
        RECT 102.410 199.110 102.730 199.170 ;
        RECT 108.850 199.110 109.170 199.170 ;
        RECT 102.410 198.970 109.170 199.110 ;
        RECT 99.650 198.910 99.970 198.970 ;
        RECT 102.410 198.910 102.730 198.970 ;
        RECT 108.850 198.910 109.170 198.970 ;
        RECT 112.990 198.910 113.310 199.170 ;
        RECT 113.910 198.910 114.230 199.170 ;
        RECT 125.870 198.910 126.190 199.170 ;
        RECT 126.330 199.110 126.650 199.170 ;
        RECT 126.805 199.110 127.095 199.155 ;
        RECT 126.330 198.970 127.095 199.110 ;
        RECT 127.340 199.110 127.480 199.310 ;
        RECT 129.550 199.310 133.510 199.450 ;
        RECT 129.550 199.265 129.840 199.310 ;
        RECT 131.120 199.265 131.410 199.310 ;
        RECT 133.220 199.265 133.510 199.310 ;
        RECT 144.730 199.110 145.050 199.170 ;
        RECT 127.340 198.970 145.050 199.110 ;
        RECT 126.330 198.910 126.650 198.970 ;
        RECT 126.805 198.925 127.095 198.970 ;
        RECT 144.730 198.910 145.050 198.970 ;
        RECT 36.100 198.290 150.180 198.770 ;
        RECT 43.530 198.090 43.850 198.150 ;
        RECT 44.005 198.090 44.295 198.135 ;
        RECT 43.530 197.950 44.295 198.090 ;
        RECT 43.530 197.890 43.850 197.950 ;
        RECT 44.005 197.905 44.295 197.950 ;
        RECT 45.830 198.090 46.150 198.150 ;
        RECT 56.425 198.090 56.715 198.135 ;
        RECT 58.710 198.090 59.030 198.150 ;
        RECT 45.830 197.950 59.030 198.090 ;
        RECT 45.830 197.890 46.150 197.950 ;
        RECT 56.425 197.905 56.715 197.950 ;
        RECT 43.620 197.410 43.760 197.890 ;
        RECT 54.570 197.750 54.890 197.810 ;
        RECT 55.965 197.750 56.255 197.795 ;
        RECT 54.570 197.610 56.255 197.750 ;
        RECT 54.570 197.550 54.890 197.610 ;
        RECT 55.965 197.565 56.255 197.610 ;
        RECT 41.320 197.270 43.760 197.410 ;
        RECT 56.500 197.410 56.640 197.905 ;
        RECT 58.710 197.890 59.030 197.950 ;
        RECT 59.170 198.090 59.490 198.150 ;
        RECT 59.645 198.090 59.935 198.135 ;
        RECT 59.170 197.950 59.935 198.090 ;
        RECT 59.170 197.890 59.490 197.950 ;
        RECT 59.645 197.905 59.935 197.950 ;
        RECT 87.690 198.090 88.010 198.150 ;
        RECT 89.545 198.090 89.835 198.135 ;
        RECT 87.690 197.950 89.835 198.090 ;
        RECT 87.690 197.890 88.010 197.950 ;
        RECT 89.545 197.905 89.835 197.950 ;
        RECT 99.650 198.090 99.970 198.150 ;
        RECT 101.045 198.090 101.335 198.135 ;
        RECT 103.790 198.090 104.110 198.150 ;
        RECT 99.650 197.950 101.335 198.090 ;
        RECT 99.650 197.890 99.970 197.950 ;
        RECT 101.045 197.905 101.335 197.950 ;
        RECT 102.500 197.950 104.110 198.090 ;
        RECT 56.870 197.750 57.190 197.810 ;
        RECT 86.770 197.750 87.090 197.810 ;
        RECT 90.910 197.750 91.230 197.810 ;
        RECT 56.870 197.610 90.220 197.750 ;
        RECT 56.870 197.550 57.190 197.610 ;
        RECT 86.770 197.550 87.090 197.610 ;
        RECT 61.025 197.410 61.315 197.455 ;
        RECT 56.500 197.270 61.315 197.410 ;
        RECT 41.320 197.115 41.460 197.270 ;
        RECT 61.025 197.225 61.315 197.270 ;
        RECT 61.930 197.210 62.250 197.470 ;
        RECT 65.610 197.410 65.930 197.470 ;
        RECT 63.860 197.270 65.930 197.410 ;
        RECT 41.245 196.885 41.535 197.115 ;
        RECT 42.150 196.870 42.470 197.130 ;
        RECT 44.910 197.070 45.230 197.130 ;
        RECT 42.700 196.930 45.230 197.070 ;
        RECT 42.700 196.450 42.840 196.930 ;
        RECT 44.910 196.870 45.230 196.930 ;
        RECT 45.845 197.070 46.135 197.115 ;
        RECT 49.510 197.070 49.830 197.130 ;
        RECT 45.845 196.930 49.830 197.070 ;
        RECT 45.845 196.885 46.135 196.930 ;
        RECT 49.510 196.870 49.830 196.930 ;
        RECT 50.890 196.870 51.210 197.130 ;
        RECT 54.570 197.070 54.890 197.130 ;
        RECT 55.045 197.070 55.335 197.115 ;
        RECT 54.570 196.930 55.335 197.070 ;
        RECT 54.570 196.870 54.890 196.930 ;
        RECT 55.045 196.885 55.335 196.930 ;
        RECT 56.870 196.870 57.190 197.130 ;
        RECT 57.345 196.885 57.635 197.115 ;
        RECT 58.725 197.070 59.015 197.115 ;
        RECT 58.725 196.930 59.400 197.070 ;
        RECT 58.725 196.885 59.015 196.930 ;
        RECT 50.980 196.730 51.120 196.870 ;
        RECT 56.960 196.730 57.100 196.870 ;
        RECT 50.980 196.590 57.100 196.730 ;
        RECT 57.420 196.730 57.560 196.885 ;
        RECT 57.420 196.590 58.940 196.730 ;
        RECT 58.800 196.450 58.940 196.590 ;
        RECT 59.260 196.450 59.400 196.930 ;
        RECT 60.550 196.870 60.870 197.130 ;
        RECT 61.485 197.070 61.775 197.115 ;
        RECT 62.850 197.070 63.170 197.130 ;
        RECT 63.860 197.070 64.000 197.270 ;
        RECT 65.610 197.210 65.930 197.270 ;
        RECT 87.690 197.210 88.010 197.470 ;
        RECT 88.150 197.210 88.470 197.470 ;
        RECT 61.485 196.930 64.000 197.070 ;
        RECT 64.245 197.070 64.535 197.115 ;
        RECT 72.970 197.070 73.290 197.130 ;
        RECT 85.865 197.070 86.155 197.115 ;
        RECT 87.245 197.070 87.535 197.115 ;
        RECT 64.245 196.930 67.680 197.070 ;
        RECT 61.485 196.885 61.775 196.930 ;
        RECT 62.850 196.870 63.170 196.930 ;
        RECT 64.245 196.885 64.535 196.930 ;
        RECT 67.540 196.790 67.680 196.930 ;
        RECT 72.970 196.930 85.620 197.070 ;
        RECT 72.970 196.870 73.290 196.930 ;
        RECT 65.610 196.730 65.930 196.790 ;
        RECT 66.545 196.730 66.835 196.775 ;
        RECT 65.610 196.590 66.835 196.730 ;
        RECT 65.610 196.530 65.930 196.590 ;
        RECT 66.545 196.545 66.835 196.590 ;
        RECT 67.450 196.530 67.770 196.790 ;
        RECT 69.290 196.730 69.610 196.790 ;
        RECT 84.025 196.730 84.315 196.775 ;
        RECT 69.290 196.590 84.315 196.730 ;
        RECT 69.290 196.530 69.610 196.590 ;
        RECT 84.025 196.545 84.315 196.590 ;
        RECT 84.470 196.730 84.790 196.790 ;
        RECT 84.945 196.730 85.235 196.775 ;
        RECT 84.470 196.590 85.235 196.730 ;
        RECT 85.480 196.730 85.620 196.930 ;
        RECT 85.865 196.930 87.535 197.070 ;
        RECT 85.865 196.885 86.155 196.930 ;
        RECT 87.245 196.885 87.535 196.930 ;
        RECT 88.610 196.870 88.930 197.130 ;
        RECT 90.080 197.070 90.220 197.610 ;
        RECT 90.910 197.610 91.600 197.750 ;
        RECT 90.910 197.550 91.230 197.610 ;
        RECT 90.450 197.210 90.770 197.470 ;
        RECT 91.460 197.455 91.600 197.610 ;
        RECT 94.130 197.550 94.450 197.810 ;
        RECT 91.385 197.225 91.675 197.455 ;
        RECT 90.925 197.070 91.215 197.115 ;
        RECT 90.080 196.930 91.215 197.070 ;
        RECT 90.925 196.885 91.215 196.930 ;
        RECT 91.830 196.870 92.150 197.130 ;
        RECT 94.220 197.070 94.360 197.550 ;
        RECT 92.380 196.930 94.360 197.070 ;
        RECT 92.380 196.730 92.520 196.930 ;
        RECT 101.950 196.870 102.270 197.130 ;
        RECT 102.500 197.115 102.640 197.950 ;
        RECT 103.790 197.890 104.110 197.950 ;
        RECT 105.645 197.905 105.935 198.135 ;
        RECT 104.725 197.565 105.015 197.795 ;
        RECT 102.425 196.885 102.715 197.115 ;
        RECT 103.790 196.870 104.110 197.130 ;
        RECT 104.265 197.070 104.555 197.115 ;
        RECT 104.800 197.070 104.940 197.565 ;
        RECT 104.265 196.930 104.940 197.070 ;
        RECT 104.265 196.885 104.555 196.930 ;
        RECT 85.480 196.590 92.520 196.730 ;
        RECT 97.810 196.730 98.130 196.790 ;
        RECT 101.490 196.730 101.810 196.790 ;
        RECT 102.885 196.730 103.175 196.775 ;
        RECT 97.810 196.590 103.175 196.730 ;
        RECT 84.470 196.530 84.790 196.590 ;
        RECT 84.945 196.545 85.235 196.590 ;
        RECT 97.810 196.530 98.130 196.590 ;
        RECT 101.490 196.530 101.810 196.590 ;
        RECT 102.885 196.545 103.175 196.590 ;
        RECT 104.710 196.730 105.030 196.790 ;
        RECT 105.720 196.730 105.860 197.905 ;
        RECT 114.370 197.890 114.690 198.150 ;
        RECT 120.350 197.890 120.670 198.150 ;
        RECT 124.950 197.890 125.270 198.150 ;
        RECT 125.870 197.890 126.190 198.150 ;
        RECT 126.790 197.890 127.110 198.150 ;
        RECT 109.785 197.410 110.075 197.455 ;
        RECT 108.020 197.270 110.075 197.410 ;
        RECT 108.020 197.130 108.160 197.270 ;
        RECT 109.785 197.225 110.075 197.270 ;
        RECT 113.910 197.210 114.230 197.470 ;
        RECT 117.605 197.410 117.895 197.455 ;
        RECT 118.970 197.410 119.290 197.470 ;
        RECT 117.605 197.270 119.290 197.410 ;
        RECT 125.960 197.410 126.100 197.890 ;
        RECT 139.710 197.750 140.000 197.795 ;
        RECT 141.810 197.750 142.100 197.795 ;
        RECT 143.380 197.750 143.670 197.795 ;
        RECT 139.710 197.610 143.670 197.750 ;
        RECT 139.710 197.565 140.000 197.610 ;
        RECT 141.810 197.565 142.100 197.610 ;
        RECT 143.380 197.565 143.670 197.610 ;
        RECT 134.610 197.410 134.930 197.470 ;
        RECT 136.450 197.410 136.770 197.470 ;
        RECT 139.225 197.410 139.515 197.455 ;
        RECT 125.960 197.270 128.860 197.410 ;
        RECT 117.605 197.225 117.895 197.270 ;
        RECT 118.970 197.210 119.290 197.270 ;
        RECT 107.930 196.870 108.250 197.130 ;
        RECT 108.865 196.885 109.155 197.115 ;
        RECT 104.710 196.590 105.860 196.730 ;
        RECT 104.710 196.530 105.030 196.590 ;
        RECT 106.550 196.530 106.870 196.790 ;
        RECT 108.940 196.730 109.080 196.885 ;
        RECT 110.230 196.870 110.550 197.130 ;
        RECT 113.005 197.070 113.295 197.115 ;
        RECT 114.000 197.070 114.140 197.210 ;
        RECT 113.005 196.930 114.140 197.070 ;
        RECT 116.225 197.070 116.515 197.115 ;
        RECT 119.430 197.070 119.750 197.130 ;
        RECT 116.225 196.930 119.750 197.070 ;
        RECT 113.005 196.885 113.295 196.930 ;
        RECT 116.225 196.885 116.515 196.930 ;
        RECT 119.430 196.870 119.750 196.930 ;
        RECT 123.110 197.070 123.430 197.130 ;
        RECT 124.045 197.070 124.335 197.115 ;
        RECT 123.110 196.930 124.335 197.070 ;
        RECT 123.110 196.870 123.430 196.930 ;
        RECT 124.045 196.885 124.335 196.930 ;
        RECT 126.330 196.870 126.650 197.130 ;
        RECT 128.720 197.115 128.860 197.270 ;
        RECT 134.610 197.270 139.515 197.410 ;
        RECT 134.610 197.210 134.930 197.270 ;
        RECT 136.450 197.210 136.770 197.270 ;
        RECT 139.225 197.225 139.515 197.270 ;
        RECT 140.105 197.410 140.395 197.455 ;
        RECT 141.295 197.410 141.585 197.455 ;
        RECT 143.815 197.410 144.105 197.455 ;
        RECT 140.105 197.270 144.105 197.410 ;
        RECT 140.105 197.225 140.395 197.270 ;
        RECT 141.295 197.225 141.585 197.270 ;
        RECT 143.815 197.225 144.105 197.270 ;
        RECT 128.185 196.885 128.475 197.115 ;
        RECT 128.645 196.885 128.935 197.115 ;
        RECT 119.905 196.730 120.195 196.775 ;
        RECT 126.420 196.730 126.560 196.870 ;
        RECT 108.020 196.590 114.140 196.730 ;
        RECT 40.770 196.390 41.090 196.450 ;
        RECT 41.705 196.390 41.995 196.435 ;
        RECT 40.770 196.250 41.995 196.390 ;
        RECT 40.770 196.190 41.090 196.250 ;
        RECT 41.705 196.205 41.995 196.250 ;
        RECT 42.610 196.190 42.930 196.450 ;
        RECT 53.190 196.390 53.510 196.450 ;
        RECT 57.805 196.390 58.095 196.435 ;
        RECT 53.190 196.250 58.095 196.390 ;
        RECT 53.190 196.190 53.510 196.250 ;
        RECT 57.805 196.205 58.095 196.250 ;
        RECT 58.710 196.190 59.030 196.450 ;
        RECT 59.170 196.190 59.490 196.450 ;
        RECT 63.785 196.390 64.075 196.435 ;
        RECT 65.150 196.390 65.470 196.450 ;
        RECT 63.785 196.250 65.470 196.390 ;
        RECT 63.785 196.205 64.075 196.250 ;
        RECT 65.150 196.190 65.470 196.250 ;
        RECT 66.990 196.190 67.310 196.450 ;
        RECT 86.325 196.390 86.615 196.435 ;
        RECT 92.750 196.390 93.070 196.450 ;
        RECT 86.325 196.250 93.070 196.390 ;
        RECT 86.325 196.205 86.615 196.250 ;
        RECT 92.750 196.190 93.070 196.250 ;
        RECT 93.670 196.390 93.990 196.450 ;
        RECT 103.330 196.390 103.650 196.450 ;
        RECT 93.670 196.250 103.650 196.390 ;
        RECT 93.670 196.190 93.990 196.250 ;
        RECT 103.330 196.190 103.650 196.250 ;
        RECT 105.565 196.390 105.855 196.435 ;
        RECT 106.090 196.390 106.410 196.450 ;
        RECT 108.020 196.390 108.160 196.590 ;
        RECT 105.565 196.250 108.160 196.390 ;
        RECT 105.565 196.205 105.855 196.250 ;
        RECT 106.090 196.190 106.410 196.250 ;
        RECT 108.390 196.190 108.710 196.450 ;
        RECT 114.000 196.435 114.140 196.590 ;
        RECT 119.905 196.590 126.560 196.730 ;
        RECT 128.260 196.730 128.400 196.885 ;
        RECT 129.090 196.870 129.410 197.130 ;
        RECT 130.025 197.070 130.315 197.115 ;
        RECT 132.770 197.070 133.090 197.130 ;
        RECT 135.070 197.070 135.390 197.130 ;
        RECT 130.025 196.930 135.390 197.070 ;
        RECT 130.025 196.885 130.315 196.930 ;
        RECT 132.770 196.870 133.090 196.930 ;
        RECT 135.070 196.870 135.390 196.930 ;
        RECT 137.385 197.070 137.675 197.115 ;
        RECT 138.750 197.070 139.070 197.130 ;
        RECT 137.385 196.930 139.070 197.070 ;
        RECT 137.385 196.885 137.675 196.930 ;
        RECT 138.750 196.870 139.070 196.930 ;
        RECT 135.530 196.730 135.850 196.790 ;
        RECT 128.260 196.590 135.850 196.730 ;
        RECT 119.905 196.545 120.195 196.590 ;
        RECT 135.530 196.530 135.850 196.590 ;
        RECT 137.830 196.730 138.150 196.790 ;
        RECT 140.450 196.730 140.740 196.775 ;
        RECT 137.830 196.590 140.740 196.730 ;
        RECT 137.830 196.530 138.150 196.590 ;
        RECT 140.450 196.545 140.740 196.590 ;
        RECT 113.925 196.390 114.215 196.435 ;
        RECT 116.685 196.390 116.975 196.435 ;
        RECT 113.925 196.250 116.975 196.390 ;
        RECT 113.925 196.205 114.215 196.250 ;
        RECT 116.685 196.205 116.975 196.250 ;
        RECT 138.290 196.190 138.610 196.450 ;
        RECT 143.810 196.390 144.130 196.450 ;
        RECT 146.125 196.390 146.415 196.435 ;
        RECT 143.810 196.250 146.415 196.390 ;
        RECT 143.810 196.190 144.130 196.250 ;
        RECT 146.125 196.205 146.415 196.250 ;
        RECT 36.100 195.570 150.180 196.050 ;
        RECT 57.790 195.170 58.110 195.430 ;
        RECT 58.710 195.370 59.030 195.430 ;
        RECT 61.025 195.370 61.315 195.415 ;
        RECT 63.325 195.370 63.615 195.415 ;
        RECT 64.230 195.370 64.550 195.430 ;
        RECT 58.710 195.230 64.550 195.370 ;
        RECT 58.710 195.170 59.030 195.230 ;
        RECT 61.025 195.185 61.315 195.230 ;
        RECT 63.325 195.185 63.615 195.230 ;
        RECT 64.230 195.170 64.550 195.230 ;
        RECT 68.845 195.370 69.135 195.415 ;
        RECT 69.290 195.370 69.610 195.430 ;
        RECT 68.845 195.230 69.610 195.370 ;
        RECT 68.845 195.185 69.135 195.230 ;
        RECT 69.290 195.170 69.610 195.230 ;
        RECT 72.510 195.370 72.830 195.430 ;
        RECT 72.985 195.370 73.275 195.415 ;
        RECT 72.510 195.230 73.275 195.370 ;
        RECT 72.510 195.170 72.830 195.230 ;
        RECT 72.985 195.185 73.275 195.230 ;
        RECT 75.730 195.370 76.050 195.430 ;
        RECT 77.090 195.370 77.380 195.415 ;
        RECT 75.730 195.230 77.380 195.370 ;
        RECT 75.730 195.170 76.050 195.230 ;
        RECT 77.090 195.185 77.380 195.230 ;
        RECT 84.470 195.370 84.790 195.430 ;
        RECT 86.325 195.370 86.615 195.415 ;
        RECT 84.470 195.230 86.615 195.370 ;
        RECT 84.470 195.170 84.790 195.230 ;
        RECT 86.325 195.185 86.615 195.230 ;
        RECT 38.470 194.490 38.790 194.750 ;
        RECT 40.770 194.735 41.090 194.750 ;
        RECT 40.740 194.690 41.090 194.735 ;
        RECT 40.575 194.550 41.090 194.690 ;
        RECT 40.740 194.505 41.090 194.550 ;
        RECT 40.770 194.490 41.090 194.505 ;
        RECT 49.970 194.690 50.290 194.750 ;
        RECT 50.445 194.690 50.735 194.735 ;
        RECT 49.970 194.550 50.735 194.690 ;
        RECT 49.970 194.490 50.290 194.550 ;
        RECT 50.445 194.505 50.735 194.550 ;
        RECT 53.205 194.690 53.495 194.735 ;
        RECT 54.110 194.690 54.430 194.750 ;
        RECT 53.205 194.550 54.430 194.690 ;
        RECT 53.205 194.505 53.495 194.550 ;
        RECT 54.110 194.490 54.430 194.550 ;
        RECT 55.045 194.690 55.335 194.735 ;
        RECT 56.870 194.690 57.190 194.750 ;
        RECT 55.045 194.550 57.190 194.690 ;
        RECT 55.045 194.505 55.335 194.550 ;
        RECT 56.870 194.490 57.190 194.550 ;
        RECT 57.345 194.505 57.635 194.735 ;
        RECT 57.880 194.690 58.020 195.170 ;
        RECT 64.705 195.030 64.995 195.075 ;
        RECT 59.260 194.890 64.995 195.030 ;
        RECT 59.260 194.690 59.400 194.890 ;
        RECT 64.705 194.845 64.995 194.890 ;
        RECT 66.530 195.030 66.850 195.090 ;
        RECT 67.005 195.030 67.295 195.075 ;
        RECT 66.530 194.890 67.295 195.030 ;
        RECT 66.530 194.830 66.850 194.890 ;
        RECT 67.005 194.845 67.295 194.890 ;
        RECT 73.905 195.030 74.195 195.075 ;
        RECT 75.270 195.030 75.590 195.090 ;
        RECT 73.905 194.890 75.590 195.030 ;
        RECT 73.905 194.845 74.195 194.890 ;
        RECT 75.270 194.830 75.590 194.890 ;
        RECT 76.665 195.030 76.955 195.075 ;
        RECT 83.090 195.030 83.410 195.090 ;
        RECT 86.400 195.030 86.540 195.185 ;
        RECT 88.610 195.170 88.930 195.430 ;
        RECT 89.530 195.370 89.850 195.430 ;
        RECT 95.970 195.370 96.290 195.430 ;
        RECT 89.530 195.230 103.560 195.370 ;
        RECT 89.530 195.170 89.850 195.230 ;
        RECT 95.970 195.170 96.290 195.230 ;
        RECT 102.410 195.030 102.730 195.090 ;
        RECT 76.665 194.890 79.640 195.030 ;
        RECT 76.665 194.845 76.955 194.890 ;
        RECT 79.500 194.750 79.640 194.890 ;
        RECT 83.090 194.890 85.620 195.030 ;
        RECT 86.400 194.890 102.730 195.030 ;
        RECT 83.090 194.830 83.410 194.890 ;
        RECT 59.645 194.690 59.935 194.735 ;
        RECT 57.880 194.550 59.935 194.690 ;
        RECT 59.645 194.505 59.935 194.550 ;
        RECT 38.560 194.350 38.700 194.490 ;
        RECT 39.405 194.350 39.695 194.395 ;
        RECT 38.560 194.210 39.695 194.350 ;
        RECT 39.405 194.165 39.695 194.210 ;
        RECT 40.285 194.350 40.575 194.395 ;
        RECT 41.475 194.350 41.765 194.395 ;
        RECT 43.995 194.350 44.285 194.395 ;
        RECT 54.570 194.350 54.890 194.410 ;
        RECT 56.425 194.350 56.715 194.395 ;
        RECT 40.285 194.210 44.285 194.350 ;
        RECT 40.285 194.165 40.575 194.210 ;
        RECT 41.475 194.165 41.765 194.210 ;
        RECT 43.995 194.165 44.285 194.210 ;
        RECT 46.380 194.210 56.715 194.350 ;
        RECT 57.420 194.350 57.560 194.505 ;
        RECT 60.090 194.490 60.410 194.750 ;
        RECT 65.165 194.690 65.455 194.735 ;
        RECT 66.070 194.690 66.390 194.750 ;
        RECT 76.205 194.690 76.495 194.735 ;
        RECT 65.165 194.550 66.390 194.690 ;
        RECT 65.165 194.505 65.455 194.550 ;
        RECT 66.070 194.490 66.390 194.550 ;
        RECT 75.820 194.550 76.495 194.690 ;
        RECT 58.250 194.350 58.570 194.410 ;
        RECT 57.420 194.210 58.570 194.350 ;
        RECT 46.380 194.055 46.520 194.210 ;
        RECT 54.570 194.150 54.890 194.210 ;
        RECT 56.425 194.165 56.715 194.210 ;
        RECT 58.250 194.150 58.570 194.210 ;
        RECT 62.405 194.350 62.695 194.395 ;
        RECT 63.325 194.350 63.615 194.395 ;
        RECT 66.530 194.350 66.850 194.410 ;
        RECT 68.385 194.350 68.675 194.395 ;
        RECT 62.405 194.210 68.675 194.350 ;
        RECT 62.405 194.165 62.695 194.210 ;
        RECT 63.325 194.165 63.615 194.210 ;
        RECT 66.530 194.150 66.850 194.210 ;
        RECT 68.385 194.165 68.675 194.210 ;
        RECT 73.890 194.350 74.210 194.410 ;
        RECT 75.820 194.395 75.960 194.550 ;
        RECT 76.205 194.505 76.495 194.550 ;
        RECT 77.570 194.490 77.890 194.750 ;
        RECT 79.410 194.490 79.730 194.750 ;
        RECT 80.330 194.690 80.650 194.750 ;
        RECT 85.480 194.735 85.620 194.890 ;
        RECT 102.410 194.830 102.730 194.890 ;
        RECT 80.805 194.690 81.095 194.735 ;
        RECT 80.330 194.550 81.095 194.690 ;
        RECT 80.330 194.490 80.650 194.550 ;
        RECT 80.805 194.505 81.095 194.550 ;
        RECT 85.405 194.505 85.695 194.735 ;
        RECT 87.690 194.690 88.010 194.750 ;
        RECT 89.545 194.690 89.835 194.735 ;
        RECT 87.690 194.550 89.835 194.690 ;
        RECT 75.745 194.350 76.035 194.395 ;
        RECT 73.890 194.210 76.035 194.350 ;
        RECT 80.880 194.350 81.020 194.505 ;
        RECT 87.690 194.490 88.010 194.550 ;
        RECT 89.545 194.505 89.835 194.550 ;
        RECT 91.385 194.690 91.675 194.735 ;
        RECT 97.350 194.690 97.670 194.750 ;
        RECT 98.745 194.690 99.035 194.735 ;
        RECT 99.190 194.690 99.510 194.750 ;
        RECT 102.870 194.690 103.190 194.750 ;
        RECT 103.420 194.735 103.560 195.230 ;
        RECT 103.790 195.170 104.110 195.430 ;
        RECT 104.710 195.170 105.030 195.430 ;
        RECT 105.630 195.170 105.950 195.430 ;
        RECT 107.930 195.170 108.250 195.430 ;
        RECT 113.910 195.370 114.230 195.430 ;
        RECT 112.620 195.230 114.230 195.370 ;
        RECT 105.720 195.030 105.860 195.170 ;
        RECT 108.020 195.030 108.160 195.170 ;
        RECT 104.340 194.890 105.860 195.030 ;
        RECT 107.560 194.890 108.160 195.030 ;
        RECT 110.230 195.030 110.550 195.090 ;
        RECT 112.620 195.075 112.760 195.230 ;
        RECT 113.910 195.170 114.230 195.230 ;
        RECT 127.725 195.370 128.015 195.415 ;
        RECT 129.090 195.370 129.410 195.430 ;
        RECT 132.770 195.370 133.090 195.430 ;
        RECT 127.725 195.230 129.410 195.370 ;
        RECT 127.725 195.185 128.015 195.230 ;
        RECT 129.090 195.170 129.410 195.230 ;
        RECT 131.940 195.230 133.090 195.370 ;
        RECT 111.625 195.030 111.915 195.075 ;
        RECT 110.230 194.890 111.915 195.030 ;
        RECT 91.385 194.550 92.060 194.690 ;
        RECT 91.385 194.505 91.675 194.550 ;
        RECT 89.070 194.350 89.390 194.410 ;
        RECT 80.880 194.210 89.390 194.350 ;
        RECT 73.890 194.150 74.210 194.210 ;
        RECT 75.745 194.165 76.035 194.210 ;
        RECT 89.070 194.150 89.390 194.210 ;
        RECT 90.925 194.165 91.215 194.395 ;
        RECT 91.920 194.350 92.060 194.550 ;
        RECT 97.350 194.550 99.510 194.690 ;
        RECT 97.350 194.490 97.670 194.550 ;
        RECT 98.745 194.505 99.035 194.550 ;
        RECT 99.190 194.490 99.510 194.550 ;
        RECT 100.200 194.550 103.190 194.690 ;
        RECT 91.460 194.210 92.060 194.350 ;
        RECT 39.890 194.010 40.180 194.055 ;
        RECT 41.990 194.010 42.280 194.055 ;
        RECT 43.560 194.010 43.850 194.055 ;
        RECT 39.890 193.870 43.850 194.010 ;
        RECT 39.890 193.825 40.180 193.870 ;
        RECT 41.990 193.825 42.280 193.870 ;
        RECT 43.560 193.825 43.850 193.870 ;
        RECT 46.305 193.825 46.595 194.055 ;
        RECT 52.730 193.810 53.050 194.070 ;
        RECT 55.030 194.010 55.350 194.070 ;
        RECT 59.170 194.010 59.490 194.070 ;
        RECT 53.280 193.870 55.350 194.010 ;
        RECT 49.510 193.670 49.830 193.730 ;
        RECT 53.280 193.670 53.420 193.870 ;
        RECT 55.030 193.810 55.350 193.870 ;
        RECT 55.580 193.870 59.490 194.010 ;
        RECT 49.510 193.530 53.420 193.670 ;
        RECT 49.510 193.470 49.830 193.530 ;
        RECT 53.650 193.470 53.970 193.730 ;
        RECT 54.570 193.670 54.890 193.730 ;
        RECT 55.580 193.715 55.720 193.870 ;
        RECT 59.170 193.810 59.490 193.870 ;
        RECT 63.785 194.010 64.075 194.055 ;
        RECT 67.925 194.010 68.215 194.055 ;
        RECT 63.785 193.870 68.215 194.010 ;
        RECT 63.785 193.825 64.075 193.870 ;
        RECT 67.925 193.825 68.215 193.870 ;
        RECT 69.765 194.010 70.055 194.055 ;
        RECT 88.610 194.010 88.930 194.070 ;
        RECT 69.765 193.870 75.500 194.010 ;
        RECT 69.765 193.825 70.055 193.870 ;
        RECT 55.505 193.670 55.795 193.715 ;
        RECT 54.570 193.530 55.795 193.670 ;
        RECT 54.570 193.470 54.890 193.530 ;
        RECT 55.505 193.485 55.795 193.530 ;
        RECT 55.965 193.670 56.255 193.715 ;
        RECT 57.330 193.670 57.650 193.730 ;
        RECT 55.965 193.530 57.650 193.670 ;
        RECT 55.965 193.485 56.255 193.530 ;
        RECT 57.330 193.470 57.650 193.530 ;
        RECT 64.245 193.670 64.535 193.715 ;
        RECT 65.625 193.670 65.915 193.715 ;
        RECT 64.245 193.530 65.915 193.670 ;
        RECT 64.245 193.485 64.535 193.530 ;
        RECT 65.625 193.485 65.915 193.530 ;
        RECT 66.545 193.670 66.835 193.715 ;
        RECT 68.845 193.670 69.135 193.715 ;
        RECT 66.545 193.530 69.135 193.670 ;
        RECT 66.545 193.485 66.835 193.530 ;
        RECT 68.845 193.485 69.135 193.530 ;
        RECT 73.905 193.670 74.195 193.715 ;
        RECT 74.350 193.670 74.670 193.730 ;
        RECT 73.905 193.530 74.670 193.670 ;
        RECT 75.360 193.670 75.500 193.870 ;
        RECT 76.280 193.870 88.930 194.010 ;
        RECT 76.280 193.670 76.420 193.870 ;
        RECT 88.610 193.810 88.930 193.870 ;
        RECT 89.530 194.010 89.850 194.070 ;
        RECT 90.465 194.010 90.755 194.055 ;
        RECT 89.530 193.870 90.755 194.010 ;
        RECT 89.530 193.810 89.850 193.870 ;
        RECT 90.465 193.825 90.755 193.870 ;
        RECT 75.360 193.530 76.420 193.670 ;
        RECT 79.410 193.670 79.730 193.730 ;
        RECT 79.885 193.670 80.175 193.715 ;
        RECT 79.410 193.530 80.175 193.670 ;
        RECT 88.700 193.670 88.840 193.810 ;
        RECT 91.000 193.670 91.140 194.165 ;
        RECT 91.460 194.070 91.600 194.210 ;
        RECT 92.750 194.150 93.070 194.410 ;
        RECT 100.200 194.395 100.340 194.550 ;
        RECT 102.870 194.490 103.190 194.550 ;
        RECT 103.345 194.505 103.635 194.735 ;
        RECT 103.790 194.690 104.110 194.750 ;
        RECT 104.340 194.735 104.480 194.890 ;
        RECT 104.265 194.690 104.555 194.735 ;
        RECT 103.790 194.550 104.555 194.690 ;
        RECT 103.790 194.490 104.110 194.550 ;
        RECT 104.265 194.505 104.555 194.550 ;
        RECT 105.645 194.690 105.935 194.735 ;
        RECT 107.560 194.720 107.700 194.890 ;
        RECT 110.230 194.830 110.550 194.890 ;
        RECT 111.625 194.845 111.915 194.890 ;
        RECT 112.545 194.845 112.835 195.075 ;
        RECT 115.290 195.030 115.610 195.090 ;
        RECT 124.490 195.030 124.810 195.090 ;
        RECT 113.540 194.890 122.880 195.030 ;
        RECT 106.640 194.690 107.700 194.720 ;
        RECT 113.540 194.690 113.680 194.890 ;
        RECT 115.290 194.830 115.610 194.890 ;
        RECT 105.645 194.580 107.700 194.690 ;
        RECT 105.645 194.550 106.780 194.580 ;
        RECT 108.480 194.550 113.680 194.690 ;
        RECT 105.645 194.505 105.935 194.550 ;
        RECT 100.125 194.165 100.415 194.395 ;
        RECT 101.490 194.350 101.810 194.410 ;
        RECT 108.480 194.350 108.620 194.550 ;
        RECT 113.910 194.490 114.230 194.750 ;
        RECT 117.130 194.490 117.450 194.750 ;
        RECT 121.270 194.490 121.590 194.750 ;
        RECT 122.740 194.735 122.880 194.890 ;
        RECT 123.660 194.890 124.810 195.030 ;
        RECT 123.660 194.735 123.800 194.890 ;
        RECT 124.490 194.830 124.810 194.890 ;
        RECT 125.885 195.030 126.175 195.075 ;
        RECT 131.940 195.030 132.080 195.230 ;
        RECT 132.770 195.170 133.090 195.230 ;
        RECT 134.625 195.370 134.915 195.415 ;
        RECT 135.990 195.370 136.310 195.430 ;
        RECT 134.625 195.230 136.310 195.370 ;
        RECT 134.625 195.185 134.915 195.230 ;
        RECT 135.990 195.170 136.310 195.230 ;
        RECT 136.450 195.170 136.770 195.430 ;
        RECT 138.290 195.370 138.610 195.430 ;
        RECT 138.290 195.230 140.360 195.370 ;
        RECT 138.290 195.170 138.610 195.230 ;
        RECT 125.885 194.890 132.080 195.030 ;
        RECT 132.310 195.030 132.630 195.090 ;
        RECT 134.165 195.030 134.455 195.075 ;
        RECT 136.540 195.030 136.680 195.170 ;
        RECT 140.220 195.030 140.360 195.230 ;
        RECT 140.910 195.030 141.200 195.075 ;
        RECT 132.310 194.890 135.300 195.030 ;
        RECT 136.540 194.890 139.900 195.030 ;
        RECT 140.220 194.890 141.200 195.030 ;
        RECT 125.885 194.845 126.175 194.890 ;
        RECT 132.310 194.830 132.630 194.890 ;
        RECT 134.165 194.845 134.455 194.890 ;
        RECT 122.665 194.505 122.955 194.735 ;
        RECT 123.585 194.505 123.875 194.735 ;
        RECT 125.410 194.690 125.730 194.750 ;
        RECT 124.120 194.550 125.730 194.690 ;
        RECT 101.490 194.210 108.620 194.350 ;
        RECT 101.490 194.150 101.810 194.210 ;
        RECT 108.850 194.150 109.170 194.410 ;
        RECT 110.230 194.350 110.550 194.410 ;
        RECT 114.385 194.350 114.675 194.395 ;
        RECT 110.230 194.210 114.675 194.350 ;
        RECT 117.220 194.350 117.360 194.490 ;
        RECT 119.905 194.350 120.195 194.395 ;
        RECT 117.220 194.210 120.195 194.350 ;
        RECT 110.230 194.150 110.550 194.210 ;
        RECT 114.385 194.165 114.675 194.210 ;
        RECT 119.905 194.165 120.195 194.210 ;
        RECT 123.110 194.150 123.430 194.410 ;
        RECT 124.120 194.395 124.260 194.550 ;
        RECT 125.410 194.490 125.730 194.550 ;
        RECT 126.805 194.690 127.095 194.735 ;
        RECT 127.250 194.690 127.570 194.750 ;
        RECT 126.805 194.550 127.570 194.690 ;
        RECT 126.805 194.505 127.095 194.550 ;
        RECT 127.250 194.490 127.570 194.550 ;
        RECT 124.045 194.165 124.335 194.395 ;
        RECT 124.965 194.350 125.255 194.395 ;
        RECT 131.850 194.350 132.170 194.410 ;
        RECT 124.965 194.210 132.170 194.350 ;
        RECT 124.965 194.165 125.255 194.210 ;
        RECT 131.850 194.150 132.170 194.210 ;
        RECT 133.245 194.350 133.535 194.395 ;
        RECT 135.160 194.350 135.300 194.890 ;
        RECT 136.450 194.690 136.770 194.750 ;
        RECT 137.845 194.690 138.135 194.735 ;
        RECT 136.450 194.550 138.135 194.690 ;
        RECT 136.450 194.490 136.770 194.550 ;
        RECT 137.845 194.505 138.135 194.550 ;
        RECT 138.750 194.490 139.070 194.750 ;
        RECT 139.760 194.735 139.900 194.890 ;
        RECT 140.910 194.845 141.200 194.890 ;
        RECT 139.685 194.505 139.975 194.735 ;
        RECT 136.925 194.350 137.215 194.395 ;
        RECT 133.245 194.210 134.380 194.350 ;
        RECT 135.160 194.210 137.215 194.350 ;
        RECT 133.245 194.165 133.535 194.210 ;
        RECT 91.370 193.810 91.690 194.070 ;
        RECT 99.650 194.010 99.970 194.070 ;
        RECT 133.690 194.010 134.010 194.070 ;
        RECT 99.650 193.870 134.010 194.010 ;
        RECT 134.240 194.010 134.380 194.210 ;
        RECT 136.925 194.165 137.215 194.210 ;
        RECT 140.565 194.350 140.855 194.395 ;
        RECT 141.755 194.350 142.045 194.395 ;
        RECT 144.275 194.350 144.565 194.395 ;
        RECT 140.565 194.210 144.565 194.350 ;
        RECT 140.565 194.165 140.855 194.210 ;
        RECT 141.755 194.165 142.045 194.210 ;
        RECT 144.275 194.165 144.565 194.210 ;
        RECT 136.465 194.010 136.755 194.055 ;
        RECT 140.170 194.010 140.460 194.055 ;
        RECT 142.270 194.010 142.560 194.055 ;
        RECT 143.840 194.010 144.130 194.055 ;
        RECT 134.240 193.870 134.840 194.010 ;
        RECT 99.650 193.810 99.970 193.870 ;
        RECT 133.690 193.810 134.010 193.870 ;
        RECT 134.700 193.730 134.840 193.870 ;
        RECT 136.465 193.870 137.140 194.010 ;
        RECT 136.465 193.825 136.755 193.870 ;
        RECT 137.000 193.730 137.140 193.870 ;
        RECT 140.170 193.870 144.130 194.010 ;
        RECT 140.170 193.825 140.460 193.870 ;
        RECT 142.270 193.825 142.560 193.870 ;
        RECT 143.840 193.825 144.130 193.870 ;
        RECT 88.700 193.530 91.140 193.670 ;
        RECT 73.905 193.485 74.195 193.530 ;
        RECT 74.350 193.470 74.670 193.530 ;
        RECT 79.410 193.470 79.730 193.530 ;
        RECT 79.885 193.485 80.175 193.530 ;
        RECT 110.690 193.470 111.010 193.730 ;
        RECT 122.190 193.670 122.510 193.730 ;
        RECT 134.610 193.670 134.930 193.730 ;
        RECT 122.190 193.530 134.930 193.670 ;
        RECT 122.190 193.470 122.510 193.530 ;
        RECT 134.610 193.470 134.930 193.530 ;
        RECT 136.910 193.470 137.230 193.730 ;
        RECT 144.730 193.670 145.050 193.730 ;
        RECT 146.585 193.670 146.875 193.715 ;
        RECT 144.730 193.530 146.875 193.670 ;
        RECT 144.730 193.470 145.050 193.530 ;
        RECT 146.585 193.485 146.875 193.530 ;
        RECT 36.100 192.850 150.180 193.330 ;
        RECT 42.150 192.650 42.470 192.710 ;
        RECT 42.625 192.650 42.915 192.695 ;
        RECT 42.150 192.510 42.915 192.650 ;
        RECT 42.150 192.450 42.470 192.510 ;
        RECT 42.625 192.465 42.915 192.510 ;
        RECT 51.810 192.650 52.130 192.710 ;
        RECT 53.205 192.650 53.495 192.695 ;
        RECT 59.630 192.650 59.950 192.710 ;
        RECT 51.810 192.510 53.495 192.650 ;
        RECT 51.810 192.450 52.130 192.510 ;
        RECT 53.205 192.465 53.495 192.510 ;
        RECT 55.120 192.510 59.950 192.650 ;
        RECT 42.150 191.770 42.470 192.030 ;
        RECT 42.610 191.630 42.930 191.690 ;
        RECT 43.085 191.630 43.375 191.675 ;
        RECT 42.610 191.490 43.375 191.630 ;
        RECT 42.610 191.430 42.930 191.490 ;
        RECT 43.085 191.445 43.375 191.490 ;
        RECT 43.545 191.630 43.835 191.675 ;
        RECT 50.890 191.630 51.210 191.690 ;
        RECT 43.545 191.490 51.210 191.630 ;
        RECT 43.545 191.445 43.835 191.490 ;
        RECT 50.890 191.430 51.210 191.490 ;
        RECT 53.205 191.630 53.495 191.675 ;
        RECT 53.650 191.630 53.970 191.690 ;
        RECT 53.205 191.490 53.970 191.630 ;
        RECT 53.205 191.445 53.495 191.490 ;
        RECT 53.650 191.430 53.970 191.490 ;
        RECT 54.110 191.630 54.430 191.690 ;
        RECT 55.120 191.675 55.260 192.510 ;
        RECT 59.630 192.450 59.950 192.510 ;
        RECT 66.530 192.650 66.850 192.710 ;
        RECT 67.005 192.650 67.295 192.695 ;
        RECT 66.530 192.510 67.295 192.650 ;
        RECT 66.530 192.450 66.850 192.510 ;
        RECT 67.005 192.465 67.295 192.510 ;
        RECT 75.270 192.450 75.590 192.710 ;
        RECT 77.570 192.650 77.890 192.710 ;
        RECT 78.505 192.650 78.795 192.695 ;
        RECT 77.570 192.510 78.795 192.650 ;
        RECT 77.570 192.450 77.890 192.510 ;
        RECT 78.505 192.465 78.795 192.510 ;
        RECT 80.790 192.450 81.110 192.710 ;
        RECT 87.690 192.450 88.010 192.710 ;
        RECT 89.990 192.650 90.310 192.710 ;
        RECT 91.845 192.650 92.135 192.695 ;
        RECT 96.430 192.650 96.750 192.710 ;
        RECT 96.905 192.650 97.195 192.695 ;
        RECT 89.990 192.510 92.135 192.650 ;
        RECT 89.990 192.450 90.310 192.510 ;
        RECT 91.845 192.465 92.135 192.510 ;
        RECT 94.220 192.510 96.200 192.650 ;
        RECT 57.330 192.310 57.650 192.370 ;
        RECT 73.890 192.310 74.210 192.370 ;
        RECT 78.965 192.310 79.255 192.355 ;
        RECT 56.960 192.170 57.650 192.310 ;
        RECT 55.045 191.630 55.335 191.675 ;
        RECT 54.110 191.490 55.335 191.630 ;
        RECT 54.110 191.430 54.430 191.490 ;
        RECT 55.045 191.445 55.335 191.490 ;
        RECT 55.505 191.630 55.795 191.675 ;
        RECT 56.425 191.630 56.715 191.675 ;
        RECT 55.505 191.490 56.715 191.630 ;
        RECT 55.505 191.445 55.795 191.490 ;
        RECT 56.425 191.445 56.715 191.490 ;
        RECT 56.960 191.290 57.100 192.170 ;
        RECT 57.330 192.110 57.650 192.170 ;
        RECT 57.880 192.170 63.080 192.310 ;
        RECT 57.880 192.015 58.020 192.170 ;
        RECT 57.805 191.785 58.095 192.015 ;
        RECT 59.170 191.970 59.490 192.030 ;
        RECT 59.645 191.970 59.935 192.015 ;
        RECT 59.170 191.830 59.935 191.970 ;
        RECT 59.170 191.770 59.490 191.830 ;
        RECT 59.645 191.785 59.935 191.830 ;
        RECT 61.010 191.970 61.330 192.030 ;
        RECT 61.010 191.830 62.620 191.970 ;
        RECT 61.010 191.770 61.330 191.830 ;
        RECT 57.330 191.430 57.650 191.690 ;
        RECT 61.485 191.630 61.775 191.675 ;
        RECT 61.485 191.490 62.160 191.630 ;
        RECT 61.485 191.445 61.775 191.490 ;
        RECT 62.020 191.350 62.160 191.490 ;
        RECT 62.480 191.350 62.620 191.830 ;
        RECT 62.940 191.630 63.080 192.170 ;
        RECT 73.890 192.170 79.255 192.310 ;
        RECT 73.890 192.110 74.210 192.170 ;
        RECT 78.965 192.125 79.255 192.170 ;
        RECT 64.705 191.970 64.995 192.015 ;
        RECT 65.610 191.970 65.930 192.030 ;
        RECT 67.450 191.970 67.770 192.030 ;
        RECT 64.705 191.830 67.770 191.970 ;
        RECT 64.705 191.785 64.995 191.830 ;
        RECT 65.610 191.770 65.930 191.830 ;
        RECT 67.450 191.770 67.770 191.830 ;
        RECT 75.820 191.830 77.340 191.970 ;
        RECT 75.820 191.690 75.960 191.830 ;
        RECT 65.150 191.630 65.470 191.690 ;
        RECT 66.085 191.630 66.375 191.675 ;
        RECT 67.910 191.630 68.230 191.690 ;
        RECT 62.940 191.490 68.230 191.630 ;
        RECT 65.150 191.430 65.470 191.490 ;
        RECT 66.085 191.445 66.375 191.490 ;
        RECT 67.910 191.430 68.230 191.490 ;
        RECT 75.730 191.430 76.050 191.690 ;
        RECT 77.200 191.675 77.340 191.830 ;
        RECT 78.030 191.770 78.350 192.030 ;
        RECT 76.435 191.630 76.725 191.675 ;
        RECT 76.435 191.445 76.780 191.630 ;
        RECT 77.125 191.445 77.415 191.675 ;
        RECT 59.185 191.290 59.475 191.335 ;
        RECT 61.930 191.290 62.250 191.350 ;
        RECT 56.960 191.150 59.475 191.290 ;
        RECT 59.185 191.105 59.475 191.150 ;
        RECT 60.180 191.150 62.250 191.290 ;
        RECT 52.270 190.750 52.590 191.010 ;
        RECT 58.725 190.950 59.015 190.995 ;
        RECT 60.180 190.950 60.320 191.150 ;
        RECT 61.930 191.090 62.250 191.150 ;
        RECT 62.390 191.290 62.710 191.350 ;
        RECT 67.465 191.290 67.755 191.335 ;
        RECT 62.390 191.150 67.755 191.290 ;
        RECT 62.390 191.090 62.710 191.150 ;
        RECT 67.465 191.105 67.755 191.150 ;
        RECT 58.725 190.810 60.320 190.950 ;
        RECT 60.565 190.950 60.855 190.995 ;
        RECT 61.010 190.950 61.330 191.010 ;
        RECT 60.565 190.810 61.330 190.950 ;
        RECT 58.725 190.765 59.015 190.810 ;
        RECT 60.565 190.765 60.855 190.810 ;
        RECT 61.010 190.750 61.330 190.810 ;
        RECT 75.730 190.950 76.050 191.010 ;
        RECT 76.640 190.950 76.780 191.445 ;
        RECT 77.570 191.430 77.890 191.690 ;
        RECT 80.880 191.675 81.020 192.450 ;
        RECT 88.610 192.310 88.930 192.370 ;
        RECT 93.685 192.310 93.975 192.355 ;
        RECT 88.610 192.170 93.975 192.310 ;
        RECT 88.610 192.110 88.930 192.170 ;
        RECT 93.685 192.125 93.975 192.170 ;
        RECT 83.090 191.970 83.410 192.030 ;
        RECT 90.005 191.970 90.295 192.015 ;
        RECT 94.220 191.970 94.360 192.510 ;
        RECT 95.525 192.125 95.815 192.355 ;
        RECT 96.060 192.310 96.200 192.510 ;
        RECT 96.430 192.510 97.195 192.650 ;
        RECT 96.430 192.450 96.750 192.510 ;
        RECT 96.905 192.465 97.195 192.510 ;
        RECT 99.190 192.650 99.510 192.710 ;
        RECT 105.185 192.650 105.475 192.695 ;
        RECT 99.190 192.510 105.475 192.650 ;
        RECT 99.190 192.450 99.510 192.510 ;
        RECT 105.185 192.465 105.475 192.510 ;
        RECT 112.530 192.650 112.850 192.710 ;
        RECT 114.845 192.650 115.135 192.695 ;
        RECT 112.530 192.510 115.135 192.650 ;
        RECT 112.530 192.450 112.850 192.510 ;
        RECT 114.845 192.465 115.135 192.510 ;
        RECT 115.290 192.650 115.610 192.710 ;
        RECT 119.905 192.650 120.195 192.695 ;
        RECT 115.290 192.510 120.195 192.650 ;
        RECT 115.290 192.450 115.610 192.510 ;
        RECT 119.905 192.465 120.195 192.510 ;
        RECT 124.490 192.650 124.810 192.710 ;
        RECT 127.725 192.650 128.015 192.695 ;
        RECT 124.490 192.510 128.015 192.650 ;
        RECT 124.490 192.450 124.810 192.510 ;
        RECT 127.725 192.465 128.015 192.510 ;
        RECT 131.405 192.650 131.695 192.695 ;
        RECT 132.310 192.650 132.630 192.710 ;
        RECT 131.405 192.510 132.630 192.650 ;
        RECT 131.405 192.465 131.695 192.510 ;
        RECT 132.310 192.450 132.630 192.510 ;
        RECT 132.770 192.450 133.090 192.710 ;
        RECT 134.625 192.650 134.915 192.695 ;
        RECT 133.320 192.510 134.915 192.650 ;
        RECT 101.045 192.310 101.335 192.355 ;
        RECT 102.870 192.310 103.190 192.370 ;
        RECT 96.060 192.170 101.335 192.310 ;
        RECT 101.045 192.125 101.335 192.170 ;
        RECT 101.580 192.170 103.190 192.310 ;
        RECT 83.090 191.830 90.295 191.970 ;
        RECT 83.090 191.770 83.410 191.830 ;
        RECT 90.005 191.785 90.295 191.830 ;
        RECT 91.030 191.830 92.520 191.970 ;
        RECT 80.805 191.630 81.095 191.675 ;
        RECT 88.625 191.630 88.915 191.675 ;
        RECT 79.420 191.350 79.710 191.565 ;
        RECT 80.805 191.490 88.915 191.630 ;
        RECT 80.805 191.445 81.095 191.490 ;
        RECT 88.625 191.445 88.915 191.490 ;
        RECT 89.070 191.630 89.390 191.690 ;
        RECT 89.545 191.630 89.835 191.675 ;
        RECT 89.070 191.490 89.835 191.630 ;
        RECT 89.070 191.430 89.390 191.490 ;
        RECT 89.545 191.445 89.835 191.490 ;
        RECT 90.450 191.430 90.770 191.690 ;
        RECT 79.410 191.090 79.730 191.350 ;
        RECT 80.330 191.290 80.650 191.350 ;
        RECT 91.030 191.290 91.170 191.830 ;
        RECT 92.380 191.690 92.520 191.830 ;
        RECT 92.840 191.830 94.360 191.970 ;
        RECT 91.385 191.630 91.675 191.675 ;
        RECT 91.385 191.490 92.060 191.630 ;
        RECT 91.385 191.445 91.675 191.490 ;
        RECT 80.330 191.150 91.170 191.290 ;
        RECT 91.920 191.290 92.060 191.490 ;
        RECT 92.290 191.430 92.610 191.690 ;
        RECT 92.840 191.675 92.980 191.830 ;
        RECT 95.600 191.690 95.740 192.125 ;
        RECT 97.350 191.770 97.670 192.030 ;
        RECT 92.765 191.445 93.055 191.675 ;
        RECT 94.130 191.430 94.450 191.690 ;
        RECT 95.510 191.630 95.830 191.690 ;
        RECT 94.680 191.490 95.830 191.630 ;
        RECT 94.680 191.290 94.820 191.490 ;
        RECT 95.510 191.430 95.830 191.490 ;
        RECT 96.445 191.630 96.735 191.675 ;
        RECT 97.440 191.630 97.580 191.770 ;
        RECT 96.445 191.490 97.580 191.630 ;
        RECT 96.445 191.445 96.735 191.490 ;
        RECT 98.270 191.430 98.590 191.690 ;
        RECT 98.745 191.445 99.035 191.675 ;
        RECT 91.920 191.150 94.820 191.290 ;
        RECT 80.330 191.090 80.650 191.150 ;
        RECT 79.885 190.950 80.175 190.995 ;
        RECT 89.990 190.950 90.310 191.010 ;
        RECT 75.730 190.810 90.310 190.950 ;
        RECT 75.730 190.750 76.050 190.810 ;
        RECT 79.885 190.765 80.175 190.810 ;
        RECT 89.990 190.750 90.310 190.810 ;
        RECT 90.450 190.950 90.770 191.010 ;
        RECT 98.820 190.950 98.960 191.445 ;
        RECT 99.190 191.430 99.510 191.690 ;
        RECT 100.125 191.445 100.415 191.675 ;
        RECT 100.200 191.290 100.340 191.445 ;
        RECT 101.580 191.290 101.720 192.170 ;
        RECT 102.870 192.110 103.190 192.170 ;
        RECT 107.945 192.310 108.235 192.355 ;
        RECT 121.285 192.310 121.575 192.355 ;
        RECT 107.945 192.170 121.575 192.310 ;
        RECT 107.945 192.125 108.235 192.170 ;
        RECT 102.410 191.970 102.730 192.030 ;
        RECT 110.230 191.970 110.550 192.030 ;
        RECT 102.410 191.830 103.560 191.970 ;
        RECT 102.410 191.770 102.730 191.830 ;
        RECT 101.950 191.430 102.270 191.690 ;
        RECT 102.870 191.430 103.190 191.690 ;
        RECT 103.420 191.675 103.560 191.830 ;
        RECT 108.940 191.830 110.550 191.970 ;
        RECT 103.345 191.445 103.635 191.675 ;
        RECT 103.790 191.430 104.110 191.690 ;
        RECT 104.250 191.580 104.570 191.690 ;
        RECT 106.090 191.630 106.410 191.690 ;
        RECT 104.725 191.580 105.015 191.625 ;
        RECT 104.250 191.440 105.015 191.580 ;
        RECT 105.895 191.490 106.410 191.630 ;
        RECT 104.250 191.430 104.570 191.440 ;
        RECT 104.725 191.395 105.015 191.440 ;
        RECT 106.090 191.430 106.410 191.490 ;
        RECT 106.550 191.630 106.870 191.690 ;
        RECT 108.940 191.675 109.080 191.830 ;
        RECT 110.230 191.770 110.550 191.830 ;
        RECT 116.685 191.970 116.975 192.015 ;
        RECT 118.510 191.970 118.830 192.030 ;
        RECT 116.685 191.830 118.830 191.970 ;
        RECT 116.685 191.785 116.975 191.830 ;
        RECT 118.510 191.770 118.830 191.830 ;
        RECT 119.060 191.690 119.200 192.170 ;
        RECT 121.285 192.125 121.575 192.170 ;
        RECT 133.320 191.970 133.460 192.510 ;
        RECT 134.625 192.465 134.915 192.510 ;
        RECT 137.830 192.450 138.150 192.710 ;
        RECT 129.180 191.830 133.460 191.970 ;
        RECT 133.780 192.170 147.720 192.310 ;
        RECT 108.405 191.630 108.695 191.675 ;
        RECT 106.550 191.490 108.695 191.630 ;
        RECT 106.550 191.430 106.870 191.490 ;
        RECT 108.405 191.445 108.695 191.490 ;
        RECT 108.865 191.445 109.155 191.675 ;
        RECT 109.770 191.430 110.090 191.690 ;
        RECT 111.625 191.630 111.915 191.675 ;
        RECT 113.910 191.630 114.230 191.690 ;
        RECT 111.625 191.490 114.230 191.630 ;
        RECT 111.625 191.445 111.915 191.490 ;
        RECT 113.910 191.430 114.230 191.490 ;
        RECT 114.370 191.630 114.690 191.690 ;
        RECT 115.765 191.630 116.055 191.675 ;
        RECT 114.370 191.490 116.055 191.630 ;
        RECT 114.370 191.430 114.690 191.490 ;
        RECT 115.765 191.445 116.055 191.490 ;
        RECT 116.225 191.445 116.515 191.675 ;
        RECT 102.410 191.290 102.730 191.350 ;
        RECT 116.300 191.290 116.440 191.445 ;
        RECT 117.130 191.430 117.450 191.690 ;
        RECT 118.970 191.430 119.290 191.690 ;
        RECT 120.365 191.630 120.655 191.675 ;
        RECT 121.270 191.630 121.590 191.690 ;
        RECT 129.180 191.675 129.320 191.830 ;
        RECT 120.365 191.490 121.590 191.630 ;
        RECT 120.365 191.445 120.655 191.490 ;
        RECT 121.270 191.430 121.590 191.490 ;
        RECT 128.645 191.445 128.935 191.675 ;
        RECT 129.105 191.445 129.395 191.675 ;
        RECT 130.010 191.630 130.330 191.690 ;
        RECT 130.485 191.630 130.775 191.675 ;
        RECT 130.010 191.490 130.775 191.630 ;
        RECT 100.200 191.150 102.730 191.290 ;
        RECT 102.410 191.090 102.730 191.150 ;
        RECT 105.260 191.150 116.440 191.290 ;
        RECT 128.720 191.290 128.860 191.445 ;
        RECT 130.010 191.430 130.330 191.490 ;
        RECT 130.485 191.445 130.775 191.490 ;
        RECT 129.565 191.290 129.855 191.335 ;
        RECT 132.555 191.290 132.845 191.505 ;
        RECT 133.780 191.335 133.920 192.170 ;
        RECT 147.580 192.030 147.720 192.170 ;
        RECT 134.610 191.970 134.930 192.030 ;
        RECT 141.065 191.970 141.355 192.015 ;
        RECT 134.610 191.830 141.355 191.970 ;
        RECT 134.610 191.770 134.930 191.830 ;
        RECT 141.065 191.785 141.355 191.830 ;
        RECT 143.810 191.970 144.130 192.030 ;
        RECT 143.810 191.830 145.420 191.970 ;
        RECT 143.810 191.770 144.130 191.830 ;
        RECT 134.165 191.445 134.455 191.675 ;
        RECT 128.720 191.150 132.080 191.290 ;
        RECT 90.450 190.810 98.960 190.950 ;
        RECT 99.190 190.950 99.510 191.010 ;
        RECT 105.260 190.950 105.400 191.150 ;
        RECT 129.565 191.105 129.855 191.150 ;
        RECT 99.190 190.810 105.400 190.950 ;
        RECT 105.630 190.950 105.950 191.010 ;
        RECT 106.105 190.950 106.395 190.995 ;
        RECT 105.630 190.810 106.395 190.950 ;
        RECT 90.450 190.750 90.770 190.810 ;
        RECT 99.190 190.750 99.510 190.810 ;
        RECT 105.630 190.750 105.950 190.810 ;
        RECT 106.105 190.765 106.395 190.810 ;
        RECT 109.785 190.950 110.075 190.995 ;
        RECT 110.230 190.950 110.550 191.010 ;
        RECT 109.785 190.810 110.550 190.950 ;
        RECT 109.785 190.765 110.075 190.810 ;
        RECT 110.230 190.750 110.550 190.810 ;
        RECT 119.430 190.950 119.750 191.010 ;
        RECT 125.870 190.950 126.190 191.010 ;
        RECT 131.940 190.995 132.080 191.150 ;
        RECT 132.400 191.275 132.845 191.290 ;
        RECT 132.400 191.150 132.770 191.275 ;
        RECT 132.400 191.010 132.540 191.150 ;
        RECT 133.705 191.105 133.995 191.335 ;
        RECT 119.430 190.810 126.190 190.950 ;
        RECT 119.430 190.750 119.750 190.810 ;
        RECT 125.870 190.750 126.190 190.810 ;
        RECT 131.865 190.765 132.155 190.995 ;
        RECT 132.310 190.750 132.630 191.010 ;
        RECT 133.230 190.950 133.550 191.010 ;
        RECT 134.240 190.950 134.380 191.445 ;
        RECT 136.910 191.430 137.230 191.690 ;
        RECT 137.370 191.430 137.690 191.690 ;
        RECT 144.360 191.675 144.500 191.830 ;
        RECT 142.445 191.630 142.735 191.675 ;
        RECT 144.285 191.630 144.575 191.675 ;
        RECT 142.445 191.490 144.575 191.630 ;
        RECT 142.445 191.445 142.735 191.490 ;
        RECT 144.285 191.445 144.575 191.490 ;
        RECT 144.730 191.430 145.050 191.690 ;
        RECT 145.280 191.630 145.420 191.830 ;
        RECT 147.490 191.770 147.810 192.030 ;
        RECT 145.280 191.490 148.180 191.630 ;
        RECT 137.460 191.290 137.600 191.430 ;
        RECT 142.905 191.290 143.195 191.335 ;
        RECT 137.460 191.150 143.195 191.290 ;
        RECT 142.905 191.105 143.195 191.150 ;
        RECT 143.825 191.290 144.115 191.335 ;
        RECT 144.820 191.290 144.960 191.430 ;
        RECT 143.825 191.150 144.960 191.290 ;
        RECT 143.825 191.105 144.115 191.150 ;
        RECT 148.040 191.010 148.180 191.490 ;
        RECT 133.230 190.810 134.380 190.950 ;
        RECT 142.430 190.950 142.750 191.010 ;
        RECT 143.365 190.950 143.655 190.995 ;
        RECT 142.430 190.810 143.655 190.950 ;
        RECT 133.230 190.750 133.550 190.810 ;
        RECT 142.430 190.750 142.750 190.810 ;
        RECT 143.365 190.765 143.655 190.810 ;
        RECT 147.950 190.750 148.270 191.010 ;
        RECT 36.100 190.130 150.180 190.610 ;
        RECT 42.150 189.930 42.470 189.990 ;
        RECT 42.625 189.930 42.915 189.975 ;
        RECT 43.990 189.930 44.310 189.990 ;
        RECT 44.925 189.930 45.215 189.975 ;
        RECT 66.990 189.930 67.310 189.990 ;
        RECT 42.150 189.790 42.915 189.930 ;
        RECT 42.150 189.730 42.470 189.790 ;
        RECT 42.625 189.745 42.915 189.790 ;
        RECT 43.160 189.790 45.215 189.930 ;
        RECT 41.245 189.250 41.535 189.295 ;
        RECT 41.690 189.250 42.010 189.310 ;
        RECT 43.160 189.295 43.300 189.790 ;
        RECT 43.990 189.730 44.310 189.790 ;
        RECT 44.925 189.745 45.215 189.790 ;
        RECT 50.520 189.790 67.310 189.930 ;
        RECT 44.540 189.450 46.520 189.590 ;
        RECT 44.540 189.295 44.680 189.450 ;
        RECT 46.380 189.310 46.520 189.450 ;
        RECT 46.750 189.390 47.070 189.650 ;
        RECT 49.510 189.635 49.830 189.650 ;
        RECT 50.520 189.635 50.660 189.790 ;
        RECT 66.990 189.730 67.310 189.790 ;
        RECT 73.890 189.930 74.210 189.990 ;
        RECT 74.365 189.930 74.655 189.975 ;
        RECT 73.890 189.790 74.655 189.930 ;
        RECT 73.890 189.730 74.210 189.790 ;
        RECT 74.365 189.745 74.655 189.790 ;
        RECT 75.730 189.730 76.050 189.990 ;
        RECT 88.610 189.930 88.930 189.990 ;
        RECT 90.450 189.930 90.770 189.990 ;
        RECT 86.400 189.790 88.930 189.930 ;
        RECT 49.445 189.405 49.830 189.635 ;
        RECT 50.445 189.405 50.735 189.635 ;
        RECT 61.010 189.590 61.330 189.650 ;
        RECT 54.200 189.450 61.330 189.590 ;
        RECT 75.820 189.590 75.960 189.730 ;
        RECT 76.205 189.590 76.495 189.635 ;
        RECT 77.570 189.590 77.890 189.650 ;
        RECT 49.510 189.390 49.830 189.405 ;
        RECT 41.245 189.110 42.010 189.250 ;
        RECT 41.245 189.065 41.535 189.110 ;
        RECT 41.690 189.050 42.010 189.110 ;
        RECT 43.085 189.065 43.375 189.295 ;
        RECT 44.005 189.065 44.295 189.295 ;
        RECT 44.465 189.065 44.755 189.295 ;
        RECT 45.845 189.065 46.135 189.295 ;
        RECT 39.390 188.710 39.710 188.970 ;
        RECT 39.480 188.570 39.620 188.710 ;
        RECT 43.085 188.570 43.375 188.615 ;
        RECT 39.480 188.430 43.375 188.570 ;
        RECT 43.085 188.385 43.375 188.430 ;
        RECT 38.930 188.230 39.250 188.290 ;
        RECT 40.325 188.230 40.615 188.275 ;
        RECT 43.530 188.230 43.850 188.290 ;
        RECT 38.930 188.090 43.850 188.230 ;
        RECT 44.080 188.230 44.220 189.065 ;
        RECT 45.920 188.570 46.060 189.065 ;
        RECT 46.290 189.050 46.610 189.310 ;
        RECT 47.455 189.065 47.745 189.295 ;
        RECT 49.970 189.250 50.290 189.310 ;
        RECT 54.200 189.250 54.340 189.450 ;
        RECT 49.970 189.110 54.340 189.250 ;
        RECT 54.570 189.250 54.890 189.310 ;
        RECT 60.180 189.295 60.320 189.450 ;
        RECT 61.010 189.390 61.330 189.450 ;
        RECT 75.055 189.420 75.345 189.465 ;
        RECT 75.820 189.450 76.495 189.590 ;
        RECT 75.055 189.310 75.420 189.420 ;
        RECT 76.205 189.405 76.495 189.450 ;
        RECT 77.200 189.450 77.890 189.590 ;
        RECT 56.425 189.250 56.715 189.295 ;
        RECT 54.570 189.110 56.715 189.250 ;
        RECT 47.530 188.910 47.670 189.065 ;
        RECT 49.970 189.050 50.290 189.110 ;
        RECT 54.570 189.050 54.890 189.110 ;
        RECT 56.425 189.065 56.715 189.110 ;
        RECT 57.345 189.065 57.635 189.295 ;
        RECT 60.105 189.065 60.395 189.295 ;
        RECT 47.530 188.770 47.900 188.910 ;
        RECT 47.760 188.630 47.900 188.770 ;
        RECT 48.145 188.725 48.435 188.955 ;
        RECT 57.420 188.910 57.560 189.065 ;
        RECT 72.510 189.050 72.830 189.310 ;
        RECT 74.810 189.110 75.420 189.310 ;
        RECT 74.810 189.050 75.130 189.110 ;
        RECT 76.650 189.050 76.970 189.310 ;
        RECT 77.200 188.955 77.340 189.450 ;
        RECT 77.570 189.390 77.890 189.450 ;
        RECT 78.490 189.050 78.810 189.310 ;
        RECT 79.425 189.065 79.715 189.295 ;
        RECT 83.090 189.250 83.410 189.310 ;
        RECT 86.400 189.295 86.540 189.790 ;
        RECT 88.610 189.730 88.930 189.790 ;
        RECT 89.620 189.790 90.770 189.930 ;
        RECT 87.245 189.590 87.535 189.635 ;
        RECT 87.245 189.450 89.300 189.590 ;
        RECT 87.245 189.405 87.535 189.450 ;
        RECT 84.485 189.250 84.775 189.295 ;
        RECT 83.090 189.110 84.775 189.250 ;
        RECT 77.125 188.910 77.415 188.955 ;
        RECT 57.420 188.770 63.540 188.910 ;
        RECT 47.210 188.570 47.530 188.630 ;
        RECT 45.920 188.430 47.530 188.570 ;
        RECT 47.210 188.370 47.530 188.430 ;
        RECT 47.670 188.370 47.990 188.630 ;
        RECT 48.220 188.570 48.360 188.725 ;
        RECT 63.400 188.630 63.540 188.770 ;
        RECT 73.060 188.770 77.415 188.910 ;
        RECT 48.605 188.570 48.895 188.615 ;
        RECT 48.220 188.430 48.895 188.570 ;
        RECT 48.605 188.385 48.895 188.430 ;
        RECT 63.310 188.570 63.630 188.630 ;
        RECT 64.230 188.570 64.550 188.630 ;
        RECT 63.310 188.430 64.550 188.570 ;
        RECT 63.310 188.370 63.630 188.430 ;
        RECT 64.230 188.370 64.550 188.430 ;
        RECT 47.760 188.230 47.900 188.370 ;
        RECT 73.060 188.290 73.200 188.770 ;
        RECT 77.125 188.725 77.415 188.770 ;
        RECT 78.045 188.910 78.335 188.955 ;
        RECT 78.580 188.910 78.720 189.050 ;
        RECT 78.045 188.770 78.720 188.910 ;
        RECT 79.500 188.910 79.640 189.065 ;
        RECT 83.090 189.050 83.410 189.110 ;
        RECT 84.485 189.065 84.775 189.110 ;
        RECT 85.865 189.065 86.155 189.295 ;
        RECT 86.325 189.065 86.615 189.295 ;
        RECT 79.870 188.910 80.190 188.970 ;
        RECT 79.500 188.770 80.190 188.910 ;
        RECT 85.940 188.910 86.080 189.065 ;
        RECT 88.150 189.050 88.470 189.310 ;
        RECT 89.160 189.295 89.300 189.450 ;
        RECT 89.620 189.310 89.760 189.790 ;
        RECT 90.450 189.730 90.770 189.790 ;
        RECT 91.385 189.930 91.675 189.975 ;
        RECT 91.830 189.930 92.150 189.990 ;
        RECT 101.950 189.930 102.270 189.990 ;
        RECT 91.385 189.790 92.150 189.930 ;
        RECT 91.385 189.745 91.675 189.790 ;
        RECT 91.830 189.730 92.150 189.790 ;
        RECT 92.380 189.790 102.270 189.930 ;
        RECT 92.380 189.590 92.520 189.790 ;
        RECT 101.950 189.730 102.270 189.790 ;
        RECT 103.790 189.930 104.110 189.990 ;
        RECT 109.770 189.930 110.090 189.990 ;
        RECT 103.790 189.790 110.090 189.930 ;
        RECT 103.790 189.730 104.110 189.790 ;
        RECT 109.770 189.730 110.090 189.790 ;
        RECT 116.685 189.930 116.975 189.975 ;
        RECT 117.130 189.930 117.450 189.990 ;
        RECT 116.685 189.790 117.450 189.930 ;
        RECT 116.685 189.745 116.975 189.790 ;
        RECT 117.130 189.730 117.450 189.790 ;
        RECT 118.970 189.930 119.290 189.990 ;
        RECT 119.445 189.930 119.735 189.975 ;
        RECT 126.790 189.930 127.110 189.990 ;
        RECT 118.970 189.790 127.110 189.930 ;
        RECT 118.970 189.730 119.290 189.790 ;
        RECT 119.445 189.745 119.735 189.790 ;
        RECT 126.790 189.730 127.110 189.790 ;
        RECT 128.185 189.930 128.475 189.975 ;
        RECT 128.630 189.930 128.950 189.990 ;
        RECT 128.185 189.790 128.950 189.930 ;
        RECT 128.185 189.745 128.475 189.790 ;
        RECT 128.630 189.730 128.950 189.790 ;
        RECT 130.010 189.930 130.330 189.990 ;
        RECT 134.150 189.930 134.470 189.990 ;
        RECT 130.010 189.790 134.470 189.930 ;
        RECT 130.010 189.730 130.330 189.790 ;
        RECT 134.150 189.730 134.470 189.790 ;
        RECT 141.050 189.730 141.370 189.990 ;
        RECT 144.270 189.730 144.590 189.990 ;
        RECT 90.540 189.450 92.520 189.590 ;
        RECT 96.430 189.590 96.750 189.650 ;
        RECT 99.665 189.590 99.955 189.635 ;
        RECT 101.045 189.590 101.335 189.635 ;
        RECT 107.010 189.590 107.330 189.650 ;
        RECT 140.145 189.590 140.435 189.635 ;
        RECT 96.430 189.450 98.960 189.590 ;
        RECT 89.085 189.065 89.375 189.295 ;
        RECT 89.530 189.050 89.850 189.310 ;
        RECT 89.990 189.295 90.310 189.310 ;
        RECT 89.990 189.250 90.395 189.295 ;
        RECT 90.540 189.250 90.680 189.450 ;
        RECT 96.430 189.390 96.750 189.450 ;
        RECT 98.270 189.250 98.590 189.310 ;
        RECT 98.820 189.295 98.960 189.450 ;
        RECT 99.665 189.450 101.335 189.590 ;
        RECT 99.665 189.405 99.955 189.450 ;
        RECT 101.045 189.405 101.335 189.450 ;
        RECT 101.580 189.450 107.330 189.590 ;
        RECT 89.990 189.110 90.680 189.250 ;
        RECT 91.920 189.110 98.590 189.250 ;
        RECT 89.990 189.065 90.395 189.110 ;
        RECT 89.990 189.050 90.310 189.065 ;
        RECT 88.610 188.910 88.930 188.970 ;
        RECT 85.940 188.770 88.930 188.910 ;
        RECT 78.045 188.725 78.335 188.770 ;
        RECT 79.870 188.710 80.190 188.770 ;
        RECT 88.610 188.710 88.930 188.770 ;
        RECT 78.505 188.570 78.795 188.615 ;
        RECT 76.740 188.430 78.795 188.570 ;
        RECT 76.740 188.290 76.880 188.430 ;
        RECT 78.505 188.385 78.795 188.430 ;
        RECT 79.410 188.570 79.730 188.630 ;
        RECT 91.920 188.570 92.060 189.110 ;
        RECT 98.270 189.050 98.590 189.110 ;
        RECT 98.745 189.065 99.035 189.295 ;
        RECT 99.190 189.250 99.510 189.310 ;
        RECT 101.580 189.295 101.720 189.450 ;
        RECT 107.010 189.390 107.330 189.450 ;
        RECT 117.680 189.450 140.435 189.590 ;
        RECT 117.680 189.310 117.820 189.450 ;
        RECT 140.145 189.405 140.435 189.450 ;
        RECT 141.140 189.450 143.810 189.590 ;
        RECT 100.125 189.250 100.415 189.295 ;
        RECT 99.190 189.110 100.415 189.250 ;
        RECT 99.190 189.050 99.510 189.110 ;
        RECT 100.125 189.065 100.415 189.110 ;
        RECT 100.585 189.065 100.875 189.295 ;
        RECT 101.505 189.065 101.795 189.295 ;
        RECT 103.330 189.250 103.650 189.310 ;
        RECT 104.710 189.250 105.030 189.310 ;
        RECT 103.330 189.110 105.030 189.250 ;
        RECT 96.890 188.710 97.210 188.970 ;
        RECT 100.660 188.910 100.800 189.065 ;
        RECT 103.330 189.050 103.650 189.110 ;
        RECT 104.710 189.050 105.030 189.110 ;
        RECT 105.630 189.050 105.950 189.310 ;
        RECT 107.485 189.250 107.775 189.295 ;
        RECT 113.450 189.250 113.770 189.310 ;
        RECT 116.670 189.250 116.990 189.310 ;
        RECT 107.485 189.110 111.380 189.250 ;
        RECT 107.485 189.065 107.775 189.110 ;
        RECT 105.720 188.910 105.860 189.050 ;
        RECT 111.240 188.970 111.380 189.110 ;
        RECT 113.450 189.110 116.990 189.250 ;
        RECT 113.450 189.050 113.770 189.110 ;
        RECT 116.670 189.050 116.990 189.110 ;
        RECT 117.590 189.050 117.910 189.310 ;
        RECT 118.755 189.250 119.045 189.295 ;
        RECT 118.755 189.110 120.580 189.250 ;
        RECT 118.755 189.065 119.045 189.110 ;
        RECT 100.660 188.770 105.860 188.910 ;
        RECT 111.150 188.710 111.470 188.970 ;
        RECT 114.370 188.910 114.690 188.970 ;
        RECT 116.210 188.910 116.530 188.970 ;
        RECT 118.065 188.910 118.355 188.955 ;
        RECT 114.370 188.770 118.355 188.910 ;
        RECT 114.370 188.710 114.690 188.770 ;
        RECT 116.210 188.710 116.530 188.770 ;
        RECT 118.065 188.725 118.355 188.770 ;
        RECT 119.890 188.710 120.210 188.970 ;
        RECT 120.440 188.910 120.580 189.110 ;
        RECT 120.810 189.050 121.130 189.310 ;
        RECT 122.190 189.050 122.510 189.310 ;
        RECT 124.950 189.250 125.270 189.310 ;
        RECT 130.945 189.250 131.235 189.295 ;
        RECT 124.950 189.110 131.235 189.250 ;
        RECT 124.950 189.050 125.270 189.110 ;
        RECT 130.945 189.065 131.235 189.110 ;
        RECT 132.310 189.250 132.630 189.310 ;
        RECT 135.545 189.250 135.835 189.295 ;
        RECT 132.310 189.110 135.835 189.250 ;
        RECT 122.280 188.910 122.420 189.050 ;
        RECT 120.440 188.770 122.420 188.910 ;
        RECT 130.010 188.710 130.330 188.970 ;
        RECT 131.020 188.910 131.160 189.065 ;
        RECT 132.310 189.050 132.630 189.110 ;
        RECT 135.545 189.065 135.835 189.110 ;
        RECT 139.685 189.065 139.975 189.295 ;
        RECT 132.770 188.910 133.090 188.970 ;
        RECT 131.020 188.770 133.090 188.910 ;
        RECT 132.770 188.710 133.090 188.770 ;
        RECT 133.690 188.910 134.010 188.970 ;
        RECT 134.625 188.910 134.915 188.955 ;
        RECT 133.690 188.770 134.915 188.910 ;
        RECT 133.690 188.710 134.010 188.770 ;
        RECT 134.625 188.725 134.915 188.770 ;
        RECT 79.410 188.430 92.060 188.570 ;
        RECT 92.290 188.570 92.610 188.630 ;
        RECT 96.980 188.570 97.120 188.710 ;
        RECT 98.745 188.570 99.035 188.615 ;
        RECT 139.210 188.570 139.530 188.630 ;
        RECT 139.760 188.570 139.900 189.065 ;
        RECT 92.290 188.430 95.280 188.570 ;
        RECT 96.980 188.430 99.035 188.570 ;
        RECT 79.410 188.370 79.730 188.430 ;
        RECT 92.290 188.370 92.610 188.430 ;
        RECT 44.080 188.090 47.900 188.230 ;
        RECT 49.050 188.230 49.370 188.290 ;
        RECT 49.525 188.230 49.815 188.275 ;
        RECT 53.650 188.230 53.970 188.290 ;
        RECT 49.050 188.090 53.970 188.230 ;
        RECT 38.930 188.030 39.250 188.090 ;
        RECT 40.325 188.045 40.615 188.090 ;
        RECT 43.530 188.030 43.850 188.090 ;
        RECT 49.050 188.030 49.370 188.090 ;
        RECT 49.525 188.045 49.815 188.090 ;
        RECT 53.650 188.030 53.970 188.090 ;
        RECT 56.870 188.030 57.190 188.290 ;
        RECT 61.010 188.230 61.330 188.290 ;
        RECT 65.610 188.230 65.930 188.290 ;
        RECT 61.010 188.090 65.930 188.230 ;
        RECT 61.010 188.030 61.330 188.090 ;
        RECT 65.610 188.030 65.930 188.090 ;
        RECT 66.085 188.230 66.375 188.275 ;
        RECT 69.750 188.230 70.070 188.290 ;
        RECT 66.085 188.090 70.070 188.230 ;
        RECT 66.085 188.045 66.375 188.090 ;
        RECT 69.750 188.030 70.070 188.090 ;
        RECT 72.970 188.030 73.290 188.290 ;
        RECT 74.810 188.230 75.130 188.290 ;
        RECT 75.285 188.230 75.575 188.275 ;
        RECT 76.650 188.230 76.970 188.290 ;
        RECT 74.810 188.090 76.970 188.230 ;
        RECT 74.810 188.030 75.130 188.090 ;
        RECT 75.285 188.045 75.575 188.090 ;
        RECT 76.650 188.030 76.970 188.090 ;
        RECT 77.570 188.030 77.890 188.290 ;
        RECT 82.170 188.230 82.490 188.290 ;
        RECT 83.090 188.230 83.410 188.290 ;
        RECT 82.170 188.090 83.410 188.230 ;
        RECT 82.170 188.030 82.490 188.090 ;
        RECT 83.090 188.030 83.410 188.090 ;
        RECT 84.945 188.230 85.235 188.275 ;
        RECT 87.690 188.230 88.010 188.290 ;
        RECT 84.945 188.090 88.010 188.230 ;
        RECT 95.140 188.230 95.280 188.430 ;
        RECT 98.745 188.385 99.035 188.430 ;
        RECT 99.740 188.430 139.900 188.570 ;
        RECT 99.740 188.230 99.880 188.430 ;
        RECT 139.210 188.370 139.530 188.430 ;
        RECT 95.140 188.090 99.880 188.230 ;
        RECT 102.870 188.230 103.190 188.290 ;
        RECT 106.550 188.230 106.870 188.290 ;
        RECT 102.870 188.090 106.870 188.230 ;
        RECT 84.945 188.045 85.235 188.090 ;
        RECT 87.690 188.030 88.010 188.090 ;
        RECT 102.870 188.030 103.190 188.090 ;
        RECT 106.550 188.030 106.870 188.090 ;
        RECT 107.010 188.230 107.330 188.290 ;
        RECT 113.910 188.230 114.230 188.290 ;
        RECT 107.010 188.090 114.230 188.230 ;
        RECT 107.010 188.030 107.330 188.090 ;
        RECT 113.910 188.030 114.230 188.090 ;
        RECT 117.130 188.230 117.450 188.290 ;
        RECT 129.550 188.230 129.870 188.290 ;
        RECT 134.610 188.230 134.930 188.290 ;
        RECT 117.130 188.090 134.930 188.230 ;
        RECT 117.130 188.030 117.450 188.090 ;
        RECT 129.550 188.030 129.870 188.090 ;
        RECT 134.610 188.030 134.930 188.090 ;
        RECT 136.450 188.030 136.770 188.290 ;
        RECT 140.220 188.230 140.360 189.405 ;
        RECT 141.140 188.970 141.280 189.450 ;
        RECT 141.510 189.250 141.830 189.310 ;
        RECT 142.905 189.250 143.195 189.295 ;
        RECT 141.510 189.110 143.195 189.250 ;
        RECT 143.670 189.250 143.810 189.450 ;
        RECT 145.205 189.250 145.495 189.295 ;
        RECT 145.650 189.250 145.970 189.310 ;
        RECT 143.670 189.110 144.960 189.250 ;
        RECT 141.510 189.050 141.830 189.110 ;
        RECT 142.905 189.065 143.195 189.110 ;
        RECT 141.050 188.710 141.370 188.970 ;
        RECT 141.970 188.710 142.290 188.970 ;
        RECT 142.445 188.725 142.735 188.955 ;
        RECT 143.365 188.910 143.655 188.955 ;
        RECT 144.270 188.910 144.590 188.970 ;
        RECT 143.365 188.770 144.590 188.910 ;
        RECT 144.820 188.910 144.960 189.110 ;
        RECT 145.205 189.110 145.970 189.250 ;
        RECT 145.205 189.065 145.495 189.110 ;
        RECT 145.650 189.050 145.970 189.110 ;
        RECT 146.125 188.910 146.415 188.955 ;
        RECT 144.820 188.770 146.415 188.910 ;
        RECT 143.365 188.725 143.655 188.770 ;
        RECT 141.140 188.570 141.280 188.710 ;
        RECT 142.520 188.570 142.660 188.725 ;
        RECT 144.270 188.710 144.590 188.770 ;
        RECT 146.125 188.725 146.415 188.770 ;
        RECT 141.140 188.430 142.660 188.570 ;
        RECT 147.030 188.230 147.350 188.290 ;
        RECT 140.220 188.090 147.350 188.230 ;
        RECT 147.030 188.030 147.350 188.090 ;
        RECT 36.100 187.410 150.180 187.890 ;
        RECT 45.845 187.210 46.135 187.255 ;
        RECT 46.290 187.210 46.610 187.270 ;
        RECT 45.845 187.070 46.610 187.210 ;
        RECT 45.845 187.025 46.135 187.070 ;
        RECT 46.290 187.010 46.610 187.070 ;
        RECT 49.510 187.010 49.830 187.270 ;
        RECT 50.445 187.025 50.735 187.255 ;
        RECT 61.010 187.210 61.330 187.270 ;
        RECT 60.180 187.070 61.330 187.210 ;
        RECT 47.225 186.870 47.515 186.915 ;
        RECT 50.520 186.870 50.660 187.025 ;
        RECT 45.000 186.730 50.660 186.870 ;
        RECT 45.000 186.250 45.140 186.730 ;
        RECT 47.225 186.685 47.515 186.730 ;
        RECT 52.730 186.530 53.050 186.590 ;
        RECT 46.840 186.390 53.050 186.530 ;
        RECT 44.910 185.990 45.230 186.250 ;
        RECT 45.370 186.190 45.690 186.250 ;
        RECT 46.840 186.235 46.980 186.390 ;
        RECT 52.730 186.330 53.050 186.390 ;
        RECT 59.185 186.530 59.475 186.575 ;
        RECT 60.180 186.530 60.320 187.070 ;
        RECT 61.010 187.010 61.330 187.070 ;
        RECT 62.865 187.210 63.155 187.255 ;
        RECT 64.245 187.210 64.535 187.255 ;
        RECT 62.865 187.070 64.535 187.210 ;
        RECT 62.865 187.025 63.155 187.070 ;
        RECT 64.245 187.025 64.535 187.070 ;
        RECT 65.165 187.210 65.455 187.255 ;
        RECT 67.465 187.210 67.755 187.255 ;
        RECT 65.165 187.070 67.755 187.210 ;
        RECT 65.165 187.025 65.455 187.070 ;
        RECT 67.465 187.025 67.755 187.070 ;
        RECT 67.910 187.210 68.230 187.270 ;
        RECT 91.370 187.210 91.690 187.270 ;
        RECT 67.910 187.070 91.690 187.210 ;
        RECT 67.910 187.010 68.230 187.070 ;
        RECT 91.370 187.010 91.690 187.070 ;
        RECT 93.210 187.210 93.530 187.270 ;
        RECT 107.010 187.210 107.330 187.270 ;
        RECT 93.210 187.070 107.330 187.210 ;
        RECT 93.210 187.010 93.530 187.070 ;
        RECT 107.010 187.010 107.330 187.070 ;
        RECT 108.020 187.070 109.080 187.210 ;
        RECT 60.550 186.670 60.870 186.930 ;
        RECT 62.405 186.870 62.695 186.915 ;
        RECT 66.545 186.870 66.835 186.915 ;
        RECT 62.405 186.730 66.835 186.870 ;
        RECT 62.405 186.685 62.695 186.730 ;
        RECT 66.545 186.685 66.835 186.730 ;
        RECT 74.365 186.870 74.655 186.915 ;
        RECT 75.770 186.870 76.060 186.915 ;
        RECT 77.870 186.870 78.160 186.915 ;
        RECT 79.440 186.870 79.730 186.915 ;
        RECT 102.195 186.870 102.485 186.915 ;
        RECT 74.365 186.730 75.445 186.870 ;
        RECT 74.365 186.685 74.655 186.730 ;
        RECT 59.185 186.390 60.320 186.530 ;
        RECT 61.025 186.530 61.315 186.575 ;
        RECT 61.945 186.530 62.235 186.575 ;
        RECT 67.005 186.530 67.295 186.575 ;
        RECT 61.025 186.390 67.295 186.530 ;
        RECT 59.185 186.345 59.475 186.390 ;
        RECT 61.025 186.345 61.315 186.390 ;
        RECT 61.945 186.345 62.235 186.390 ;
        RECT 46.765 186.190 47.055 186.235 ;
        RECT 45.370 186.050 47.055 186.190 ;
        RECT 45.370 185.990 45.690 186.050 ;
        RECT 46.765 186.005 47.055 186.050 ;
        RECT 47.685 186.005 47.975 186.235 ;
        RECT 48.145 186.190 48.435 186.235 ;
        RECT 49.050 186.190 49.370 186.250 ;
        RECT 48.145 186.050 49.370 186.190 ;
        RECT 48.145 186.005 48.435 186.050 ;
        RECT 47.760 185.850 47.900 186.005 ;
        RECT 49.050 185.990 49.370 186.050 ;
        RECT 49.510 185.990 49.830 186.250 ;
        RECT 50.445 186.005 50.735 186.235 ;
        RECT 49.600 185.850 49.740 185.990 ;
        RECT 47.760 185.710 49.740 185.850 ;
        RECT 50.520 185.850 50.660 186.005 ;
        RECT 50.890 185.990 51.210 186.250 ;
        RECT 54.110 186.190 54.430 186.250 ;
        RECT 56.870 186.190 57.190 186.250 ;
        RECT 51.440 186.050 57.190 186.190 ;
        RECT 51.440 185.850 51.580 186.050 ;
        RECT 54.110 185.990 54.430 186.050 ;
        RECT 56.870 185.990 57.190 186.050 ;
        RECT 58.250 185.990 58.570 186.250 ;
        RECT 58.725 186.005 59.015 186.235 ;
        RECT 50.520 185.710 51.580 185.850 ;
        RECT 51.825 185.850 52.115 185.895 ;
        RECT 52.730 185.850 53.050 185.910 ;
        RECT 51.825 185.710 53.050 185.850 ;
        RECT 51.825 185.665 52.115 185.710 ;
        RECT 52.730 185.650 53.050 185.710 ;
        RECT 44.450 185.510 44.770 185.570 ;
        RECT 49.050 185.510 49.370 185.570 ;
        RECT 44.450 185.370 49.370 185.510 ;
        RECT 58.800 185.510 58.940 186.005 ;
        RECT 59.630 185.990 59.950 186.250 ;
        RECT 62.480 186.190 62.620 186.390 ;
        RECT 67.005 186.345 67.295 186.390 ;
        RECT 69.750 186.530 70.070 186.590 ;
        RECT 75.305 186.530 75.445 186.730 ;
        RECT 75.770 186.730 79.730 186.870 ;
        RECT 75.770 186.685 76.060 186.730 ;
        RECT 77.870 186.685 78.160 186.730 ;
        RECT 79.440 186.685 79.730 186.730 ;
        RECT 94.220 186.730 102.485 186.870 ;
        RECT 94.220 186.590 94.360 186.730 ;
        RECT 102.195 186.685 102.485 186.730 ;
        RECT 76.165 186.530 76.455 186.575 ;
        RECT 77.355 186.530 77.645 186.575 ;
        RECT 79.875 186.530 80.165 186.575 ;
        RECT 69.750 186.390 74.580 186.530 ;
        RECT 75.305 186.390 75.960 186.530 ;
        RECT 69.750 186.330 70.070 186.390 ;
        RECT 60.180 186.050 62.620 186.190 ;
        RECT 60.180 185.910 60.320 186.050 ;
        RECT 62.850 185.990 63.170 186.250 ;
        RECT 65.610 185.990 65.930 186.250 ;
        RECT 73.445 186.190 73.735 186.235 ;
        RECT 73.890 186.190 74.210 186.250 ;
        RECT 60.090 185.650 60.410 185.910 ;
        RECT 61.945 185.850 62.235 185.895 ;
        RECT 62.940 185.850 63.080 185.990 ;
        RECT 73.000 185.910 73.290 186.125 ;
        RECT 73.445 186.050 74.210 186.190 ;
        RECT 74.440 186.190 74.580 186.390 ;
        RECT 75.285 186.190 75.575 186.235 ;
        RECT 74.440 186.050 75.575 186.190 ;
        RECT 75.820 186.190 75.960 186.390 ;
        RECT 76.165 186.390 80.165 186.530 ;
        RECT 76.165 186.345 76.455 186.390 ;
        RECT 77.355 186.345 77.645 186.390 ;
        RECT 79.875 186.345 80.165 186.390 ;
        RECT 94.130 186.330 94.450 186.590 ;
        RECT 95.510 186.530 95.830 186.590 ;
        RECT 94.680 186.390 95.830 186.530 ;
        RECT 76.565 186.190 76.855 186.235 ;
        RECT 75.820 186.050 76.855 186.190 ;
        RECT 73.445 186.005 73.735 186.050 ;
        RECT 73.890 185.990 74.210 186.050 ;
        RECT 75.285 186.005 75.575 186.050 ;
        RECT 76.565 186.005 76.855 186.050 ;
        RECT 78.030 186.190 78.350 186.250 ;
        RECT 81.710 186.190 82.030 186.250 ;
        RECT 78.030 186.050 82.030 186.190 ;
        RECT 78.030 185.990 78.350 186.050 ;
        RECT 81.710 185.990 82.030 186.050 ;
        RECT 84.470 186.190 84.790 186.250 ;
        RECT 94.680 186.235 94.820 186.390 ;
        RECT 95.510 186.330 95.830 186.390 ;
        RECT 95.985 186.530 96.275 186.575 ;
        RECT 97.810 186.530 98.130 186.590 ;
        RECT 98.730 186.530 99.050 186.590 ;
        RECT 95.985 186.390 99.050 186.530 ;
        RECT 95.985 186.345 96.275 186.390 ;
        RECT 97.810 186.330 98.130 186.390 ;
        RECT 98.730 186.330 99.050 186.390 ;
        RECT 99.190 186.530 99.510 186.590 ;
        RECT 100.570 186.530 100.890 186.590 ;
        RECT 99.190 186.390 100.890 186.530 ;
        RECT 99.190 186.330 99.510 186.390 ;
        RECT 100.570 186.330 100.890 186.390 ;
        RECT 101.045 186.530 101.335 186.575 ;
        RECT 103.330 186.530 103.650 186.590 ;
        RECT 101.045 186.390 103.650 186.530 ;
        RECT 101.045 186.345 101.335 186.390 ;
        RECT 103.330 186.330 103.650 186.390 ;
        RECT 88.625 186.190 88.915 186.235 ;
        RECT 94.605 186.190 94.895 186.235 ;
        RECT 101.950 186.190 102.270 186.250 ;
        RECT 108.020 186.190 108.160 187.070 ;
        RECT 108.390 186.670 108.710 186.930 ;
        RECT 108.940 186.870 109.080 187.070 ;
        RECT 117.130 187.010 117.450 187.270 ;
        RECT 118.510 187.210 118.830 187.270 ;
        RECT 120.365 187.210 120.655 187.255 ;
        RECT 118.510 187.070 120.655 187.210 ;
        RECT 118.510 187.010 118.830 187.070 ;
        RECT 120.365 187.025 120.655 187.070 ;
        RECT 121.730 187.210 122.050 187.270 ;
        RECT 127.725 187.210 128.015 187.255 ;
        RECT 121.730 187.070 128.015 187.210 ;
        RECT 121.730 187.010 122.050 187.070 ;
        RECT 127.725 187.025 128.015 187.070 ;
        RECT 128.645 187.210 128.935 187.255 ;
        RECT 132.325 187.210 132.615 187.255 ;
        RECT 136.450 187.210 136.770 187.270 ;
        RECT 128.645 187.070 132.080 187.210 ;
        RECT 128.645 187.025 128.935 187.070 ;
        RECT 124.950 186.870 125.270 186.930 ;
        RECT 131.940 186.870 132.080 187.070 ;
        RECT 132.325 187.070 136.770 187.210 ;
        RECT 132.325 187.025 132.615 187.070 ;
        RECT 136.450 187.010 136.770 187.070 ;
        RECT 139.210 187.010 139.530 187.270 ;
        RECT 140.130 187.210 140.450 187.270 ;
        RECT 141.985 187.210 142.275 187.255 ;
        RECT 140.130 187.070 142.275 187.210 ;
        RECT 140.130 187.010 140.450 187.070 ;
        RECT 141.985 187.025 142.275 187.070 ;
        RECT 143.810 187.010 144.130 187.270 ;
        RECT 144.270 187.210 144.590 187.270 ;
        RECT 145.650 187.210 145.970 187.270 ;
        RECT 146.125 187.210 146.415 187.255 ;
        RECT 144.270 187.070 145.420 187.210 ;
        RECT 144.270 187.010 144.590 187.070 ;
        RECT 132.770 186.870 133.090 186.930 ;
        RECT 108.940 186.730 113.220 186.870 ;
        RECT 108.480 186.530 108.620 186.670 ;
        RECT 113.080 186.590 113.220 186.730 ;
        RECT 116.300 186.730 124.720 186.870 ;
        RECT 109.785 186.530 110.075 186.575 ;
        RECT 108.480 186.390 110.075 186.530 ;
        RECT 109.785 186.345 110.075 186.390 ;
        RECT 111.625 186.345 111.915 186.575 ;
        RECT 84.470 186.050 87.920 186.190 ;
        RECT 84.470 185.990 84.790 186.050 ;
        RECT 61.945 185.710 63.080 185.850 ;
        RECT 61.945 185.665 62.235 185.710 ;
        RECT 63.310 185.650 63.630 185.910 ;
        RECT 63.785 185.850 64.075 185.895 ;
        RECT 66.070 185.850 66.390 185.910 ;
        RECT 63.785 185.710 66.390 185.850 ;
        RECT 63.785 185.665 64.075 185.710 ;
        RECT 66.070 185.650 66.390 185.710 ;
        RECT 72.970 185.650 73.290 185.910 ;
        RECT 74.365 185.850 74.655 185.895 ;
        RECT 77.570 185.850 77.890 185.910 ;
        RECT 87.230 185.850 87.550 185.910 ;
        RECT 74.365 185.710 77.890 185.850 ;
        RECT 74.365 185.665 74.655 185.710 ;
        RECT 77.570 185.650 77.890 185.710 ;
        RECT 81.800 185.710 87.550 185.850 ;
        RECT 87.780 185.850 87.920 186.050 ;
        RECT 88.625 186.050 94.895 186.190 ;
        RECT 88.625 186.005 88.915 186.050 ;
        RECT 94.605 186.005 94.895 186.050 ;
        RECT 95.370 186.050 102.270 186.190 ;
        RECT 95.370 185.850 95.510 186.050 ;
        RECT 101.950 185.990 102.270 186.050 ;
        RECT 102.500 186.050 108.160 186.190 ;
        RECT 87.780 185.710 95.510 185.850 ;
        RECT 98.730 185.850 99.050 185.910 ;
        RECT 102.500 185.850 102.640 186.050 ;
        RECT 108.405 186.005 108.695 186.235 ;
        RECT 110.245 186.190 110.535 186.235 ;
        RECT 111.150 186.190 111.470 186.250 ;
        RECT 110.245 186.050 111.470 186.190 ;
        RECT 110.245 186.005 110.535 186.050 ;
        RECT 98.730 185.710 102.640 185.850 ;
        RECT 104.250 185.850 104.570 185.910 ;
        RECT 108.480 185.850 108.620 186.005 ;
        RECT 111.150 185.990 111.470 186.050 ;
        RECT 111.700 185.910 111.840 186.345 ;
        RECT 112.990 186.330 113.310 186.590 ;
        RECT 116.300 186.235 116.440 186.730 ;
        RECT 124.580 186.530 124.720 186.730 ;
        RECT 124.950 186.730 131.160 186.870 ;
        RECT 131.940 186.730 133.090 186.870 ;
        RECT 124.950 186.670 125.270 186.730 ;
        RECT 126.330 186.530 126.650 186.590 ;
        RECT 124.580 186.390 126.650 186.530 ;
        RECT 115.305 186.005 115.595 186.235 ;
        RECT 116.225 186.005 116.515 186.235 ;
        RECT 116.670 186.190 116.990 186.250 ;
        RECT 117.145 186.190 117.435 186.235 ;
        RECT 116.670 186.050 117.435 186.190 ;
        RECT 104.250 185.710 108.620 185.850 ;
        RECT 62.850 185.510 63.170 185.570 ;
        RECT 67.465 185.510 67.755 185.555 ;
        RECT 58.800 185.370 67.755 185.510 ;
        RECT 44.450 185.310 44.770 185.370 ;
        RECT 49.050 185.310 49.370 185.370 ;
        RECT 62.850 185.310 63.170 185.370 ;
        RECT 67.465 185.325 67.755 185.370 ;
        RECT 68.385 185.510 68.675 185.555 ;
        RECT 81.800 185.510 81.940 185.710 ;
        RECT 87.230 185.650 87.550 185.710 ;
        RECT 98.730 185.650 99.050 185.710 ;
        RECT 104.250 185.650 104.570 185.710 ;
        RECT 111.610 185.650 111.930 185.910 ;
        RECT 68.385 185.370 81.940 185.510 ;
        RECT 68.385 185.325 68.675 185.370 ;
        RECT 82.170 185.310 82.490 185.570 ;
        RECT 87.705 185.510 87.995 185.555 ;
        RECT 88.150 185.510 88.470 185.570 ;
        RECT 87.705 185.370 88.470 185.510 ;
        RECT 87.705 185.325 87.995 185.370 ;
        RECT 88.150 185.310 88.470 185.370 ;
        RECT 89.990 185.510 90.310 185.570 ;
        RECT 112.530 185.510 112.850 185.570 ;
        RECT 89.990 185.370 112.850 185.510 ;
        RECT 115.380 185.510 115.520 186.005 ;
        RECT 116.670 185.990 116.990 186.050 ;
        RECT 117.145 186.005 117.435 186.050 ;
        RECT 118.985 186.175 119.275 186.235 ;
        RECT 122.650 186.190 122.970 186.250 ;
        RECT 124.580 186.235 124.720 186.390 ;
        RECT 126.330 186.330 126.650 186.390 ;
        RECT 129.090 186.330 129.410 186.590 ;
        RECT 131.020 186.575 131.160 186.730 ;
        RECT 132.770 186.670 133.090 186.730 ;
        RECT 133.245 186.870 133.535 186.915 ;
        RECT 135.990 186.870 136.310 186.930 ;
        RECT 143.350 186.870 143.670 186.930 ;
        RECT 133.245 186.730 136.310 186.870 ;
        RECT 133.245 186.685 133.535 186.730 ;
        RECT 135.990 186.670 136.310 186.730 ;
        RECT 139.760 186.730 143.670 186.870 ;
        RECT 130.945 186.345 131.235 186.575 ;
        RECT 133.690 186.330 134.010 186.590 ;
        RECT 139.760 186.575 139.900 186.730 ;
        RECT 143.350 186.670 143.670 186.730 ;
        RECT 139.685 186.345 139.975 186.575 ;
        RECT 143.900 186.530 144.040 187.010 ;
        RECT 145.280 186.915 145.420 187.070 ;
        RECT 145.650 187.070 146.415 187.210 ;
        RECT 145.650 187.010 145.970 187.070 ;
        RECT 146.125 187.025 146.415 187.070 ;
        RECT 145.205 186.685 145.495 186.915 ;
        RECT 140.680 186.390 144.040 186.530 ;
        RECT 144.745 186.530 145.035 186.575 ;
        RECT 145.740 186.530 145.880 187.010 ;
        RECT 144.745 186.390 145.880 186.530 ;
        RECT 119.520 186.175 123.340 186.190 ;
        RECT 118.985 186.050 123.340 186.175 ;
        RECT 118.985 186.035 119.660 186.050 ;
        RECT 118.985 186.005 119.275 186.035 ;
        RECT 122.650 185.990 122.970 186.050 ;
        RECT 117.590 185.850 117.910 185.910 ;
        RECT 123.200 185.895 123.340 186.050 ;
        RECT 124.505 186.005 124.795 186.235 ;
        RECT 130.025 186.005 130.315 186.235 ;
        RECT 133.780 186.115 133.920 186.330 ;
        RECT 137.370 186.190 137.690 186.250 ;
        RECT 138.305 186.190 138.595 186.235 ;
        RECT 132.770 186.065 133.090 186.080 ;
        RECT 130.100 185.930 130.310 186.005 ;
        RECT 117.590 185.710 122.880 185.850 ;
        RECT 117.590 185.650 117.910 185.710 ;
        RECT 117.130 185.510 117.450 185.570 ;
        RECT 115.380 185.370 117.450 185.510 ;
        RECT 89.990 185.310 90.310 185.370 ;
        RECT 112.530 185.310 112.850 185.370 ;
        RECT 117.130 185.310 117.450 185.370 ;
        RECT 119.430 185.510 119.750 185.570 ;
        RECT 121.285 185.510 121.575 185.555 ;
        RECT 119.430 185.370 121.575 185.510 ;
        RECT 119.430 185.310 119.750 185.370 ;
        RECT 121.285 185.325 121.575 185.370 ;
        RECT 121.730 185.310 122.050 185.570 ;
        RECT 122.190 185.310 122.510 185.570 ;
        RECT 122.740 185.510 122.880 185.710 ;
        RECT 123.125 185.665 123.415 185.895 ;
        RECT 123.585 185.665 123.875 185.895 ;
        RECT 123.660 185.510 123.800 185.665 ;
        RECT 126.790 185.650 127.110 185.910 ;
        RECT 122.740 185.370 123.800 185.510 ;
        RECT 124.030 185.510 124.350 185.570 ;
        RECT 125.425 185.510 125.715 185.555 ;
        RECT 127.250 185.510 127.570 185.570 ;
        RECT 124.030 185.370 127.570 185.510 ;
        RECT 124.030 185.310 124.350 185.370 ;
        RECT 125.425 185.325 125.715 185.370 ;
        RECT 127.250 185.310 127.570 185.370 ;
        RECT 127.710 185.555 128.030 185.570 ;
        RECT 127.710 185.325 128.095 185.555 ;
        RECT 130.170 185.510 130.310 185.930 ;
        RECT 130.930 185.850 131.250 185.910 ;
        RECT 131.405 185.850 131.695 185.895 ;
        RECT 130.930 185.710 131.695 185.850 ;
        RECT 132.555 185.835 133.090 186.065 ;
        RECT 133.705 185.885 133.995 186.115 ;
        RECT 137.370 186.050 138.595 186.190 ;
        RECT 137.370 185.990 137.690 186.050 ;
        RECT 138.305 186.005 138.595 186.050 ;
        RECT 138.750 185.990 139.070 186.250 ;
        RECT 140.680 186.235 140.820 186.390 ;
        RECT 144.745 186.345 145.035 186.390 ;
        RECT 140.435 186.050 140.820 186.235 ;
        RECT 140.435 186.005 140.725 186.050 ;
        RECT 141.065 186.005 141.355 186.235 ;
        RECT 141.510 186.190 141.830 186.250 ;
        RECT 142.445 186.190 142.735 186.235 ;
        RECT 141.510 186.050 142.735 186.190 ;
        RECT 132.770 185.820 133.090 185.835 ;
        RECT 130.930 185.650 131.250 185.710 ;
        RECT 131.405 185.665 131.695 185.710 ;
        RECT 133.230 185.510 133.550 185.570 ;
        RECT 134.625 185.510 134.915 185.555 ;
        RECT 130.170 185.370 134.915 185.510 ;
        RECT 127.710 185.310 128.030 185.325 ;
        RECT 133.230 185.310 133.550 185.370 ;
        RECT 134.625 185.325 134.915 185.370 ;
        RECT 136.910 185.310 137.230 185.570 ;
        RECT 141.140 185.510 141.280 186.005 ;
        RECT 141.510 185.990 141.830 186.050 ;
        RECT 142.445 186.005 142.735 186.050 ;
        RECT 142.905 186.005 143.195 186.235 ;
        RECT 143.365 186.190 143.655 186.235 ;
        RECT 144.270 186.190 144.590 186.250 ;
        RECT 147.490 186.190 147.810 186.250 ;
        RECT 143.365 186.050 147.810 186.190 ;
        RECT 143.365 186.005 143.655 186.050 ;
        RECT 142.980 185.850 143.120 186.005 ;
        RECT 144.270 185.990 144.590 186.050 ;
        RECT 147.490 185.990 147.810 186.050 ;
        RECT 143.810 185.850 144.130 185.910 ;
        RECT 142.980 185.710 144.130 185.850 ;
        RECT 143.810 185.650 144.130 185.710 ;
        RECT 147.030 185.650 147.350 185.910 ;
        RECT 141.510 185.510 141.830 185.570 ;
        RECT 141.140 185.370 141.830 185.510 ;
        RECT 141.510 185.310 141.830 185.370 ;
        RECT 143.350 185.510 143.670 185.570 ;
        RECT 145.995 185.510 146.285 185.555 ;
        RECT 143.350 185.370 146.285 185.510 ;
        RECT 143.350 185.310 143.670 185.370 ;
        RECT 145.995 185.325 146.285 185.370 ;
        RECT 36.100 184.690 150.180 185.170 ;
        RECT 44.465 184.305 44.755 184.535 ;
        RECT 50.890 184.490 51.210 184.550 ;
        RECT 47.070 184.350 51.210 184.490 ;
        RECT 44.540 184.150 44.680 184.305 ;
        RECT 47.070 184.150 47.210 184.350 ;
        RECT 50.890 184.290 51.210 184.350 ;
        RECT 52.745 184.305 53.035 184.535 ;
        RECT 59.630 184.490 59.950 184.550 ;
        RECT 60.105 184.490 60.395 184.535 ;
        RECT 78.030 184.490 78.350 184.550 ;
        RECT 59.630 184.350 60.395 184.490 ;
        RECT 51.350 184.150 51.670 184.210 ;
        RECT 44.540 184.010 47.210 184.150 ;
        RECT 48.680 184.010 51.670 184.150 ;
        RECT 43.085 183.625 43.375 183.855 ;
        RECT 43.160 183.470 43.300 183.625 ;
        RECT 43.990 183.610 44.310 183.870 ;
        RECT 44.450 183.610 44.770 183.870 ;
        RECT 44.925 183.810 45.215 183.855 ;
        RECT 45.370 183.810 45.690 183.870 ;
        RECT 44.925 183.670 45.690 183.810 ;
        RECT 44.925 183.625 45.215 183.670 ;
        RECT 45.000 183.470 45.140 183.625 ;
        RECT 45.370 183.610 45.690 183.670 ;
        RECT 45.845 183.625 46.135 183.855 ;
        RECT 46.290 183.810 46.610 183.870 ;
        RECT 48.680 183.855 48.820 184.010 ;
        RECT 51.350 183.950 51.670 184.010 ;
        RECT 48.145 183.810 48.435 183.855 ;
        RECT 46.290 183.670 48.435 183.810 ;
        RECT 43.160 183.330 45.140 183.470 ;
        RECT 45.920 183.130 46.060 183.625 ;
        RECT 46.290 183.610 46.610 183.670 ;
        RECT 48.145 183.625 48.435 183.670 ;
        RECT 48.605 183.625 48.895 183.855 ;
        RECT 49.510 183.810 49.830 183.870 ;
        RECT 50.905 183.810 51.195 183.855 ;
        RECT 52.820 183.810 52.960 184.305 ;
        RECT 59.630 184.290 59.950 184.350 ;
        RECT 60.105 184.305 60.395 184.350 ;
        RECT 62.480 184.350 78.350 184.490 ;
        RECT 62.480 184.210 62.620 184.350 ;
        RECT 78.030 184.290 78.350 184.350 ;
        RECT 78.950 184.290 79.270 184.550 ;
        RECT 80.805 184.490 81.095 184.535 ;
        RECT 80.805 184.350 84.700 184.490 ;
        RECT 80.805 184.305 81.095 184.350 ;
        RECT 62.390 183.950 62.710 184.210 ;
        RECT 81.710 184.150 82.030 184.210 ;
        RECT 80.420 184.010 81.480 184.150 ;
        RECT 80.420 183.870 80.560 184.010 ;
        RECT 53.205 183.810 53.495 183.855 ;
        RECT 49.510 183.670 50.660 183.810 ;
        RECT 46.765 183.470 47.055 183.515 ;
        RECT 48.680 183.470 48.820 183.625 ;
        RECT 49.510 183.610 49.830 183.670 ;
        RECT 46.765 183.330 48.820 183.470 ;
        RECT 46.765 183.285 47.055 183.330 ;
        RECT 49.970 183.130 50.290 183.190 ;
        RECT 45.920 182.990 50.290 183.130 ;
        RECT 50.520 183.130 50.660 183.670 ;
        RECT 50.905 183.670 52.500 183.810 ;
        RECT 52.820 183.670 53.495 183.810 ;
        RECT 50.905 183.625 51.195 183.670 ;
        RECT 51.350 183.270 51.670 183.530 ;
        RECT 52.360 183.470 52.500 183.670 ;
        RECT 53.205 183.625 53.495 183.670 ;
        RECT 53.650 183.610 53.970 183.870 ;
        RECT 58.250 183.610 58.570 183.870 ;
        RECT 58.710 183.810 59.030 183.870 ;
        RECT 59.185 183.810 59.475 183.855 ;
        RECT 58.710 183.670 59.475 183.810 ;
        RECT 58.710 183.610 59.030 183.670 ;
        RECT 59.185 183.625 59.475 183.670 ;
        RECT 61.010 183.810 61.330 183.870 ;
        RECT 64.245 183.810 64.535 183.855 ;
        RECT 67.450 183.810 67.770 183.870 ;
        RECT 77.585 183.810 77.875 183.855 ;
        RECT 61.010 183.670 67.770 183.810 ;
        RECT 61.010 183.610 61.330 183.670 ;
        RECT 64.245 183.625 64.535 183.670 ;
        RECT 67.450 183.610 67.770 183.670 ;
        RECT 76.740 183.670 77.875 183.810 ;
        RECT 54.570 183.470 54.890 183.530 ;
        RECT 52.360 183.330 54.890 183.470 ;
        RECT 54.570 183.270 54.890 183.330 ;
        RECT 59.630 183.470 59.950 183.530 ;
        RECT 66.530 183.470 66.850 183.530 ;
        RECT 59.630 183.330 66.850 183.470 ;
        RECT 59.630 183.270 59.950 183.330 ;
        RECT 66.530 183.270 66.850 183.330 ;
        RECT 55.045 183.130 55.335 183.175 ;
        RECT 50.520 182.990 55.335 183.130 ;
        RECT 46.840 182.850 46.980 182.990 ;
        RECT 49.970 182.930 50.290 182.990 ;
        RECT 55.045 182.945 55.335 182.990 ;
        RECT 61.470 183.130 61.790 183.190 ;
        RECT 63.770 183.130 64.090 183.190 ;
        RECT 61.470 182.990 64.090 183.130 ;
        RECT 61.470 182.930 61.790 182.990 ;
        RECT 63.770 182.930 64.090 182.990 ;
        RECT 76.740 183.130 76.880 183.670 ;
        RECT 77.585 183.625 77.875 183.670 ;
        RECT 79.885 183.625 80.175 183.855 ;
        RECT 79.960 183.470 80.100 183.625 ;
        RECT 80.330 183.610 80.650 183.870 ;
        RECT 81.340 183.855 81.480 184.010 ;
        RECT 81.710 184.010 82.860 184.150 ;
        RECT 81.710 183.950 82.030 184.010 ;
        RECT 82.720 183.855 82.860 184.010 ;
        RECT 81.265 183.625 81.555 183.855 ;
        RECT 82.645 183.625 82.935 183.855 ;
        RECT 81.725 183.470 82.015 183.515 ;
        RECT 79.960 183.330 82.015 183.470 ;
        RECT 81.725 183.285 82.015 183.330 ;
        RECT 83.565 183.285 83.855 183.515 ;
        RECT 82.170 183.130 82.490 183.190 ;
        RECT 83.640 183.130 83.780 183.285 ;
        RECT 84.560 183.190 84.700 184.350 ;
        RECT 84.930 184.290 85.250 184.550 ;
        RECT 87.230 184.490 87.550 184.550 ;
        RECT 100.125 184.490 100.415 184.535 ;
        RECT 100.570 184.490 100.890 184.550 ;
        RECT 87.230 184.350 92.980 184.490 ;
        RECT 87.230 184.290 87.550 184.350 ;
        RECT 85.020 183.855 85.160 184.290 ;
        RECT 91.845 184.150 92.135 184.195 ;
        RECT 89.160 184.010 92.135 184.150 ;
        RECT 84.945 183.625 85.235 183.855 ;
        RECT 88.150 183.610 88.470 183.870 ;
        RECT 89.160 183.855 89.300 184.010 ;
        RECT 91.845 183.965 92.135 184.010 ;
        RECT 89.085 183.625 89.375 183.855 ;
        RECT 89.530 183.610 89.850 183.870 ;
        RECT 90.005 183.810 90.295 183.855 ;
        RECT 92.290 183.810 92.610 183.870 ;
        RECT 92.840 183.855 92.980 184.350 ;
        RECT 94.680 184.350 99.880 184.490 ;
        RECT 90.005 183.670 92.610 183.810 ;
        RECT 90.005 183.625 90.295 183.670 ;
        RECT 89.620 183.470 89.760 183.610 ;
        RECT 91.370 183.470 91.690 183.530 ;
        RECT 89.620 183.330 91.690 183.470 ;
        RECT 91.370 183.270 91.690 183.330 ;
        RECT 76.740 182.990 83.780 183.130 ;
        RECT 76.740 182.850 76.880 182.990 ;
        RECT 82.170 182.930 82.490 182.990 ;
        RECT 84.470 182.930 84.790 183.190 ;
        RECT 91.920 183.130 92.060 183.670 ;
        RECT 92.290 183.610 92.610 183.670 ;
        RECT 92.765 183.625 93.055 183.855 ;
        RECT 90.080 182.990 92.060 183.130 ;
        RECT 92.840 183.130 92.980 183.625 ;
        RECT 93.210 183.610 93.530 183.870 ;
        RECT 94.680 183.855 94.820 184.350 ;
        RECT 95.050 184.150 95.370 184.210 ;
        RECT 98.270 184.150 98.590 184.210 ;
        RECT 99.740 184.150 99.880 184.350 ;
        RECT 100.125 184.350 100.890 184.490 ;
        RECT 100.125 184.305 100.415 184.350 ;
        RECT 100.570 184.290 100.890 184.350 ;
        RECT 101.950 184.490 102.270 184.550 ;
        RECT 110.690 184.490 111.010 184.550 ;
        RECT 101.950 184.350 111.010 184.490 ;
        RECT 101.950 184.290 102.270 184.350 ;
        RECT 110.690 184.290 111.010 184.350 ;
        RECT 111.150 184.490 111.470 184.550 ;
        RECT 111.150 184.350 114.600 184.490 ;
        RECT 111.150 184.290 111.470 184.350 ;
        RECT 114.460 184.195 114.600 184.350 ;
        RECT 122.190 184.290 122.510 184.550 ;
        RECT 123.585 184.305 123.875 184.535 ;
        RECT 127.250 184.490 127.570 184.550 ;
        RECT 134.165 184.490 134.455 184.535 ;
        RECT 135.530 184.490 135.850 184.550 ;
        RECT 127.250 184.350 133.920 184.490 ;
        RECT 95.050 184.010 98.040 184.150 ;
        RECT 95.050 183.950 95.370 184.010 ;
        RECT 94.605 183.625 94.895 183.855 ;
        RECT 95.510 183.810 95.830 183.870 ;
        RECT 95.985 183.810 96.275 183.855 ;
        RECT 95.510 183.670 96.275 183.810 ;
        RECT 95.510 183.610 95.830 183.670 ;
        RECT 95.985 183.625 96.275 183.670 ;
        RECT 96.445 183.810 96.735 183.855 ;
        RECT 96.890 183.810 97.210 183.870 ;
        RECT 96.445 183.670 97.210 183.810 ;
        RECT 96.445 183.625 96.735 183.670 ;
        RECT 96.890 183.610 97.210 183.670 ;
        RECT 97.350 183.610 97.670 183.870 ;
        RECT 97.900 183.855 98.040 184.010 ;
        RECT 98.270 184.010 99.420 184.150 ;
        RECT 99.740 184.010 112.300 184.150 ;
        RECT 98.270 183.950 98.590 184.010 ;
        RECT 97.825 183.625 98.115 183.855 ;
        RECT 98.730 183.610 99.050 183.870 ;
        RECT 99.280 183.855 99.420 184.010 ;
        RECT 99.205 183.625 99.495 183.855 ;
        RECT 101.490 183.610 101.810 183.870 ;
        RECT 102.870 183.855 103.190 183.870 ;
        RECT 102.195 183.625 102.485 183.855 ;
        RECT 102.870 183.810 103.205 183.855 ;
        RECT 102.705 183.670 103.205 183.810 ;
        RECT 102.870 183.625 103.205 183.670 ;
        RECT 103.405 183.820 103.695 183.865 ;
        RECT 104.265 183.820 104.555 183.855 ;
        RECT 104.710 183.820 105.030 183.870 ;
        RECT 105.720 183.855 105.860 184.010 ;
        RECT 103.405 183.680 103.975 183.820 ;
        RECT 103.405 183.635 103.695 183.680 ;
        RECT 93.670 183.470 93.990 183.530 ;
        RECT 98.285 183.470 98.575 183.515 ;
        RECT 98.820 183.470 98.960 183.610 ;
        RECT 93.670 183.330 98.960 183.470 ;
        RECT 93.670 183.270 93.990 183.330 ;
        RECT 98.285 183.285 98.575 183.330 ;
        RECT 102.270 183.130 102.410 183.625 ;
        RECT 102.870 183.610 103.190 183.625 ;
        RECT 102.870 183.130 103.190 183.190 ;
        RECT 103.835 183.130 103.975 183.680 ;
        RECT 104.265 183.680 105.030 183.820 ;
        RECT 104.265 183.625 104.555 183.680 ;
        RECT 104.710 183.610 105.030 183.680 ;
        RECT 105.645 183.625 105.935 183.855 ;
        RECT 107.025 183.810 107.315 183.855 ;
        RECT 106.640 183.670 107.315 183.810 ;
        RECT 106.640 183.530 106.780 183.670 ;
        RECT 107.025 183.625 107.315 183.670 ;
        RECT 107.945 183.625 108.235 183.855 ;
        RECT 106.550 183.270 106.870 183.530 ;
        RECT 108.020 183.470 108.160 183.625 ;
        RECT 109.770 183.610 110.090 183.870 ;
        RECT 108.390 183.470 108.710 183.530 ;
        RECT 108.020 183.330 108.710 183.470 ;
        RECT 108.390 183.270 108.710 183.330 ;
        RECT 107.930 183.130 108.250 183.190 ;
        RECT 92.840 182.990 101.720 183.130 ;
        RECT 102.270 182.990 103.190 183.130 ;
        RECT 46.750 182.590 47.070 182.850 ;
        RECT 47.210 182.590 47.530 182.850 ;
        RECT 49.050 182.590 49.370 182.850 ;
        RECT 51.825 182.790 52.115 182.835 ;
        RECT 52.270 182.790 52.590 182.850 ;
        RECT 51.825 182.650 52.590 182.790 ;
        RECT 51.825 182.605 52.115 182.650 ;
        RECT 52.270 182.590 52.590 182.650 ;
        RECT 52.730 182.790 53.050 182.850 ;
        RECT 53.205 182.790 53.495 182.835 ;
        RECT 52.730 182.650 53.495 182.790 ;
        RECT 52.730 182.590 53.050 182.650 ;
        RECT 53.205 182.605 53.495 182.650 ;
        RECT 62.850 182.790 63.170 182.850 ;
        RECT 63.325 182.790 63.615 182.835 ;
        RECT 62.850 182.650 63.615 182.790 ;
        RECT 62.850 182.590 63.170 182.650 ;
        RECT 63.325 182.605 63.615 182.650 ;
        RECT 76.650 182.590 76.970 182.850 ;
        RECT 78.505 182.790 78.795 182.835 ;
        RECT 79.870 182.790 80.190 182.850 ;
        RECT 90.080 182.790 90.220 182.990 ;
        RECT 78.505 182.650 90.220 182.790 ;
        RECT 90.450 182.790 90.770 182.850 ;
        RECT 91.385 182.790 91.675 182.835 ;
        RECT 90.450 182.650 91.675 182.790 ;
        RECT 78.505 182.605 78.795 182.650 ;
        RECT 79.870 182.590 80.190 182.650 ;
        RECT 90.450 182.590 90.770 182.650 ;
        RECT 91.385 182.605 91.675 182.650 ;
        RECT 92.290 182.790 92.610 182.850 ;
        RECT 94.145 182.790 94.435 182.835 ;
        RECT 94.590 182.790 94.910 182.850 ;
        RECT 92.290 182.650 94.910 182.790 ;
        RECT 92.290 182.590 92.610 182.650 ;
        RECT 94.145 182.605 94.435 182.650 ;
        RECT 94.590 182.590 94.910 182.650 ;
        RECT 95.050 182.590 95.370 182.850 ;
        RECT 99.190 182.790 99.510 182.850 ;
        RECT 100.585 182.790 100.875 182.835 ;
        RECT 99.190 182.650 100.875 182.790 ;
        RECT 101.580 182.790 101.720 182.990 ;
        RECT 102.870 182.930 103.190 182.990 ;
        RECT 103.420 182.990 108.250 183.130 ;
        RECT 103.420 182.790 103.560 182.990 ;
        RECT 107.930 182.930 108.250 182.990 ;
        RECT 101.580 182.650 103.560 182.790 ;
        RECT 104.725 182.790 105.015 182.835 ;
        RECT 105.630 182.790 105.950 182.850 ;
        RECT 104.725 182.650 105.950 182.790 ;
        RECT 99.190 182.590 99.510 182.650 ;
        RECT 100.585 182.605 100.875 182.650 ;
        RECT 104.725 182.605 105.015 182.650 ;
        RECT 105.630 182.590 105.950 182.650 ;
        RECT 107.470 182.590 107.790 182.850 ;
        RECT 109.860 182.790 110.000 183.610 ;
        RECT 112.160 183.130 112.300 184.010 ;
        RECT 114.385 183.965 114.675 184.195 ;
        RECT 117.130 184.150 117.450 184.210 ;
        RECT 121.270 184.150 121.590 184.210 ;
        RECT 121.745 184.150 122.035 184.195 ;
        RECT 117.130 184.010 122.035 184.150 ;
        RECT 117.130 183.950 117.450 184.010 ;
        RECT 121.270 183.950 121.590 184.010 ;
        RECT 121.745 183.965 122.035 184.010 ;
        RECT 117.220 183.775 117.360 183.950 ;
        RECT 118.525 183.810 118.815 183.855 ;
        RECT 122.280 183.810 122.420 184.290 ;
        RECT 122.650 184.195 122.970 184.210 ;
        RECT 122.650 183.965 123.035 184.195 ;
        RECT 123.660 184.150 123.800 184.305 ;
        RECT 127.250 184.290 127.570 184.350 ;
        RECT 133.780 184.210 133.920 184.350 ;
        RECT 134.165 184.350 135.850 184.490 ;
        RECT 134.165 184.305 134.455 184.350 ;
        RECT 135.530 184.290 135.850 184.350 ;
        RECT 141.970 184.490 142.290 184.550 ;
        RECT 142.445 184.490 142.735 184.535 ;
        RECT 141.970 184.350 142.735 184.490 ;
        RECT 141.970 184.290 142.290 184.350 ;
        RECT 142.445 184.305 142.735 184.350 ;
        RECT 144.270 184.290 144.590 184.550 ;
        RECT 127.710 184.150 128.030 184.210 ;
        RECT 123.660 184.010 129.780 184.150 ;
        RECT 122.650 183.950 122.970 183.965 ;
        RECT 127.710 183.950 128.030 184.010 ;
        RECT 117.145 183.545 117.435 183.775 ;
        RECT 118.525 183.670 122.420 183.810 ;
        RECT 118.525 183.625 118.815 183.670 ;
        RECT 124.950 183.610 125.270 183.870 ;
        RECT 125.870 183.810 126.190 183.870 ;
        RECT 127.265 183.810 127.555 183.855 ;
        RECT 129.090 183.810 129.410 183.870 ;
        RECT 129.640 183.855 129.780 184.010 ;
        RECT 133.690 183.950 134.010 184.210 ;
        RECT 140.590 184.150 140.910 184.210 ;
        RECT 140.590 184.010 141.740 184.150 ;
        RECT 140.590 183.950 140.910 184.010 ;
        RECT 125.870 183.670 129.410 183.810 ;
        RECT 125.870 183.610 126.190 183.670 ;
        RECT 127.265 183.625 127.555 183.670 ;
        RECT 129.090 183.610 129.410 183.670 ;
        RECT 129.565 183.625 129.855 183.855 ;
        RECT 130.010 183.810 130.330 183.870 ;
        RECT 131.405 183.810 131.695 183.855 ;
        RECT 130.010 183.670 131.695 183.810 ;
        RECT 130.010 183.610 130.330 183.670 ;
        RECT 131.405 183.625 131.695 183.670 ;
        RECT 132.310 183.610 132.630 183.870 ;
        RECT 132.785 183.810 133.075 183.855 ;
        RECT 133.230 183.810 133.550 183.870 ;
        RECT 135.085 183.810 135.375 183.855 ;
        RECT 132.785 183.670 135.375 183.810 ;
        RECT 132.785 183.625 133.075 183.670 ;
        RECT 133.230 183.610 133.550 183.670 ;
        RECT 135.085 183.625 135.375 183.670 ;
        RECT 138.290 183.810 138.610 183.870 ;
        RECT 141.600 183.855 141.740 184.010 ;
        RECT 140.080 183.810 140.370 183.855 ;
        RECT 138.290 183.670 140.650 183.810 ;
        RECT 138.290 183.610 138.610 183.670 ;
        RECT 140.080 183.625 140.370 183.670 ;
        RECT 119.430 183.470 119.750 183.530 ;
        RECT 119.905 183.470 120.195 183.515 ;
        RECT 118.140 183.330 120.195 183.470 ;
        RECT 118.140 183.175 118.280 183.330 ;
        RECT 119.430 183.270 119.750 183.330 ;
        RECT 119.905 183.285 120.195 183.330 ;
        RECT 118.065 183.130 118.355 183.175 ;
        RECT 124.030 183.130 124.350 183.190 ;
        RECT 125.960 183.175 126.100 183.610 ;
        RECT 131.850 183.470 132.170 183.530 ;
        RECT 134.150 183.470 134.470 183.530 ;
        RECT 129.870 183.330 132.170 183.470 ;
        RECT 112.160 182.990 118.355 183.130 ;
        RECT 118.065 182.945 118.355 182.990 ;
        RECT 120.440 182.990 124.350 183.130 ;
        RECT 112.070 182.790 112.390 182.850 ;
        RECT 109.860 182.650 112.390 182.790 ;
        RECT 112.070 182.590 112.390 182.650 ;
        RECT 112.990 182.790 113.310 182.850 ;
        RECT 114.845 182.790 115.135 182.835 ;
        RECT 112.990 182.650 115.135 182.790 ;
        RECT 112.990 182.590 113.310 182.650 ;
        RECT 114.845 182.605 115.135 182.650 ;
        RECT 116.670 182.790 116.990 182.850 ;
        RECT 120.440 182.835 120.580 182.990 ;
        RECT 124.030 182.930 124.350 182.990 ;
        RECT 125.885 182.945 126.175 183.175 ;
        RECT 127.250 183.130 127.570 183.190 ;
        RECT 128.185 183.130 128.475 183.175 ;
        RECT 127.250 182.990 128.475 183.130 ;
        RECT 127.250 182.930 127.570 182.990 ;
        RECT 128.185 182.945 128.475 182.990 ;
        RECT 128.630 182.930 128.950 183.190 ;
        RECT 129.870 183.130 130.010 183.330 ;
        RECT 131.850 183.270 132.170 183.330 ;
        RECT 133.320 183.330 134.470 183.470 ;
        RECT 133.320 183.175 133.460 183.330 ;
        RECT 134.150 183.270 134.470 183.330 ;
        RECT 137.830 183.470 138.150 183.530 ;
        RECT 140.510 183.470 140.650 183.670 ;
        RECT 141.525 183.625 141.815 183.855 ;
        RECT 143.825 183.810 144.115 183.855 ;
        RECT 144.360 183.810 144.500 184.290 ;
        RECT 143.825 183.670 144.500 183.810 ;
        RECT 143.825 183.625 144.115 183.670 ;
        RECT 137.830 183.330 140.360 183.470 ;
        RECT 140.510 183.330 143.120 183.470 ;
        RECT 137.830 183.270 138.150 183.330 ;
        RECT 133.245 183.130 133.535 183.175 ;
        RECT 129.180 182.990 130.010 183.130 ;
        RECT 131.940 182.990 133.535 183.130 ;
        RECT 140.220 183.130 140.360 183.330 ;
        RECT 142.980 183.175 143.120 183.330 ;
        RECT 140.605 183.130 140.895 183.175 ;
        RECT 140.220 182.990 140.895 183.130 ;
        RECT 120.365 182.790 120.655 182.835 ;
        RECT 116.670 182.650 120.655 182.790 ;
        RECT 116.670 182.590 116.990 182.650 ;
        RECT 120.365 182.605 120.655 182.650 ;
        RECT 121.285 182.790 121.575 182.835 ;
        RECT 121.730 182.790 122.050 182.850 ;
        RECT 121.285 182.650 122.050 182.790 ;
        RECT 121.285 182.605 121.575 182.650 ;
        RECT 121.730 182.590 122.050 182.650 ;
        RECT 122.190 182.790 122.510 182.850 ;
        RECT 122.665 182.790 122.955 182.835 ;
        RECT 129.180 182.790 129.320 182.990 ;
        RECT 122.190 182.650 129.320 182.790 ;
        RECT 130.010 182.790 130.330 182.850 ;
        RECT 131.940 182.790 132.080 182.990 ;
        RECT 133.245 182.945 133.535 182.990 ;
        RECT 140.605 182.945 140.895 182.990 ;
        RECT 141.065 182.945 141.355 183.175 ;
        RECT 142.905 182.945 143.195 183.175 ;
        RECT 130.010 182.650 132.080 182.790 ;
        RECT 132.325 182.790 132.615 182.835 ;
        RECT 132.770 182.790 133.090 182.850 ;
        RECT 132.325 182.650 133.090 182.790 ;
        RECT 122.190 182.590 122.510 182.650 ;
        RECT 122.665 182.605 122.955 182.650 ;
        RECT 130.010 182.590 130.330 182.650 ;
        RECT 132.325 182.605 132.615 182.650 ;
        RECT 132.770 182.590 133.090 182.650 ;
        RECT 134.610 182.790 134.930 182.850 ;
        RECT 138.290 182.790 138.610 182.850 ;
        RECT 141.140 182.790 141.280 182.945 ;
        RECT 134.610 182.650 141.280 182.790 ;
        RECT 134.610 182.590 134.930 182.650 ;
        RECT 138.290 182.590 138.610 182.650 ;
        RECT 36.100 181.970 150.180 182.450 ;
        RECT 44.910 181.770 45.230 181.830 ;
        RECT 46.290 181.770 46.610 181.830 ;
        RECT 46.765 181.770 47.055 181.815 ;
        RECT 44.910 181.630 46.015 181.770 ;
        RECT 44.910 181.570 45.230 181.630 ;
        RECT 45.385 181.245 45.675 181.475 ;
        RECT 45.875 181.430 46.015 181.630 ;
        RECT 46.290 181.630 47.055 181.770 ;
        RECT 46.290 181.570 46.610 181.630 ;
        RECT 46.765 181.585 47.055 181.630 ;
        RECT 48.590 181.770 48.910 181.830 ;
        RECT 49.525 181.770 49.815 181.815 ;
        RECT 48.590 181.630 49.815 181.770 ;
        RECT 48.590 181.570 48.910 181.630 ;
        RECT 49.525 181.585 49.815 181.630 ;
        RECT 50.430 181.770 50.750 181.830 ;
        RECT 51.810 181.770 52.130 181.830 ;
        RECT 50.430 181.630 52.130 181.770 ;
        RECT 50.430 181.570 50.750 181.630 ;
        RECT 51.810 181.570 52.130 181.630 ;
        RECT 63.785 181.770 64.075 181.815 ;
        RECT 65.165 181.770 65.455 181.815 ;
        RECT 63.785 181.630 65.455 181.770 ;
        RECT 63.785 181.585 64.075 181.630 ;
        RECT 65.165 181.585 65.455 181.630 ;
        RECT 66.085 181.770 66.375 181.815 ;
        RECT 68.385 181.770 68.675 181.815 ;
        RECT 66.085 181.630 68.675 181.770 ;
        RECT 66.085 181.585 66.375 181.630 ;
        RECT 68.385 181.585 68.675 181.630 ;
        RECT 75.285 181.770 75.575 181.815 ;
        RECT 76.205 181.770 76.495 181.815 ;
        RECT 75.285 181.630 76.495 181.770 ;
        RECT 75.285 181.585 75.575 181.630 ;
        RECT 76.205 181.585 76.495 181.630 ;
        RECT 87.690 181.770 88.010 181.830 ;
        RECT 90.465 181.770 90.755 181.815 ;
        RECT 92.290 181.770 92.610 181.830 ;
        RECT 87.690 181.630 92.610 181.770 ;
        RECT 87.690 181.570 88.010 181.630 ;
        RECT 90.465 181.585 90.755 181.630 ;
        RECT 92.290 181.570 92.610 181.630 ;
        RECT 94.590 181.770 94.910 181.830 ;
        RECT 97.810 181.770 98.130 181.830 ;
        RECT 94.590 181.630 98.130 181.770 ;
        RECT 94.590 181.570 94.910 181.630 ;
        RECT 97.810 181.570 98.130 181.630 ;
        RECT 99.665 181.770 99.955 181.815 ;
        RECT 108.390 181.770 108.710 181.830 ;
        RECT 112.530 181.770 112.850 181.830 ;
        RECT 114.845 181.770 115.135 181.815 ;
        RECT 99.665 181.630 110.000 181.770 ;
        RECT 99.665 181.585 99.955 181.630 ;
        RECT 108.390 181.570 108.710 181.630 ;
        RECT 47.685 181.430 47.975 181.475 ;
        RECT 63.325 181.430 63.615 181.475 ;
        RECT 67.465 181.430 67.755 181.475 ;
        RECT 45.875 181.290 47.975 181.430 ;
        RECT 47.685 181.245 47.975 181.290 ;
        RECT 49.140 181.290 61.240 181.430 ;
        RECT 44.465 180.565 44.755 180.795 ;
        RECT 45.460 180.750 45.600 181.245 ;
        RECT 45.845 180.750 46.135 180.795 ;
        RECT 48.605 180.750 48.895 180.795 ;
        RECT 49.140 180.750 49.280 181.290 ;
        RECT 61.100 181.150 61.240 181.290 ;
        RECT 63.325 181.290 67.755 181.430 ;
        RECT 63.325 181.245 63.615 181.290 ;
        RECT 67.465 181.245 67.755 181.290 ;
        RECT 69.305 181.430 69.595 181.475 ;
        RECT 83.090 181.430 83.410 181.490 ;
        RECT 69.305 181.290 83.410 181.430 ;
        RECT 69.305 181.245 69.595 181.290 ;
        RECT 83.090 181.230 83.410 181.290 ;
        RECT 88.610 181.230 88.930 181.490 ;
        RECT 90.910 181.430 91.230 181.490 ;
        RECT 106.550 181.430 106.870 181.490 ;
        RECT 90.910 181.290 106.870 181.430 ;
        RECT 90.910 181.230 91.230 181.290 ;
        RECT 49.510 181.090 49.830 181.150 ;
        RECT 55.030 181.090 55.350 181.150 ;
        RECT 49.510 180.950 55.350 181.090 ;
        RECT 49.510 180.890 49.830 180.950 ;
        RECT 45.460 180.610 49.280 180.750 ;
        RECT 49.970 180.750 50.290 180.810 ;
        RECT 50.980 180.795 51.120 180.950 ;
        RECT 55.030 180.890 55.350 180.950 ;
        RECT 61.010 180.890 61.330 181.150 ;
        RECT 61.470 181.090 61.790 181.150 ;
        RECT 61.945 181.090 62.235 181.135 ;
        RECT 62.865 181.090 63.155 181.135 ;
        RECT 67.925 181.090 68.215 181.135 ;
        RECT 61.470 180.950 68.215 181.090 ;
        RECT 61.470 180.890 61.790 180.950 ;
        RECT 61.945 180.905 62.235 180.950 ;
        RECT 62.865 180.905 63.155 180.950 ;
        RECT 67.925 180.905 68.215 180.950 ;
        RECT 76.650 180.890 76.970 181.150 ;
        RECT 81.710 181.090 82.030 181.150 ;
        RECT 81.570 180.890 82.030 181.090 ;
        RECT 50.445 180.750 50.735 180.795 ;
        RECT 49.970 180.610 50.735 180.750 ;
        RECT 45.845 180.565 46.135 180.610 ;
        RECT 48.605 180.565 48.895 180.610 ;
        RECT 44.540 180.130 44.680 180.565 ;
        RECT 49.970 180.550 50.290 180.610 ;
        RECT 50.445 180.565 50.735 180.610 ;
        RECT 50.905 180.565 51.195 180.795 ;
        RECT 56.885 180.750 57.175 180.795 ;
        RECT 58.710 180.750 59.030 180.810 ;
        RECT 54.660 180.610 59.030 180.750 ;
        RECT 46.750 180.410 47.070 180.470 ;
        RECT 47.225 180.410 47.515 180.455 ;
        RECT 46.750 180.270 47.515 180.410 ;
        RECT 46.750 180.210 47.070 180.270 ;
        RECT 47.225 180.225 47.515 180.270 ;
        RECT 48.145 180.410 48.435 180.455 ;
        RECT 49.525 180.410 49.815 180.455 ;
        RECT 54.110 180.410 54.430 180.470 ;
        RECT 48.145 180.270 49.280 180.410 ;
        RECT 48.145 180.225 48.435 180.270 ;
        RECT 44.450 179.870 44.770 180.130 ;
        RECT 49.140 180.070 49.280 180.270 ;
        RECT 49.525 180.270 54.430 180.410 ;
        RECT 49.525 180.225 49.815 180.270 ;
        RECT 54.110 180.210 54.430 180.270 ;
        RECT 49.970 180.070 50.290 180.130 ;
        RECT 49.140 179.930 50.290 180.070 ;
        RECT 49.970 179.870 50.290 179.930 ;
        RECT 51.825 180.070 52.115 180.115 ;
        RECT 52.270 180.070 52.590 180.130 ;
        RECT 51.825 179.930 52.590 180.070 ;
        RECT 51.825 179.885 52.115 179.930 ;
        RECT 52.270 179.870 52.590 179.930 ;
        RECT 53.650 180.070 53.970 180.130 ;
        RECT 54.660 180.070 54.800 180.610 ;
        RECT 56.885 180.565 57.175 180.610 ;
        RECT 58.710 180.550 59.030 180.610 ;
        RECT 59.170 180.750 59.490 180.810 ;
        RECT 64.245 180.750 64.535 180.795 ;
        RECT 59.170 180.610 64.535 180.750 ;
        RECT 59.170 180.550 59.490 180.610 ;
        RECT 64.245 180.565 64.535 180.610 ;
        RECT 64.690 180.750 65.010 180.810 ;
        RECT 66.990 180.750 67.310 180.810 ;
        RECT 78.980 180.795 79.240 180.840 ;
        RECT 64.690 180.610 67.310 180.750 ;
        RECT 64.690 180.550 65.010 180.610 ;
        RECT 66.990 180.550 67.310 180.610 ;
        RECT 76.205 180.750 76.495 180.795 ;
        RECT 78.965 180.750 79.255 180.795 ;
        RECT 81.570 180.750 81.710 180.890 ;
        RECT 76.205 180.610 81.710 180.750 ;
        RECT 83.180 180.750 83.320 181.230 ;
        RECT 88.700 181.090 88.840 181.230 ;
        RECT 93.210 181.090 93.530 181.150 ;
        RECT 88.700 180.950 93.530 181.090 ;
        RECT 89.620 180.795 89.760 180.950 ;
        RECT 93.210 180.890 93.530 180.950 ;
        RECT 89.085 180.750 89.375 180.795 ;
        RECT 83.180 180.610 89.375 180.750 ;
        RECT 76.205 180.565 76.495 180.610 ;
        RECT 78.965 180.565 79.255 180.610 ;
        RECT 89.085 180.565 89.375 180.610 ;
        RECT 89.545 180.565 89.835 180.795 ;
        RECT 89.990 180.750 90.310 180.810 ;
        RECT 90.910 180.750 91.230 180.810 ;
        RECT 89.990 180.610 91.230 180.750 ;
        RECT 78.980 180.520 79.240 180.565 ;
        RECT 62.850 180.210 63.170 180.470 ;
        RECT 65.610 180.410 65.930 180.470 ;
        RECT 66.545 180.410 66.835 180.455 ;
        RECT 65.610 180.270 66.835 180.410 ;
        RECT 65.610 180.210 65.930 180.270 ;
        RECT 66.545 180.225 66.835 180.270 ;
        RECT 79.425 180.410 79.715 180.455 ;
        RECT 79.870 180.410 80.190 180.470 ;
        RECT 79.425 180.270 80.190 180.410 ;
        RECT 79.425 180.225 79.715 180.270 ;
        RECT 79.870 180.210 80.190 180.270 ;
        RECT 88.165 180.410 88.455 180.455 ;
        RECT 88.610 180.410 88.930 180.470 ;
        RECT 88.165 180.270 88.930 180.410 ;
        RECT 89.160 180.410 89.300 180.565 ;
        RECT 89.990 180.550 90.310 180.610 ;
        RECT 90.910 180.550 91.230 180.610 ;
        RECT 91.385 180.565 91.675 180.795 ;
        RECT 91.845 180.565 92.135 180.795 ;
        RECT 91.460 180.410 91.600 180.565 ;
        RECT 89.160 180.270 91.600 180.410 ;
        RECT 91.920 180.410 92.060 180.565 ;
        RECT 92.750 180.550 93.070 180.810 ;
        RECT 95.140 180.795 95.280 181.290 ;
        RECT 106.550 181.230 106.870 181.290 ;
        RECT 107.470 181.230 107.790 181.490 ;
        RECT 107.930 181.430 108.250 181.490 ;
        RECT 109.860 181.430 110.000 181.630 ;
        RECT 112.530 181.630 115.135 181.770 ;
        RECT 112.530 181.570 112.850 181.630 ;
        RECT 114.845 181.585 115.135 181.630 ;
        RECT 117.130 181.770 117.450 181.830 ;
        RECT 117.605 181.770 117.895 181.815 ;
        RECT 117.130 181.630 117.895 181.770 ;
        RECT 117.130 181.570 117.450 181.630 ;
        RECT 117.605 181.585 117.895 181.630 ;
        RECT 119.430 181.570 119.750 181.830 ;
        RECT 119.890 181.570 120.210 181.830 ;
        RECT 121.270 181.570 121.590 181.830 ;
        RECT 125.410 181.770 125.730 181.830 ;
        RECT 127.710 181.770 128.030 181.830 ;
        RECT 128.630 181.770 128.950 181.830 ;
        RECT 125.410 181.630 128.950 181.770 ;
        RECT 125.410 181.570 125.730 181.630 ;
        RECT 127.710 181.570 128.030 181.630 ;
        RECT 128.630 181.570 128.950 181.630 ;
        RECT 129.550 181.570 129.870 181.830 ;
        RECT 132.310 181.770 132.630 181.830 ;
        RECT 132.785 181.770 133.075 181.815 ;
        RECT 132.310 181.630 133.075 181.770 ;
        RECT 132.310 181.570 132.630 181.630 ;
        RECT 132.785 181.585 133.075 181.630 ;
        RECT 133.690 181.770 134.010 181.830 ;
        RECT 135.085 181.770 135.375 181.815 ;
        RECT 136.465 181.770 136.755 181.815 ;
        RECT 133.690 181.630 136.755 181.770 ;
        RECT 133.690 181.570 134.010 181.630 ;
        RECT 135.085 181.585 135.375 181.630 ;
        RECT 136.465 181.585 136.755 181.630 ;
        RECT 136.910 181.570 137.230 181.830 ;
        RECT 140.130 181.570 140.450 181.830 ;
        RECT 141.525 181.770 141.815 181.815 ;
        RECT 143.350 181.770 143.670 181.830 ;
        RECT 141.525 181.630 143.670 181.770 ;
        RECT 141.525 181.585 141.815 181.630 ;
        RECT 143.350 181.570 143.670 181.630 ;
        RECT 113.005 181.430 113.295 181.475 ;
        RECT 119.520 181.430 119.660 181.570 ;
        RECT 121.360 181.430 121.500 181.570 ;
        RECT 107.930 181.290 109.540 181.430 ;
        RECT 109.860 181.290 113.295 181.430 ;
        RECT 107.930 181.230 108.250 181.290 ;
        RECT 95.970 180.890 96.290 181.150 ;
        RECT 99.190 181.090 99.510 181.150 ;
        RECT 98.820 180.950 99.510 181.090 ;
        RECT 95.065 180.565 95.355 180.795 ;
        RECT 96.060 180.750 96.200 180.890 ;
        RECT 98.820 180.795 98.960 180.950 ;
        RECT 99.190 180.890 99.510 180.950 ;
        RECT 100.110 181.090 100.430 181.150 ;
        RECT 103.790 181.090 104.110 181.150 ;
        RECT 105.630 181.090 105.950 181.150 ;
        RECT 100.110 180.950 105.950 181.090 ;
        RECT 107.560 181.090 107.700 181.230 ;
        RECT 109.400 181.135 109.540 181.290 ;
        RECT 113.005 181.245 113.295 181.290 ;
        RECT 115.840 181.290 119.660 181.430 ;
        RECT 120.900 181.290 121.500 181.430 ;
        RECT 108.865 181.090 109.155 181.135 ;
        RECT 107.560 180.950 109.155 181.090 ;
        RECT 100.110 180.890 100.430 180.950 ;
        RECT 103.790 180.890 104.110 180.950 ;
        RECT 105.630 180.890 105.950 180.950 ;
        RECT 108.865 180.905 109.155 180.950 ;
        RECT 109.325 180.905 109.615 181.135 ;
        RECT 110.230 181.090 110.550 181.150 ;
        RECT 110.230 180.950 114.600 181.090 ;
        RECT 110.230 180.890 110.550 180.950 ;
        RECT 96.060 180.610 98.500 180.750 ;
        RECT 96.060 180.410 96.200 180.610 ;
        RECT 91.920 180.270 96.200 180.410 ;
        RECT 88.165 180.225 88.455 180.270 ;
        RECT 88.610 180.210 88.930 180.270 ;
        RECT 97.810 180.210 98.130 180.470 ;
        RECT 98.360 180.410 98.500 180.610 ;
        RECT 98.745 180.565 99.035 180.795 ;
        RECT 107.485 180.750 107.775 180.795 ;
        RECT 109.785 180.750 110.075 180.795 ;
        RECT 101.580 180.610 110.075 180.750 ;
        RECT 101.580 180.410 101.720 180.610 ;
        RECT 107.485 180.565 107.775 180.610 ;
        RECT 109.785 180.565 110.075 180.610 ;
        RECT 110.690 180.550 111.010 180.810 ;
        RECT 112.085 180.750 112.375 180.795 ;
        RECT 113.450 180.750 113.770 180.810 ;
        RECT 114.460 180.795 114.600 180.950 ;
        RECT 115.840 180.795 115.980 181.290 ;
        RECT 117.590 181.090 117.910 181.150 ;
        RECT 120.900 181.090 121.040 181.290 ;
        RECT 128.645 181.090 128.935 181.135 ;
        RECT 129.640 181.090 129.780 181.570 ;
        RECT 133.230 181.430 133.550 181.490 ;
        RECT 135.545 181.430 135.835 181.475 ;
        RECT 137.000 181.430 137.140 181.570 ;
        RECT 140.590 181.430 140.910 181.490 ;
        RECT 147.045 181.430 147.335 181.475 ;
        RECT 116.300 180.950 117.910 181.090 ;
        RECT 116.300 180.810 116.440 180.950 ;
        RECT 117.590 180.890 117.910 180.950 ;
        RECT 119.060 180.950 121.040 181.090 ;
        RECT 121.360 180.950 128.400 181.090 ;
        RECT 112.085 180.610 113.770 180.750 ;
        RECT 112.085 180.565 112.375 180.610 ;
        RECT 113.450 180.550 113.770 180.610 ;
        RECT 114.385 180.565 114.675 180.795 ;
        RECT 115.765 180.565 116.055 180.795 ;
        RECT 98.360 180.270 101.720 180.410 ;
        RECT 101.950 180.410 102.270 180.470 ;
        RECT 103.330 180.410 103.650 180.470 ;
        RECT 101.950 180.270 103.650 180.410 ;
        RECT 101.950 180.210 102.270 180.270 ;
        RECT 103.330 180.210 103.650 180.270 ;
        RECT 105.630 180.410 105.950 180.470 ;
        RECT 111.625 180.410 111.915 180.455 ;
        RECT 105.630 180.270 111.915 180.410 ;
        RECT 105.630 180.210 105.950 180.270 ;
        RECT 111.625 180.225 111.915 180.270 ;
        RECT 53.650 179.930 54.800 180.070 ;
        RECT 55.030 180.070 55.350 180.130 ;
        RECT 57.805 180.070 58.095 180.115 ;
        RECT 55.030 179.930 58.095 180.070 ;
        RECT 53.650 179.870 53.970 179.930 ;
        RECT 55.030 179.870 55.350 179.930 ;
        RECT 57.805 179.885 58.095 179.930 ;
        RECT 63.310 180.070 63.630 180.130 ;
        RECT 68.370 180.070 68.690 180.130 ;
        RECT 63.310 179.930 68.690 180.070 ;
        RECT 63.310 179.870 63.630 179.930 ;
        RECT 68.370 179.870 68.690 179.930 ;
        RECT 91.830 180.070 92.150 180.130 ;
        RECT 93.685 180.070 93.975 180.115 ;
        RECT 91.830 179.930 93.975 180.070 ;
        RECT 91.830 179.870 92.150 179.930 ;
        RECT 93.685 179.885 93.975 179.930 ;
        RECT 94.145 180.070 94.435 180.115 ;
        RECT 95.970 180.070 96.290 180.130 ;
        RECT 94.145 179.930 96.290 180.070 ;
        RECT 94.145 179.885 94.435 179.930 ;
        RECT 95.970 179.870 96.290 179.930 ;
        RECT 97.350 180.070 97.670 180.130 ;
        RECT 98.730 180.070 99.050 180.130 ;
        RECT 97.350 179.930 99.050 180.070 ;
        RECT 97.350 179.870 97.670 179.930 ;
        RECT 98.730 179.870 99.050 179.930 ;
        RECT 99.190 180.070 99.510 180.130 ;
        RECT 104.250 180.070 104.570 180.130 ;
        RECT 99.190 179.930 104.570 180.070 ;
        RECT 99.190 179.870 99.510 179.930 ;
        RECT 104.250 179.870 104.570 179.930 ;
        RECT 109.770 180.070 110.090 180.130 ;
        RECT 113.465 180.070 113.755 180.115 ;
        RECT 109.770 179.930 113.755 180.070 ;
        RECT 115.840 180.070 115.980 180.565 ;
        RECT 116.210 180.550 116.530 180.810 ;
        RECT 116.670 180.750 116.990 180.810 ;
        RECT 119.060 180.795 119.200 180.950 ;
        RECT 118.525 180.750 118.815 180.795 ;
        RECT 116.670 180.610 117.820 180.750 ;
        RECT 116.670 180.550 116.990 180.610 ;
        RECT 117.680 180.455 117.820 180.610 ;
        RECT 118.140 180.610 118.815 180.750 ;
        RECT 117.605 180.225 117.895 180.455 ;
        RECT 117.145 180.070 117.435 180.115 ;
        RECT 115.840 179.930 117.435 180.070 ;
        RECT 118.140 180.070 118.280 180.610 ;
        RECT 118.525 180.565 118.815 180.610 ;
        RECT 118.985 180.565 119.275 180.795 ;
        RECT 119.890 180.750 120.210 180.810 ;
        RECT 120.365 180.750 120.655 180.795 ;
        RECT 121.360 180.750 121.500 180.950 ;
        RECT 119.890 180.610 121.500 180.750 ;
        RECT 119.890 180.550 120.210 180.610 ;
        RECT 120.365 180.565 120.655 180.610 ;
        RECT 121.730 180.550 122.050 180.810 ;
        RECT 122.650 180.750 122.970 180.810 ;
        RECT 127.725 180.750 128.015 180.795 ;
        RECT 122.650 180.610 128.015 180.750 ;
        RECT 128.260 180.750 128.400 180.950 ;
        RECT 128.645 180.950 129.780 181.090 ;
        RECT 130.560 181.290 133.550 181.430 ;
        RECT 128.645 180.905 128.935 180.950 ;
        RECT 130.010 180.750 130.330 180.810 ;
        RECT 130.560 180.795 130.700 181.290 ;
        RECT 133.230 181.230 133.550 181.290 ;
        RECT 133.780 181.290 135.835 181.430 ;
        RECT 133.780 181.090 133.920 181.290 ;
        RECT 135.545 181.245 135.835 181.290 ;
        RECT 136.080 181.290 137.600 181.430 ;
        RECT 131.480 180.950 133.920 181.090 ;
        RECT 134.625 181.090 134.915 181.135 ;
        RECT 136.080 181.090 136.220 181.290 ;
        RECT 137.460 181.135 137.600 181.290 ;
        RECT 140.590 181.290 147.335 181.430 ;
        RECT 140.590 181.230 140.910 181.290 ;
        RECT 147.045 181.245 147.335 181.290 ;
        RECT 134.625 180.950 136.220 181.090 ;
        RECT 131.480 180.795 131.620 180.950 ;
        RECT 134.625 180.905 134.915 180.950 ;
        RECT 137.385 180.905 137.675 181.135 ;
        RECT 139.670 180.890 139.990 181.150 ;
        RECT 141.510 181.090 141.830 181.150 ;
        RECT 143.365 181.090 143.655 181.135 ;
        RECT 147.950 181.090 148.270 181.150 ;
        RECT 141.510 180.950 143.655 181.090 ;
        RECT 141.510 180.890 141.830 180.950 ;
        RECT 143.365 180.905 143.655 180.950 ;
        RECT 146.660 180.950 148.270 181.090 ;
        RECT 128.260 180.610 130.330 180.750 ;
        RECT 122.650 180.550 122.970 180.610 ;
        RECT 127.725 180.565 128.015 180.610 ;
        RECT 130.010 180.550 130.330 180.610 ;
        RECT 130.485 180.565 130.775 180.795 ;
        RECT 131.405 180.565 131.695 180.795 ;
        RECT 133.705 180.750 133.995 180.795 ;
        RECT 135.990 180.750 136.310 180.810 ;
        RECT 136.465 180.750 136.755 180.795 ;
        RECT 133.705 180.610 136.755 180.750 ;
        RECT 133.705 180.565 133.995 180.610 ;
        RECT 135.990 180.550 136.310 180.610 ;
        RECT 136.465 180.565 136.755 180.610 ;
        RECT 137.845 180.750 138.135 180.795 ;
        RECT 140.130 180.750 140.450 180.810 ;
        RECT 146.660 180.795 146.800 180.950 ;
        RECT 147.950 180.890 148.270 180.950 ;
        RECT 140.605 180.750 140.895 180.795 ;
        RECT 141.985 180.750 142.275 180.795 ;
        RECT 137.845 180.610 139.900 180.750 ;
        RECT 137.845 180.565 138.135 180.610 ;
        RECT 121.820 180.410 121.960 180.550 ;
        RECT 139.760 180.470 139.900 180.610 ;
        RECT 140.130 180.610 142.275 180.750 ;
        RECT 140.130 180.550 140.450 180.610 ;
        RECT 140.605 180.565 140.895 180.610 ;
        RECT 141.985 180.565 142.275 180.610 ;
        RECT 146.585 180.565 146.875 180.795 ;
        RECT 147.505 180.565 147.795 180.795 ;
        RECT 133.230 180.410 133.550 180.470 ;
        RECT 121.820 180.270 133.550 180.410 ;
        RECT 133.230 180.210 133.550 180.270 ;
        RECT 134.610 180.410 134.930 180.470 ;
        RECT 135.085 180.410 135.375 180.455 ;
        RECT 134.610 180.270 135.375 180.410 ;
        RECT 134.610 180.210 134.930 180.270 ;
        RECT 135.085 180.225 135.375 180.270 ;
        RECT 139.210 180.210 139.530 180.470 ;
        RECT 139.670 180.210 139.990 180.470 ;
        RECT 142.060 180.410 142.200 180.565 ;
        RECT 147.580 180.410 147.720 180.565 ;
        RECT 142.060 180.270 147.720 180.410 ;
        RECT 121.270 180.070 121.590 180.130 ;
        RECT 118.140 179.930 121.590 180.070 ;
        RECT 109.770 179.870 110.090 179.930 ;
        RECT 113.465 179.885 113.755 179.930 ;
        RECT 117.145 179.885 117.435 179.930 ;
        RECT 121.270 179.870 121.590 179.930 ;
        RECT 126.790 179.870 127.110 180.130 ;
        RECT 130.945 180.070 131.235 180.115 ;
        RECT 132.310 180.070 132.630 180.130 ;
        RECT 130.945 179.930 132.630 180.070 ;
        RECT 130.945 179.885 131.235 179.930 ;
        RECT 132.310 179.870 132.630 179.930 ;
        RECT 36.100 179.250 150.180 179.730 ;
        RECT 44.450 179.050 44.770 179.110 ;
        RECT 44.450 178.910 49.740 179.050 ;
        RECT 44.450 178.850 44.770 178.910 ;
        RECT 38.930 178.415 39.250 178.430 ;
        RECT 38.900 178.185 39.250 178.415 ;
        RECT 38.930 178.170 39.250 178.185 ;
        RECT 46.750 178.370 47.070 178.430 ;
        RECT 49.600 178.415 49.740 178.910 ;
        RECT 50.430 178.850 50.750 179.110 ;
        RECT 50.890 179.050 51.210 179.110 ;
        RECT 52.745 179.050 53.035 179.095 ;
        RECT 53.650 179.050 53.970 179.110 ;
        RECT 50.890 178.910 53.970 179.050 ;
        RECT 50.890 178.850 51.210 178.910 ;
        RECT 52.745 178.865 53.035 178.910 ;
        RECT 53.650 178.850 53.970 178.910 ;
        RECT 58.250 178.850 58.570 179.110 ;
        RECT 58.710 178.850 59.030 179.110 ;
        RECT 59.170 179.050 59.490 179.110 ;
        RECT 63.310 179.050 63.630 179.110 ;
        RECT 59.170 178.910 63.630 179.050 ;
        RECT 59.170 178.850 59.490 178.910 ;
        RECT 63.310 178.850 63.630 178.910 ;
        RECT 63.770 179.050 64.090 179.110 ;
        RECT 68.845 179.050 69.135 179.095 ;
        RECT 63.770 178.910 69.135 179.050 ;
        RECT 63.770 178.850 64.090 178.910 ;
        RECT 68.845 178.865 69.135 178.910 ;
        RECT 89.085 179.050 89.375 179.095 ;
        RECT 92.750 179.050 93.070 179.110 ;
        RECT 89.085 178.910 93.070 179.050 ;
        RECT 89.085 178.865 89.375 178.910 ;
        RECT 92.750 178.850 93.070 178.910 ;
        RECT 95.510 179.050 95.830 179.110 ;
        RECT 101.950 179.050 102.270 179.110 ;
        RECT 95.510 178.910 102.270 179.050 ;
        RECT 95.510 178.850 95.830 178.910 ;
        RECT 101.950 178.850 102.270 178.910 ;
        RECT 102.410 179.050 102.730 179.110 ;
        RECT 102.410 178.910 105.400 179.050 ;
        RECT 102.410 178.850 102.730 178.910 ;
        RECT 49.970 178.710 50.290 178.770 ;
        RECT 58.340 178.710 58.480 178.850 ;
        RECT 49.970 178.570 58.480 178.710 ;
        RECT 49.970 178.510 50.290 178.570 ;
        RECT 47.225 178.370 47.515 178.415 ;
        RECT 49.525 178.370 49.815 178.415 ;
        RECT 50.890 178.370 51.210 178.430 ;
        RECT 58.340 178.415 58.480 178.570 ;
        RECT 46.750 178.230 49.280 178.370 ;
        RECT 46.750 178.170 47.070 178.230 ;
        RECT 47.225 178.185 47.515 178.230 ;
        RECT 37.550 177.830 37.870 178.090 ;
        RECT 38.445 178.030 38.735 178.075 ;
        RECT 39.635 178.030 39.925 178.075 ;
        RECT 42.155 178.030 42.445 178.075 ;
        RECT 38.445 177.890 42.445 178.030 ;
        RECT 38.445 177.845 38.735 177.890 ;
        RECT 39.635 177.845 39.925 177.890 ;
        RECT 42.155 177.845 42.445 177.890 ;
        RECT 48.590 177.830 48.910 178.090 ;
        RECT 49.140 178.030 49.280 178.230 ;
        RECT 49.525 178.230 51.210 178.370 ;
        RECT 49.525 178.185 49.815 178.230 ;
        RECT 50.890 178.170 51.210 178.230 ;
        RECT 51.825 178.370 52.115 178.415 ;
        RECT 51.825 178.230 53.420 178.370 ;
        RECT 51.825 178.185 52.115 178.230 ;
        RECT 49.140 177.890 52.040 178.030 ;
        RECT 38.050 177.690 38.340 177.735 ;
        RECT 40.150 177.690 40.440 177.735 ;
        RECT 41.720 177.690 42.010 177.735 ;
        RECT 38.050 177.550 42.010 177.690 ;
        RECT 38.050 177.505 38.340 177.550 ;
        RECT 40.150 177.505 40.440 177.550 ;
        RECT 41.720 177.505 42.010 177.550 ;
        RECT 49.050 177.690 49.370 177.750 ;
        RECT 51.365 177.690 51.655 177.735 ;
        RECT 49.050 177.550 51.655 177.690 ;
        RECT 49.050 177.490 49.370 177.550 ;
        RECT 49.600 177.395 49.740 177.550 ;
        RECT 51.365 177.505 51.655 177.550 ;
        RECT 49.525 177.165 49.815 177.395 ;
        RECT 51.900 177.350 52.040 177.890 ;
        RECT 53.280 177.750 53.420 178.230 ;
        RECT 53.665 178.185 53.955 178.415 ;
        RECT 58.265 178.185 58.555 178.415 ;
        RECT 58.800 178.370 58.940 178.850 ;
        RECT 64.230 178.540 64.550 178.770 ;
        RECT 64.230 178.510 64.920 178.540 ;
        RECT 66.530 178.510 66.850 178.770 ;
        RECT 90.910 178.710 91.230 178.770 ;
        RECT 95.970 178.710 96.290 178.770 ;
        RECT 90.910 178.570 91.600 178.710 ;
        RECT 90.910 178.510 91.230 178.570 ;
        RECT 64.320 178.415 64.920 178.510 ;
        RECT 59.645 178.370 59.935 178.415 ;
        RECT 64.320 178.400 64.960 178.415 ;
        RECT 58.800 178.230 59.935 178.370 ;
        RECT 59.645 178.185 59.935 178.230 ;
        RECT 64.670 178.185 64.960 178.400 ;
        RECT 65.105 178.380 65.395 178.415 ;
        RECT 65.105 178.370 65.840 178.380 ;
        RECT 66.620 178.370 66.760 178.510 ;
        RECT 65.105 178.240 66.760 178.370 ;
        RECT 65.105 178.185 65.395 178.240 ;
        RECT 65.700 178.230 66.760 178.240 ;
        RECT 67.005 178.370 67.295 178.415 ;
        RECT 67.450 178.370 67.770 178.430 ;
        RECT 67.005 178.230 67.770 178.370 ;
        RECT 67.005 178.185 67.295 178.230 ;
        RECT 53.190 177.490 53.510 177.750 ;
        RECT 53.740 177.350 53.880 178.185 ;
        RECT 67.450 178.170 67.770 178.230 ;
        RECT 79.870 178.170 80.190 178.430 ;
        RECT 81.265 178.370 81.555 178.415 ;
        RECT 84.470 178.370 84.790 178.430 ;
        RECT 81.265 178.230 84.790 178.370 ;
        RECT 81.265 178.185 81.555 178.230 ;
        RECT 84.470 178.170 84.790 178.230 ;
        RECT 89.070 178.170 89.390 178.430 ;
        RECT 89.530 178.370 89.850 178.430 ;
        RECT 91.460 178.415 91.600 178.570 ;
        RECT 91.920 178.570 96.290 178.710 ;
        RECT 91.920 178.415 92.060 178.570 ;
        RECT 95.970 178.510 96.290 178.570 ;
        RECT 96.980 178.570 102.640 178.710 ;
        RECT 96.980 178.430 97.120 178.570 ;
        RECT 90.005 178.370 90.295 178.415 ;
        RECT 89.530 178.230 90.295 178.370 ;
        RECT 89.530 178.170 89.850 178.230 ;
        RECT 90.005 178.185 90.295 178.230 ;
        RECT 91.385 178.185 91.675 178.415 ;
        RECT 91.845 178.185 92.135 178.415 ;
        RECT 92.765 178.370 93.055 178.415 ;
        RECT 95.050 178.370 95.370 178.430 ;
        RECT 96.890 178.370 97.210 178.430 ;
        RECT 92.765 178.230 97.210 178.370 ;
        RECT 92.765 178.185 93.055 178.230 ;
        RECT 95.050 178.170 95.370 178.230 ;
        RECT 96.890 178.170 97.210 178.230 ;
        RECT 99.650 178.370 99.970 178.430 ;
        RECT 102.500 178.415 102.640 178.570 ;
        RECT 101.965 178.370 102.255 178.415 ;
        RECT 99.650 178.230 102.255 178.370 ;
        RECT 99.650 178.170 99.970 178.230 ;
        RECT 101.965 178.185 102.255 178.230 ;
        RECT 102.425 178.185 102.715 178.415 ;
        RECT 103.330 178.170 103.650 178.430 ;
        RECT 103.790 178.170 104.110 178.430 ;
        RECT 104.250 178.170 104.570 178.430 ;
        RECT 105.260 178.415 105.400 178.910 ;
        RECT 107.470 178.850 107.790 179.110 ;
        RECT 107.930 179.050 108.250 179.110 ;
        RECT 111.165 179.050 111.455 179.095 ;
        RECT 107.930 178.910 111.455 179.050 ;
        RECT 107.930 178.850 108.250 178.910 ;
        RECT 111.165 178.865 111.455 178.910 ;
        RECT 118.510 178.850 118.830 179.110 ;
        RECT 119.445 179.050 119.735 179.095 ;
        RECT 135.085 179.050 135.375 179.095 ;
        RECT 137.385 179.050 137.675 179.095 ;
        RECT 119.445 178.910 126.100 179.050 ;
        RECT 119.445 178.865 119.735 178.910 ;
        RECT 107.560 178.710 107.700 178.850 ;
        RECT 118.600 178.710 118.740 178.850 ;
        RECT 105.720 178.570 107.240 178.710 ;
        RECT 107.560 178.570 110.460 178.710 ;
        RECT 105.185 178.185 105.475 178.415 ;
        RECT 61.470 178.030 61.790 178.090 ;
        RECT 62.405 178.030 62.695 178.075 ;
        RECT 63.325 178.030 63.615 178.075 ;
        RECT 68.385 178.030 68.675 178.075 ;
        RECT 61.470 177.890 68.675 178.030 ;
        RECT 61.470 177.830 61.790 177.890 ;
        RECT 62.405 177.845 62.695 177.890 ;
        RECT 63.325 177.845 63.615 177.890 ;
        RECT 68.385 177.845 68.675 177.890 ;
        RECT 77.570 177.830 77.890 178.090 ;
        RECT 89.160 178.030 89.300 178.170 ;
        RECT 90.925 178.030 91.215 178.075 ;
        RECT 99.190 178.030 99.510 178.090 ;
        RECT 89.160 177.890 99.510 178.030 ;
        RECT 103.880 178.030 104.020 178.170 ;
        RECT 105.720 178.030 105.860 178.570 ;
        RECT 106.550 178.170 106.870 178.430 ;
        RECT 107.100 178.370 107.240 178.570 ;
        RECT 107.485 178.370 107.775 178.415 ;
        RECT 107.100 178.230 107.775 178.370 ;
        RECT 107.485 178.185 107.775 178.230 ;
        RECT 109.770 178.170 110.090 178.430 ;
        RECT 110.320 178.415 110.460 178.570 ;
        RECT 118.140 178.570 118.740 178.710 ;
        RECT 119.905 178.710 120.195 178.755 ;
        RECT 120.810 178.710 121.130 178.770 ;
        RECT 119.905 178.570 121.130 178.710 ;
        RECT 125.960 178.710 126.100 178.910 ;
        RECT 135.085 178.910 137.675 179.050 ;
        RECT 135.085 178.865 135.375 178.910 ;
        RECT 137.385 178.865 137.675 178.910 ;
        RECT 136.925 178.710 137.215 178.755 ;
        RECT 125.960 178.570 137.215 178.710 ;
        RECT 118.140 178.415 118.280 178.570 ;
        RECT 119.905 178.525 120.195 178.570 ;
        RECT 120.810 178.510 121.130 178.570 ;
        RECT 136.925 178.525 137.215 178.570 ;
        RECT 110.245 178.185 110.535 178.415 ;
        RECT 117.605 178.370 117.895 178.415 ;
        RECT 116.760 178.230 117.895 178.370 ;
        RECT 103.880 177.890 105.860 178.030 ;
        RECT 106.105 178.030 106.395 178.075 ;
        RECT 110.690 178.030 111.010 178.090 ;
        RECT 106.105 177.890 111.010 178.030 ;
        RECT 90.925 177.845 91.215 177.890 ;
        RECT 99.190 177.830 99.510 177.890 ;
        RECT 106.105 177.845 106.395 177.890 ;
        RECT 110.690 177.830 111.010 177.890 ;
        RECT 63.785 177.690 64.075 177.735 ;
        RECT 67.925 177.690 68.215 177.735 ;
        RECT 89.070 177.690 89.390 177.750 ;
        RECT 91.370 177.690 91.690 177.750 ;
        RECT 108.865 177.690 109.155 177.735 ;
        RECT 63.785 177.550 68.215 177.690 ;
        RECT 63.785 177.505 64.075 177.550 ;
        RECT 67.925 177.505 68.215 177.550 ;
        RECT 69.380 177.550 88.840 177.690 ;
        RECT 69.380 177.410 69.520 177.550 ;
        RECT 51.900 177.210 53.880 177.350 ;
        RECT 54.110 177.350 54.430 177.410 ;
        RECT 60.090 177.350 60.410 177.410 ;
        RECT 54.110 177.210 60.410 177.350 ;
        RECT 54.110 177.150 54.430 177.210 ;
        RECT 60.090 177.150 60.410 177.210 ;
        RECT 60.565 177.350 60.855 177.395 ;
        RECT 63.310 177.350 63.630 177.410 ;
        RECT 60.565 177.210 63.630 177.350 ;
        RECT 60.565 177.165 60.855 177.210 ;
        RECT 63.310 177.150 63.630 177.210 ;
        RECT 64.245 177.350 64.535 177.395 ;
        RECT 65.625 177.350 65.915 177.395 ;
        RECT 64.245 177.210 65.915 177.350 ;
        RECT 64.245 177.165 64.535 177.210 ;
        RECT 65.625 177.165 65.915 177.210 ;
        RECT 66.545 177.350 66.835 177.395 ;
        RECT 68.845 177.350 69.135 177.395 ;
        RECT 66.545 177.210 69.135 177.350 ;
        RECT 66.545 177.165 66.835 177.210 ;
        RECT 68.845 177.165 69.135 177.210 ;
        RECT 69.290 177.150 69.610 177.410 ;
        RECT 69.750 177.150 70.070 177.410 ;
        RECT 79.405 177.350 79.695 177.395 ;
        RECT 80.325 177.350 80.615 177.395 ;
        RECT 79.405 177.210 80.615 177.350 ;
        RECT 88.700 177.350 88.840 177.550 ;
        RECT 89.070 177.550 93.900 177.690 ;
        RECT 89.070 177.490 89.390 177.550 ;
        RECT 91.370 177.490 91.690 177.550 ;
        RECT 93.210 177.350 93.530 177.410 ;
        RECT 88.700 177.210 93.530 177.350 ;
        RECT 93.760 177.350 93.900 177.550 ;
        RECT 104.340 177.550 109.155 177.690 ;
        RECT 116.760 177.690 116.900 178.230 ;
        RECT 117.605 178.185 117.895 178.230 ;
        RECT 118.065 178.185 118.355 178.415 ;
        RECT 118.525 178.370 118.815 178.415 ;
        RECT 126.790 178.370 127.110 178.430 ;
        RECT 131.865 178.370 132.155 178.415 ;
        RECT 118.525 178.230 132.155 178.370 ;
        RECT 118.525 178.185 118.815 178.230 ;
        RECT 126.790 178.170 127.110 178.230 ;
        RECT 131.865 178.185 132.155 178.230 ;
        RECT 132.310 178.370 132.630 178.430 ;
        RECT 134.165 178.370 134.455 178.415 ;
        RECT 135.990 178.370 136.310 178.430 ;
        RECT 132.310 178.230 133.920 178.370 ;
        RECT 132.310 178.170 132.630 178.230 ;
        RECT 117.130 178.030 117.450 178.090 ;
        RECT 122.190 178.030 122.510 178.090 ;
        RECT 117.130 177.890 122.510 178.030 ;
        RECT 117.130 177.830 117.450 177.890 ;
        RECT 122.190 177.830 122.510 177.890 ;
        RECT 133.230 177.830 133.550 178.090 ;
        RECT 133.780 178.030 133.920 178.230 ;
        RECT 134.165 178.230 136.310 178.370 ;
        RECT 134.165 178.185 134.455 178.230 ;
        RECT 135.990 178.170 136.310 178.230 ;
        RECT 137.370 178.370 137.690 178.430 ;
        RECT 141.425 178.370 141.715 178.415 ;
        RECT 137.370 178.230 141.715 178.370 ;
        RECT 137.370 178.170 137.690 178.230 ;
        RECT 141.425 178.185 141.715 178.230 ;
        RECT 134.610 178.030 134.930 178.090 ;
        RECT 135.545 178.030 135.835 178.075 ;
        RECT 133.780 177.890 135.835 178.030 ;
        RECT 134.610 177.830 134.930 177.890 ;
        RECT 135.545 177.845 135.835 177.890 ;
        RECT 136.910 178.030 137.230 178.090 ;
        RECT 137.970 178.030 138.260 178.075 ;
        RECT 136.910 177.890 138.260 178.030 ;
        RECT 136.910 177.830 137.230 177.890 ;
        RECT 137.970 177.845 138.260 177.890 ;
        RECT 140.145 177.845 140.435 178.075 ;
        RECT 141.025 178.030 141.315 178.075 ;
        RECT 142.215 178.030 142.505 178.075 ;
        RECT 144.735 178.030 145.025 178.075 ;
        RECT 141.025 177.890 145.025 178.030 ;
        RECT 141.025 177.845 141.315 177.890 ;
        RECT 142.215 177.845 142.505 177.890 ;
        RECT 144.735 177.845 145.025 177.890 ;
        RECT 140.220 177.690 140.360 177.845 ;
        RECT 116.760 177.550 117.360 177.690 ;
        RECT 104.340 177.350 104.480 177.550 ;
        RECT 108.865 177.505 109.155 177.550 ;
        RECT 117.220 177.410 117.360 177.550 ;
        RECT 127.340 177.550 140.360 177.690 ;
        RECT 140.630 177.690 140.920 177.735 ;
        RECT 142.730 177.690 143.020 177.735 ;
        RECT 144.300 177.690 144.590 177.735 ;
        RECT 140.630 177.550 144.590 177.690 ;
        RECT 127.340 177.410 127.480 177.550 ;
        RECT 140.630 177.505 140.920 177.550 ;
        RECT 142.730 177.505 143.020 177.550 ;
        RECT 144.300 177.505 144.590 177.550 ;
        RECT 93.760 177.210 104.480 177.350 ;
        RECT 108.405 177.350 108.695 177.395 ;
        RECT 110.690 177.350 111.010 177.410 ;
        RECT 108.405 177.210 111.010 177.350 ;
        RECT 79.405 177.165 79.695 177.210 ;
        RECT 80.325 177.165 80.615 177.210 ;
        RECT 93.210 177.150 93.530 177.210 ;
        RECT 108.405 177.165 108.695 177.210 ;
        RECT 110.690 177.150 111.010 177.210 ;
        RECT 117.130 177.150 117.450 177.410 ;
        RECT 118.970 177.350 119.290 177.410 ;
        RECT 123.110 177.350 123.430 177.410 ;
        RECT 118.970 177.210 123.430 177.350 ;
        RECT 118.970 177.150 119.290 177.210 ;
        RECT 123.110 177.150 123.430 177.210 ;
        RECT 127.250 177.150 127.570 177.410 ;
        RECT 130.485 177.350 130.775 177.395 ;
        RECT 133.230 177.350 133.550 177.410 ;
        RECT 130.485 177.210 133.550 177.350 ;
        RECT 130.485 177.165 130.775 177.210 ;
        RECT 133.230 177.150 133.550 177.210 ;
        RECT 138.750 177.150 139.070 177.410 ;
        RECT 140.130 177.350 140.450 177.410 ;
        RECT 147.045 177.350 147.335 177.395 ;
        RECT 140.130 177.210 147.335 177.350 ;
        RECT 140.130 177.150 140.450 177.210 ;
        RECT 147.045 177.165 147.335 177.210 ;
        RECT 36.100 176.530 150.180 177.010 ;
        RECT 38.930 176.330 39.250 176.390 ;
        RECT 40.325 176.330 40.615 176.375 ;
        RECT 38.930 176.190 40.615 176.330 ;
        RECT 38.930 176.130 39.250 176.190 ;
        RECT 40.325 176.145 40.615 176.190 ;
        RECT 47.670 176.330 47.990 176.390 ;
        RECT 49.525 176.330 49.815 176.375 ;
        RECT 47.670 176.190 49.815 176.330 ;
        RECT 47.670 176.130 47.990 176.190 ;
        RECT 49.525 176.145 49.815 176.190 ;
        RECT 49.970 176.130 50.290 176.390 ;
        RECT 51.825 176.145 52.115 176.375 ;
        RECT 55.045 176.330 55.335 176.375 ;
        RECT 57.345 176.330 57.635 176.375 ;
        RECT 55.045 176.190 57.635 176.330 ;
        RECT 55.045 176.145 55.335 176.190 ;
        RECT 57.345 176.145 57.635 176.190 ;
        RECT 58.265 176.330 58.555 176.375 ;
        RECT 59.645 176.330 59.935 176.375 ;
        RECT 58.265 176.190 59.935 176.330 ;
        RECT 58.265 176.145 58.555 176.190 ;
        RECT 59.645 176.145 59.935 176.190 ;
        RECT 60.550 176.330 60.870 176.390 ;
        RECT 69.290 176.330 69.610 176.390 ;
        RECT 60.550 176.190 69.610 176.330 ;
        RECT 46.290 175.650 46.610 175.710 ;
        RECT 48.130 175.650 48.450 175.710 ;
        RECT 48.605 175.650 48.895 175.695 ;
        RECT 46.290 175.510 48.895 175.650 ;
        RECT 50.060 175.650 50.200 176.130 ;
        RECT 51.900 175.990 52.040 176.145 ;
        RECT 60.550 176.130 60.870 176.190 ;
        RECT 69.290 176.130 69.610 176.190 ;
        RECT 69.750 176.330 70.070 176.390 ;
        RECT 97.350 176.330 97.670 176.390 ;
        RECT 101.030 176.330 101.350 176.390 ;
        RECT 69.750 176.190 97.120 176.330 ;
        RECT 69.750 176.130 70.070 176.190 ;
        RECT 53.205 175.990 53.495 176.035 ;
        RECT 53.650 175.990 53.970 176.050 ;
        RECT 51.900 175.850 53.970 175.990 ;
        RECT 53.205 175.805 53.495 175.850 ;
        RECT 53.650 175.790 53.970 175.850 ;
        RECT 54.110 175.790 54.430 176.050 ;
        RECT 55.965 175.990 56.255 176.035 ;
        RECT 60.105 175.990 60.395 176.035 ;
        RECT 55.965 175.850 60.395 175.990 ;
        RECT 55.965 175.805 56.255 175.850 ;
        RECT 60.105 175.805 60.395 175.850 ;
        RECT 87.690 175.990 88.010 176.050 ;
        RECT 92.750 175.990 93.070 176.050 ;
        RECT 87.690 175.850 93.070 175.990 ;
        RECT 96.980 175.990 97.120 176.190 ;
        RECT 97.350 176.190 101.350 176.330 ;
        RECT 97.350 176.130 97.670 176.190 ;
        RECT 101.030 176.130 101.350 176.190 ;
        RECT 101.950 176.330 102.270 176.390 ;
        RECT 110.705 176.330 110.995 176.375 ;
        RECT 111.610 176.330 111.930 176.390 ;
        RECT 101.950 176.190 110.460 176.330 ;
        RECT 101.950 176.130 102.270 176.190 ;
        RECT 107.010 175.990 107.330 176.050 ;
        RECT 96.980 175.850 107.330 175.990 ;
        RECT 87.690 175.790 88.010 175.850 ;
        RECT 92.750 175.790 93.070 175.850 ;
        RECT 61.500 175.695 61.760 175.740 ;
        RECT 55.505 175.650 55.795 175.695 ;
        RECT 60.565 175.650 60.855 175.695 ;
        RECT 61.485 175.650 61.775 175.695 ;
        RECT 72.510 175.650 72.830 175.710 ;
        RECT 95.510 175.650 95.830 175.710 ;
        RECT 50.060 175.510 52.500 175.650 ;
        RECT 46.290 175.450 46.610 175.510 ;
        RECT 48.130 175.450 48.450 175.510 ;
        RECT 48.605 175.465 48.895 175.510 ;
        RECT 52.360 175.370 52.500 175.510 ;
        RECT 55.505 175.510 61.775 175.650 ;
        RECT 55.505 175.465 55.795 175.510 ;
        RECT 60.565 175.465 60.855 175.510 ;
        RECT 61.485 175.465 61.775 175.510 ;
        RECT 70.760 175.510 95.830 175.650 ;
        RECT 61.500 175.420 61.760 175.465 ;
        RECT 40.310 175.110 40.630 175.370 ;
        RECT 41.245 175.310 41.535 175.355 ;
        RECT 42.610 175.310 42.930 175.370 ;
        RECT 45.370 175.310 45.690 175.370 ;
        RECT 41.245 175.170 45.690 175.310 ;
        RECT 41.245 175.125 41.535 175.170 ;
        RECT 42.610 175.110 42.930 175.170 ;
        RECT 45.370 175.110 45.690 175.170 ;
        RECT 47.225 175.310 47.515 175.355 ;
        RECT 47.225 175.170 49.740 175.310 ;
        RECT 47.225 175.125 47.515 175.170 ;
        RECT 49.600 175.030 49.740 175.170 ;
        RECT 50.445 175.125 50.735 175.355 ;
        RECT 49.510 174.770 49.830 175.030 ;
        RECT 50.520 174.970 50.660 175.125 ;
        RECT 50.890 175.110 51.210 175.370 ;
        RECT 51.810 175.110 52.130 175.370 ;
        RECT 52.270 175.110 52.590 175.370 ;
        RECT 53.650 175.310 53.970 175.370 ;
        RECT 52.820 175.170 53.970 175.310 ;
        RECT 52.820 174.970 52.960 175.170 ;
        RECT 53.650 175.110 53.970 175.170 ;
        RECT 54.570 175.310 54.890 175.370 ;
        RECT 56.885 175.310 57.175 175.355 ;
        RECT 58.250 175.310 58.570 175.370 ;
        RECT 54.570 175.170 58.570 175.310 ;
        RECT 54.570 175.110 54.890 175.170 ;
        RECT 56.885 175.125 57.175 175.170 ;
        RECT 58.250 175.110 58.570 175.170 ;
        RECT 59.170 175.110 59.490 175.370 ;
        RECT 70.760 175.355 70.900 175.510 ;
        RECT 72.510 175.450 72.830 175.510 ;
        RECT 95.510 175.450 95.830 175.510 ;
        RECT 95.970 175.650 96.290 175.710 ;
        RECT 99.190 175.650 99.510 175.710 ;
        RECT 95.970 175.510 99.510 175.650 ;
        RECT 95.970 175.450 96.290 175.510 ;
        RECT 99.190 175.450 99.510 175.510 ;
        RECT 99.650 175.650 99.970 175.710 ;
        RECT 100.125 175.650 100.415 175.695 ;
        RECT 99.650 175.510 100.415 175.650 ;
        RECT 99.650 175.450 99.970 175.510 ;
        RECT 100.125 175.465 100.415 175.510 ;
        RECT 70.685 175.125 70.975 175.355 ;
        RECT 83.090 175.110 83.410 175.370 ;
        RECT 84.025 175.125 84.315 175.355 ;
        RECT 84.945 175.310 85.235 175.355 ;
        RECT 86.770 175.310 87.090 175.370 ;
        RECT 84.945 175.170 87.090 175.310 ;
        RECT 84.945 175.125 85.235 175.170 ;
        RECT 50.520 174.830 52.960 174.970 ;
        RECT 58.725 174.970 59.015 175.015 ;
        RECT 59.630 174.970 59.950 175.030 ;
        RECT 58.725 174.830 59.950 174.970 ;
        RECT 58.725 174.785 59.015 174.830 ;
        RECT 59.630 174.770 59.950 174.830 ;
        RECT 61.010 174.970 61.330 175.030 ;
        RECT 84.100 174.970 84.240 175.125 ;
        RECT 86.770 175.110 87.090 175.170 ;
        RECT 87.245 175.125 87.535 175.355 ;
        RECT 87.705 175.310 87.995 175.355 ;
        RECT 88.150 175.310 88.470 175.370 ;
        RECT 87.705 175.170 88.470 175.310 ;
        RECT 87.705 175.125 87.995 175.170 ;
        RECT 84.470 174.970 84.790 175.030 ;
        RECT 61.010 174.830 83.780 174.970 ;
        RECT 84.100 174.830 84.790 174.970 ;
        RECT 61.010 174.770 61.330 174.830 ;
        RECT 54.570 174.630 54.890 174.690 ;
        RECT 55.045 174.630 55.335 174.675 ;
        RECT 54.570 174.490 55.335 174.630 ;
        RECT 54.570 174.430 54.890 174.490 ;
        RECT 55.045 174.445 55.335 174.490 ;
        RECT 60.550 174.430 60.870 174.690 ;
        RECT 64.245 174.630 64.535 174.675 ;
        RECT 65.610 174.630 65.930 174.690 ;
        RECT 64.245 174.490 65.930 174.630 ;
        RECT 83.640 174.630 83.780 174.830 ;
        RECT 84.470 174.770 84.790 174.830 ;
        RECT 85.405 174.785 85.695 175.015 ;
        RECT 86.325 174.785 86.615 175.015 ;
        RECT 87.320 174.970 87.460 175.125 ;
        RECT 88.150 175.110 88.470 175.170 ;
        RECT 88.610 175.110 88.930 175.370 ;
        RECT 89.070 175.110 89.390 175.370 ;
        RECT 89.530 175.110 89.850 175.370 ;
        RECT 91.830 175.110 92.150 175.370 ;
        RECT 92.290 175.110 92.610 175.370 ;
        RECT 92.750 175.110 93.070 175.370 ;
        RECT 93.225 175.125 93.515 175.355 ;
        RECT 97.350 175.310 97.670 175.370 ;
        RECT 98.270 175.310 98.590 175.370 ;
        RECT 97.350 175.170 98.590 175.310 ;
        RECT 93.300 174.970 93.440 175.125 ;
        RECT 97.350 175.110 97.670 175.170 ;
        RECT 98.270 175.110 98.590 175.170 ;
        RECT 98.745 175.125 99.035 175.355 ;
        RECT 95.970 174.970 96.290 175.030 ;
        RECT 98.820 174.970 98.960 175.125 ;
        RECT 101.030 175.110 101.350 175.370 ;
        RECT 102.040 175.355 102.180 175.850 ;
        RECT 107.010 175.790 107.330 175.850 ;
        RECT 107.470 175.990 107.790 176.050 ;
        RECT 108.850 175.990 109.170 176.050 ;
        RECT 110.320 175.990 110.460 176.190 ;
        RECT 110.705 176.190 111.930 176.330 ;
        RECT 110.705 176.145 110.995 176.190 ;
        RECT 111.610 176.130 111.930 176.190 ;
        RECT 121.285 176.330 121.575 176.375 ;
        RECT 126.790 176.330 127.110 176.390 ;
        RECT 121.285 176.190 127.110 176.330 ;
        RECT 121.285 176.145 121.575 176.190 ;
        RECT 107.470 175.850 110.000 175.990 ;
        RECT 110.320 175.850 115.980 175.990 ;
        RECT 107.470 175.790 107.790 175.850 ;
        RECT 108.850 175.790 109.170 175.850 ;
        RECT 102.410 175.450 102.730 175.710 ;
        RECT 102.870 175.450 103.190 175.710 ;
        RECT 105.630 175.450 105.950 175.710 ;
        RECT 107.100 175.650 107.240 175.790 ;
        RECT 107.100 175.510 109.540 175.650 ;
        RECT 101.965 175.125 102.255 175.355 ;
        RECT 103.805 175.125 104.095 175.355 ;
        RECT 104.250 175.310 104.570 175.370 ;
        RECT 109.400 175.355 109.540 175.510 ;
        RECT 109.860 175.355 110.000 175.850 ;
        RECT 110.690 175.450 111.010 175.710 ;
        RECT 112.530 175.650 112.850 175.710 ;
        RECT 115.840 175.695 115.980 175.850 ;
        RECT 120.350 175.790 120.670 176.050 ;
        RECT 114.385 175.650 114.675 175.695 ;
        RECT 112.530 175.510 114.675 175.650 ;
        RECT 112.530 175.450 112.850 175.510 ;
        RECT 114.385 175.465 114.675 175.510 ;
        RECT 115.765 175.650 116.055 175.695 ;
        RECT 117.130 175.650 117.450 175.710 ;
        RECT 121.360 175.650 121.500 176.145 ;
        RECT 126.790 176.130 127.110 176.190 ;
        RECT 127.250 176.130 127.570 176.390 ;
        RECT 130.010 176.330 130.330 176.390 ;
        RECT 135.070 176.330 135.390 176.390 ;
        RECT 130.010 176.190 135.390 176.330 ;
        RECT 130.010 176.130 130.330 176.190 ;
        RECT 135.070 176.130 135.390 176.190 ;
        RECT 137.370 176.130 137.690 176.390 ;
        RECT 138.750 176.130 139.070 176.390 ;
        RECT 127.340 175.990 127.480 176.130 ;
        RECT 128.670 175.990 128.960 176.035 ;
        RECT 130.770 175.990 131.060 176.035 ;
        RECT 132.340 175.990 132.630 176.035 ;
        RECT 127.340 175.850 128.400 175.990 ;
        RECT 128.260 175.695 128.400 175.850 ;
        RECT 128.670 175.850 132.630 175.990 ;
        RECT 128.670 175.805 128.960 175.850 ;
        RECT 130.770 175.805 131.060 175.850 ;
        RECT 132.340 175.805 132.630 175.850 ;
        RECT 135.990 175.990 136.310 176.050 ;
        RECT 138.305 175.990 138.595 176.035 ;
        RECT 135.990 175.850 138.595 175.990 ;
        RECT 135.990 175.790 136.310 175.850 ;
        RECT 138.305 175.805 138.595 175.850 ;
        RECT 122.205 175.650 122.495 175.695 ;
        RECT 115.765 175.510 117.450 175.650 ;
        RECT 115.765 175.465 116.055 175.510 ;
        RECT 117.130 175.450 117.450 175.510 ;
        RECT 119.060 175.510 121.500 175.650 ;
        RECT 121.820 175.510 122.495 175.650 ;
        RECT 106.105 175.310 106.395 175.355 ;
        RECT 104.250 175.170 106.395 175.310 ;
        RECT 100.570 174.970 100.890 175.030 ;
        RECT 87.320 174.830 93.440 174.970 ;
        RECT 93.760 174.830 94.820 174.970 ;
        RECT 85.480 174.630 85.620 174.785 ;
        RECT 83.640 174.490 85.620 174.630 ;
        RECT 86.400 174.630 86.540 174.785 ;
        RECT 89.990 174.630 90.310 174.690 ;
        RECT 86.400 174.490 90.310 174.630 ;
        RECT 64.245 174.445 64.535 174.490 ;
        RECT 65.610 174.430 65.930 174.490 ;
        RECT 89.990 174.430 90.310 174.490 ;
        RECT 90.910 174.430 91.230 174.690 ;
        RECT 91.370 174.630 91.690 174.690 ;
        RECT 93.760 174.630 93.900 174.830 ;
        RECT 91.370 174.490 93.900 174.630 ;
        RECT 91.370 174.430 91.690 174.490 ;
        RECT 94.130 174.430 94.450 174.690 ;
        RECT 94.680 174.630 94.820 174.830 ;
        RECT 95.970 174.830 100.890 174.970 ;
        RECT 95.970 174.770 96.290 174.830 ;
        RECT 100.570 174.770 100.890 174.830 ;
        RECT 101.490 174.970 101.810 175.030 ;
        RECT 103.880 174.970 104.020 175.125 ;
        RECT 104.250 175.110 104.570 175.170 ;
        RECT 106.105 175.125 106.395 175.170 ;
        RECT 106.565 175.125 106.855 175.355 ;
        RECT 107.025 175.310 107.315 175.355 ;
        RECT 107.025 175.170 109.080 175.310 ;
        RECT 107.025 175.125 107.315 175.170 ;
        RECT 101.490 174.830 104.020 174.970 ;
        RECT 105.630 174.970 105.950 175.030 ;
        RECT 106.640 174.970 106.780 175.125 ;
        RECT 108.405 174.970 108.695 175.015 ;
        RECT 105.630 174.830 106.780 174.970 ;
        RECT 107.100 174.830 108.695 174.970 ;
        RECT 108.940 174.970 109.080 175.170 ;
        RECT 109.325 175.125 109.615 175.355 ;
        RECT 109.785 175.125 110.075 175.355 ;
        RECT 110.780 174.970 110.920 175.450 ;
        RECT 111.165 175.310 111.455 175.355 ;
        RECT 117.590 175.310 117.910 175.370 ;
        RECT 119.060 175.355 119.200 175.510 ;
        RECT 121.820 175.370 121.960 175.510 ;
        RECT 122.205 175.465 122.495 175.510 ;
        RECT 123.200 175.510 127.480 175.650 ;
        RECT 111.165 175.170 117.910 175.310 ;
        RECT 111.165 175.125 111.455 175.170 ;
        RECT 117.590 175.110 117.910 175.170 ;
        RECT 118.985 175.125 119.275 175.355 ;
        RECT 120.825 175.310 121.115 175.355 ;
        RECT 119.520 175.170 121.115 175.310 ;
        RECT 108.940 174.830 110.920 174.970 ;
        RECT 101.490 174.770 101.810 174.830 ;
        RECT 105.630 174.770 105.950 174.830 ;
        RECT 101.950 174.630 102.270 174.690 ;
        RECT 94.680 174.490 102.270 174.630 ;
        RECT 101.950 174.430 102.270 174.490 ;
        RECT 102.410 174.630 102.730 174.690 ;
        RECT 104.725 174.630 105.015 174.675 ;
        RECT 102.410 174.490 105.015 174.630 ;
        RECT 102.410 174.430 102.730 174.490 ;
        RECT 104.725 174.445 105.015 174.490 ;
        RECT 106.550 174.630 106.870 174.690 ;
        RECT 107.100 174.630 107.240 174.830 ;
        RECT 108.405 174.785 108.695 174.830 ;
        RECT 119.520 174.690 119.660 175.170 ;
        RECT 120.825 175.125 121.115 175.170 ;
        RECT 121.730 175.110 122.050 175.370 ;
        RECT 123.200 175.355 123.340 175.510 ;
        RECT 123.125 175.125 123.415 175.355 ;
        RECT 124.030 175.110 124.350 175.370 ;
        RECT 124.950 175.110 125.270 175.370 ;
        RECT 126.790 175.110 127.110 175.370 ;
        RECT 127.340 175.355 127.480 175.510 ;
        RECT 128.185 175.465 128.475 175.695 ;
        RECT 129.065 175.650 129.355 175.695 ;
        RECT 130.255 175.650 130.545 175.695 ;
        RECT 132.775 175.650 133.065 175.695 ;
        RECT 138.840 175.650 138.980 176.130 ;
        RECT 129.065 175.510 133.065 175.650 ;
        RECT 129.065 175.465 129.355 175.510 ;
        RECT 130.255 175.465 130.545 175.510 ;
        RECT 132.775 175.465 133.065 175.510 ;
        RECT 136.540 175.510 138.980 175.650 ;
        RECT 127.265 175.125 127.555 175.355 ;
        RECT 127.710 175.110 128.030 175.370 ;
        RECT 128.260 175.310 128.400 175.465 ;
        RECT 132.310 175.310 132.630 175.370 ;
        RECT 136.540 175.355 136.680 175.510 ;
        RECT 128.260 175.170 132.630 175.310 ;
        RECT 132.310 175.110 132.630 175.170 ;
        RECT 136.465 175.125 136.755 175.355 ;
        RECT 138.765 175.310 139.055 175.355 ;
        RECT 140.130 175.310 140.450 175.370 ;
        RECT 138.765 175.170 140.450 175.310 ;
        RECT 138.765 175.125 139.055 175.170 ;
        RECT 140.130 175.110 140.450 175.170 ;
        RECT 120.365 174.970 120.655 175.015 ;
        RECT 122.205 174.970 122.495 175.015 ;
        RECT 124.505 174.970 124.795 175.015 ;
        RECT 129.410 174.970 129.700 175.015 ;
        RECT 120.365 174.830 122.495 174.970 ;
        RECT 120.365 174.785 120.655 174.830 ;
        RECT 122.205 174.785 122.495 174.830 ;
        RECT 123.200 174.830 124.795 174.970 ;
        RECT 123.200 174.690 123.340 174.830 ;
        RECT 124.505 174.785 124.795 174.830 ;
        RECT 125.960 174.830 129.700 174.970 ;
        RECT 106.550 174.490 107.240 174.630 ;
        RECT 107.945 174.630 108.235 174.675 ;
        RECT 118.510 174.630 118.830 174.690 ;
        RECT 107.945 174.490 118.830 174.630 ;
        RECT 106.550 174.430 106.870 174.490 ;
        RECT 107.945 174.445 108.235 174.490 ;
        RECT 118.510 174.430 118.830 174.490 ;
        RECT 119.430 174.430 119.750 174.690 ;
        RECT 123.110 174.430 123.430 174.690 ;
        RECT 125.960 174.675 126.100 174.830 ;
        RECT 129.410 174.785 129.700 174.830 ;
        RECT 125.885 174.445 126.175 174.675 ;
        RECT 36.100 173.810 150.180 174.290 ;
        RECT 40.310 173.610 40.630 173.670 ;
        RECT 42.165 173.610 42.455 173.655 ;
        RECT 40.310 173.470 42.455 173.610 ;
        RECT 40.310 173.410 40.630 173.470 ;
        RECT 42.165 173.425 42.455 173.470 ;
        RECT 43.990 173.410 44.310 173.670 ;
        RECT 45.370 173.410 45.690 173.670 ;
        RECT 49.985 173.610 50.275 173.655 ;
        RECT 50.890 173.610 51.210 173.670 ;
        RECT 45.920 173.470 49.740 173.610 ;
        RECT 44.080 173.270 44.220 173.410 ;
        RECT 45.920 173.270 46.060 173.470 ;
        RECT 46.290 173.315 46.610 173.330 ;
        RECT 44.080 173.130 46.060 173.270 ;
        RECT 46.225 173.085 46.610 173.315 ;
        RECT 47.225 173.270 47.515 173.315 ;
        RECT 48.130 173.270 48.450 173.330 ;
        RECT 49.600 173.270 49.740 173.470 ;
        RECT 49.985 173.470 51.210 173.610 ;
        RECT 49.985 173.425 50.275 173.470 ;
        RECT 50.890 173.410 51.210 173.470 ;
        RECT 51.365 173.425 51.655 173.655 ;
        RECT 51.440 173.270 51.580 173.425 ;
        RECT 52.270 173.410 52.590 173.670 ;
        RECT 53.650 173.610 53.970 173.670 ;
        RECT 59.630 173.610 59.950 173.670 ;
        RECT 53.650 173.470 59.950 173.610 ;
        RECT 53.650 173.410 53.970 173.470 ;
        RECT 59.630 173.410 59.950 173.470 ;
        RECT 63.770 173.610 64.090 173.670 ;
        RECT 65.150 173.610 65.470 173.670 ;
        RECT 70.225 173.610 70.515 173.655 ;
        RECT 83.090 173.610 83.410 173.670 ;
        RECT 84.470 173.610 84.790 173.670 ;
        RECT 63.770 173.470 64.460 173.610 ;
        RECT 63.770 173.410 64.090 173.470 ;
        RECT 60.550 173.270 60.870 173.330 ;
        RECT 47.225 173.130 49.280 173.270 ;
        RECT 49.600 173.130 60.870 173.270 ;
        RECT 64.320 173.270 64.460 173.470 ;
        RECT 65.150 173.470 78.720 173.610 ;
        RECT 65.150 173.410 65.470 173.470 ;
        RECT 70.225 173.425 70.515 173.470 ;
        RECT 78.580 173.330 78.720 173.470 ;
        RECT 83.090 173.470 84.790 173.610 ;
        RECT 83.090 173.410 83.410 173.470 ;
        RECT 84.470 173.410 84.790 173.470 ;
        RECT 89.070 173.410 89.390 173.670 ;
        RECT 89.990 173.610 90.310 173.670 ;
        RECT 91.830 173.610 92.150 173.670 ;
        RECT 93.670 173.610 93.990 173.670 ;
        RECT 89.990 173.470 93.990 173.610 ;
        RECT 89.990 173.410 90.310 173.470 ;
        RECT 91.830 173.410 92.150 173.470 ;
        RECT 93.670 173.410 93.990 173.470 ;
        RECT 95.050 173.610 95.370 173.670 ;
        RECT 95.050 173.470 96.660 173.610 ;
        RECT 95.050 173.410 95.370 173.470 ;
        RECT 64.705 173.270 64.995 173.315 ;
        RECT 64.320 173.130 64.995 173.270 ;
        RECT 47.225 173.085 47.515 173.130 ;
        RECT 46.290 173.070 46.610 173.085 ;
        RECT 48.130 173.070 48.450 173.130 ;
        RECT 43.545 172.930 43.835 172.975 ;
        RECT 43.545 172.790 47.210 172.930 ;
        RECT 43.545 172.745 43.835 172.790 ;
        RECT 42.150 172.390 42.470 172.650 ;
        RECT 47.070 172.590 47.210 172.790 ;
        RECT 47.670 172.730 47.990 172.990 ;
        RECT 49.140 172.975 49.280 173.130 ;
        RECT 60.550 173.070 60.870 173.130 ;
        RECT 64.705 173.085 64.995 173.130 ;
        RECT 65.610 173.270 65.930 173.330 ;
        RECT 74.810 173.270 75.130 173.330 ;
        RECT 76.190 173.270 76.510 173.330 ;
        RECT 65.610 173.130 69.015 173.270 ;
        RECT 65.610 173.070 65.930 173.130 ;
        RECT 49.065 172.745 49.355 172.975 ;
        RECT 49.985 172.745 50.275 172.975 ;
        RECT 50.445 172.930 50.735 172.975 ;
        RECT 51.350 172.930 51.670 172.990 ;
        RECT 50.445 172.790 51.670 172.930 ;
        RECT 50.445 172.745 50.735 172.790 ;
        RECT 49.510 172.590 49.830 172.650 ;
        RECT 47.070 172.450 49.830 172.590 ;
        RECT 49.510 172.390 49.830 172.450 ;
        RECT 50.060 172.250 50.200 172.745 ;
        RECT 51.350 172.730 51.670 172.790 ;
        RECT 51.810 172.930 52.130 172.990 ;
        RECT 53.190 172.930 53.510 172.990 ;
        RECT 51.810 172.790 53.510 172.930 ;
        RECT 51.810 172.730 52.130 172.790 ;
        RECT 53.190 172.730 53.510 172.790 ;
        RECT 54.125 172.745 54.415 172.975 ;
        RECT 56.425 172.930 56.715 172.975 ;
        RECT 57.330 172.930 57.650 172.990 ;
        RECT 54.660 172.790 57.650 172.930 ;
        RECT 51.440 172.590 51.580 172.730 ;
        RECT 54.200 172.590 54.340 172.745 ;
        RECT 54.660 172.650 54.800 172.790 ;
        RECT 56.425 172.745 56.715 172.790 ;
        RECT 57.330 172.730 57.650 172.790 ;
        RECT 62.850 172.930 63.170 172.990 ;
        RECT 63.400 172.930 64.460 172.960 ;
        RECT 66.085 172.930 66.375 172.975 ;
        RECT 62.850 172.820 66.375 172.930 ;
        RECT 62.850 172.790 63.540 172.820 ;
        RECT 64.320 172.790 66.375 172.820 ;
        RECT 62.850 172.730 63.170 172.790 ;
        RECT 66.085 172.745 66.375 172.790 ;
        RECT 66.545 172.930 66.835 172.975 ;
        RECT 66.990 172.930 67.310 172.990 ;
        RECT 66.545 172.790 67.310 172.930 ;
        RECT 66.545 172.745 66.835 172.790 ;
        RECT 66.990 172.730 67.310 172.790 ;
        RECT 68.370 172.730 68.690 172.990 ;
        RECT 68.875 172.930 69.015 173.130 ;
        RECT 72.600 173.130 76.510 173.270 ;
        RECT 72.600 172.975 72.740 173.130 ;
        RECT 74.810 173.070 75.130 173.130 ;
        RECT 76.190 173.070 76.510 173.130 ;
        RECT 78.490 173.070 78.810 173.330 ;
        RECT 86.770 173.270 87.090 173.330 ;
        RECT 89.160 173.270 89.300 173.410 ;
        RECT 96.520 173.330 96.660 173.470 ;
        RECT 99.190 173.410 99.510 173.670 ;
        RECT 100.570 173.410 100.890 173.670 ;
        RECT 103.345 173.610 103.635 173.655 ;
        RECT 117.130 173.610 117.450 173.670 ;
        RECT 103.345 173.470 107.700 173.610 ;
        RECT 103.345 173.425 103.635 173.470 ;
        RECT 86.770 173.130 88.380 173.270 ;
        RECT 89.160 173.130 91.140 173.270 ;
        RECT 86.770 173.070 87.090 173.130 ;
        RECT 68.875 172.790 70.440 172.930 ;
        RECT 51.440 172.450 54.340 172.590 ;
        RECT 54.200 172.250 54.340 172.450 ;
        RECT 54.570 172.390 54.890 172.650 ;
        RECT 61.470 172.590 61.790 172.650 ;
        RECT 63.785 172.590 64.075 172.635 ;
        RECT 64.705 172.590 64.995 172.635 ;
        RECT 69.765 172.590 70.055 172.635 ;
        RECT 61.470 172.450 70.055 172.590 ;
        RECT 70.300 172.590 70.440 172.790 ;
        RECT 72.525 172.745 72.815 172.975 ;
        RECT 75.240 172.930 75.530 172.975 ;
        RECT 81.250 172.930 81.570 172.990 ;
        RECT 88.240 172.975 88.380 173.130 ;
        RECT 75.240 172.790 81.570 172.930 ;
        RECT 75.240 172.745 75.530 172.790 ;
        RECT 81.250 172.730 81.570 172.790 ;
        RECT 86.325 172.745 86.615 172.975 ;
        RECT 87.245 172.745 87.535 172.975 ;
        RECT 88.165 172.745 88.455 172.975 ;
        RECT 88.610 172.930 88.930 172.990 ;
        RECT 89.085 172.930 89.375 172.975 ;
        RECT 88.610 172.790 89.375 172.930 ;
        RECT 73.905 172.590 74.195 172.635 ;
        RECT 70.300 172.450 74.195 172.590 ;
        RECT 61.470 172.390 61.790 172.450 ;
        RECT 63.785 172.405 64.075 172.450 ;
        RECT 64.705 172.405 64.995 172.450 ;
        RECT 69.765 172.405 70.055 172.450 ;
        RECT 73.905 172.405 74.195 172.450 ;
        RECT 74.785 172.590 75.075 172.635 ;
        RECT 75.975 172.590 76.265 172.635 ;
        RECT 78.495 172.590 78.785 172.635 ;
        RECT 74.785 172.450 78.785 172.590 ;
        RECT 74.785 172.405 75.075 172.450 ;
        RECT 75.975 172.405 76.265 172.450 ;
        RECT 78.495 172.405 78.785 172.450 ;
        RECT 80.330 172.390 80.650 172.650 ;
        RECT 55.505 172.250 55.795 172.295 ;
        RECT 50.060 172.110 52.960 172.250 ;
        RECT 54.200 172.110 55.795 172.250 ;
        RECT 43.070 171.710 43.390 171.970 ;
        RECT 46.305 171.910 46.595 171.955 ;
        RECT 47.670 171.910 47.990 171.970 ;
        RECT 46.305 171.770 47.990 171.910 ;
        RECT 46.305 171.725 46.595 171.770 ;
        RECT 47.670 171.710 47.990 171.770 ;
        RECT 48.605 171.910 48.895 171.955 ;
        RECT 52.270 171.910 52.590 171.970 ;
        RECT 48.605 171.770 52.590 171.910 ;
        RECT 52.820 171.910 52.960 172.110 ;
        RECT 55.505 172.065 55.795 172.110 ;
        RECT 65.165 172.250 65.455 172.295 ;
        RECT 69.305 172.250 69.595 172.295 ;
        RECT 65.165 172.110 69.595 172.250 ;
        RECT 65.165 172.065 65.455 172.110 ;
        RECT 69.305 172.065 69.595 172.110 ;
        RECT 71.145 172.250 71.435 172.295 ;
        RECT 74.390 172.250 74.680 172.295 ;
        RECT 76.490 172.250 76.780 172.295 ;
        RECT 78.060 172.250 78.350 172.295 ;
        RECT 71.145 172.110 74.120 172.250 ;
        RECT 71.145 172.065 71.435 172.110 ;
        RECT 54.110 171.910 54.430 171.970 ;
        RECT 52.820 171.770 54.430 171.910 ;
        RECT 48.605 171.725 48.895 171.770 ;
        RECT 52.270 171.710 52.590 171.770 ;
        RECT 54.110 171.710 54.430 171.770 ;
        RECT 55.045 171.910 55.335 171.955 ;
        RECT 58.710 171.910 59.030 171.970 ;
        RECT 64.690 171.910 65.010 171.970 ;
        RECT 55.045 171.770 65.010 171.910 ;
        RECT 55.045 171.725 55.335 171.770 ;
        RECT 58.710 171.710 59.030 171.770 ;
        RECT 64.690 171.710 65.010 171.770 ;
        RECT 65.625 171.910 65.915 171.955 ;
        RECT 67.005 171.910 67.295 171.955 ;
        RECT 65.625 171.770 67.295 171.910 ;
        RECT 65.625 171.725 65.915 171.770 ;
        RECT 67.005 171.725 67.295 171.770 ;
        RECT 67.925 171.910 68.215 171.955 ;
        RECT 70.225 171.910 70.515 171.955 ;
        RECT 67.925 171.770 70.515 171.910 ;
        RECT 67.925 171.725 68.215 171.770 ;
        RECT 70.225 171.725 70.515 171.770 ;
        RECT 73.430 171.710 73.750 171.970 ;
        RECT 73.980 171.910 74.120 172.110 ;
        RECT 74.390 172.110 78.350 172.250 ;
        RECT 80.420 172.250 80.560 172.390 ;
        RECT 80.805 172.250 81.095 172.295 ;
        RECT 80.420 172.110 81.095 172.250 ;
        RECT 74.390 172.065 74.680 172.110 ;
        RECT 76.490 172.065 76.780 172.110 ;
        RECT 78.060 172.065 78.350 172.110 ;
        RECT 80.805 172.065 81.095 172.110 ;
        RECT 86.400 171.970 86.540 172.745 ;
        RECT 87.320 172.590 87.460 172.745 ;
        RECT 88.610 172.730 88.930 172.790 ;
        RECT 89.085 172.745 89.375 172.790 ;
        RECT 89.545 172.745 89.835 172.975 ;
        RECT 89.620 172.590 89.760 172.745 ;
        RECT 89.990 172.730 90.310 172.990 ;
        RECT 91.000 172.975 91.140 173.130 ;
        RECT 96.430 173.070 96.750 173.330 ;
        RECT 99.280 173.270 99.420 173.410 ;
        RECT 100.660 173.270 100.800 173.410 ;
        RECT 99.280 173.130 100.340 173.270 ;
        RECT 100.660 173.130 104.940 173.270 ;
        RECT 90.925 172.745 91.215 172.975 ;
        RECT 91.370 172.730 91.690 172.990 ;
        RECT 92.750 172.930 93.070 172.990 ;
        RECT 94.605 172.930 94.895 172.975 ;
        RECT 92.750 172.790 94.895 172.930 ;
        RECT 92.750 172.730 93.070 172.790 ;
        RECT 94.605 172.745 94.895 172.790 ;
        RECT 99.665 172.745 99.955 172.975 ;
        RECT 100.200 172.930 100.340 173.130 ;
        RECT 100.585 172.930 100.875 172.975 ;
        RECT 100.200 172.790 100.875 172.930 ;
        RECT 100.585 172.745 100.875 172.790 ;
        RECT 101.950 172.930 102.270 172.990 ;
        RECT 102.425 172.930 102.715 172.975 ;
        RECT 101.950 172.790 102.715 172.930 ;
        RECT 91.460 172.590 91.600 172.730 ;
        RECT 93.225 172.590 93.515 172.635 ;
        RECT 87.320 172.450 91.600 172.590 ;
        RECT 92.840 172.450 93.515 172.590 ;
        RECT 86.785 172.250 87.075 172.295 ;
        RECT 87.690 172.250 88.010 172.310 ;
        RECT 86.785 172.110 88.010 172.250 ;
        RECT 86.785 172.065 87.075 172.110 ;
        RECT 87.690 172.050 88.010 172.110 ;
        RECT 88.700 172.110 92.520 172.250 ;
        RECT 80.330 171.910 80.650 171.970 ;
        RECT 73.980 171.770 80.650 171.910 ;
        RECT 80.330 171.710 80.650 171.770 ;
        RECT 86.310 171.710 86.630 171.970 ;
        RECT 87.230 171.910 87.550 171.970 ;
        RECT 88.700 171.910 88.840 172.110 ;
        RECT 87.230 171.770 88.840 171.910 ;
        RECT 89.530 171.910 89.850 171.970 ;
        RECT 92.380 171.955 92.520 172.110 ;
        RECT 92.840 171.970 92.980 172.450 ;
        RECT 93.225 172.405 93.515 172.450 ;
        RECT 93.670 172.390 93.990 172.650 ;
        RECT 94.145 172.405 94.435 172.635 ;
        RECT 96.890 172.590 97.210 172.650 ;
        RECT 99.740 172.590 99.880 172.745 ;
        RECT 101.950 172.730 102.270 172.790 ;
        RECT 102.425 172.745 102.715 172.790 ;
        RECT 103.330 172.730 103.650 172.990 ;
        RECT 103.790 172.730 104.110 172.990 ;
        RECT 104.800 172.975 104.940 173.130 ;
        RECT 104.725 172.745 105.015 172.975 ;
        RECT 106.105 172.930 106.395 172.975 ;
        RECT 107.010 172.930 107.330 172.990 ;
        RECT 107.560 172.975 107.700 173.470 ;
        RECT 116.300 173.470 117.450 173.610 ;
        RECT 111.610 173.270 111.930 173.330 ;
        RECT 113.910 173.270 114.230 173.330 ;
        RECT 111.610 173.130 114.230 173.270 ;
        RECT 111.610 173.070 111.930 173.130 ;
        RECT 113.910 173.070 114.230 173.130 ;
        RECT 116.300 172.975 116.440 173.470 ;
        RECT 117.130 173.410 117.450 173.470 ;
        RECT 118.510 173.610 118.830 173.670 ;
        RECT 120.350 173.610 120.670 173.670 ;
        RECT 118.510 173.470 120.670 173.610 ;
        RECT 118.510 173.410 118.830 173.470 ;
        RECT 120.350 173.410 120.670 173.470 ;
        RECT 139.670 173.410 139.990 173.670 ;
        RECT 123.110 173.270 123.430 173.330 ;
        RECT 119.980 173.130 123.430 173.270 ;
        RECT 119.980 172.975 120.120 173.130 ;
        RECT 123.110 173.070 123.430 173.130 ;
        RECT 138.380 173.130 140.360 173.270 ;
        RECT 106.105 172.790 107.330 172.930 ;
        RECT 106.105 172.745 106.395 172.790 ;
        RECT 96.890 172.450 99.880 172.590 ;
        RECT 91.845 171.910 92.135 171.955 ;
        RECT 89.530 171.770 92.135 171.910 ;
        RECT 87.230 171.710 87.550 171.770 ;
        RECT 89.530 171.710 89.850 171.770 ;
        RECT 91.845 171.725 92.135 171.770 ;
        RECT 92.305 171.725 92.595 171.955 ;
        RECT 92.750 171.710 93.070 171.970 ;
        RECT 94.220 171.910 94.360 172.405 ;
        RECT 96.890 172.390 97.210 172.450 ;
        RECT 101.045 172.405 101.335 172.635 ;
        RECT 101.505 172.590 101.795 172.635 ;
        RECT 103.420 172.590 103.560 172.730 ;
        RECT 101.505 172.450 103.560 172.590 ;
        RECT 104.800 172.590 104.940 172.745 ;
        RECT 107.010 172.730 107.330 172.790 ;
        RECT 107.485 172.745 107.775 172.975 ;
        RECT 116.225 172.745 116.515 172.975 ;
        RECT 119.905 172.930 120.195 172.975 ;
        RECT 116.760 172.790 120.195 172.930 ;
        RECT 116.760 172.590 116.900 172.790 ;
        RECT 119.905 172.745 120.195 172.790 ;
        RECT 120.825 172.745 121.115 172.975 ;
        RECT 121.285 172.930 121.575 172.975 ;
        RECT 122.650 172.930 122.970 172.990 ;
        RECT 121.285 172.790 122.970 172.930 ;
        RECT 121.285 172.745 121.575 172.790 ;
        RECT 119.430 172.590 119.750 172.650 ;
        RECT 120.900 172.590 121.040 172.745 ;
        RECT 122.650 172.730 122.970 172.790 ;
        RECT 135.070 172.930 135.390 172.990 ;
        RECT 138.380 172.930 138.520 173.130 ;
        RECT 135.070 172.790 138.520 172.930 ;
        RECT 135.070 172.730 135.390 172.790 ;
        RECT 138.765 172.745 139.055 172.975 ;
        RECT 140.220 172.930 140.360 173.130 ;
        RECT 141.065 172.930 141.355 172.975 ;
        RECT 140.220 172.790 141.355 172.930 ;
        RECT 141.065 172.745 141.355 172.790 ;
        RECT 141.985 172.930 142.275 172.975 ;
        RECT 142.430 172.930 142.750 172.990 ;
        RECT 141.985 172.790 142.750 172.930 ;
        RECT 141.985 172.745 142.275 172.790 ;
        RECT 104.800 172.450 116.900 172.590 ;
        RECT 117.220 172.450 121.040 172.590 ;
        RECT 101.505 172.405 101.795 172.450 ;
        RECT 98.730 172.250 99.050 172.310 ;
        RECT 100.570 172.250 100.890 172.310 ;
        RECT 98.730 172.110 100.890 172.250 ;
        RECT 101.120 172.250 101.260 172.405 ;
        RECT 102.870 172.250 103.190 172.310 ;
        RECT 117.220 172.295 117.360 172.450 ;
        RECT 119.430 172.390 119.750 172.450 ;
        RECT 126.790 172.390 127.110 172.650 ;
        RECT 138.840 172.590 138.980 172.745 ;
        RECT 142.430 172.730 142.750 172.790 ;
        RECT 142.890 172.930 143.210 172.990 ;
        RECT 143.365 172.930 143.655 172.975 ;
        RECT 142.890 172.790 143.655 172.930 ;
        RECT 142.890 172.730 143.210 172.790 ;
        RECT 143.365 172.745 143.655 172.790 ;
        RECT 138.840 172.450 142.200 172.590 ;
        RECT 117.145 172.250 117.435 172.295 ;
        RECT 101.120 172.110 103.190 172.250 ;
        RECT 98.730 172.050 99.050 172.110 ;
        RECT 100.570 172.050 100.890 172.110 ;
        RECT 102.870 172.050 103.190 172.110 ;
        RECT 103.880 172.110 117.435 172.250 ;
        RECT 103.880 171.910 104.020 172.110 ;
        RECT 117.145 172.065 117.435 172.110 ;
        RECT 119.905 172.250 120.195 172.295 ;
        RECT 126.880 172.250 127.020 172.390 ;
        RECT 119.905 172.110 127.020 172.250 ;
        RECT 119.905 172.065 120.195 172.110 ;
        RECT 142.060 171.970 142.200 172.450 ;
        RECT 94.220 171.770 104.020 171.910 ;
        RECT 104.265 171.910 104.555 171.955 ;
        RECT 105.630 171.910 105.950 171.970 ;
        RECT 104.265 171.770 105.950 171.910 ;
        RECT 104.265 171.725 104.555 171.770 ;
        RECT 105.630 171.710 105.950 171.770 ;
        RECT 106.550 171.910 106.870 171.970 ;
        RECT 107.930 171.910 108.250 171.970 ;
        RECT 106.550 171.770 108.250 171.910 ;
        RECT 106.550 171.710 106.870 171.770 ;
        RECT 107.930 171.710 108.250 171.770 ;
        RECT 108.405 171.910 108.695 171.955 ;
        RECT 108.850 171.910 109.170 171.970 ;
        RECT 108.405 171.770 109.170 171.910 ;
        RECT 108.405 171.725 108.695 171.770 ;
        RECT 108.850 171.710 109.170 171.770 ;
        RECT 136.910 171.910 137.230 171.970 ;
        RECT 137.845 171.910 138.135 171.955 ;
        RECT 136.910 171.770 138.135 171.910 ;
        RECT 136.910 171.710 137.230 171.770 ;
        RECT 137.845 171.725 138.135 171.770 ;
        RECT 141.510 171.710 141.830 171.970 ;
        RECT 141.970 171.910 142.290 171.970 ;
        RECT 142.445 171.910 142.735 171.955 ;
        RECT 141.970 171.770 142.735 171.910 ;
        RECT 141.970 171.710 142.290 171.770 ;
        RECT 142.445 171.725 142.735 171.770 ;
        RECT 36.100 171.090 150.180 171.570 ;
        RECT 43.070 170.890 43.390 170.950 ;
        RECT 44.465 170.890 44.755 170.935 ;
        RECT 43.070 170.750 44.755 170.890 ;
        RECT 43.070 170.690 43.390 170.750 ;
        RECT 44.465 170.705 44.755 170.750 ;
        RECT 45.370 170.890 45.690 170.950 ;
        RECT 46.290 170.890 46.610 170.950 ;
        RECT 45.370 170.750 46.610 170.890 ;
        RECT 41.245 170.550 41.535 170.595 ;
        RECT 41.690 170.550 42.010 170.610 ;
        RECT 41.245 170.410 43.760 170.550 ;
        RECT 41.245 170.365 41.535 170.410 ;
        RECT 41.690 170.350 42.010 170.410 ;
        RECT 42.150 170.010 42.470 170.270 ;
        RECT 40.785 169.685 41.075 169.915 ;
        RECT 40.860 169.190 41.000 169.685 ;
        RECT 43.070 169.670 43.390 169.930 ;
        RECT 43.620 169.915 43.760 170.410 ;
        RECT 44.540 170.210 44.680 170.705 ;
        RECT 45.370 170.690 45.690 170.750 ;
        RECT 46.290 170.690 46.610 170.750 ;
        RECT 47.225 170.890 47.515 170.935 ;
        RECT 51.350 170.890 51.670 170.950 ;
        RECT 47.225 170.750 51.670 170.890 ;
        RECT 47.225 170.705 47.515 170.750 ;
        RECT 51.350 170.690 51.670 170.750 ;
        RECT 61.010 170.890 61.330 170.950 ;
        RECT 63.310 170.890 63.630 170.950 ;
        RECT 61.010 170.750 63.630 170.890 ;
        RECT 61.010 170.690 61.330 170.750 ;
        RECT 63.310 170.690 63.630 170.750 ;
        RECT 64.245 170.890 64.535 170.935 ;
        RECT 65.625 170.890 65.915 170.935 ;
        RECT 64.245 170.750 65.915 170.890 ;
        RECT 64.245 170.705 64.535 170.750 ;
        RECT 65.625 170.705 65.915 170.750 ;
        RECT 66.545 170.890 66.835 170.935 ;
        RECT 68.845 170.890 69.135 170.935 ;
        RECT 66.545 170.750 69.135 170.890 ;
        RECT 66.545 170.705 66.835 170.750 ;
        RECT 68.845 170.705 69.135 170.750 ;
        RECT 76.190 170.690 76.510 170.950 ;
        RECT 85.850 170.890 86.170 170.950 ;
        RECT 81.570 170.750 86.170 170.890 ;
        RECT 63.785 170.550 64.075 170.595 ;
        RECT 67.925 170.550 68.215 170.595 ;
        RECT 63.785 170.410 68.215 170.550 ;
        RECT 63.785 170.365 64.075 170.410 ;
        RECT 67.925 170.365 68.215 170.410 ;
        RECT 73.430 170.550 73.750 170.610 ;
        RECT 78.045 170.550 78.335 170.595 ;
        RECT 73.430 170.410 78.335 170.550 ;
        RECT 73.430 170.350 73.750 170.410 ;
        RECT 78.045 170.365 78.335 170.410 ;
        RECT 78.490 170.550 78.810 170.610 ;
        RECT 81.570 170.550 81.710 170.750 ;
        RECT 85.850 170.690 86.170 170.750 ;
        RECT 86.310 170.890 86.630 170.950 ;
        RECT 93.670 170.890 93.990 170.950 ;
        RECT 86.310 170.750 93.990 170.890 ;
        RECT 86.310 170.690 86.630 170.750 ;
        RECT 93.670 170.690 93.990 170.750 ;
        RECT 97.350 170.890 97.670 170.950 ;
        RECT 121.270 170.890 121.590 170.950 ;
        RECT 136.910 170.890 137.230 170.950 ;
        RECT 137.845 170.890 138.135 170.935 ;
        RECT 97.350 170.750 102.180 170.890 ;
        RECT 97.350 170.690 97.670 170.750 ;
        RECT 102.040 170.610 102.180 170.750 ;
        RECT 121.270 170.750 138.135 170.890 ;
        RECT 121.270 170.690 121.590 170.750 ;
        RECT 136.910 170.690 137.230 170.750 ;
        RECT 137.845 170.705 138.135 170.750 ;
        RECT 142.430 170.890 142.750 170.950 ;
        RECT 147.505 170.890 147.795 170.935 ;
        RECT 142.430 170.750 147.795 170.890 ;
        RECT 142.430 170.690 142.750 170.750 ;
        RECT 147.505 170.705 147.795 170.750 ;
        RECT 90.910 170.550 91.230 170.610 ;
        RECT 101.950 170.550 102.270 170.610 ;
        RECT 102.885 170.550 103.175 170.595 ;
        RECT 78.490 170.410 81.710 170.550 ;
        RECT 87.780 170.410 89.300 170.550 ;
        RECT 78.490 170.350 78.810 170.410 ;
        RECT 87.780 170.270 87.920 170.410 ;
        RECT 52.270 170.210 52.590 170.270 ;
        RECT 61.930 170.210 62.250 170.270 ;
        RECT 62.405 170.210 62.695 170.255 ;
        RECT 63.325 170.210 63.615 170.255 ;
        RECT 68.385 170.210 68.675 170.255 ;
        RECT 44.540 170.070 45.140 170.210 ;
        RECT 43.545 169.870 43.835 169.915 ;
        RECT 44.450 169.870 44.770 169.930 ;
        RECT 45.000 169.915 45.140 170.070 ;
        RECT 52.270 170.070 61.700 170.210 ;
        RECT 52.270 170.010 52.590 170.070 ;
        RECT 43.545 169.730 44.770 169.870 ;
        RECT 43.545 169.685 43.835 169.730 ;
        RECT 44.450 169.670 44.770 169.730 ;
        RECT 44.925 169.685 45.215 169.915 ;
        RECT 45.845 169.685 46.135 169.915 ;
        RECT 42.165 169.530 42.455 169.575 ;
        RECT 45.920 169.530 46.060 169.685 ;
        RECT 61.010 169.670 61.330 169.930 ;
        RECT 61.560 169.870 61.700 170.070 ;
        RECT 61.930 170.070 68.675 170.210 ;
        RECT 61.930 170.010 62.250 170.070 ;
        RECT 62.405 170.025 62.695 170.070 ;
        RECT 63.325 170.025 63.615 170.070 ;
        RECT 68.385 170.025 68.675 170.070 ;
        RECT 68.830 170.210 69.150 170.270 ;
        RECT 87.690 170.210 88.010 170.270 ;
        RECT 89.160 170.255 89.300 170.410 ;
        RECT 89.620 170.410 91.230 170.550 ;
        RECT 89.620 170.255 89.760 170.410 ;
        RECT 90.910 170.350 91.230 170.410 ;
        RECT 91.920 170.410 101.720 170.550 ;
        RECT 68.830 170.070 88.010 170.210 ;
        RECT 68.830 170.010 69.150 170.070 ;
        RECT 87.690 170.010 88.010 170.070 ;
        RECT 89.085 170.025 89.375 170.255 ;
        RECT 89.545 170.025 89.835 170.255 ;
        RECT 90.005 170.210 90.295 170.255 ;
        RECT 90.450 170.210 90.770 170.270 ;
        RECT 91.920 170.255 92.060 170.410 ;
        RECT 90.005 170.070 90.770 170.210 ;
        RECT 90.005 170.025 90.295 170.070 ;
        RECT 90.450 170.010 90.770 170.070 ;
        RECT 91.840 170.025 92.130 170.255 ;
        RECT 92.750 170.010 93.070 170.270 ;
        RECT 101.580 170.210 101.720 170.410 ;
        RECT 101.950 170.410 103.175 170.550 ;
        RECT 101.950 170.350 102.270 170.410 ;
        RECT 102.885 170.365 103.175 170.410 ;
        RECT 104.250 170.550 104.570 170.610 ;
        RECT 108.390 170.550 108.710 170.610 ;
        RECT 104.250 170.410 108.710 170.550 ;
        RECT 104.250 170.350 104.570 170.410 ;
        RECT 108.390 170.350 108.710 170.410 ;
        RECT 141.090 170.550 141.380 170.595 ;
        RECT 143.190 170.550 143.480 170.595 ;
        RECT 144.760 170.550 145.050 170.595 ;
        RECT 141.090 170.410 145.050 170.550 ;
        RECT 141.090 170.365 141.380 170.410 ;
        RECT 143.190 170.365 143.480 170.410 ;
        RECT 144.760 170.365 145.050 170.410 ;
        RECT 101.580 170.070 108.620 170.210 ;
        RECT 108.480 169.930 108.620 170.070 ;
        RECT 109.770 170.010 110.090 170.270 ;
        RECT 127.250 170.210 127.570 170.270 ;
        RECT 122.740 170.070 124.260 170.210 ;
        RECT 122.740 169.930 122.880 170.070 ;
        RECT 64.230 169.870 64.550 169.930 ;
        RECT 64.705 169.870 64.995 169.915 ;
        RECT 61.560 169.730 64.000 169.870 ;
        RECT 42.165 169.390 46.060 169.530 ;
        RECT 48.145 169.530 48.435 169.575 ;
        RECT 58.250 169.530 58.570 169.590 ;
        RECT 48.145 169.390 58.570 169.530 ;
        RECT 42.165 169.345 42.455 169.390 ;
        RECT 48.145 169.345 48.435 169.390 ;
        RECT 58.250 169.330 58.570 169.390 ;
        RECT 60.550 169.530 60.870 169.590 ;
        RECT 63.325 169.530 63.615 169.575 ;
        RECT 60.550 169.390 63.615 169.530 ;
        RECT 63.860 169.530 64.000 169.730 ;
        RECT 64.230 169.730 64.995 169.870 ;
        RECT 64.230 169.670 64.550 169.730 ;
        RECT 64.705 169.685 64.995 169.730 ;
        RECT 65.165 169.870 65.455 169.915 ;
        RECT 66.070 169.870 66.390 169.930 ;
        RECT 86.310 169.870 86.630 169.930 ;
        RECT 65.165 169.730 66.390 169.870 ;
        RECT 65.165 169.685 65.455 169.730 ;
        RECT 66.070 169.670 66.390 169.730 ;
        RECT 66.620 169.730 86.630 169.870 ;
        RECT 66.620 169.530 66.760 169.730 ;
        RECT 86.310 169.670 86.630 169.730 ;
        RECT 88.625 169.870 88.915 169.915 ;
        RECT 90.910 169.870 91.230 169.930 ;
        RECT 88.625 169.730 91.230 169.870 ;
        RECT 88.625 169.685 88.915 169.730 ;
        RECT 90.910 169.670 91.230 169.730 ;
        RECT 91.370 169.670 91.690 169.930 ;
        RECT 92.355 169.685 92.645 169.915 ;
        RECT 101.965 169.870 102.255 169.915 ;
        RECT 102.410 169.870 102.730 169.930 ;
        RECT 93.760 169.730 101.720 169.870 ;
        RECT 63.860 169.390 66.760 169.530 ;
        RECT 60.550 169.330 60.870 169.390 ;
        RECT 63.325 169.345 63.615 169.390 ;
        RECT 66.990 169.330 67.310 169.590 ;
        RECT 89.990 169.530 90.310 169.590 ;
        RECT 68.460 169.390 90.310 169.530 ;
        RECT 43.070 169.190 43.390 169.250 ;
        RECT 40.860 169.050 43.390 169.190 ;
        RECT 43.070 168.990 43.390 169.050 ;
        RECT 45.370 168.990 45.690 169.250 ;
        RECT 47.210 169.235 47.530 169.250 ;
        RECT 47.095 169.005 47.530 169.235 ;
        RECT 47.210 168.990 47.530 169.005 ;
        RECT 61.930 169.190 62.250 169.250 ;
        RECT 68.460 169.190 68.600 169.390 ;
        RECT 89.990 169.330 90.310 169.390 ;
        RECT 61.930 169.050 68.600 169.190 ;
        RECT 68.845 169.190 69.135 169.235 ;
        RECT 69.290 169.190 69.610 169.250 ;
        RECT 68.845 169.050 69.610 169.190 ;
        RECT 61.930 168.990 62.250 169.050 ;
        RECT 68.845 169.005 69.135 169.050 ;
        RECT 69.290 168.990 69.610 169.050 ;
        RECT 69.750 168.990 70.070 169.250 ;
        RECT 74.810 169.190 75.130 169.250 ;
        RECT 75.285 169.190 75.575 169.235 ;
        RECT 74.810 169.050 75.575 169.190 ;
        RECT 74.810 168.990 75.130 169.050 ;
        RECT 75.285 169.005 75.575 169.050 ;
        RECT 76.190 168.990 76.510 169.250 ;
        RECT 84.470 169.190 84.790 169.250 ;
        RECT 87.705 169.190 87.995 169.235 ;
        RECT 84.470 169.050 87.995 169.190 ;
        RECT 92.380 169.190 92.520 169.685 ;
        RECT 93.760 169.530 93.900 169.730 ;
        RECT 93.300 169.390 93.900 169.530 ;
        RECT 93.300 169.250 93.440 169.390 ;
        RECT 94.130 169.330 94.450 169.590 ;
        RECT 95.065 169.530 95.355 169.575 ;
        RECT 97.350 169.530 97.670 169.590 ;
        RECT 95.065 169.390 97.670 169.530 ;
        RECT 101.580 169.530 101.720 169.730 ;
        RECT 101.965 169.730 102.730 169.870 ;
        RECT 101.965 169.685 102.255 169.730 ;
        RECT 102.410 169.670 102.730 169.730 ;
        RECT 102.870 169.870 103.190 169.930 ;
        RECT 103.345 169.870 103.635 169.915 ;
        RECT 102.870 169.730 103.635 169.870 ;
        RECT 102.870 169.670 103.190 169.730 ;
        RECT 103.345 169.685 103.635 169.730 ;
        RECT 107.485 169.685 107.775 169.915 ;
        RECT 107.560 169.530 107.700 169.685 ;
        RECT 108.390 169.670 108.710 169.930 ;
        RECT 108.850 169.870 109.170 169.930 ;
        RECT 109.325 169.870 109.615 169.915 ;
        RECT 108.850 169.730 109.615 169.870 ;
        RECT 108.850 169.670 109.170 169.730 ;
        RECT 109.325 169.685 109.615 169.730 ;
        RECT 110.245 169.685 110.535 169.915 ;
        RECT 110.705 169.870 110.995 169.915 ;
        RECT 113.925 169.870 114.215 169.915 ;
        RECT 110.705 169.730 114.215 169.870 ;
        RECT 110.705 169.685 110.995 169.730 ;
        RECT 113.925 169.685 114.215 169.730 ;
        RECT 115.305 169.870 115.595 169.915 ;
        RECT 117.590 169.870 117.910 169.930 ;
        RECT 115.305 169.730 122.420 169.870 ;
        RECT 115.305 169.685 115.595 169.730 ;
        RECT 101.580 169.390 107.700 169.530 ;
        RECT 95.065 169.345 95.355 169.390 ;
        RECT 97.350 169.330 97.670 169.390 ;
        RECT 93.210 169.190 93.530 169.250 ;
        RECT 92.380 169.050 93.530 169.190 ;
        RECT 84.470 168.990 84.790 169.050 ;
        RECT 87.705 169.005 87.995 169.050 ;
        RECT 93.210 168.990 93.530 169.050 ;
        RECT 93.685 169.190 93.975 169.235 ;
        RECT 94.590 169.190 94.910 169.250 ;
        RECT 93.685 169.050 94.910 169.190 ;
        RECT 93.685 169.005 93.975 169.050 ;
        RECT 94.590 168.990 94.910 169.050 ;
        RECT 95.970 168.990 96.290 169.250 ;
        RECT 98.270 169.190 98.590 169.250 ;
        RECT 101.045 169.190 101.335 169.235 ;
        RECT 98.270 169.050 101.335 169.190 ;
        RECT 107.560 169.190 107.700 169.390 ;
        RECT 107.945 169.530 108.235 169.575 ;
        RECT 110.320 169.530 110.460 169.685 ;
        RECT 117.590 169.670 117.910 169.730 ;
        RECT 122.280 169.590 122.420 169.730 ;
        RECT 122.650 169.670 122.970 169.930 ;
        RECT 123.110 169.670 123.430 169.930 ;
        RECT 124.120 169.915 124.260 170.070 ;
        RECT 125.040 170.070 128.860 170.210 ;
        RECT 125.040 169.930 125.180 170.070 ;
        RECT 127.250 170.010 127.570 170.070 ;
        RECT 124.045 169.685 124.335 169.915 ;
        RECT 124.950 169.670 125.270 169.930 ;
        RECT 128.720 169.915 128.860 170.070 ;
        RECT 138.290 170.010 138.610 170.270 ;
        RECT 139.670 170.210 139.990 170.270 ;
        RECT 140.605 170.210 140.895 170.255 ;
        RECT 138.840 170.070 140.895 170.210 ;
        RECT 126.805 169.685 127.095 169.915 ;
        RECT 128.645 169.685 128.935 169.915 ;
        RECT 132.310 169.870 132.630 169.930 ;
        RECT 138.840 169.870 138.980 170.070 ;
        RECT 139.670 170.010 139.990 170.070 ;
        RECT 140.605 170.025 140.895 170.070 ;
        RECT 141.485 170.210 141.775 170.255 ;
        RECT 142.675 170.210 142.965 170.255 ;
        RECT 145.195 170.210 145.485 170.255 ;
        RECT 141.485 170.070 145.485 170.210 ;
        RECT 141.485 170.025 141.775 170.070 ;
        RECT 142.675 170.025 142.965 170.070 ;
        RECT 145.195 170.025 145.485 170.070 ;
        RECT 132.310 169.730 138.980 169.870 ;
        RECT 112.085 169.530 112.375 169.575 ;
        RECT 107.945 169.390 110.460 169.530 ;
        RECT 110.780 169.390 112.375 169.530 ;
        RECT 107.945 169.345 108.235 169.390 ;
        RECT 110.780 169.190 110.920 169.390 ;
        RECT 112.085 169.345 112.375 169.390 ;
        RECT 112.990 169.530 113.310 169.590 ;
        RECT 112.990 169.390 114.600 169.530 ;
        RECT 112.990 169.330 113.310 169.390 ;
        RECT 107.560 169.050 110.920 169.190 ;
        RECT 111.625 169.190 111.915 169.235 ;
        RECT 113.910 169.190 114.230 169.250 ;
        RECT 114.460 169.235 114.600 169.390 ;
        RECT 122.190 169.330 122.510 169.590 ;
        RECT 123.585 169.530 123.875 169.575 ;
        RECT 126.880 169.530 127.020 169.685 ;
        RECT 132.310 169.670 132.630 169.730 ;
        RECT 139.225 169.685 139.515 169.915 ;
        RECT 123.585 169.390 127.020 169.530 ;
        RECT 123.585 169.345 123.875 169.390 ;
        RECT 127.725 169.345 128.015 169.575 ;
        RECT 128.185 169.345 128.475 169.575 ;
        RECT 111.625 169.050 114.230 169.190 ;
        RECT 98.270 168.990 98.590 169.050 ;
        RECT 101.045 169.005 101.335 169.050 ;
        RECT 111.625 169.005 111.915 169.050 ;
        RECT 113.910 168.990 114.230 169.050 ;
        RECT 114.385 169.005 114.675 169.235 ;
        RECT 124.030 169.190 124.350 169.250 ;
        RECT 127.800 169.190 127.940 169.345 ;
        RECT 124.030 169.050 127.940 169.190 ;
        RECT 128.260 169.190 128.400 169.345 ;
        RECT 137.830 169.330 138.150 169.590 ;
        RECT 138.290 169.530 138.610 169.590 ;
        RECT 139.300 169.530 139.440 169.685 ;
        RECT 141.830 169.530 142.120 169.575 ;
        RECT 138.290 169.390 139.440 169.530 ;
        RECT 139.760 169.390 142.120 169.530 ;
        RECT 138.290 169.330 138.610 169.390 ;
        RECT 128.630 169.190 128.950 169.250 ;
        RECT 128.260 169.050 128.950 169.190 ;
        RECT 124.030 168.990 124.350 169.050 ;
        RECT 128.630 168.990 128.950 169.050 ;
        RECT 129.565 169.190 129.855 169.235 ;
        RECT 139.760 169.190 139.900 169.390 ;
        RECT 141.830 169.345 142.120 169.390 ;
        RECT 129.565 169.050 139.900 169.190 ;
        RECT 140.145 169.190 140.435 169.235 ;
        RECT 141.050 169.190 141.370 169.250 ;
        RECT 140.145 169.050 141.370 169.190 ;
        RECT 129.565 169.005 129.855 169.050 ;
        RECT 140.145 169.005 140.435 169.050 ;
        RECT 141.050 168.990 141.370 169.050 ;
        RECT 36.100 168.370 150.180 168.850 ;
        RECT 43.070 168.170 43.390 168.230 ;
        RECT 52.270 168.170 52.590 168.230 ;
        RECT 43.070 168.030 52.590 168.170 ;
        RECT 43.070 167.970 43.390 168.030 ;
        RECT 52.270 167.970 52.590 168.030 ;
        RECT 60.550 168.170 60.870 168.230 ;
        RECT 66.990 168.170 67.310 168.230 ;
        RECT 60.550 168.030 67.310 168.170 ;
        RECT 60.550 167.970 60.870 168.030 ;
        RECT 66.990 167.970 67.310 168.030 ;
        RECT 68.370 168.170 68.690 168.230 ;
        RECT 69.290 168.170 69.610 168.230 ;
        RECT 68.370 168.030 69.610 168.170 ;
        RECT 68.370 167.970 68.690 168.030 ;
        RECT 69.290 167.970 69.610 168.030 ;
        RECT 73.905 168.170 74.195 168.215 ;
        RECT 74.350 168.170 74.670 168.230 ;
        RECT 73.905 168.030 74.670 168.170 ;
        RECT 73.905 167.985 74.195 168.030 ;
        RECT 74.350 167.970 74.670 168.030 ;
        RECT 75.270 167.970 75.590 168.230 ;
        RECT 75.745 168.170 76.035 168.215 ;
        RECT 76.190 168.170 76.510 168.230 ;
        RECT 81.710 168.170 82.030 168.230 ;
        RECT 75.745 168.030 76.510 168.170 ;
        RECT 75.745 167.985 76.035 168.030 ;
        RECT 76.190 167.970 76.510 168.030 ;
        RECT 76.740 168.030 82.030 168.170 ;
        RECT 43.530 167.630 43.850 167.890 ;
        RECT 66.530 167.830 66.850 167.890 ;
        RECT 73.445 167.830 73.735 167.875 ;
        RECT 76.740 167.830 76.880 168.030 ;
        RECT 81.710 167.970 82.030 168.030 ;
        RECT 91.370 167.970 91.690 168.230 ;
        RECT 93.670 168.170 93.990 168.230 ;
        RECT 94.590 168.170 94.910 168.230 ;
        RECT 93.670 168.030 94.910 168.170 ;
        RECT 93.670 167.970 93.990 168.030 ;
        RECT 94.590 167.970 94.910 168.030 ;
        RECT 95.970 167.970 96.290 168.230 ;
        RECT 97.350 167.970 97.670 168.230 ;
        RECT 107.930 168.170 108.250 168.230 ;
        RECT 103.420 168.030 108.250 168.170 ;
        RECT 90.910 167.830 91.230 167.890 ;
        RECT 93.210 167.830 93.530 167.890 ;
        RECT 45.000 167.690 47.210 167.830 ;
        RECT 37.550 167.490 37.870 167.550 ;
        RECT 45.000 167.535 45.140 167.690 ;
        RECT 44.925 167.490 45.215 167.535 ;
        RECT 37.550 167.350 45.215 167.490 ;
        RECT 37.550 167.290 37.870 167.350 ;
        RECT 44.925 167.305 45.215 167.350 ;
        RECT 45.370 167.490 45.690 167.550 ;
        RECT 46.205 167.490 46.495 167.535 ;
        RECT 45.370 167.350 46.495 167.490 ;
        RECT 47.070 167.490 47.210 167.690 ;
        RECT 62.480 167.690 65.840 167.830 ;
        RECT 58.250 167.490 58.570 167.550 ;
        RECT 62.480 167.535 62.620 167.690 ;
        RECT 65.700 167.550 65.840 167.690 ;
        RECT 66.530 167.690 76.880 167.830 ;
        RECT 78.580 167.690 90.220 167.830 ;
        RECT 66.530 167.630 66.850 167.690 ;
        RECT 73.445 167.645 73.735 167.690 ;
        RECT 78.580 167.550 78.720 167.690 ;
        RECT 62.405 167.490 62.695 167.535 ;
        RECT 47.070 167.350 62.695 167.490 ;
        RECT 45.370 167.290 45.690 167.350 ;
        RECT 46.205 167.305 46.495 167.350 ;
        RECT 58.250 167.290 58.570 167.350 ;
        RECT 62.405 167.305 62.695 167.350 ;
        RECT 62.850 167.490 63.170 167.550 ;
        RECT 63.685 167.490 63.975 167.535 ;
        RECT 62.850 167.350 63.975 167.490 ;
        RECT 62.850 167.290 63.170 167.350 ;
        RECT 63.685 167.305 63.975 167.350 ;
        RECT 65.610 167.290 65.930 167.550 ;
        RECT 68.830 167.290 69.150 167.550 ;
        RECT 71.145 167.490 71.435 167.535 ;
        RECT 72.525 167.490 72.815 167.535 ;
        RECT 74.365 167.490 74.655 167.535 ;
        RECT 76.665 167.490 76.955 167.535 ;
        RECT 71.145 167.350 72.815 167.490 ;
        RECT 71.145 167.305 71.435 167.350 ;
        RECT 72.525 167.305 72.815 167.350 ;
        RECT 73.060 167.350 76.955 167.490 ;
        RECT 78.490 167.480 78.810 167.550 ;
        RECT 41.690 166.950 42.010 167.210 ;
        RECT 45.805 167.150 46.095 167.195 ;
        RECT 46.995 167.150 47.285 167.195 ;
        RECT 49.515 167.150 49.805 167.195 ;
        RECT 45.805 167.010 49.805 167.150 ;
        RECT 45.805 166.965 46.095 167.010 ;
        RECT 46.995 166.965 47.285 167.010 ;
        RECT 49.515 166.965 49.805 167.010 ;
        RECT 49.970 167.150 50.290 167.210 ;
        RECT 49.970 167.010 58.480 167.150 ;
        RECT 49.970 166.950 50.290 167.010 ;
        RECT 45.410 166.810 45.700 166.855 ;
        RECT 47.510 166.810 47.800 166.855 ;
        RECT 49.080 166.810 49.370 166.855 ;
        RECT 43.620 166.670 45.140 166.810 ;
        RECT 43.620 166.515 43.760 166.670 ;
        RECT 43.545 166.285 43.835 166.515 ;
        RECT 44.450 166.270 44.770 166.530 ;
        RECT 45.000 166.470 45.140 166.670 ;
        RECT 45.410 166.670 49.370 166.810 ;
        RECT 45.410 166.625 45.700 166.670 ;
        RECT 47.510 166.625 47.800 166.670 ;
        RECT 49.080 166.625 49.370 166.670 ;
        RECT 51.440 166.670 58.020 166.810 ;
        RECT 51.440 166.470 51.580 166.670 ;
        RECT 45.000 166.330 51.580 166.470 ;
        RECT 51.810 166.270 52.130 166.530 ;
        RECT 57.880 166.515 58.020 166.670 ;
        RECT 57.805 166.285 58.095 166.515 ;
        RECT 58.340 166.470 58.480 167.010 ;
        RECT 58.710 166.950 59.030 167.210 ;
        RECT 59.185 166.965 59.475 167.195 ;
        RECT 59.260 166.810 59.400 166.965 ;
        RECT 59.630 166.950 59.950 167.210 ;
        RECT 60.105 167.150 60.395 167.195 ;
        RECT 61.930 167.150 62.250 167.210 ;
        RECT 60.105 167.010 62.250 167.150 ;
        RECT 60.105 166.965 60.395 167.010 ;
        RECT 61.930 166.950 62.250 167.010 ;
        RECT 63.285 167.150 63.575 167.195 ;
        RECT 64.475 167.150 64.765 167.195 ;
        RECT 66.995 167.150 67.285 167.195 ;
        RECT 63.285 167.010 67.285 167.150 ;
        RECT 63.285 166.965 63.575 167.010 ;
        RECT 64.475 166.965 64.765 167.010 ;
        RECT 66.995 166.965 67.285 167.010 ;
        RECT 61.470 166.810 61.790 166.870 ;
        RECT 59.260 166.670 61.790 166.810 ;
        RECT 61.470 166.610 61.790 166.670 ;
        RECT 62.890 166.810 63.180 166.855 ;
        RECT 64.990 166.810 65.280 166.855 ;
        RECT 66.560 166.810 66.850 166.855 ;
        RECT 68.920 166.810 69.060 167.290 ;
        RECT 71.220 167.150 71.360 167.305 ;
        RECT 73.060 167.210 73.200 167.350 ;
        RECT 74.365 167.305 74.655 167.350 ;
        RECT 76.665 167.305 76.955 167.350 ;
        RECT 77.660 167.340 78.810 167.480 ;
        RECT 62.890 166.670 66.850 166.810 ;
        RECT 62.890 166.625 63.180 166.670 ;
        RECT 64.990 166.625 65.280 166.670 ;
        RECT 66.560 166.625 66.850 166.670 ;
        RECT 67.080 166.670 69.060 166.810 ;
        RECT 69.380 167.010 71.360 167.150 ;
        RECT 67.080 166.470 67.220 166.670 ;
        RECT 69.380 166.530 69.520 167.010 ;
        RECT 72.970 166.950 73.290 167.210 ;
        RECT 75.270 167.150 75.590 167.210 ;
        RECT 77.660 167.195 77.800 167.340 ;
        RECT 78.490 167.290 78.810 167.340 ;
        RECT 78.965 167.490 79.255 167.535 ;
        RECT 79.870 167.490 80.190 167.550 ;
        RECT 78.965 167.350 80.190 167.490 ;
        RECT 78.965 167.305 79.255 167.350 ;
        RECT 79.870 167.290 80.190 167.350 ;
        RECT 81.250 167.290 81.570 167.550 ;
        RECT 84.010 167.490 84.330 167.550 ;
        RECT 87.245 167.490 87.535 167.535 ;
        RECT 84.010 167.350 87.535 167.490 ;
        RECT 84.010 167.290 84.330 167.350 ;
        RECT 87.245 167.305 87.535 167.350 ;
        RECT 87.690 167.290 88.010 167.550 ;
        RECT 88.150 167.290 88.470 167.550 ;
        RECT 90.080 167.535 90.220 167.690 ;
        RECT 90.910 167.690 93.530 167.830 ;
        RECT 90.910 167.630 91.230 167.690 ;
        RECT 93.210 167.630 93.530 167.690 ;
        RECT 89.085 167.305 89.375 167.535 ;
        RECT 89.545 167.305 89.835 167.535 ;
        RECT 90.005 167.305 90.295 167.535 ;
        RECT 92.290 167.490 92.610 167.550 ;
        RECT 94.605 167.490 94.895 167.535 ;
        RECT 92.290 167.350 94.895 167.490 ;
        RECT 77.125 167.150 77.415 167.195 ;
        RECT 75.270 167.010 77.415 167.150 ;
        RECT 75.270 166.950 75.590 167.010 ;
        RECT 77.125 166.965 77.415 167.010 ;
        RECT 77.585 166.965 77.875 167.195 ;
        RECT 78.045 166.965 78.335 167.195 ;
        RECT 79.410 167.150 79.730 167.210 ;
        RECT 81.340 167.150 81.480 167.290 ;
        RECT 79.410 167.010 81.480 167.150 ;
        RECT 87.780 167.150 87.920 167.290 ;
        RECT 89.160 167.150 89.300 167.305 ;
        RECT 87.780 167.010 89.300 167.150 ;
        RECT 72.065 166.810 72.355 166.855 ;
        RECT 78.120 166.810 78.260 166.965 ;
        RECT 79.410 166.950 79.730 167.010 ;
        RECT 89.070 166.810 89.390 166.870 ;
        RECT 72.065 166.670 89.390 166.810 ;
        RECT 72.065 166.625 72.355 166.670 ;
        RECT 89.070 166.610 89.390 166.670 ;
        RECT 58.340 166.330 67.220 166.470 ;
        RECT 69.290 166.270 69.610 166.530 ;
        RECT 72.970 166.470 73.290 166.530 ;
        RECT 78.490 166.470 78.810 166.530 ;
        RECT 72.970 166.330 78.810 166.470 ;
        RECT 72.970 166.270 73.290 166.330 ;
        RECT 78.490 166.270 78.810 166.330 ;
        RECT 86.325 166.470 86.615 166.515 ;
        RECT 87.230 166.470 87.550 166.530 ;
        RECT 86.325 166.330 87.550 166.470 ;
        RECT 89.620 166.470 89.760 167.305 ;
        RECT 92.290 167.290 92.610 167.350 ;
        RECT 94.605 167.305 94.895 167.350 ;
        RECT 95.525 167.490 95.815 167.535 ;
        RECT 96.060 167.490 96.200 167.970 ;
        RECT 97.440 167.830 97.580 167.970 ;
        RECT 103.420 167.890 103.560 168.030 ;
        RECT 107.930 167.970 108.250 168.030 ;
        RECT 108.390 168.170 108.710 168.230 ;
        RECT 110.705 168.170 110.995 168.215 ;
        RECT 108.390 168.030 110.995 168.170 ;
        RECT 108.390 167.970 108.710 168.030 ;
        RECT 110.705 167.985 110.995 168.030 ;
        RECT 112.990 167.970 113.310 168.230 ;
        RECT 118.510 168.170 118.830 168.230 ;
        RECT 121.270 168.170 121.590 168.230 ;
        RECT 118.510 168.030 121.590 168.170 ;
        RECT 118.510 167.970 118.830 168.030 ;
        RECT 121.270 167.970 121.590 168.030 ;
        RECT 121.745 168.170 122.035 168.215 ;
        RECT 123.110 168.170 123.430 168.230 ;
        RECT 121.745 168.030 123.430 168.170 ;
        RECT 121.745 167.985 122.035 168.030 ;
        RECT 123.110 167.970 123.430 168.030 ;
        RECT 127.725 168.170 128.015 168.215 ;
        RECT 138.765 168.170 139.055 168.215 ;
        RECT 127.725 168.030 130.700 168.170 ;
        RECT 127.725 167.985 128.015 168.030 ;
        RECT 103.330 167.830 103.650 167.890 ;
        RECT 112.070 167.830 112.390 167.890 ;
        RECT 97.440 167.690 103.650 167.830 ;
        RECT 95.525 167.350 96.200 167.490 ;
        RECT 95.525 167.305 95.815 167.350 ;
        RECT 96.890 167.290 97.210 167.550 ;
        RECT 94.215 166.965 94.505 167.195 ;
        RECT 94.220 166.810 94.360 166.965 ;
        RECT 95.050 166.950 95.370 167.210 ;
        RECT 97.440 167.150 97.580 167.690 ;
        RECT 103.330 167.630 103.650 167.690 ;
        RECT 108.020 167.690 112.390 167.830 ;
        RECT 97.825 167.490 98.115 167.535 ;
        RECT 99.190 167.490 99.510 167.550 ;
        RECT 97.825 167.350 99.510 167.490 ;
        RECT 97.825 167.305 98.115 167.350 ;
        RECT 99.190 167.290 99.510 167.350 ;
        RECT 99.650 167.290 99.970 167.550 ;
        RECT 100.585 167.490 100.875 167.535 ;
        RECT 101.965 167.490 102.255 167.535 ;
        RECT 108.020 167.490 108.160 167.690 ;
        RECT 112.070 167.630 112.390 167.690 ;
        RECT 100.585 167.350 102.255 167.490 ;
        RECT 100.585 167.305 100.875 167.350 ;
        RECT 101.965 167.305 102.255 167.350 ;
        RECT 102.500 167.350 108.160 167.490 ;
        RECT 98.285 167.150 98.575 167.195 ;
        RECT 97.440 167.010 98.575 167.150 ;
        RECT 98.285 166.965 98.575 167.010 ;
        RECT 98.745 167.150 99.035 167.195 ;
        RECT 102.500 167.150 102.640 167.350 ;
        RECT 108.390 167.290 108.710 167.550 ;
        RECT 110.245 167.490 110.535 167.535 ;
        RECT 111.150 167.490 111.470 167.550 ;
        RECT 110.245 167.350 111.470 167.490 ;
        RECT 110.245 167.305 110.535 167.350 ;
        RECT 111.150 167.290 111.470 167.350 ;
        RECT 111.625 167.490 111.915 167.535 ;
        RECT 113.080 167.490 113.220 167.970 ;
        RECT 119.430 167.830 119.750 167.890 ;
        RECT 125.885 167.830 126.175 167.875 ;
        RECT 128.645 167.830 128.935 167.875 ;
        RECT 117.680 167.690 119.200 167.830 ;
        RECT 117.680 167.550 117.820 167.690 ;
        RECT 111.625 167.350 113.220 167.490 ;
        RECT 111.625 167.305 111.915 167.350 ;
        RECT 117.590 167.290 117.910 167.550 ;
        RECT 118.510 167.290 118.830 167.550 ;
        RECT 119.060 167.535 119.200 167.690 ;
        RECT 119.430 167.690 125.640 167.830 ;
        RECT 119.430 167.630 119.750 167.690 ;
        RECT 118.985 167.305 119.275 167.535 ;
        RECT 121.285 167.305 121.575 167.535 ;
        RECT 122.205 167.490 122.495 167.535 ;
        RECT 123.585 167.490 123.875 167.535 ;
        RECT 122.205 167.350 123.875 167.490 ;
        RECT 122.205 167.305 122.495 167.350 ;
        RECT 123.585 167.305 123.875 167.350 ;
        RECT 124.030 167.490 124.350 167.550 ;
        RECT 124.965 167.490 125.255 167.535 ;
        RECT 124.030 167.350 125.255 167.490 ;
        RECT 125.500 167.490 125.640 167.690 ;
        RECT 125.885 167.690 128.935 167.830 ;
        RECT 130.560 167.830 130.700 168.030 ;
        RECT 138.765 168.030 141.280 168.170 ;
        RECT 138.765 167.985 139.055 168.030 ;
        RECT 133.090 167.830 133.380 167.875 ;
        RECT 130.560 167.690 133.380 167.830 ;
        RECT 125.885 167.645 126.175 167.690 ;
        RECT 128.645 167.645 128.935 167.690 ;
        RECT 133.090 167.645 133.380 167.690 ;
        RECT 141.140 167.830 141.280 168.030 ;
        RECT 143.810 167.970 144.130 168.230 ;
        RECT 141.140 167.690 144.500 167.830 ;
        RECT 126.345 167.490 126.635 167.535 ;
        RECT 125.500 167.350 126.635 167.490 ;
        RECT 98.745 167.010 102.640 167.150 ;
        RECT 102.870 167.150 103.190 167.210 ;
        RECT 103.345 167.150 103.635 167.195 ;
        RECT 102.870 167.010 103.635 167.150 ;
        RECT 98.745 166.965 99.035 167.010 ;
        RECT 102.870 166.950 103.190 167.010 ;
        RECT 103.345 166.965 103.635 167.010 ;
        RECT 106.550 166.950 106.870 167.210 ;
        RECT 107.930 166.950 108.250 167.210 ;
        RECT 108.480 167.150 108.620 167.290 ;
        RECT 121.360 167.150 121.500 167.305 ;
        RECT 108.480 167.010 121.500 167.150 ;
        RECT 101.045 166.810 101.335 166.855 ;
        RECT 94.220 166.670 101.335 166.810 ;
        RECT 101.045 166.625 101.335 166.670 ;
        RECT 95.970 166.470 96.290 166.530 ;
        RECT 89.620 166.330 96.290 166.470 ;
        RECT 86.325 166.285 86.615 166.330 ;
        RECT 87.230 166.270 87.550 166.330 ;
        RECT 95.970 166.270 96.290 166.330 ;
        RECT 96.445 166.470 96.735 166.515 ;
        RECT 99.190 166.470 99.510 166.530 ;
        RECT 96.445 166.330 99.510 166.470 ;
        RECT 96.445 166.285 96.735 166.330 ;
        RECT 99.190 166.270 99.510 166.330 ;
        RECT 102.885 166.470 103.175 166.515 ;
        RECT 105.630 166.470 105.950 166.530 ;
        RECT 106.640 166.470 106.780 166.950 ;
        RECT 108.020 166.810 108.160 166.950 ;
        RECT 108.020 166.670 110.000 166.810 ;
        RECT 102.885 166.330 106.780 166.470 ;
        RECT 102.885 166.285 103.175 166.330 ;
        RECT 105.630 166.270 105.950 166.330 ;
        RECT 109.310 166.270 109.630 166.530 ;
        RECT 109.860 166.470 110.000 166.670 ;
        RECT 119.430 166.610 119.750 166.870 ;
        RECT 117.590 166.470 117.910 166.530 ;
        RECT 109.860 166.330 117.910 166.470 ;
        RECT 119.520 166.470 119.660 166.610 ;
        RECT 119.905 166.470 120.195 166.515 ;
        RECT 119.520 166.330 120.195 166.470 ;
        RECT 121.360 166.470 121.500 167.010 ;
        RECT 122.650 166.950 122.970 167.210 ;
        RECT 123.660 166.810 123.800 167.305 ;
        RECT 124.030 167.290 124.350 167.350 ;
        RECT 124.965 167.305 125.255 167.350 ;
        RECT 126.345 167.305 126.635 167.350 ;
        RECT 126.805 167.490 127.095 167.535 ;
        RECT 127.250 167.490 127.570 167.550 ;
        RECT 126.805 167.350 127.570 167.490 ;
        RECT 126.805 167.305 127.095 167.350 ;
        RECT 127.250 167.290 127.570 167.350 ;
        RECT 127.710 167.490 128.030 167.550 ;
        RECT 128.185 167.490 128.475 167.535 ;
        RECT 127.710 167.350 128.475 167.490 ;
        RECT 127.710 167.290 128.030 167.350 ;
        RECT 128.185 167.305 128.475 167.350 ;
        RECT 129.090 167.290 129.410 167.550 ;
        RECT 131.865 167.490 132.155 167.535 ;
        RECT 132.310 167.490 132.630 167.550 ;
        RECT 141.140 167.535 141.280 167.690 ;
        RECT 131.865 167.350 132.630 167.490 ;
        RECT 131.865 167.305 132.155 167.350 ;
        RECT 132.310 167.290 132.630 167.350 ;
        RECT 141.065 167.305 141.355 167.535 ;
        RECT 142.430 167.290 142.750 167.550 ;
        RECT 142.890 167.290 143.210 167.550 ;
        RECT 144.360 167.535 144.500 167.690 ;
        RECT 144.285 167.305 144.575 167.535 ;
        RECT 124.490 166.950 124.810 167.210 ;
        RECT 127.800 166.810 127.940 167.290 ;
        RECT 132.745 167.150 133.035 167.195 ;
        RECT 133.935 167.150 134.225 167.195 ;
        RECT 136.455 167.150 136.745 167.195 ;
        RECT 132.745 167.010 136.745 167.150 ;
        RECT 132.745 166.965 133.035 167.010 ;
        RECT 133.935 166.965 134.225 167.010 ;
        RECT 136.455 166.965 136.745 167.010 ;
        RECT 140.605 167.150 140.895 167.195 ;
        RECT 142.520 167.150 142.660 167.290 ;
        RECT 140.605 167.010 142.660 167.150 ;
        RECT 140.605 166.965 140.895 167.010 ;
        RECT 123.660 166.670 127.940 166.810 ;
        RECT 132.350 166.810 132.640 166.855 ;
        RECT 134.450 166.810 134.740 166.855 ;
        RECT 136.020 166.810 136.310 166.855 ;
        RECT 132.350 166.670 136.310 166.810 ;
        RECT 132.350 166.625 132.640 166.670 ;
        RECT 134.450 166.625 134.740 166.670 ;
        RECT 136.020 166.625 136.310 166.670 ;
        RECT 140.130 166.810 140.450 166.870 ;
        RECT 141.970 166.810 142.290 166.870 ;
        RECT 145.205 166.810 145.495 166.855 ;
        RECT 140.130 166.670 145.495 166.810 ;
        RECT 140.130 166.610 140.450 166.670 ;
        RECT 141.970 166.610 142.290 166.670 ;
        RECT 145.205 166.625 145.495 166.670 ;
        RECT 128.630 166.470 128.950 166.530 ;
        RECT 121.360 166.330 128.950 166.470 ;
        RECT 117.590 166.270 117.910 166.330 ;
        RECT 119.905 166.285 120.195 166.330 ;
        RECT 128.630 166.270 128.950 166.330 ;
        RECT 142.905 166.470 143.195 166.515 ;
        RECT 143.810 166.470 144.130 166.530 ;
        RECT 142.905 166.330 144.130 166.470 ;
        RECT 142.905 166.285 143.195 166.330 ;
        RECT 143.810 166.270 144.130 166.330 ;
        RECT 36.100 165.650 150.180 166.130 ;
        RECT 42.150 165.250 42.470 165.510 ;
        RECT 60.105 165.450 60.395 165.495 ;
        RECT 62.850 165.450 63.170 165.510 ;
        RECT 60.105 165.310 63.170 165.450 ;
        RECT 60.105 165.265 60.395 165.310 ;
        RECT 62.850 165.250 63.170 165.310 ;
        RECT 66.315 165.450 66.605 165.495 ;
        RECT 67.910 165.450 68.230 165.510 ;
        RECT 72.970 165.450 73.290 165.510 ;
        RECT 66.315 165.310 73.290 165.450 ;
        RECT 66.315 165.265 66.605 165.310 ;
        RECT 67.910 165.250 68.230 165.310 ;
        RECT 72.970 165.250 73.290 165.310 ;
        RECT 74.810 165.250 75.130 165.510 ;
        RECT 76.190 165.450 76.510 165.510 ;
        RECT 79.870 165.450 80.190 165.510 ;
        RECT 88.610 165.450 88.930 165.510 ;
        RECT 76.190 165.310 80.190 165.450 ;
        RECT 76.190 165.250 76.510 165.310 ;
        RECT 79.870 165.250 80.190 165.310 ;
        RECT 88.240 165.310 88.930 165.450 ;
        RECT 42.240 164.770 42.380 165.250 ;
        RECT 44.005 165.110 44.295 165.155 ;
        RECT 47.210 165.110 47.530 165.170 ;
        RECT 74.900 165.110 75.040 165.250 ;
        RECT 44.005 164.970 47.530 165.110 ;
        RECT 44.005 164.925 44.295 164.970 ;
        RECT 47.210 164.910 47.530 164.970 ;
        RECT 59.260 164.970 75.040 165.110 ;
        RECT 88.240 165.110 88.380 165.310 ;
        RECT 88.610 165.250 88.930 165.310 ;
        RECT 89.070 165.450 89.390 165.510 ;
        RECT 91.830 165.450 92.150 165.510 ;
        RECT 89.070 165.310 92.150 165.450 ;
        RECT 89.070 165.250 89.390 165.310 ;
        RECT 91.830 165.250 92.150 165.310 ;
        RECT 92.290 165.450 92.610 165.510 ;
        RECT 95.065 165.450 95.355 165.495 ;
        RECT 92.290 165.310 95.355 165.450 ;
        RECT 92.290 165.250 92.610 165.310 ;
        RECT 95.065 165.265 95.355 165.310 ;
        RECT 101.950 165.450 102.270 165.510 ;
        RECT 107.470 165.450 107.790 165.510 ;
        RECT 101.950 165.310 107.790 165.450 ;
        RECT 101.950 165.250 102.270 165.310 ;
        RECT 107.470 165.250 107.790 165.310 ;
        RECT 111.150 165.450 111.470 165.510 ;
        RECT 112.070 165.450 112.390 165.510 ;
        RECT 111.150 165.310 112.390 165.450 ;
        RECT 111.150 165.250 111.470 165.310 ;
        RECT 112.070 165.250 112.390 165.310 ;
        RECT 114.370 165.450 114.690 165.510 ;
        RECT 121.270 165.450 121.590 165.510 ;
        RECT 114.370 165.310 121.590 165.450 ;
        RECT 114.370 165.250 114.690 165.310 ;
        RECT 121.270 165.250 121.590 165.310 ;
        RECT 125.885 165.450 126.175 165.495 ;
        RECT 129.090 165.450 129.410 165.510 ;
        RECT 125.885 165.310 129.410 165.450 ;
        RECT 125.885 165.265 126.175 165.310 ;
        RECT 129.090 165.250 129.410 165.310 ;
        RECT 137.830 165.450 138.150 165.510 ;
        RECT 138.765 165.450 139.055 165.495 ;
        RECT 137.830 165.310 139.055 165.450 ;
        RECT 137.830 165.250 138.150 165.310 ;
        RECT 138.765 165.265 139.055 165.310 ;
        RECT 140.605 165.450 140.895 165.495 ;
        RECT 141.050 165.450 141.370 165.510 ;
        RECT 140.605 165.310 141.370 165.450 ;
        RECT 140.605 165.265 140.895 165.310 ;
        RECT 141.050 165.250 141.370 165.310 ;
        RECT 141.510 165.450 141.830 165.510 ;
        RECT 143.365 165.450 143.655 165.495 ;
        RECT 141.510 165.310 143.655 165.450 ;
        RECT 141.510 165.250 141.830 165.310 ;
        RECT 143.365 165.265 143.655 165.310 ;
        RECT 89.990 165.110 90.310 165.170 ;
        RECT 92.750 165.110 93.070 165.170 ;
        RECT 88.240 164.970 90.310 165.110 ;
        RECT 43.085 164.770 43.375 164.815 ;
        RECT 42.240 164.630 43.375 164.770 ;
        RECT 43.085 164.585 43.375 164.630 ;
        RECT 44.910 164.770 45.230 164.830 ;
        RECT 57.345 164.770 57.635 164.815 ;
        RECT 58.710 164.770 59.030 164.830 ;
        RECT 44.910 164.630 46.060 164.770 ;
        RECT 44.910 164.570 45.230 164.630 ;
        RECT 44.450 164.430 44.770 164.490 ;
        RECT 45.920 164.475 46.060 164.630 ;
        RECT 57.345 164.630 59.030 164.770 ;
        RECT 57.345 164.585 57.635 164.630 ;
        RECT 58.710 164.570 59.030 164.630 ;
        RECT 59.260 164.475 59.400 164.970 ;
        RECT 61.470 164.770 61.790 164.830 ;
        RECT 61.945 164.770 62.235 164.815 ;
        RECT 61.470 164.630 62.235 164.770 ;
        RECT 61.470 164.570 61.790 164.630 ;
        RECT 61.945 164.585 62.235 164.630 ;
        RECT 65.165 164.770 65.455 164.815 ;
        RECT 66.530 164.770 66.850 164.830 ;
        RECT 65.165 164.630 66.850 164.770 ;
        RECT 65.165 164.585 65.455 164.630 ;
        RECT 44.450 164.290 45.600 164.430 ;
        RECT 44.450 164.230 44.770 164.290 ;
        RECT 45.460 164.090 45.600 164.290 ;
        RECT 45.845 164.245 46.135 164.475 ;
        RECT 55.965 164.245 56.255 164.475 ;
        RECT 59.185 164.245 59.475 164.475 ;
        RECT 56.040 164.090 56.180 164.245 ;
        RECT 60.550 164.230 60.870 164.490 ;
        RECT 62.020 164.430 62.160 164.585 ;
        RECT 66.530 164.570 66.850 164.630 ;
        RECT 71.590 164.770 71.910 164.830 ;
        RECT 71.590 164.630 75.500 164.770 ;
        RECT 71.590 164.570 71.910 164.630 ;
        RECT 75.360 164.475 75.500 164.630 ;
        RECT 71.145 164.430 71.435 164.475 ;
        RECT 62.020 164.290 67.680 164.430 ;
        RECT 45.460 163.950 64.000 164.090 ;
        RECT 63.860 163.810 64.000 163.950 ;
        RECT 67.540 163.810 67.680 164.290 ;
        RECT 71.145 164.290 75.040 164.430 ;
        RECT 71.145 164.245 71.435 164.290 ;
        RECT 43.070 163.550 43.390 163.810 ;
        RECT 44.910 163.550 45.230 163.810 ;
        RECT 50.890 163.750 51.210 163.810 ;
        RECT 62.390 163.750 62.710 163.810 ;
        RECT 50.890 163.610 62.710 163.750 ;
        RECT 50.890 163.550 51.210 163.610 ;
        RECT 62.390 163.550 62.710 163.610 ;
        RECT 63.770 163.550 64.090 163.810 ;
        RECT 67.450 163.550 67.770 163.810 ;
        RECT 72.970 163.550 73.290 163.810 ;
        RECT 74.900 163.750 75.040 164.290 ;
        RECT 75.285 164.245 75.575 164.475 ;
        RECT 76.650 164.230 76.970 164.490 ;
        RECT 79.410 164.230 79.730 164.490 ;
        RECT 80.330 164.430 80.650 164.490 ;
        RECT 88.240 164.475 88.380 164.970 ;
        RECT 89.990 164.910 90.310 164.970 ;
        RECT 91.000 164.970 119.660 165.110 ;
        RECT 88.625 164.770 88.915 164.815 ;
        RECT 91.000 164.770 91.140 164.970 ;
        RECT 92.750 164.910 93.070 164.970 ;
        RECT 119.520 164.830 119.660 164.970 ;
        RECT 123.660 164.970 126.100 165.110 ;
        RECT 88.625 164.630 91.140 164.770 ;
        RECT 88.625 164.585 88.915 164.630 ;
        RECT 84.945 164.430 85.235 164.475 ;
        RECT 80.330 164.290 85.235 164.430 ;
        RECT 80.330 164.230 80.650 164.290 ;
        RECT 84.945 164.245 85.235 164.290 ;
        RECT 86.785 164.430 87.075 164.475 ;
        RECT 87.245 164.430 87.535 164.475 ;
        RECT 86.785 164.290 87.535 164.430 ;
        RECT 86.785 164.245 87.075 164.290 ;
        RECT 87.245 164.245 87.535 164.290 ;
        RECT 88.165 164.245 88.455 164.475 ;
        RECT 89.070 164.230 89.390 164.490 ;
        RECT 90.005 164.430 90.295 164.475 ;
        RECT 90.450 164.430 90.770 164.490 ;
        RECT 90.005 164.290 90.770 164.430 ;
        RECT 91.000 164.430 91.140 164.630 ;
        RECT 91.830 164.570 92.150 164.830 ;
        RECT 110.230 164.770 110.550 164.830 ;
        RECT 96.060 164.630 107.240 164.770 ;
        RECT 96.060 164.490 96.200 164.630 ;
        RECT 92.305 164.430 92.595 164.475 ;
        RECT 91.000 164.290 92.595 164.430 ;
        RECT 90.005 164.245 90.295 164.290 ;
        RECT 90.450 164.230 90.770 164.290 ;
        RECT 92.305 164.245 92.595 164.290 ;
        RECT 92.765 164.245 93.055 164.475 ;
        RECT 75.745 164.090 76.035 164.135 ;
        RECT 79.500 164.090 79.640 164.230 ;
        RECT 75.745 163.950 79.640 164.090 ;
        RECT 83.090 164.090 83.410 164.150 ;
        RECT 85.865 164.090 86.155 164.135 ;
        RECT 91.370 164.090 91.690 164.150 ;
        RECT 92.840 164.090 92.980 164.245 ;
        RECT 93.210 164.230 93.530 164.490 ;
        RECT 94.130 164.230 94.450 164.490 ;
        RECT 95.510 164.230 95.830 164.490 ;
        RECT 95.970 164.230 96.290 164.490 ;
        RECT 96.430 164.230 96.750 164.490 ;
        RECT 96.980 164.475 97.120 164.630 ;
        RECT 96.905 164.245 97.195 164.475 ;
        RECT 97.350 164.230 97.670 164.490 ;
        RECT 98.285 164.245 98.575 164.475 ;
        RECT 101.045 164.245 101.335 164.475 ;
        RECT 101.490 164.430 101.810 164.490 ;
        RECT 102.410 164.430 102.730 164.490 ;
        RECT 101.490 164.290 102.730 164.430 ;
        RECT 83.090 163.950 91.690 164.090 ;
        RECT 75.745 163.905 76.035 163.950 ;
        RECT 83.090 163.890 83.410 163.950 ;
        RECT 85.865 163.905 86.155 163.950 ;
        RECT 91.370 163.890 91.690 163.950 ;
        RECT 91.920 163.950 92.980 164.090 ;
        RECT 94.220 164.090 94.360 164.230 ;
        RECT 95.600 164.090 95.740 164.230 ;
        RECT 98.360 164.090 98.500 164.245 ;
        RECT 94.220 163.950 95.280 164.090 ;
        RECT 95.600 163.950 98.500 164.090 ;
        RECT 101.120 164.090 101.260 164.245 ;
        RECT 101.490 164.230 101.810 164.290 ;
        RECT 102.410 164.230 102.730 164.290 ;
        RECT 104.250 164.230 104.570 164.490 ;
        RECT 104.340 164.090 104.480 164.230 ;
        RECT 106.090 164.090 106.410 164.150 ;
        RECT 101.120 163.950 106.410 164.090 ;
        RECT 91.920 163.810 92.060 163.950 ;
        RECT 76.190 163.750 76.510 163.810 ;
        RECT 74.900 163.610 76.510 163.750 ;
        RECT 76.190 163.550 76.510 163.610 ;
        RECT 77.585 163.750 77.875 163.795 ;
        RECT 78.490 163.750 78.810 163.810 ;
        RECT 77.585 163.610 78.810 163.750 ;
        RECT 77.585 163.565 77.875 163.610 ;
        RECT 78.490 163.550 78.810 163.610 ;
        RECT 90.910 163.550 91.230 163.810 ;
        RECT 91.830 163.550 92.150 163.810 ;
        RECT 94.130 163.550 94.450 163.810 ;
        RECT 95.140 163.750 95.280 163.950 ;
        RECT 106.090 163.890 106.410 163.950 ;
        RECT 99.190 163.750 99.510 163.810 ;
        RECT 107.100 163.795 107.240 164.630 ;
        RECT 108.020 164.630 110.550 164.770 ;
        RECT 108.020 164.475 108.160 164.630 ;
        RECT 110.230 164.570 110.550 164.630 ;
        RECT 110.690 164.770 111.010 164.830 ;
        RECT 112.545 164.770 112.835 164.815 ;
        RECT 110.690 164.630 112.835 164.770 ;
        RECT 110.690 164.570 111.010 164.630 ;
        RECT 112.545 164.585 112.835 164.630 ;
        RECT 112.990 164.570 113.310 164.830 ;
        RECT 113.450 164.770 113.770 164.830 ;
        RECT 114.370 164.770 114.690 164.830 ;
        RECT 113.450 164.630 114.690 164.770 ;
        RECT 113.450 164.570 113.770 164.630 ;
        RECT 114.370 164.570 114.690 164.630 ;
        RECT 119.430 164.570 119.750 164.830 ;
        RECT 107.945 164.245 108.235 164.475 ;
        RECT 109.310 164.230 109.630 164.490 ;
        RECT 109.785 164.245 110.075 164.475 ;
        RECT 111.165 164.430 111.455 164.475 ;
        RECT 111.610 164.430 111.930 164.490 ;
        RECT 111.165 164.290 111.930 164.430 ;
        RECT 111.165 164.245 111.455 164.290 ;
        RECT 107.470 164.090 107.790 164.150 ;
        RECT 109.860 164.090 110.000 164.245 ;
        RECT 111.610 164.230 111.930 164.290 ;
        RECT 118.510 164.430 118.830 164.490 ;
        RECT 121.745 164.430 122.035 164.475 ;
        RECT 123.660 164.430 123.800 164.970 ;
        RECT 124.045 164.770 124.335 164.815 ;
        RECT 125.960 164.770 126.100 164.970 ;
        RECT 127.710 164.910 128.030 165.170 ;
        RECT 135.070 165.110 135.390 165.170 ;
        RECT 141.600 165.110 141.740 165.250 ;
        RECT 135.070 164.970 141.740 165.110 ;
        RECT 135.070 164.910 135.390 164.970 ;
        RECT 141.065 164.770 141.355 164.815 ;
        RECT 124.045 164.630 125.640 164.770 ;
        RECT 125.960 164.630 141.355 164.770 ;
        RECT 124.045 164.585 124.335 164.630 ;
        RECT 125.500 164.490 125.640 164.630 ;
        RECT 141.065 164.585 141.355 164.630 ;
        RECT 143.810 164.570 144.130 164.830 ;
        RECT 124.490 164.430 124.810 164.490 ;
        RECT 118.510 164.290 124.810 164.430 ;
        RECT 118.510 164.230 118.830 164.290 ;
        RECT 121.745 164.245 122.035 164.290 ;
        RECT 124.490 164.230 124.810 164.290 ;
        RECT 124.965 164.245 125.255 164.475 ;
        RECT 125.410 164.430 125.730 164.490 ;
        RECT 126.805 164.430 127.095 164.475 ;
        RECT 125.410 164.290 127.095 164.430 ;
        RECT 125.040 164.090 125.180 164.245 ;
        RECT 125.410 164.230 125.730 164.290 ;
        RECT 126.805 164.245 127.095 164.290 ;
        RECT 127.725 164.430 128.015 164.475 ;
        RECT 135.070 164.430 135.390 164.490 ;
        RECT 127.725 164.290 135.390 164.430 ;
        RECT 127.725 164.245 128.015 164.290 ;
        RECT 127.800 164.090 127.940 164.245 ;
        RECT 135.070 164.230 135.390 164.290 ;
        RECT 140.130 164.230 140.450 164.490 ;
        RECT 140.590 164.230 140.910 164.490 ;
        RECT 141.985 164.430 142.275 164.475 ;
        RECT 142.430 164.430 142.750 164.490 ;
        RECT 141.985 164.290 142.750 164.430 ;
        RECT 141.985 164.245 142.275 164.290 ;
        RECT 142.430 164.230 142.750 164.290 ;
        RECT 142.890 164.230 143.210 164.490 ;
        RECT 143.900 164.425 144.040 164.570 ;
        RECT 143.825 164.195 144.115 164.425 ;
        RECT 107.470 163.950 123.340 164.090 ;
        RECT 125.040 163.950 127.940 164.090 ;
        RECT 133.230 164.090 133.550 164.150 ;
        RECT 138.750 164.090 139.070 164.150 ;
        RECT 133.230 163.950 139.070 164.090 ;
        RECT 107.470 163.890 107.790 163.950 ;
        RECT 95.140 163.610 99.510 163.750 ;
        RECT 99.190 163.550 99.510 163.610 ;
        RECT 107.025 163.750 107.315 163.795 ;
        RECT 107.930 163.750 108.250 163.810 ;
        RECT 107.025 163.610 108.250 163.750 ;
        RECT 107.025 163.565 107.315 163.610 ;
        RECT 107.930 163.550 108.250 163.610 ;
        RECT 108.405 163.750 108.695 163.795 ;
        RECT 109.310 163.750 109.630 163.810 ;
        RECT 108.405 163.610 109.630 163.750 ;
        RECT 108.405 163.565 108.695 163.610 ;
        RECT 109.310 163.550 109.630 163.610 ;
        RECT 111.610 163.550 111.930 163.810 ;
        RECT 114.845 163.750 115.135 163.795 ;
        RECT 117.590 163.750 117.910 163.810 ;
        RECT 114.845 163.610 117.910 163.750 ;
        RECT 114.845 163.565 115.135 163.610 ;
        RECT 117.590 163.550 117.910 163.610 ;
        RECT 122.650 163.550 122.970 163.810 ;
        RECT 123.200 163.750 123.340 163.950 ;
        RECT 133.230 163.890 133.550 163.950 ;
        RECT 138.750 163.890 139.070 163.950 ;
        RECT 141.050 163.750 141.370 163.810 ;
        RECT 123.200 163.610 141.370 163.750 ;
        RECT 141.050 163.550 141.370 163.610 ;
        RECT 36.100 162.930 150.180 163.410 ;
        RECT 44.910 162.530 45.230 162.790 ;
        RECT 46.750 162.530 47.070 162.790 ;
        RECT 50.445 162.730 50.735 162.775 ;
        RECT 54.110 162.730 54.430 162.790 ;
        RECT 60.550 162.730 60.870 162.790 ;
        RECT 50.445 162.590 60.870 162.730 ;
        RECT 50.445 162.545 50.735 162.590 ;
        RECT 54.110 162.530 54.430 162.590 ;
        RECT 60.550 162.530 60.870 162.590 ;
        RECT 61.025 162.730 61.315 162.775 ;
        RECT 66.530 162.730 66.850 162.790 ;
        RECT 61.025 162.590 66.850 162.730 ;
        RECT 61.025 162.545 61.315 162.590 ;
        RECT 66.530 162.530 66.850 162.590 ;
        RECT 72.065 162.730 72.355 162.775 ;
        RECT 76.650 162.730 76.970 162.790 ;
        RECT 72.065 162.590 76.970 162.730 ;
        RECT 72.065 162.545 72.355 162.590 ;
        RECT 76.650 162.530 76.970 162.590 ;
        RECT 80.330 162.730 80.650 162.790 ;
        RECT 92.765 162.730 93.055 162.775 ;
        RECT 95.050 162.730 95.370 162.790 ;
        RECT 80.330 162.590 91.140 162.730 ;
        RECT 80.330 162.530 80.650 162.590 ;
        RECT 41.200 162.390 41.490 162.435 ;
        RECT 45.000 162.390 45.140 162.530 ;
        RECT 41.200 162.250 45.140 162.390 ;
        RECT 51.810 162.390 52.130 162.450 ;
        RECT 63.770 162.390 64.090 162.450 ;
        RECT 91.000 162.390 91.140 162.590 ;
        RECT 92.765 162.590 95.370 162.730 ;
        RECT 92.765 162.545 93.055 162.590 ;
        RECT 95.050 162.530 95.370 162.590 ;
        RECT 97.350 162.730 97.670 162.790 ;
        RECT 101.045 162.730 101.335 162.775 ;
        RECT 97.350 162.590 101.335 162.730 ;
        RECT 97.350 162.530 97.670 162.590 ;
        RECT 101.045 162.545 101.335 162.590 ;
        RECT 107.010 162.530 107.330 162.790 ;
        RECT 117.590 162.530 117.910 162.790 ;
        RECT 125.885 162.730 126.175 162.775 ;
        RECT 137.370 162.730 137.690 162.790 ;
        RECT 125.885 162.590 137.690 162.730 ;
        RECT 125.885 162.545 126.175 162.590 ;
        RECT 137.370 162.530 137.690 162.590 ;
        RECT 138.765 162.730 139.055 162.775 ;
        RECT 139.210 162.730 139.530 162.790 ;
        RECT 138.765 162.590 139.530 162.730 ;
        RECT 138.765 162.545 139.055 162.590 ;
        RECT 139.210 162.530 139.530 162.590 ;
        RECT 142.890 162.730 143.210 162.790 ;
        RECT 144.730 162.730 145.050 162.790 ;
        RECT 146.585 162.730 146.875 162.775 ;
        RECT 142.890 162.590 146.875 162.730 ;
        RECT 142.890 162.530 143.210 162.590 ;
        RECT 144.730 162.530 145.050 162.590 ;
        RECT 146.585 162.545 146.875 162.590 ;
        RECT 102.870 162.390 103.190 162.450 ;
        RECT 51.810 162.250 63.540 162.390 ;
        RECT 41.200 162.205 41.490 162.250 ;
        RECT 51.810 162.190 52.130 162.250 ;
        RECT 37.550 162.050 37.870 162.110 ;
        RECT 39.865 162.050 40.155 162.095 ;
        RECT 37.550 161.910 40.155 162.050 ;
        RECT 37.550 161.850 37.870 161.910 ;
        RECT 39.865 161.865 40.155 161.910 ;
        RECT 51.350 161.850 51.670 162.110 ;
        RECT 55.030 162.050 55.350 162.110 ;
        RECT 57.345 162.050 57.635 162.095 ;
        RECT 55.030 161.910 57.635 162.050 ;
        RECT 55.030 161.850 55.350 161.910 ;
        RECT 57.345 161.865 57.635 161.910 ;
        RECT 60.105 161.865 60.395 162.095 ;
        RECT 62.405 161.865 62.695 162.095 ;
        RECT 40.745 161.710 41.035 161.755 ;
        RECT 41.935 161.710 42.225 161.755 ;
        RECT 44.455 161.710 44.745 161.755 ;
        RECT 40.745 161.570 44.745 161.710 ;
        RECT 40.745 161.525 41.035 161.570 ;
        RECT 41.935 161.525 42.225 161.570 ;
        RECT 44.455 161.525 44.745 161.570 ;
        RECT 51.825 161.710 52.115 161.755 ;
        RECT 52.270 161.710 52.590 161.770 ;
        RECT 51.825 161.570 52.590 161.710 ;
        RECT 51.825 161.525 52.115 161.570 ;
        RECT 52.270 161.510 52.590 161.570 ;
        RECT 53.205 161.525 53.495 161.755 ;
        RECT 54.110 161.710 54.430 161.770 ;
        RECT 56.425 161.710 56.715 161.755 ;
        RECT 60.180 161.710 60.320 161.865 ;
        RECT 54.110 161.570 60.320 161.710 ;
        RECT 40.350 161.370 40.640 161.415 ;
        RECT 42.450 161.370 42.740 161.415 ;
        RECT 44.020 161.370 44.310 161.415 ;
        RECT 40.350 161.230 44.310 161.370 ;
        RECT 53.280 161.370 53.420 161.525 ;
        RECT 54.110 161.510 54.430 161.570 ;
        RECT 56.425 161.525 56.715 161.570 ;
        RECT 62.480 161.370 62.620 161.865 ;
        RECT 62.850 161.510 63.170 161.770 ;
        RECT 63.400 161.710 63.540 162.250 ;
        RECT 63.770 162.250 88.840 162.390 ;
        RECT 91.000 162.250 103.190 162.390 ;
        RECT 63.770 162.190 64.090 162.250 ;
        RECT 67.925 162.050 68.215 162.095 ;
        RECT 69.290 162.060 69.610 162.110 ;
        RECT 70.225 162.060 70.515 162.095 ;
        RECT 69.290 162.050 70.515 162.060 ;
        RECT 67.925 161.920 70.515 162.050 ;
        RECT 67.925 161.910 69.610 161.920 ;
        RECT 67.925 161.865 68.215 161.910 ;
        RECT 69.290 161.850 69.610 161.910 ;
        RECT 70.225 161.865 70.515 161.920 ;
        RECT 70.670 162.050 70.990 162.110 ;
        RECT 71.145 162.050 71.435 162.095 ;
        RECT 70.670 161.910 71.435 162.050 ;
        RECT 70.670 161.850 70.990 161.910 ;
        RECT 71.145 161.865 71.435 161.910 ;
        RECT 86.325 162.060 86.615 162.095 ;
        RECT 86.325 162.050 87.000 162.060 ;
        RECT 87.230 162.050 87.550 162.110 ;
        RECT 86.325 161.920 87.550 162.050 ;
        RECT 86.325 161.865 86.615 161.920 ;
        RECT 86.860 161.910 87.550 161.920 ;
        RECT 88.700 162.050 88.840 162.250 ;
        RECT 91.830 162.050 92.150 162.110 ;
        RECT 88.700 161.910 92.150 162.050 ;
        RECT 87.230 161.850 87.550 161.910 ;
        RECT 91.830 161.850 92.150 161.910 ;
        RECT 92.750 161.850 93.070 162.110 ;
        RECT 98.730 161.850 99.050 162.110 ;
        RECT 102.040 162.095 102.180 162.250 ;
        RECT 102.870 162.190 103.190 162.250 ;
        RECT 103.330 162.190 103.650 162.450 ;
        RECT 107.100 162.390 107.240 162.530 ;
        RECT 112.990 162.390 113.310 162.450 ;
        RECT 114.370 162.390 114.690 162.450 ;
        RECT 123.585 162.390 123.875 162.435 ;
        RECT 124.490 162.390 124.810 162.450 ;
        RECT 132.310 162.390 132.630 162.450 ;
        RECT 135.530 162.390 135.850 162.450 ;
        RECT 107.100 162.250 114.140 162.390 ;
        RECT 101.965 161.865 102.255 162.095 ;
        RECT 102.410 161.850 102.730 162.110 ;
        RECT 103.420 162.050 103.560 162.190 ;
        RECT 103.805 162.050 104.095 162.095 ;
        RECT 103.420 161.910 104.095 162.050 ;
        RECT 103.805 161.865 104.095 161.910 ;
        RECT 104.250 162.050 104.570 162.110 ;
        RECT 105.185 162.050 105.475 162.095 ;
        RECT 108.850 162.050 109.170 162.110 ;
        RECT 109.400 162.095 109.540 162.250 ;
        RECT 112.990 162.190 113.310 162.250 ;
        RECT 104.250 161.910 109.170 162.050 ;
        RECT 104.250 161.850 104.570 161.910 ;
        RECT 105.185 161.865 105.475 161.910 ;
        RECT 108.850 161.850 109.170 161.910 ;
        RECT 109.325 161.865 109.615 162.095 ;
        RECT 110.230 161.850 110.550 162.110 ;
        RECT 111.150 161.850 111.470 162.110 ;
        RECT 112.070 161.850 112.390 162.110 ;
        RECT 114.000 162.095 114.140 162.250 ;
        RECT 114.370 162.250 115.980 162.390 ;
        RECT 114.370 162.190 114.690 162.250 ;
        RECT 115.840 162.095 115.980 162.250 ;
        RECT 122.280 162.250 132.630 162.390 ;
        RECT 113.925 161.865 114.215 162.095 ;
        RECT 114.845 161.865 115.135 162.095 ;
        RECT 115.305 161.865 115.595 162.095 ;
        RECT 115.765 161.865 116.055 162.095 ;
        RECT 116.685 162.050 116.975 162.095 ;
        RECT 119.430 162.050 119.750 162.110 ;
        RECT 116.685 161.910 119.750 162.050 ;
        RECT 116.685 161.865 116.975 161.910 ;
        RECT 68.385 161.710 68.675 161.755 ;
        RECT 72.050 161.710 72.370 161.770 ;
        RECT 85.850 161.710 86.170 161.770 ;
        RECT 63.400 161.570 69.520 161.710 ;
        RECT 68.385 161.525 68.675 161.570 ;
        RECT 69.380 161.430 69.520 161.570 ;
        RECT 72.050 161.570 86.170 161.710 ;
        RECT 72.050 161.510 72.370 161.570 ;
        RECT 85.850 161.510 86.170 161.570 ;
        RECT 92.290 161.710 92.610 161.770 ;
        RECT 92.290 161.570 93.900 161.710 ;
        RECT 92.290 161.510 92.610 161.570 ;
        RECT 63.770 161.370 64.090 161.430 ;
        RECT 53.280 161.230 59.860 161.370 ;
        RECT 62.480 161.230 64.090 161.370 ;
        RECT 40.350 161.185 40.640 161.230 ;
        RECT 42.450 161.185 42.740 161.230 ;
        RECT 44.020 161.185 44.310 161.230 ;
        RECT 59.720 161.090 59.860 161.230 ;
        RECT 63.770 161.170 64.090 161.230 ;
        RECT 69.290 161.170 69.610 161.430 ;
        RECT 69.765 161.370 70.055 161.415 ;
        RECT 71.590 161.370 71.910 161.430 ;
        RECT 69.765 161.230 71.910 161.370 ;
        RECT 69.765 161.185 70.055 161.230 ;
        RECT 71.590 161.170 71.910 161.230 ;
        RECT 87.245 161.370 87.535 161.415 ;
        RECT 93.210 161.370 93.530 161.430 ;
        RECT 87.245 161.230 93.530 161.370 ;
        RECT 93.760 161.370 93.900 161.570 ;
        RECT 97.350 161.510 97.670 161.770 ;
        RECT 97.825 161.710 98.115 161.755 ;
        RECT 103.345 161.710 103.635 161.755 ;
        RECT 109.770 161.710 110.090 161.770 ;
        RECT 97.825 161.570 110.090 161.710 ;
        RECT 97.825 161.525 98.115 161.570 ;
        RECT 98.820 161.430 98.960 161.570 ;
        RECT 103.345 161.525 103.635 161.570 ;
        RECT 109.770 161.510 110.090 161.570 ;
        RECT 110.705 161.525 110.995 161.755 ;
        RECT 114.920 161.710 115.060 161.865 ;
        RECT 112.160 161.570 115.060 161.710 ;
        RECT 115.380 161.710 115.520 161.865 ;
        RECT 119.430 161.850 119.750 161.910 ;
        RECT 122.280 161.710 122.420 162.250 ;
        RECT 123.585 162.205 123.875 162.250 ;
        RECT 124.490 162.190 124.810 162.250 ;
        RECT 122.650 162.050 122.970 162.110 ;
        RECT 131.020 162.095 131.160 162.250 ;
        RECT 132.310 162.190 132.630 162.250 ;
        RECT 132.860 162.250 135.850 162.390 ;
        RECT 124.965 162.050 125.255 162.095 ;
        RECT 122.650 161.910 125.255 162.050 ;
        RECT 122.650 161.850 122.970 161.910 ;
        RECT 124.965 161.865 125.255 161.910 ;
        RECT 128.645 161.865 128.935 162.095 ;
        RECT 130.945 161.865 131.235 162.095 ;
        RECT 131.405 162.050 131.695 162.095 ;
        RECT 132.860 162.050 133.000 162.250 ;
        RECT 135.530 162.190 135.850 162.250 ;
        RECT 136.465 162.390 136.755 162.435 ;
        RECT 141.510 162.390 141.830 162.450 ;
        RECT 136.465 162.250 141.830 162.390 ;
        RECT 136.465 162.205 136.755 162.250 ;
        RECT 141.510 162.190 141.830 162.250 ;
        RECT 131.405 161.910 133.000 162.050 ;
        RECT 131.405 161.865 131.695 161.910 ;
        RECT 115.380 161.570 122.420 161.710 ;
        RECT 93.760 161.230 98.040 161.370 ;
        RECT 87.245 161.185 87.535 161.230 ;
        RECT 93.210 161.170 93.530 161.230 ;
        RECT 97.900 161.090 98.040 161.230 ;
        RECT 98.730 161.170 99.050 161.430 ;
        RECT 107.470 161.370 107.790 161.430 ;
        RECT 110.780 161.370 110.920 161.525 ;
        RECT 107.470 161.230 110.920 161.370 ;
        RECT 107.470 161.170 107.790 161.230 ;
        RECT 58.265 161.030 58.555 161.075 ;
        RECT 59.170 161.030 59.490 161.090 ;
        RECT 58.265 160.890 59.490 161.030 ;
        RECT 58.265 160.845 58.555 160.890 ;
        RECT 59.170 160.830 59.490 160.890 ;
        RECT 59.630 161.030 59.950 161.090 ;
        RECT 95.050 161.030 95.370 161.090 ;
        RECT 59.630 160.890 95.370 161.030 ;
        RECT 59.630 160.830 59.950 160.890 ;
        RECT 95.050 160.830 95.370 160.890 ;
        RECT 97.810 160.830 98.130 161.090 ;
        RECT 99.650 160.830 99.970 161.090 ;
        RECT 104.250 160.830 104.570 161.090 ;
        RECT 106.090 161.030 106.410 161.090 ;
        RECT 112.160 161.030 112.300 161.570 ;
        RECT 124.505 161.525 124.795 161.755 ;
        RECT 126.790 161.710 127.110 161.770 ;
        RECT 128.720 161.710 128.860 161.865 ;
        RECT 133.230 161.850 133.550 162.110 ;
        RECT 137.845 162.050 138.135 162.095 ;
        RECT 138.290 162.050 138.610 162.110 ;
        RECT 137.845 161.910 138.610 162.050 ;
        RECT 137.845 161.865 138.135 161.910 ;
        RECT 138.290 161.850 138.610 161.910 ;
        RECT 139.670 161.850 139.990 162.110 ;
        RECT 140.965 162.050 141.255 162.095 ;
        RECT 140.220 161.910 141.255 162.050 ;
        RECT 126.790 161.570 128.860 161.710 ;
        RECT 132.325 161.710 132.615 161.755 ;
        RECT 133.320 161.710 133.460 161.850 ;
        RECT 132.325 161.570 133.460 161.710 ;
        RECT 137.385 161.710 137.675 161.755 ;
        RECT 138.750 161.710 139.070 161.770 ;
        RECT 140.220 161.710 140.360 161.910 ;
        RECT 140.965 161.865 141.255 161.910 ;
        RECT 137.385 161.570 139.070 161.710 ;
        RECT 115.290 161.370 115.610 161.430 ;
        RECT 124.580 161.370 124.720 161.525 ;
        RECT 126.790 161.510 127.110 161.570 ;
        RECT 132.325 161.525 132.615 161.570 ;
        RECT 137.385 161.525 137.675 161.570 ;
        RECT 138.750 161.510 139.070 161.570 ;
        RECT 139.300 161.570 140.360 161.710 ;
        RECT 140.565 161.710 140.855 161.755 ;
        RECT 141.755 161.710 142.045 161.755 ;
        RECT 144.275 161.710 144.565 161.755 ;
        RECT 140.565 161.570 144.565 161.710 ;
        RECT 131.390 161.370 131.710 161.430 ;
        RECT 115.290 161.230 131.710 161.370 ;
        RECT 115.290 161.170 115.610 161.230 ;
        RECT 131.390 161.170 131.710 161.230 ;
        RECT 134.150 161.370 134.470 161.430 ;
        RECT 134.625 161.370 134.915 161.415 ;
        RECT 138.290 161.370 138.610 161.430 ;
        RECT 134.150 161.230 138.610 161.370 ;
        RECT 134.150 161.170 134.470 161.230 ;
        RECT 134.625 161.185 134.915 161.230 ;
        RECT 138.290 161.170 138.610 161.230 ;
        RECT 106.090 160.890 112.300 161.030 ;
        RECT 113.005 161.030 113.295 161.075 ;
        RECT 114.370 161.030 114.690 161.090 ;
        RECT 113.005 160.890 114.690 161.030 ;
        RECT 106.090 160.830 106.410 160.890 ;
        RECT 113.005 160.845 113.295 160.890 ;
        RECT 114.370 160.830 114.690 160.890 ;
        RECT 124.965 161.030 125.255 161.075 ;
        RECT 125.410 161.030 125.730 161.090 ;
        RECT 124.965 160.890 125.730 161.030 ;
        RECT 124.965 160.845 125.255 160.890 ;
        RECT 125.410 160.830 125.730 160.890 ;
        RECT 127.710 160.830 128.030 161.090 ;
        RECT 131.865 161.030 132.155 161.075 ;
        RECT 133.230 161.030 133.550 161.090 ;
        RECT 131.865 160.890 133.550 161.030 ;
        RECT 131.865 160.845 132.155 160.890 ;
        RECT 133.230 160.830 133.550 160.890 ;
        RECT 136.910 160.830 137.230 161.090 ;
        RECT 137.370 161.030 137.690 161.090 ;
        RECT 139.300 161.030 139.440 161.570 ;
        RECT 140.565 161.525 140.855 161.570 ;
        RECT 141.755 161.525 142.045 161.570 ;
        RECT 144.275 161.525 144.565 161.570 ;
        RECT 140.170 161.370 140.460 161.415 ;
        RECT 142.270 161.370 142.560 161.415 ;
        RECT 143.840 161.370 144.130 161.415 ;
        RECT 140.170 161.230 144.130 161.370 ;
        RECT 140.170 161.185 140.460 161.230 ;
        RECT 142.270 161.185 142.560 161.230 ;
        RECT 143.840 161.185 144.130 161.230 ;
        RECT 137.370 160.890 139.440 161.030 ;
        RECT 137.370 160.830 137.690 160.890 ;
        RECT 36.100 160.210 150.180 160.690 ;
        RECT 46.765 160.010 47.055 160.055 ;
        RECT 47.210 160.010 47.530 160.070 ;
        RECT 46.765 159.870 47.530 160.010 ;
        RECT 46.765 159.825 47.055 159.870 ;
        RECT 46.840 159.330 46.980 159.825 ;
        RECT 47.210 159.810 47.530 159.870 ;
        RECT 52.270 160.010 52.590 160.070 ;
        RECT 68.370 160.010 68.690 160.070 ;
        RECT 52.270 159.870 68.690 160.010 ;
        RECT 52.270 159.810 52.590 159.870 ;
        RECT 68.370 159.810 68.690 159.870 ;
        RECT 78.505 160.010 78.795 160.055 ;
        RECT 79.425 160.010 79.715 160.055 ;
        RECT 78.505 159.870 79.715 160.010 ;
        RECT 78.505 159.825 78.795 159.870 ;
        RECT 79.425 159.825 79.715 159.870 ;
        RECT 91.370 160.010 91.690 160.070 ;
        RECT 91.370 159.870 101.260 160.010 ;
        RECT 91.370 159.810 91.690 159.870 ;
        RECT 62.850 159.670 63.170 159.730 ;
        RECT 100.570 159.670 100.890 159.730 ;
        RECT 61.100 159.530 100.890 159.670 ;
        RECT 43.620 159.190 46.980 159.330 ;
        RECT 47.210 159.330 47.530 159.390 ;
        RECT 55.030 159.330 55.350 159.390 ;
        RECT 47.210 159.190 55.350 159.330 ;
        RECT 42.165 158.990 42.455 159.035 ;
        RECT 43.070 158.990 43.390 159.050 ;
        RECT 43.620 159.035 43.760 159.190 ;
        RECT 47.210 159.130 47.530 159.190 ;
        RECT 55.030 159.130 55.350 159.190 ;
        RECT 56.425 159.330 56.715 159.375 ;
        RECT 61.100 159.330 61.240 159.530 ;
        RECT 62.850 159.470 63.170 159.530 ;
        RECT 100.570 159.470 100.890 159.530 ;
        RECT 56.425 159.190 58.480 159.330 ;
        RECT 56.425 159.145 56.715 159.190 ;
        RECT 42.165 158.850 43.390 158.990 ;
        RECT 42.165 158.805 42.455 158.850 ;
        RECT 43.070 158.790 43.390 158.850 ;
        RECT 43.545 158.805 43.835 159.035 ;
        RECT 44.450 158.790 44.770 159.050 ;
        RECT 44.910 158.790 45.230 159.050 ;
        RECT 45.845 158.990 46.135 159.035 ;
        RECT 51.350 158.990 51.670 159.050 ;
        RECT 45.845 158.850 51.670 158.990 ;
        RECT 45.845 158.805 46.135 158.850 ;
        RECT 51.350 158.790 51.670 158.850 ;
        RECT 54.110 158.990 54.430 159.050 ;
        RECT 58.340 159.035 58.480 159.190 ;
        RECT 58.800 159.190 61.240 159.330 ;
        RECT 71.605 159.330 71.895 159.375 ;
        RECT 72.970 159.330 73.290 159.390 ;
        RECT 71.605 159.190 76.420 159.330 ;
        RECT 58.800 159.035 58.940 159.190 ;
        RECT 71.605 159.145 71.895 159.190 ;
        RECT 72.970 159.130 73.290 159.190 ;
        RECT 54.585 158.990 54.875 159.035 ;
        RECT 54.110 158.850 54.875 158.990 ;
        RECT 54.110 158.790 54.430 158.850 ;
        RECT 54.585 158.805 54.875 158.850 ;
        RECT 58.265 158.805 58.555 159.035 ;
        RECT 58.725 158.805 59.015 159.035 ;
        RECT 59.170 158.990 59.490 159.050 ;
        RECT 59.645 158.990 59.935 159.035 ;
        RECT 59.170 158.850 59.935 158.990 ;
        RECT 42.610 158.355 42.930 158.370 ;
        RECT 42.610 158.125 42.945 158.355 ;
        RECT 43.085 158.310 43.375 158.355 ;
        RECT 44.540 158.310 44.680 158.790 ;
        RECT 58.340 158.650 58.480 158.805 ;
        RECT 59.170 158.790 59.490 158.850 ;
        RECT 59.645 158.805 59.935 158.850 ;
        RECT 72.525 158.990 72.815 159.035 ;
        RECT 75.285 158.990 75.575 159.035 ;
        RECT 72.525 158.850 75.575 158.990 ;
        RECT 72.525 158.805 72.815 158.850 ;
        RECT 75.285 158.805 75.575 158.850 ;
        RECT 60.565 158.650 60.855 158.695 ;
        RECT 72.600 158.650 72.740 158.805 ;
        RECT 75.730 158.790 76.050 159.050 ;
        RECT 76.280 159.035 76.420 159.190 ;
        RECT 77.570 159.130 77.890 159.390 ;
        RECT 78.490 159.330 78.810 159.390 ;
        RECT 79.870 159.330 80.190 159.390 ;
        RECT 78.490 159.190 80.190 159.330 ;
        RECT 78.490 159.130 78.810 159.190 ;
        RECT 76.205 158.805 76.495 159.035 ;
        RECT 77.660 158.990 77.800 159.130 ;
        RECT 79.500 159.035 79.640 159.190 ;
        RECT 79.870 159.130 80.190 159.190 ;
        RECT 81.250 159.330 81.570 159.390 ;
        RECT 82.630 159.330 82.950 159.390 ;
        RECT 81.250 159.190 82.950 159.330 ;
        RECT 81.250 159.130 81.570 159.190 ;
        RECT 82.630 159.130 82.950 159.190 ;
        RECT 95.970 159.330 96.290 159.390 ;
        RECT 95.970 159.190 98.500 159.330 ;
        RECT 95.970 159.130 96.290 159.190 ;
        RECT 78.965 158.990 79.255 159.035 ;
        RECT 77.660 158.850 79.255 158.990 ;
        RECT 78.965 158.805 79.255 158.850 ;
        RECT 79.425 158.990 79.715 159.035 ;
        RECT 82.185 158.990 82.475 159.035 ;
        RECT 79.425 158.850 82.475 158.990 ;
        RECT 79.425 158.805 79.715 158.850 ;
        RECT 82.185 158.805 82.475 158.850 ;
        RECT 95.510 158.990 95.830 159.050 ;
        RECT 96.905 158.990 97.195 159.035 ;
        RECT 95.510 158.850 97.195 158.990 ;
        RECT 95.510 158.790 95.830 158.850 ;
        RECT 96.905 158.805 97.195 158.850 ;
        RECT 58.340 158.510 60.320 158.650 ;
        RECT 60.180 158.370 60.320 158.510 ;
        RECT 60.565 158.510 72.740 158.650 ;
        RECT 78.490 158.650 78.810 158.710 ;
        RECT 84.025 158.650 84.315 158.695 ;
        RECT 87.690 158.650 88.010 158.710 ;
        RECT 78.490 158.510 88.010 158.650 ;
        RECT 60.565 158.465 60.855 158.510 ;
        RECT 78.490 158.450 78.810 158.510 ;
        RECT 84.025 158.465 84.315 158.510 ;
        RECT 87.690 158.450 88.010 158.510 ;
        RECT 43.085 158.170 44.680 158.310 ;
        RECT 43.085 158.125 43.375 158.170 ;
        RECT 42.610 158.110 42.930 158.125 ;
        RECT 60.090 158.110 60.410 158.370 ;
        RECT 73.430 158.110 73.750 158.370 ;
        RECT 75.270 158.310 75.590 158.370 ;
        RECT 90.450 158.310 90.770 158.370 ;
        RECT 75.270 158.170 90.770 158.310 ;
        RECT 96.980 158.310 97.120 158.805 ;
        RECT 97.350 158.790 97.670 159.050 ;
        RECT 97.810 158.790 98.130 159.050 ;
        RECT 98.360 159.035 98.500 159.190 ;
        RECT 100.110 159.130 100.430 159.390 ;
        RECT 101.120 159.330 101.260 159.870 ;
        RECT 106.090 159.810 106.410 160.070 ;
        RECT 108.850 160.010 109.170 160.070 ;
        RECT 108.850 159.870 111.840 160.010 ;
        RECT 108.850 159.810 109.170 159.870 ;
        RECT 106.180 159.670 106.320 159.810 ;
        RECT 102.960 159.530 106.320 159.670 ;
        RECT 102.960 159.375 103.100 159.530 ;
        RECT 110.230 159.470 110.550 159.730 ;
        RECT 111.700 159.670 111.840 159.870 ;
        RECT 121.730 159.810 122.050 160.070 ;
        RECT 124.490 160.010 124.810 160.070 ;
        RECT 124.965 160.010 125.255 160.055 ;
        RECT 124.490 159.870 125.255 160.010 ;
        RECT 124.490 159.810 124.810 159.870 ;
        RECT 124.965 159.825 125.255 159.870 ;
        RECT 125.870 160.010 126.190 160.070 ;
        RECT 134.150 160.010 134.470 160.070 ;
        RECT 125.870 159.870 134.470 160.010 ;
        RECT 125.870 159.810 126.190 159.870 ;
        RECT 134.150 159.810 134.470 159.870 ;
        RECT 140.130 160.010 140.450 160.070 ;
        RECT 143.350 160.010 143.670 160.070 ;
        RECT 140.130 159.870 143.670 160.010 ;
        RECT 140.130 159.810 140.450 159.870 ;
        RECT 143.350 159.810 143.670 159.870 ;
        RECT 143.810 160.010 144.130 160.070 ;
        RECT 143.810 159.870 147.260 160.010 ;
        RECT 143.810 159.810 144.130 159.870 ;
        RECT 121.820 159.670 121.960 159.810 ;
        RECT 133.690 159.670 134.010 159.730 ;
        RECT 136.450 159.670 136.770 159.730 ;
        RECT 141.050 159.670 141.370 159.730 ;
        RECT 141.525 159.670 141.815 159.715 ;
        RECT 146.125 159.670 146.415 159.715 ;
        RECT 111.700 159.530 115.520 159.670 ;
        RECT 121.820 159.530 128.400 159.670 ;
        RECT 102.425 159.330 102.715 159.375 ;
        RECT 101.120 159.190 102.715 159.330 ;
        RECT 102.425 159.145 102.715 159.190 ;
        RECT 102.885 159.145 103.175 159.375 ;
        RECT 105.185 159.330 105.475 159.375 ;
        RECT 103.420 159.190 105.475 159.330 ;
        RECT 98.285 158.805 98.575 159.035 ;
        RECT 98.745 158.805 99.035 159.035 ;
        RECT 97.440 158.650 97.580 158.790 ;
        RECT 98.820 158.650 98.960 158.805 ;
        RECT 99.190 158.790 99.510 159.050 ;
        RECT 99.650 158.990 99.970 159.050 ;
        RECT 101.045 158.990 101.335 159.035 ;
        RECT 99.650 158.850 101.335 158.990 ;
        RECT 99.650 158.790 99.970 158.850 ;
        RECT 101.045 158.805 101.335 158.850 ;
        RECT 101.965 158.990 102.255 159.035 ;
        RECT 103.420 158.990 103.560 159.190 ;
        RECT 105.185 159.145 105.475 159.190 ;
        RECT 105.630 159.330 105.950 159.390 ;
        RECT 110.320 159.330 110.460 159.470 ;
        RECT 111.700 159.375 111.840 159.530 ;
        RECT 115.380 159.390 115.520 159.530 ;
        RECT 105.630 159.190 110.000 159.330 ;
        RECT 110.320 159.190 110.920 159.330 ;
        RECT 105.630 159.130 105.950 159.190 ;
        RECT 101.965 158.850 103.560 158.990 ;
        RECT 103.805 158.990 104.095 159.035 ;
        RECT 104.250 158.990 104.570 159.050 ;
        RECT 103.805 158.850 104.570 158.990 ;
        RECT 101.965 158.805 102.255 158.850 ;
        RECT 103.805 158.805 104.095 158.850 ;
        RECT 97.440 158.510 98.960 158.650 ;
        RECT 99.280 158.650 99.420 158.790 ;
        RECT 102.040 158.650 102.180 158.805 ;
        RECT 104.250 158.790 104.570 158.850 ;
        RECT 106.565 158.990 106.855 159.035 ;
        RECT 109.325 158.990 109.615 159.035 ;
        RECT 106.565 158.850 109.615 158.990 ;
        RECT 106.565 158.805 106.855 158.850 ;
        RECT 109.325 158.805 109.615 158.850 ;
        RECT 99.280 158.510 102.180 158.650 ;
        RECT 104.725 158.650 105.015 158.695 ;
        RECT 108.850 158.650 109.170 158.710 ;
        RECT 104.725 158.510 109.170 158.650 ;
        RECT 104.725 158.465 105.015 158.510 ;
        RECT 108.850 158.450 109.170 158.510 ;
        RECT 105.630 158.310 105.950 158.370 ;
        RECT 96.980 158.170 105.950 158.310 ;
        RECT 75.270 158.110 75.590 158.170 ;
        RECT 90.450 158.110 90.770 158.170 ;
        RECT 105.630 158.110 105.950 158.170 ;
        RECT 107.470 158.110 107.790 158.370 ;
        RECT 109.860 158.310 110.000 159.190 ;
        RECT 110.230 158.790 110.550 159.050 ;
        RECT 110.780 158.650 110.920 159.190 ;
        RECT 111.625 159.145 111.915 159.375 ;
        RECT 112.990 159.130 113.310 159.390 ;
        RECT 113.450 159.130 113.770 159.390 ;
        RECT 115.290 159.130 115.610 159.390 ;
        RECT 126.790 159.130 127.110 159.390 ;
        RECT 111.150 158.790 111.470 159.050 ;
        RECT 112.085 158.805 112.375 159.035 ;
        RECT 113.080 158.985 113.220 159.130 ;
        RECT 112.160 158.650 112.300 158.805 ;
        RECT 113.005 158.755 113.295 158.985 ;
        RECT 113.925 158.805 114.215 159.035 ;
        RECT 114.370 158.990 114.690 159.050 ;
        RECT 128.260 159.035 128.400 159.530 ;
        RECT 133.690 159.530 135.715 159.670 ;
        RECT 133.690 159.470 134.010 159.530 ;
        RECT 133.780 159.330 133.920 159.470 ;
        RECT 135.070 159.330 135.390 159.390 ;
        RECT 132.860 159.190 133.920 159.330 ;
        RECT 134.240 159.190 135.390 159.330 ;
        RECT 135.575 159.330 135.715 159.530 ;
        RECT 136.450 159.530 138.060 159.670 ;
        RECT 136.450 159.470 136.770 159.530 ;
        RECT 135.575 159.190 136.220 159.330 ;
        RECT 132.860 159.035 133.000 159.190 ;
        RECT 114.845 158.990 115.135 159.035 ;
        RECT 114.370 158.850 115.135 158.990 ;
        RECT 110.780 158.510 112.300 158.650 ;
        RECT 114.000 158.310 114.140 158.805 ;
        RECT 114.370 158.790 114.690 158.850 ;
        RECT 114.845 158.805 115.135 158.850 ;
        RECT 125.885 158.805 126.175 159.035 ;
        RECT 128.185 158.805 128.475 159.035 ;
        RECT 132.785 158.805 133.075 159.035 ;
        RECT 133.230 158.990 133.550 159.050 ;
        RECT 134.240 159.035 134.380 159.190 ;
        RECT 135.070 159.130 135.390 159.190 ;
        RECT 133.705 158.990 133.995 159.035 ;
        RECT 133.230 158.850 133.995 158.990 ;
        RECT 125.960 158.650 126.100 158.805 ;
        RECT 133.230 158.790 133.550 158.850 ;
        RECT 133.705 158.805 133.995 158.850 ;
        RECT 134.165 158.805 134.455 159.035 ;
        RECT 134.625 158.990 134.915 159.035 ;
        RECT 135.530 158.990 135.850 159.050 ;
        RECT 134.625 158.850 135.850 158.990 ;
        RECT 136.080 158.990 136.220 159.190 ;
        RECT 136.450 158.990 136.770 159.050 ;
        RECT 136.080 158.850 136.770 158.990 ;
        RECT 134.625 158.805 134.915 158.850 ;
        RECT 126.330 158.650 126.650 158.710 ;
        RECT 125.960 158.510 126.650 158.650 ;
        RECT 126.330 158.450 126.650 158.510 ;
        RECT 131.390 158.650 131.710 158.710 ;
        RECT 134.700 158.650 134.840 158.805 ;
        RECT 135.530 158.790 135.850 158.850 ;
        RECT 136.450 158.790 136.770 158.850 ;
        RECT 136.910 158.790 137.230 159.050 ;
        RECT 137.370 158.790 137.690 159.050 ;
        RECT 137.920 159.035 138.060 159.530 ;
        RECT 141.050 159.530 141.815 159.670 ;
        RECT 141.050 159.470 141.370 159.530 ;
        RECT 141.525 159.485 141.815 159.530 ;
        RECT 142.520 159.530 146.415 159.670 ;
        RECT 137.845 158.805 138.135 159.035 ;
        RECT 138.305 158.990 138.595 159.035 ;
        RECT 138.305 158.850 140.360 158.990 ;
        RECT 138.305 158.805 138.595 158.850 ;
        RECT 131.390 158.510 134.840 158.650 ;
        RECT 136.005 158.650 136.295 158.695 ;
        RECT 137.000 158.650 137.140 158.790 ;
        RECT 136.005 158.510 137.140 158.650 ;
        RECT 131.390 158.450 131.710 158.510 ;
        RECT 136.005 158.465 136.295 158.510 ;
        RECT 109.860 158.170 114.140 158.310 ;
        RECT 114.830 158.310 115.150 158.370 ;
        RECT 115.765 158.310 116.055 158.355 ;
        RECT 114.830 158.170 116.055 158.310 ;
        RECT 114.830 158.110 115.150 158.170 ;
        RECT 115.765 158.125 116.055 158.170 ;
        RECT 117.130 158.310 117.450 158.370 ;
        RECT 138.380 158.310 138.520 158.805 ;
        RECT 117.130 158.170 138.520 158.310 ;
        RECT 139.210 158.310 139.530 158.370 ;
        RECT 140.220 158.355 140.360 158.850 ;
        RECT 140.590 158.790 140.910 159.050 ;
        RECT 141.140 159.035 141.280 159.470 ;
        RECT 141.065 158.805 141.355 159.035 ;
        RECT 141.510 158.990 141.830 159.050 ;
        RECT 142.520 159.035 142.660 159.530 ;
        RECT 146.125 159.485 146.415 159.530 ;
        RECT 142.445 158.990 142.735 159.035 ;
        RECT 141.510 158.850 142.735 158.990 ;
        RECT 141.510 158.790 141.830 158.850 ;
        RECT 142.445 158.805 142.735 158.850 ;
        RECT 143.825 158.990 144.115 159.035 ;
        RECT 144.730 158.990 145.050 159.050 ;
        RECT 147.120 159.035 147.260 159.870 ;
        RECT 143.825 158.850 145.050 158.990 ;
        RECT 143.825 158.805 144.115 158.850 ;
        RECT 144.730 158.790 145.050 158.850 ;
        RECT 145.665 158.805 145.955 159.035 ;
        RECT 147.045 158.990 147.335 159.035 ;
        RECT 147.490 158.990 147.810 159.050 ;
        RECT 147.045 158.850 147.810 158.990 ;
        RECT 147.045 158.805 147.335 158.850 ;
        RECT 139.685 158.310 139.975 158.355 ;
        RECT 139.210 158.170 139.975 158.310 ;
        RECT 117.130 158.110 117.450 158.170 ;
        RECT 139.210 158.110 139.530 158.170 ;
        RECT 139.685 158.125 139.975 158.170 ;
        RECT 140.145 158.125 140.435 158.355 ;
        RECT 140.680 158.310 140.820 158.790 ;
        RECT 143.350 158.650 143.670 158.710 ;
        RECT 144.270 158.650 144.590 158.710 ;
        RECT 145.740 158.650 145.880 158.805 ;
        RECT 147.490 158.790 147.810 158.850 ;
        RECT 143.350 158.510 145.880 158.650 ;
        RECT 143.350 158.450 143.670 158.510 ;
        RECT 144.270 158.450 144.590 158.510 ;
        RECT 144.745 158.310 145.035 158.355 ;
        RECT 140.680 158.170 145.035 158.310 ;
        RECT 144.745 158.125 145.035 158.170 ;
        RECT 36.100 157.490 150.180 157.970 ;
        RECT 44.910 157.290 45.230 157.350 ;
        RECT 51.365 157.290 51.655 157.335 ;
        RECT 54.110 157.290 54.430 157.350 ;
        RECT 44.910 157.150 47.440 157.290 ;
        RECT 44.910 157.090 45.230 157.150 ;
        RECT 47.300 156.995 47.440 157.150 ;
        RECT 51.365 157.150 54.430 157.290 ;
        RECT 51.365 157.105 51.655 157.150 ;
        RECT 54.110 157.090 54.430 157.150 ;
        RECT 65.165 157.290 65.455 157.335 ;
        RECT 67.910 157.290 68.230 157.350 ;
        RECT 65.165 157.150 68.600 157.290 ;
        RECT 65.165 157.105 65.455 157.150 ;
        RECT 67.910 157.090 68.230 157.150 ;
        RECT 47.225 156.765 47.515 156.995 ;
        RECT 48.145 156.950 48.435 156.995 ;
        RECT 50.430 156.950 50.750 157.010 ;
        RECT 52.270 156.950 52.590 157.010 ;
        RECT 48.145 156.810 52.590 156.950 ;
        RECT 48.145 156.765 48.435 156.810 ;
        RECT 50.430 156.750 50.750 156.810 ;
        RECT 52.270 156.750 52.590 156.810 ;
        RECT 57.040 156.950 57.330 156.995 ;
        RECT 66.085 156.950 66.375 156.995 ;
        RECT 57.040 156.810 66.375 156.950 ;
        RECT 57.040 156.765 57.330 156.810 ;
        RECT 66.085 156.765 66.375 156.810 ;
        RECT 66.620 156.810 68.140 156.950 ;
        RECT 37.550 156.610 37.870 156.670 ;
        RECT 39.390 156.655 39.710 156.670 ;
        RECT 38.025 156.610 38.315 156.655 ;
        RECT 37.550 156.470 38.315 156.610 ;
        RECT 37.550 156.410 37.870 156.470 ;
        RECT 38.025 156.425 38.315 156.470 ;
        RECT 39.360 156.425 39.710 156.655 ;
        RECT 39.390 156.410 39.710 156.425 ;
        RECT 58.250 156.410 58.570 156.670 ;
        RECT 60.565 156.610 60.855 156.655 ;
        RECT 63.770 156.610 64.090 156.670 ;
        RECT 60.565 156.470 64.090 156.610 ;
        RECT 60.565 156.425 60.855 156.470 ;
        RECT 63.770 156.410 64.090 156.470 ;
        RECT 65.625 156.610 65.915 156.655 ;
        RECT 66.620 156.610 66.760 156.810 ;
        RECT 65.625 156.470 66.760 156.610 ;
        RECT 65.625 156.425 65.915 156.470 ;
        RECT 67.005 156.425 67.295 156.655 ;
        RECT 38.905 156.270 39.195 156.315 ;
        RECT 40.095 156.270 40.385 156.315 ;
        RECT 42.615 156.270 42.905 156.315 ;
        RECT 38.905 156.130 42.905 156.270 ;
        RECT 38.905 156.085 39.195 156.130 ;
        RECT 40.095 156.085 40.385 156.130 ;
        RECT 42.615 156.085 42.905 156.130 ;
        RECT 53.675 156.270 53.965 156.315 ;
        RECT 56.195 156.270 56.485 156.315 ;
        RECT 57.385 156.270 57.675 156.315 ;
        RECT 53.675 156.130 57.675 156.270 ;
        RECT 53.675 156.085 53.965 156.130 ;
        RECT 56.195 156.085 56.485 156.130 ;
        RECT 57.385 156.085 57.675 156.130 ;
        RECT 60.090 156.070 60.410 156.330 ;
        RECT 63.325 156.085 63.615 156.315 ;
        RECT 64.245 156.270 64.535 156.315 ;
        RECT 67.080 156.270 67.220 156.425 ;
        RECT 64.245 156.130 67.220 156.270 ;
        RECT 64.245 156.085 64.535 156.130 ;
        RECT 38.510 155.930 38.800 155.975 ;
        RECT 40.610 155.930 40.900 155.975 ;
        RECT 42.180 155.930 42.470 155.975 ;
        RECT 38.510 155.790 42.470 155.930 ;
        RECT 38.510 155.745 38.800 155.790 ;
        RECT 40.610 155.745 40.900 155.790 ;
        RECT 42.180 155.745 42.470 155.790 ;
        RECT 54.110 155.930 54.400 155.975 ;
        RECT 55.680 155.930 55.970 155.975 ;
        RECT 57.780 155.930 58.070 155.975 ;
        RECT 54.110 155.790 58.070 155.930 ;
        RECT 54.110 155.745 54.400 155.790 ;
        RECT 55.680 155.745 55.970 155.790 ;
        RECT 57.780 155.745 58.070 155.790 ;
        RECT 58.710 155.730 59.030 155.990 ;
        RECT 63.400 155.930 63.540 156.085 ;
        RECT 66.530 155.930 66.850 155.990 ;
        RECT 63.400 155.790 66.850 155.930 ;
        RECT 66.530 155.730 66.850 155.790 ;
        RECT 68.000 155.635 68.140 156.810 ;
        RECT 68.460 156.655 68.600 157.150 ;
        RECT 75.730 157.090 76.050 157.350 ;
        RECT 77.570 157.290 77.890 157.350 ;
        RECT 78.505 157.290 78.795 157.335 ;
        RECT 80.790 157.290 81.110 157.350 ;
        RECT 76.280 157.150 77.340 157.290 ;
        RECT 73.430 156.750 73.750 157.010 ;
        RECT 75.820 156.950 75.960 157.090 ;
        RECT 73.980 156.810 75.960 156.950 ;
        RECT 68.385 156.425 68.675 156.655 ;
        RECT 71.605 156.425 71.895 156.655 ;
        RECT 72.985 156.610 73.275 156.655 ;
        RECT 73.520 156.610 73.660 156.750 ;
        RECT 73.980 156.655 74.120 156.810 ;
        RECT 76.280 156.655 76.420 157.150 ;
        RECT 72.985 156.470 73.660 156.610 ;
        RECT 72.985 156.425 73.275 156.470 ;
        RECT 73.905 156.425 74.195 156.655 ;
        RECT 74.365 156.425 74.655 156.655 ;
        RECT 76.205 156.425 76.495 156.655 ;
        RECT 77.200 156.610 77.340 157.150 ;
        RECT 77.570 157.150 78.260 157.290 ;
        RECT 77.570 157.090 77.890 157.150 ;
        RECT 78.120 156.950 78.260 157.150 ;
        RECT 78.505 157.150 81.110 157.290 ;
        RECT 78.505 157.105 78.795 157.150 ;
        RECT 80.790 157.090 81.110 157.150 ;
        RECT 83.550 157.090 83.870 157.350 ;
        RECT 86.310 157.290 86.630 157.350 ;
        RECT 92.290 157.290 92.610 157.350 ;
        RECT 97.810 157.290 98.130 157.350 ;
        RECT 98.745 157.290 99.035 157.335 ;
        RECT 84.100 157.150 86.630 157.290 ;
        RECT 84.100 156.950 84.240 157.150 ;
        RECT 86.310 157.090 86.630 157.150 ;
        RECT 86.860 157.150 92.610 157.290 ;
        RECT 85.390 156.950 85.710 157.010 ;
        RECT 86.860 156.950 87.000 157.150 ;
        RECT 92.290 157.090 92.610 157.150 ;
        RECT 93.760 157.150 95.510 157.290 ;
        RECT 78.120 156.810 80.560 156.950 ;
        RECT 78.965 156.610 79.255 156.655 ;
        RECT 77.200 156.470 79.255 156.610 ;
        RECT 78.965 156.425 79.255 156.470 ;
        RECT 69.750 155.930 70.070 155.990 ;
        RECT 71.680 155.930 71.820 156.425 ;
        RECT 73.445 156.270 73.735 156.315 ;
        RECT 74.440 156.270 74.580 156.425 ;
        RECT 79.870 156.410 80.190 156.670 ;
        RECT 80.420 156.655 80.560 156.810 ;
        RECT 81.800 156.810 84.240 156.950 ;
        RECT 84.560 156.810 85.710 156.950 ;
        RECT 80.345 156.425 80.635 156.655 ;
        RECT 73.445 156.130 75.960 156.270 ;
        RECT 73.445 156.085 73.735 156.130 ;
        RECT 73.890 155.930 74.210 155.990 ;
        RECT 69.750 155.790 74.210 155.930 ;
        RECT 69.750 155.730 70.070 155.790 ;
        RECT 73.890 155.730 74.210 155.790 ;
        RECT 74.810 155.730 75.130 155.990 ;
        RECT 75.820 155.930 75.960 156.130 ;
        RECT 76.650 156.070 76.970 156.330 ;
        RECT 77.125 156.085 77.415 156.315 ;
        RECT 77.585 156.270 77.875 156.315 ;
        RECT 78.490 156.270 78.810 156.330 ;
        RECT 81.800 156.270 81.940 156.810 ;
        RECT 82.185 156.610 82.475 156.655 ;
        RECT 84.560 156.610 84.700 156.810 ;
        RECT 85.390 156.750 85.710 156.810 ;
        RECT 85.940 156.810 87.000 156.950 ;
        RECT 82.185 156.470 82.860 156.610 ;
        RECT 82.185 156.425 82.475 156.470 ;
        RECT 82.720 156.315 82.860 156.470 ;
        RECT 84.100 156.470 84.700 156.610 ;
        RECT 84.945 156.610 85.235 156.655 ;
        RECT 85.940 156.610 86.080 156.810 ;
        RECT 90.450 156.750 90.770 157.010 ;
        RECT 93.145 156.950 93.435 156.995 ;
        RECT 93.760 156.950 93.900 157.150 ;
        RECT 93.145 156.810 93.900 156.950 ;
        RECT 93.145 156.765 93.435 156.810 ;
        RECT 94.145 156.765 94.435 156.995 ;
        RECT 95.370 156.950 95.510 157.150 ;
        RECT 97.810 157.150 99.035 157.290 ;
        RECT 97.810 157.090 98.130 157.150 ;
        RECT 98.745 157.105 99.035 157.150 ;
        RECT 99.280 157.150 105.400 157.290 ;
        RECT 99.280 156.950 99.420 157.150 ;
        RECT 95.370 156.810 99.420 156.950 ;
        RECT 84.945 156.470 86.080 156.610 ;
        RECT 77.585 156.130 78.810 156.270 ;
        RECT 77.585 156.085 77.875 156.130 ;
        RECT 77.200 155.930 77.340 156.085 ;
        RECT 78.490 156.070 78.810 156.130 ;
        RECT 79.040 156.130 81.940 156.270 ;
        RECT 79.040 155.990 79.180 156.130 ;
        RECT 82.645 156.085 82.935 156.315 ;
        RECT 83.105 156.270 83.395 156.315 ;
        RECT 84.100 156.270 84.240 156.470 ;
        RECT 84.945 156.425 85.235 156.470 ;
        RECT 86.310 156.410 86.630 156.670 ;
        RECT 87.245 156.610 87.535 156.655 ;
        RECT 87.690 156.610 88.010 156.670 ;
        RECT 87.245 156.470 88.010 156.610 ;
        RECT 90.540 156.610 90.680 156.750 ;
        RECT 94.220 156.610 94.360 156.765 ;
        RECT 100.570 156.750 100.890 157.010 ;
        RECT 104.250 156.950 104.570 157.010 ;
        RECT 102.960 156.810 104.570 156.950 ;
        RECT 90.540 156.470 94.360 156.610 ;
        RECT 94.605 156.610 94.895 156.655 ;
        RECT 95.050 156.610 95.370 156.670 ;
        RECT 94.605 156.470 95.370 156.610 ;
        RECT 87.245 156.425 87.535 156.470 ;
        RECT 87.690 156.410 88.010 156.470 ;
        RECT 94.605 156.425 94.895 156.470 ;
        RECT 95.050 156.410 95.370 156.470 ;
        RECT 99.190 156.610 99.510 156.670 ;
        RECT 99.665 156.610 99.955 156.655 ;
        RECT 99.190 156.470 99.955 156.610 ;
        RECT 99.190 156.410 99.510 156.470 ;
        RECT 99.665 156.425 99.955 156.470 ;
        RECT 100.125 156.610 100.415 156.655 ;
        RECT 100.660 156.610 100.800 156.750 ;
        RECT 102.960 156.670 103.100 156.810 ;
        RECT 104.250 156.750 104.570 156.810 ;
        RECT 101.490 156.655 101.810 156.670 ;
        RECT 100.125 156.470 100.800 156.610 ;
        RECT 100.125 156.425 100.415 156.470 ;
        RECT 101.415 156.425 101.810 156.655 ;
        RECT 101.965 156.610 102.255 156.655 ;
        RECT 101.965 156.470 102.640 156.610 ;
        RECT 101.965 156.425 102.255 156.470 ;
        RECT 101.490 156.410 101.810 156.425 ;
        RECT 102.500 156.330 102.640 156.470 ;
        RECT 102.870 156.410 103.190 156.670 ;
        RECT 83.105 156.130 84.240 156.270 ;
        RECT 84.485 156.270 84.775 156.315 ;
        RECT 85.850 156.270 86.170 156.330 ;
        RECT 84.485 156.130 86.170 156.270 ;
        RECT 83.105 156.085 83.395 156.130 ;
        RECT 84.485 156.085 84.775 156.130 ;
        RECT 75.820 155.790 77.340 155.930 ;
        RECT 78.950 155.730 79.270 155.990 ;
        RECT 82.170 155.930 82.490 155.990 ;
        RECT 80.420 155.790 82.490 155.930 ;
        RECT 82.720 155.930 82.860 156.085 ;
        RECT 85.850 156.070 86.170 156.130 ;
        RECT 91.385 156.085 91.675 156.315 ;
        RECT 86.785 155.930 87.075 155.975 ;
        RECT 82.720 155.790 87.075 155.930 ;
        RECT 67.925 155.590 68.215 155.635 ;
        RECT 68.370 155.590 68.690 155.650 ;
        RECT 67.925 155.450 68.690 155.590 ;
        RECT 67.925 155.405 68.215 155.450 ;
        RECT 68.370 155.390 68.690 155.450 ;
        RECT 72.525 155.590 72.815 155.635 ;
        RECT 72.970 155.590 73.290 155.650 ;
        RECT 74.900 155.590 75.040 155.730 ;
        RECT 72.525 155.450 75.040 155.590 ;
        RECT 75.285 155.590 75.575 155.635 ;
        RECT 80.420 155.590 80.560 155.790 ;
        RECT 82.170 155.730 82.490 155.790 ;
        RECT 86.785 155.745 87.075 155.790 ;
        RECT 88.610 155.930 88.930 155.990 ;
        RECT 89.545 155.930 89.835 155.975 ;
        RECT 88.610 155.790 89.835 155.930 ;
        RECT 91.460 155.930 91.600 156.085 ;
        RECT 102.410 156.070 102.730 156.330 ;
        RECT 105.260 156.270 105.400 157.150 ;
        RECT 107.930 157.090 108.250 157.350 ;
        RECT 110.230 157.290 110.550 157.350 ;
        RECT 110.230 157.150 124.720 157.290 ;
        RECT 110.230 157.090 110.550 157.150 ;
        RECT 108.020 156.950 108.160 157.090 ;
        RECT 117.130 156.950 117.450 157.010 ;
        RECT 123.585 156.950 123.875 156.995 ;
        RECT 108.020 156.810 110.460 156.950 ;
        RECT 105.630 156.610 105.950 156.670 ;
        RECT 108.865 156.610 109.155 156.655 ;
        RECT 105.630 156.470 109.155 156.610 ;
        RECT 105.630 156.410 105.950 156.470 ;
        RECT 108.865 156.425 109.155 156.470 ;
        RECT 109.770 156.410 110.090 156.670 ;
        RECT 110.320 156.655 110.460 156.810 ;
        RECT 114.000 156.810 117.450 156.950 ;
        RECT 110.245 156.425 110.535 156.655 ;
        RECT 110.705 156.425 110.995 156.655 ;
        RECT 109.310 156.270 109.630 156.330 ;
        RECT 105.260 156.130 109.630 156.270 ;
        RECT 110.780 156.270 110.920 156.425 ;
        RECT 112.070 156.410 112.390 156.670 ;
        RECT 113.450 156.610 113.770 156.670 ;
        RECT 114.000 156.655 114.140 156.810 ;
        RECT 117.130 156.750 117.450 156.810 ;
        RECT 119.980 156.810 123.875 156.950 ;
        RECT 113.925 156.610 114.215 156.655 ;
        RECT 113.450 156.470 114.215 156.610 ;
        RECT 113.450 156.410 113.770 156.470 ;
        RECT 113.925 156.425 114.215 156.470 ;
        RECT 114.845 156.610 115.135 156.655 ;
        RECT 115.290 156.610 115.610 156.670 ;
        RECT 114.845 156.470 115.610 156.610 ;
        RECT 114.845 156.425 115.135 156.470 ;
        RECT 115.290 156.410 115.610 156.470 ;
        RECT 119.430 156.610 119.750 156.670 ;
        RECT 119.980 156.655 120.120 156.810 ;
        RECT 123.585 156.765 123.875 156.810 ;
        RECT 124.580 156.950 124.720 157.150 ;
        RECT 126.330 157.090 126.650 157.350 ;
        RECT 129.235 157.290 129.525 157.335 ;
        RECT 132.770 157.290 133.090 157.350 ;
        RECT 129.235 157.150 133.090 157.290 ;
        RECT 129.235 157.105 129.525 157.150 ;
        RECT 132.770 157.090 133.090 157.150 ;
        RECT 133.245 157.290 133.535 157.335 ;
        RECT 137.370 157.290 137.690 157.350 ;
        RECT 133.245 157.150 137.690 157.290 ;
        RECT 133.245 157.105 133.535 157.150 ;
        RECT 137.370 157.090 137.690 157.150 ;
        RECT 139.210 157.090 139.530 157.350 ;
        RECT 146.585 157.290 146.875 157.335 ;
        RECT 147.490 157.290 147.810 157.350 ;
        RECT 146.585 157.150 147.810 157.290 ;
        RECT 146.585 157.105 146.875 157.150 ;
        RECT 147.490 157.090 147.810 157.150 ;
        RECT 128.185 156.950 128.475 156.995 ;
        RECT 137.830 156.950 138.150 157.010 ;
        RECT 124.580 156.810 138.150 156.950 ;
        RECT 139.300 156.950 139.440 157.090 ;
        RECT 140.910 156.950 141.200 156.995 ;
        RECT 139.300 156.810 141.200 156.950 ;
        RECT 119.905 156.610 120.195 156.655 ;
        RECT 119.430 156.470 120.195 156.610 ;
        RECT 119.430 156.410 119.750 156.470 ;
        RECT 119.905 156.425 120.195 156.470 ;
        RECT 120.825 156.610 121.115 156.655 ;
        RECT 123.110 156.610 123.430 156.670 ;
        RECT 124.580 156.655 124.720 156.810 ;
        RECT 128.185 156.765 128.475 156.810 ;
        RECT 137.830 156.750 138.150 156.810 ;
        RECT 140.910 156.765 141.200 156.810 ;
        RECT 120.825 156.470 123.430 156.610 ;
        RECT 120.825 156.425 121.115 156.470 ;
        RECT 123.110 156.410 123.430 156.470 ;
        RECT 124.045 156.425 124.335 156.655 ;
        RECT 124.505 156.425 124.795 156.655 ;
        RECT 126.805 156.425 127.095 156.655 ;
        RECT 112.160 156.270 112.300 156.410 ;
        RECT 124.120 156.270 124.260 156.425 ;
        RECT 110.780 156.130 123.800 156.270 ;
        RECT 124.120 156.130 126.560 156.270 ;
        RECT 109.310 156.070 109.630 156.130 ;
        RECT 95.525 155.930 95.815 155.975 ;
        RECT 110.690 155.930 111.010 155.990 ;
        RECT 117.590 155.930 117.910 155.990 ;
        RECT 91.460 155.790 110.000 155.930 ;
        RECT 88.610 155.730 88.930 155.790 ;
        RECT 89.545 155.745 89.835 155.790 ;
        RECT 95.525 155.745 95.815 155.790 ;
        RECT 75.285 155.450 80.560 155.590 ;
        RECT 80.790 155.590 81.110 155.650 ;
        RECT 85.865 155.590 86.155 155.635 ;
        RECT 80.790 155.450 86.155 155.590 ;
        RECT 72.525 155.405 72.815 155.450 ;
        RECT 72.970 155.390 73.290 155.450 ;
        RECT 75.285 155.405 75.575 155.450 ;
        RECT 80.790 155.390 81.110 155.450 ;
        RECT 85.865 155.405 86.155 155.450 ;
        RECT 86.310 155.590 86.630 155.650 ;
        RECT 89.085 155.590 89.375 155.635 ;
        RECT 86.310 155.450 89.375 155.590 ;
        RECT 86.310 155.390 86.630 155.450 ;
        RECT 89.085 155.405 89.375 155.450 ;
        RECT 92.290 155.390 92.610 155.650 ;
        RECT 93.225 155.590 93.515 155.635 ;
        RECT 97.350 155.590 97.670 155.650 ;
        RECT 93.225 155.450 97.670 155.590 ;
        RECT 93.225 155.405 93.515 155.450 ;
        RECT 97.350 155.390 97.670 155.450 ;
        RECT 98.730 155.590 99.050 155.650 ;
        RECT 101.045 155.590 101.335 155.635 ;
        RECT 98.730 155.450 101.335 155.590 ;
        RECT 98.730 155.390 99.050 155.450 ;
        RECT 101.045 155.405 101.335 155.450 ;
        RECT 102.425 155.590 102.715 155.635 ;
        RECT 105.630 155.590 105.950 155.650 ;
        RECT 102.425 155.450 105.950 155.590 ;
        RECT 109.860 155.590 110.000 155.790 ;
        RECT 110.690 155.790 117.910 155.930 ;
        RECT 123.660 155.930 123.800 156.130 ;
        RECT 124.950 155.930 125.270 155.990 ;
        RECT 123.660 155.790 125.270 155.930 ;
        RECT 110.690 155.730 111.010 155.790 ;
        RECT 117.590 155.730 117.910 155.790 ;
        RECT 124.950 155.730 125.270 155.790 ;
        RECT 111.150 155.590 111.470 155.650 ;
        RECT 109.860 155.450 111.470 155.590 ;
        RECT 102.425 155.405 102.715 155.450 ;
        RECT 105.630 155.390 105.950 155.450 ;
        RECT 111.150 155.390 111.470 155.450 ;
        RECT 112.070 155.390 112.390 155.650 ;
        RECT 114.370 155.390 114.690 155.650 ;
        RECT 119.890 155.390 120.210 155.650 ;
        RECT 125.425 155.590 125.715 155.635 ;
        RECT 125.870 155.590 126.190 155.650 ;
        RECT 125.425 155.450 126.190 155.590 ;
        RECT 126.420 155.590 126.560 156.130 ;
        RECT 126.880 155.990 127.020 156.425 ;
        RECT 131.390 156.410 131.710 156.670 ;
        RECT 132.310 156.410 132.630 156.670 ;
        RECT 134.625 156.610 134.915 156.655 ;
        RECT 137.370 156.610 137.690 156.670 ;
        RECT 134.625 156.470 137.690 156.610 ;
        RECT 134.625 156.425 134.915 156.470 ;
        RECT 133.230 156.270 133.550 156.330 ;
        RECT 128.720 156.130 133.550 156.270 ;
        RECT 126.790 155.930 127.110 155.990 ;
        RECT 128.720 155.930 128.860 156.130 ;
        RECT 133.230 156.070 133.550 156.130 ;
        RECT 134.700 155.930 134.840 156.425 ;
        RECT 137.370 156.410 137.690 156.470 ;
        RECT 139.670 156.410 139.990 156.670 ;
        RECT 140.565 156.270 140.855 156.315 ;
        RECT 141.755 156.270 142.045 156.315 ;
        RECT 144.275 156.270 144.565 156.315 ;
        RECT 140.565 156.130 144.565 156.270 ;
        RECT 140.565 156.085 140.855 156.130 ;
        RECT 141.755 156.085 142.045 156.130 ;
        RECT 144.275 156.085 144.565 156.130 ;
        RECT 126.790 155.790 128.860 155.930 ;
        RECT 129.180 155.790 134.840 155.930 ;
        RECT 140.170 155.930 140.460 155.975 ;
        RECT 142.270 155.930 142.560 155.975 ;
        RECT 143.840 155.930 144.130 155.975 ;
        RECT 140.170 155.790 144.130 155.930 ;
        RECT 126.790 155.730 127.110 155.790 ;
        RECT 128.630 155.590 128.950 155.650 ;
        RECT 129.180 155.635 129.320 155.790 ;
        RECT 140.170 155.745 140.460 155.790 ;
        RECT 142.270 155.745 142.560 155.790 ;
        RECT 143.840 155.745 144.130 155.790 ;
        RECT 129.105 155.590 129.395 155.635 ;
        RECT 126.420 155.450 129.395 155.590 ;
        RECT 125.425 155.405 125.715 155.450 ;
        RECT 125.870 155.390 126.190 155.450 ;
        RECT 128.630 155.390 128.950 155.450 ;
        RECT 129.105 155.405 129.395 155.450 ;
        RECT 130.025 155.590 130.315 155.635 ;
        RECT 132.770 155.590 133.090 155.650 ;
        RECT 130.025 155.450 133.090 155.590 ;
        RECT 130.025 155.405 130.315 155.450 ;
        RECT 132.770 155.390 133.090 155.450 ;
        RECT 133.690 155.390 134.010 155.650 ;
        RECT 36.100 154.770 150.180 155.250 ;
        RECT 39.390 154.570 39.710 154.630 ;
        RECT 40.325 154.570 40.615 154.615 ;
        RECT 39.390 154.430 40.615 154.570 ;
        RECT 39.390 154.370 39.710 154.430 ;
        RECT 40.325 154.385 40.615 154.430 ;
        RECT 47.225 154.570 47.515 154.615 ;
        RECT 49.525 154.570 49.815 154.615 ;
        RECT 52.730 154.570 53.050 154.630 ;
        RECT 47.225 154.430 53.050 154.570 ;
        RECT 47.225 154.385 47.515 154.430 ;
        RECT 49.525 154.385 49.815 154.430 ;
        RECT 52.730 154.370 53.050 154.430 ;
        RECT 66.085 154.570 66.375 154.615 ;
        RECT 66.530 154.570 66.850 154.630 ;
        RECT 68.370 154.570 68.690 154.630 ;
        RECT 96.905 154.570 97.195 154.615 ;
        RECT 98.270 154.570 98.590 154.630 ;
        RECT 66.085 154.430 66.850 154.570 ;
        RECT 66.085 154.385 66.375 154.430 ;
        RECT 45.385 154.230 45.675 154.275 ;
        RECT 48.590 154.230 48.910 154.290 ;
        RECT 45.385 154.090 48.910 154.230 ;
        RECT 45.385 154.045 45.675 154.090 ;
        RECT 48.590 154.030 48.910 154.090 ;
        RECT 41.230 153.350 41.550 153.610 ;
        RECT 43.085 153.365 43.375 153.595 ;
        RECT 43.160 153.210 43.300 153.365 ;
        RECT 44.910 153.350 45.230 153.610 ;
        RECT 45.830 153.350 46.150 153.610 ;
        RECT 48.590 153.550 48.910 153.610 ;
        RECT 47.070 153.425 48.910 153.550 ;
        RECT 46.995 153.410 48.910 153.425 ;
        RECT 43.160 153.070 46.520 153.210 ;
        RECT 46.995 153.195 47.285 153.410 ;
        RECT 48.590 153.350 48.910 153.410 ;
        RECT 50.430 153.350 50.750 153.610 ;
        RECT 51.350 153.350 51.670 153.610 ;
        RECT 48.145 153.210 48.435 153.255 ;
        RECT 66.160 153.210 66.300 154.385 ;
        RECT 66.530 154.370 66.850 154.430 ;
        RECT 67.540 154.430 80.560 154.570 ;
        RECT 67.540 154.230 67.680 154.430 ;
        RECT 68.370 154.370 68.690 154.430 ;
        RECT 67.080 154.090 67.680 154.230 ;
        RECT 78.490 154.230 78.810 154.290 ;
        RECT 80.420 154.230 80.560 154.430 ;
        RECT 96.905 154.430 98.590 154.570 ;
        RECT 96.905 154.385 97.195 154.430 ;
        RECT 98.270 154.370 98.590 154.430 ;
        RECT 100.125 154.570 100.415 154.615 ;
        RECT 103.330 154.570 103.650 154.630 ;
        RECT 100.125 154.430 103.650 154.570 ;
        RECT 100.125 154.385 100.415 154.430 ;
        RECT 103.330 154.370 103.650 154.430 ;
        RECT 107.010 154.570 107.330 154.630 ;
        RECT 109.785 154.570 110.075 154.615 ;
        RECT 107.010 154.430 110.075 154.570 ;
        RECT 107.010 154.370 107.330 154.430 ;
        RECT 109.785 154.385 110.075 154.430 ;
        RECT 112.070 154.370 112.390 154.630 ;
        RECT 114.370 154.370 114.690 154.630 ;
        RECT 114.830 154.370 115.150 154.630 ;
        RECT 119.890 154.370 120.210 154.630 ;
        RECT 127.710 154.570 128.030 154.630 ;
        RECT 131.865 154.570 132.155 154.615 ;
        RECT 127.710 154.430 132.155 154.570 ;
        RECT 127.710 154.370 128.030 154.430 ;
        RECT 131.865 154.385 132.155 154.430 ;
        RECT 137.830 154.570 138.150 154.630 ;
        RECT 141.970 154.570 142.290 154.630 ;
        RECT 137.830 154.430 142.290 154.570 ;
        RECT 137.830 154.370 138.150 154.430 ;
        RECT 141.970 154.370 142.290 154.430 ;
        RECT 80.790 154.230 81.110 154.290 ;
        RECT 82.170 154.230 82.490 154.290 ;
        RECT 78.490 154.090 80.100 154.230 ;
        RECT 80.420 154.090 81.110 154.230 ;
        RECT 67.080 153.550 67.220 154.090 ;
        RECT 78.490 154.030 78.810 154.090 ;
        RECT 67.450 153.890 67.770 153.950 ;
        RECT 76.190 153.890 76.510 153.950 ;
        RECT 67.450 153.750 76.510 153.890 ;
        RECT 67.450 153.690 67.770 153.750 ;
        RECT 76.190 153.690 76.510 153.750 ;
        RECT 78.950 153.690 79.270 153.950 ;
        RECT 67.925 153.550 68.215 153.595 ;
        RECT 67.080 153.410 68.215 153.550 ;
        RECT 67.925 153.365 68.215 153.410 ;
        RECT 71.605 153.550 71.895 153.595 ;
        RECT 72.970 153.550 73.290 153.610 ;
        RECT 78.045 153.550 78.335 153.595 ;
        RECT 71.605 153.410 73.290 153.550 ;
        RECT 71.605 153.365 71.895 153.410 ;
        RECT 72.970 153.350 73.290 153.410 ;
        RECT 76.740 153.410 78.335 153.550 ;
        RECT 79.040 153.550 79.180 153.690 ;
        RECT 79.960 153.595 80.100 154.090 ;
        RECT 80.790 154.030 81.110 154.090 ;
        RECT 81.270 154.090 82.490 154.230 ;
        RECT 81.270 153.595 81.410 154.090 ;
        RECT 82.170 154.030 82.490 154.090 ;
        RECT 85.850 154.030 86.170 154.290 ;
        RECT 101.120 154.090 108.160 154.230 ;
        RECT 85.940 153.890 86.080 154.030 ;
        RECT 87.245 153.890 87.535 153.935 ;
        RECT 101.120 153.890 101.260 154.090 ;
        RECT 85.940 153.750 101.260 153.890 ;
        RECT 87.245 153.705 87.535 153.750 ;
        RECT 101.490 153.690 101.810 153.950 ;
        RECT 101.950 153.690 102.270 153.950 ;
        RECT 102.960 153.935 103.100 154.090 ;
        RECT 102.885 153.705 103.175 153.935 ;
        RECT 105.630 153.690 105.950 153.950 ;
        RECT 106.090 153.690 106.410 153.950 ;
        RECT 106.565 153.890 106.855 153.935 ;
        RECT 107.470 153.890 107.790 153.950 ;
        RECT 106.565 153.750 107.790 153.890 ;
        RECT 106.565 153.705 106.855 153.750 ;
        RECT 107.470 153.690 107.790 153.750 ;
        RECT 79.425 153.550 79.715 153.595 ;
        RECT 79.040 153.410 79.715 153.550 ;
        RECT 42.150 152.670 42.470 152.930 ;
        RECT 46.380 152.915 46.520 153.070 ;
        RECT 48.145 153.070 66.300 153.210 ;
        RECT 48.145 153.025 48.435 153.070 ;
        RECT 72.510 153.010 72.830 153.270 ;
        RECT 76.740 152.930 76.880 153.410 ;
        RECT 78.045 153.365 78.335 153.410 ;
        RECT 79.425 153.365 79.715 153.410 ;
        RECT 79.885 153.365 80.175 153.595 ;
        RECT 80.440 153.550 80.730 153.595 ;
        RECT 80.420 153.365 80.730 153.550 ;
        RECT 81.265 153.365 81.555 153.595 ;
        RECT 80.420 153.210 80.560 153.365 ;
        RECT 81.710 153.350 82.030 153.610 ;
        RECT 82.170 153.550 82.490 153.610 ;
        RECT 83.105 153.550 83.395 153.595 ;
        RECT 82.170 153.410 83.395 153.550 ;
        RECT 82.170 153.350 82.490 153.410 ;
        RECT 83.105 153.365 83.395 153.410 ;
        RECT 83.550 153.550 83.870 153.610 ;
        RECT 84.025 153.550 84.315 153.595 ;
        RECT 83.550 153.410 84.315 153.550 ;
        RECT 83.550 153.350 83.870 153.410 ;
        RECT 84.025 153.365 84.315 153.410 ;
        RECT 84.470 153.550 84.790 153.610 ;
        RECT 85.865 153.550 86.155 153.595 ;
        RECT 84.470 153.410 86.155 153.550 ;
        RECT 84.470 153.350 84.790 153.410 ;
        RECT 85.865 153.365 86.155 153.410 ;
        RECT 97.810 153.350 98.130 153.610 ;
        RECT 102.410 153.550 102.730 153.610 ;
        RECT 98.360 153.410 102.730 153.550 ;
        RECT 79.960 153.070 80.560 153.210 ;
        RECT 81.800 153.210 81.940 153.350 ;
        RECT 86.310 153.210 86.630 153.270 ;
        RECT 98.360 153.255 98.500 153.410 ;
        RECT 102.410 153.350 102.730 153.410 ;
        RECT 103.330 153.550 103.650 153.610 ;
        RECT 105.185 153.550 105.475 153.595 ;
        RECT 103.330 153.410 105.475 153.550 ;
        RECT 103.330 153.350 103.650 153.410 ;
        RECT 105.185 153.365 105.475 153.410 ;
        RECT 98.285 153.210 98.575 153.255 ;
        RECT 81.800 153.070 86.630 153.210 ;
        RECT 46.305 152.685 46.595 152.915 ;
        RECT 59.170 152.870 59.490 152.930 ;
        RECT 65.165 152.870 65.455 152.915 ;
        RECT 59.170 152.730 65.455 152.870 ;
        RECT 59.170 152.670 59.490 152.730 ;
        RECT 65.165 152.685 65.455 152.730 ;
        RECT 66.085 152.870 66.375 152.915 ;
        RECT 70.685 152.870 70.975 152.915 ;
        RECT 66.085 152.730 70.975 152.870 ;
        RECT 66.085 152.685 66.375 152.730 ;
        RECT 70.685 152.685 70.975 152.730 ;
        RECT 76.650 152.670 76.970 152.930 ;
        RECT 78.490 152.870 78.810 152.930 ;
        RECT 78.965 152.870 79.255 152.915 ;
        RECT 79.960 152.870 80.100 153.070 ;
        RECT 86.310 153.010 86.630 153.070 ;
        RECT 92.380 153.070 98.575 153.210 ;
        RECT 92.380 152.930 92.520 153.070 ;
        RECT 98.285 153.025 98.575 153.070 ;
        RECT 99.205 153.025 99.495 153.255 ;
        RECT 78.490 152.730 80.100 152.870 ;
        RECT 78.490 152.670 78.810 152.730 ;
        RECT 78.965 152.685 79.255 152.730 ;
        RECT 82.170 152.670 82.490 152.930 ;
        RECT 84.945 152.870 85.235 152.915 ;
        RECT 88.610 152.870 88.930 152.930 ;
        RECT 84.945 152.730 88.930 152.870 ;
        RECT 84.945 152.685 85.235 152.730 ;
        RECT 88.610 152.670 88.930 152.730 ;
        RECT 92.290 152.670 92.610 152.930 ;
        RECT 95.050 152.870 95.370 152.930 ;
        RECT 98.730 152.870 99.050 152.930 ;
        RECT 95.050 152.730 99.050 152.870 ;
        RECT 99.280 152.870 99.420 153.025 ;
        RECT 107.470 153.010 107.790 153.270 ;
        RECT 108.020 153.210 108.160 154.090 ;
        RECT 112.160 153.935 112.300 154.370 ;
        RECT 108.480 153.750 111.840 153.890 ;
        RECT 108.480 153.595 108.620 153.750 ;
        RECT 108.405 153.365 108.695 153.595 ;
        RECT 110.690 153.550 111.010 153.610 ;
        RECT 108.940 153.410 111.010 153.550 ;
        RECT 108.940 153.210 109.080 153.410 ;
        RECT 110.690 153.350 111.010 153.410 ;
        RECT 111.150 153.350 111.470 153.610 ;
        RECT 111.700 153.595 111.840 153.750 ;
        RECT 112.085 153.705 112.375 153.935 ;
        RECT 113.450 153.690 113.770 153.950 ;
        RECT 114.460 153.935 114.600 154.370 ;
        RECT 114.920 154.230 115.060 154.370 ;
        RECT 119.980 154.230 120.120 154.370 ;
        RECT 114.920 154.090 115.520 154.230 ;
        RECT 114.385 153.705 114.675 153.935 ;
        RECT 114.830 153.690 115.150 153.950 ;
        RECT 115.380 153.935 115.520 154.090 ;
        RECT 118.140 154.090 120.120 154.230 ;
        RECT 125.870 154.230 126.190 154.290 ;
        RECT 130.470 154.230 130.790 154.290 ;
        RECT 125.870 154.090 130.790 154.230 ;
        RECT 115.305 153.705 115.595 153.935 ;
        RECT 111.625 153.550 111.915 153.595 ;
        RECT 113.540 153.550 113.680 153.690 ;
        RECT 111.625 153.410 113.680 153.550 ;
        RECT 111.625 153.365 111.915 153.410 ;
        RECT 113.925 153.365 114.215 153.595 ;
        RECT 108.020 153.070 109.080 153.210 ;
        RECT 109.325 153.210 109.615 153.255 ;
        RECT 114.000 153.210 114.140 153.365 ;
        RECT 116.210 153.350 116.530 153.610 ;
        RECT 118.140 153.595 118.280 154.090 ;
        RECT 125.870 154.030 126.190 154.090 ;
        RECT 130.470 154.030 130.790 154.090 ;
        RECT 132.785 154.045 133.075 154.275 ;
        RECT 124.950 153.890 125.270 153.950 ;
        RECT 124.950 153.750 127.940 153.890 ;
        RECT 124.950 153.690 125.270 153.750 ;
        RECT 118.065 153.365 118.355 153.595 ;
        RECT 118.510 153.550 118.830 153.610 ;
        RECT 118.985 153.550 119.275 153.595 ;
        RECT 118.510 153.410 127.020 153.550 ;
        RECT 109.325 153.070 114.140 153.210 ;
        RECT 116.685 153.210 116.975 153.255 ;
        RECT 117.130 153.210 117.450 153.270 ;
        RECT 116.685 153.070 117.450 153.210 ;
        RECT 109.325 153.025 109.615 153.070 ;
        RECT 116.685 153.025 116.975 153.070 ;
        RECT 117.130 153.010 117.450 153.070 ;
        RECT 101.030 152.870 101.350 152.930 ;
        RECT 99.280 152.730 101.350 152.870 ;
        RECT 95.050 152.670 95.370 152.730 ;
        RECT 98.730 152.670 99.050 152.730 ;
        RECT 101.030 152.670 101.350 152.730 ;
        RECT 103.790 152.670 104.110 152.930 ;
        RECT 104.265 152.870 104.555 152.915 ;
        RECT 111.150 152.870 111.470 152.930 ;
        RECT 104.265 152.730 111.470 152.870 ;
        RECT 104.265 152.685 104.555 152.730 ;
        RECT 111.150 152.670 111.470 152.730 ;
        RECT 112.990 152.670 113.310 152.930 ;
        RECT 114.370 152.870 114.690 152.930 ;
        RECT 118.140 152.870 118.280 153.365 ;
        RECT 118.510 153.350 118.830 153.410 ;
        RECT 118.985 153.365 119.275 153.410 ;
        RECT 126.880 152.930 127.020 153.410 ;
        RECT 127.250 153.350 127.570 153.610 ;
        RECT 114.370 152.730 118.280 152.870 ;
        RECT 126.790 152.870 127.110 152.930 ;
        RECT 127.265 152.870 127.555 152.915 ;
        RECT 126.790 152.730 127.555 152.870 ;
        RECT 127.800 152.870 127.940 153.750 ;
        RECT 128.185 153.550 128.475 153.595 ;
        RECT 128.630 153.550 128.950 153.610 ;
        RECT 128.185 153.410 128.950 153.550 ;
        RECT 128.185 153.365 128.475 153.410 ;
        RECT 128.630 153.350 128.950 153.410 ;
        RECT 130.010 153.350 130.330 153.610 ;
        RECT 132.860 153.550 133.000 154.045 ;
        RECT 138.765 153.550 139.055 153.595 ;
        RECT 132.860 153.410 139.055 153.550 ;
        RECT 138.765 153.365 139.055 153.410 ;
        RECT 131.865 153.210 132.155 153.255 ;
        RECT 133.245 153.210 133.535 153.255 ;
        RECT 131.865 153.070 133.535 153.210 ;
        RECT 131.865 153.025 132.155 153.070 ;
        RECT 133.245 153.025 133.535 153.070 ;
        RECT 133.690 153.210 134.010 153.270 ;
        RECT 134.165 153.210 134.455 153.255 ;
        RECT 133.690 153.070 134.455 153.210 ;
        RECT 133.690 153.010 134.010 153.070 ;
        RECT 134.165 153.025 134.455 153.070 ;
        RECT 134.610 153.210 134.930 153.270 ;
        RECT 135.085 153.210 135.375 153.255 ;
        RECT 134.610 153.070 135.375 153.210 ;
        RECT 134.240 152.870 134.380 153.025 ;
        RECT 134.610 153.010 134.930 153.070 ;
        RECT 135.085 153.025 135.375 153.070 ;
        RECT 127.800 152.730 134.380 152.870 ;
        RECT 114.370 152.670 114.690 152.730 ;
        RECT 126.790 152.670 127.110 152.730 ;
        RECT 127.265 152.685 127.555 152.730 ;
        RECT 139.670 152.670 139.990 152.930 ;
        RECT 36.100 152.050 150.180 152.530 ;
        RECT 45.830 151.850 46.150 151.910 ;
        RECT 53.650 151.850 53.970 151.910 ;
        RECT 45.830 151.710 53.970 151.850 ;
        RECT 45.830 151.650 46.150 151.710 ;
        RECT 40.280 151.510 40.570 151.555 ;
        RECT 42.150 151.510 42.470 151.570 ;
        RECT 40.280 151.370 42.470 151.510 ;
        RECT 40.280 151.325 40.570 151.370 ;
        RECT 42.150 151.310 42.470 151.370 ;
        RECT 38.945 151.170 39.235 151.215 ;
        RECT 39.390 151.170 39.710 151.230 ;
        RECT 47.760 151.215 47.900 151.710 ;
        RECT 53.650 151.650 53.970 151.710 ;
        RECT 78.030 151.850 78.350 151.910 ;
        RECT 82.185 151.850 82.475 151.895 ;
        RECT 83.090 151.850 83.410 151.910 ;
        RECT 78.030 151.710 81.020 151.850 ;
        RECT 78.030 151.650 78.350 151.710 ;
        RECT 51.350 151.510 51.670 151.570 ;
        RECT 51.350 151.370 79.180 151.510 ;
        RECT 51.350 151.310 51.670 151.370 ;
        RECT 38.945 151.030 39.710 151.170 ;
        RECT 38.945 150.985 39.235 151.030 ;
        RECT 39.390 150.970 39.710 151.030 ;
        RECT 47.685 150.985 47.975 151.215 ;
        RECT 49.065 151.170 49.355 151.215 ;
        RECT 51.440 151.170 51.580 151.310 ;
        RECT 49.065 151.030 51.580 151.170 ;
        RECT 53.205 151.170 53.495 151.215 ;
        RECT 59.170 151.170 59.490 151.230 ;
        RECT 53.205 151.030 59.490 151.170 ;
        RECT 49.065 150.985 49.355 151.030 ;
        RECT 53.205 150.985 53.495 151.030 ;
        RECT 59.170 150.970 59.490 151.030 ;
        RECT 39.825 150.830 40.115 150.875 ;
        RECT 41.015 150.830 41.305 150.875 ;
        RECT 43.535 150.830 43.825 150.875 ;
        RECT 39.825 150.690 43.825 150.830 ;
        RECT 39.825 150.645 40.115 150.690 ;
        RECT 41.015 150.645 41.305 150.690 ;
        RECT 43.535 150.645 43.825 150.690 ;
        RECT 52.730 150.830 53.050 150.890 ;
        RECT 55.505 150.830 55.795 150.875 ;
        RECT 52.730 150.690 55.795 150.830 ;
        RECT 52.730 150.630 53.050 150.690 ;
        RECT 55.505 150.645 55.795 150.690 ;
        RECT 56.885 150.830 57.175 150.875 ;
        RECT 69.750 150.830 70.070 150.890 ;
        RECT 56.885 150.690 70.070 150.830 ;
        RECT 56.885 150.645 57.175 150.690 ;
        RECT 69.750 150.630 70.070 150.690 ;
        RECT 39.430 150.490 39.720 150.535 ;
        RECT 41.530 150.490 41.820 150.535 ;
        RECT 43.100 150.490 43.390 150.535 ;
        RECT 78.490 150.490 78.810 150.550 ;
        RECT 39.430 150.350 43.390 150.490 ;
        RECT 39.430 150.305 39.720 150.350 ;
        RECT 41.530 150.305 41.820 150.350 ;
        RECT 43.100 150.305 43.390 150.350 ;
        RECT 51.900 150.350 78.810 150.490 ;
        RECT 51.900 150.210 52.040 150.350 ;
        RECT 78.490 150.290 78.810 150.350 ;
        RECT 51.810 149.950 52.130 150.210 ;
        RECT 52.270 149.950 52.590 150.210 ;
        RECT 69.750 150.150 70.070 150.210 ;
        RECT 77.110 150.150 77.430 150.210 ;
        RECT 69.750 150.010 77.430 150.150 ;
        RECT 79.040 150.150 79.180 151.370 ;
        RECT 79.410 151.310 79.730 151.570 ;
        RECT 80.880 151.555 81.020 151.710 ;
        RECT 82.185 151.710 83.410 151.850 ;
        RECT 82.185 151.665 82.475 151.710 ;
        RECT 83.090 151.650 83.410 151.710 ;
        RECT 84.470 151.850 84.790 151.910 ;
        RECT 87.230 151.850 87.550 151.910 ;
        RECT 91.830 151.850 92.150 151.910 ;
        RECT 97.350 151.850 97.670 151.910 ;
        RECT 84.470 151.710 90.680 151.850 ;
        RECT 84.470 151.650 84.790 151.710 ;
        RECT 87.230 151.650 87.550 151.710 ;
        RECT 80.805 151.325 81.095 151.555 ;
        RECT 81.725 151.510 82.015 151.555 ;
        RECT 82.630 151.510 82.950 151.570 ;
        RECT 81.725 151.370 82.950 151.510 ;
        RECT 81.725 151.325 82.015 151.370 ;
        RECT 82.630 151.310 82.950 151.370 ;
        RECT 83.550 151.510 83.870 151.570 ;
        RECT 88.610 151.510 88.930 151.570 ;
        RECT 83.550 151.370 84.700 151.510 ;
        RECT 83.550 151.310 83.870 151.370 ;
        RECT 79.500 151.170 79.640 151.310 ;
        RECT 82.170 151.170 82.490 151.230 ;
        RECT 79.500 151.030 82.490 151.170 ;
        RECT 82.720 151.170 82.860 151.310 ;
        RECT 84.560 151.215 84.700 151.370 ;
        RECT 88.610 151.370 90.220 151.510 ;
        RECT 88.610 151.310 88.930 151.370 ;
        RECT 90.080 151.215 90.220 151.370 ;
        RECT 83.105 151.170 83.395 151.215 ;
        RECT 82.720 151.030 83.395 151.170 ;
        RECT 82.170 150.970 82.490 151.030 ;
        RECT 83.105 150.985 83.395 151.030 ;
        RECT 84.025 150.985 84.315 151.215 ;
        RECT 84.485 150.985 84.775 151.215 ;
        RECT 89.545 151.170 89.835 151.215 ;
        RECT 86.400 151.030 89.835 151.170 ;
        RECT 80.790 150.830 81.110 150.890 ;
        RECT 82.260 150.830 82.400 150.970 ;
        RECT 84.100 150.830 84.240 150.985 ;
        RECT 80.790 150.690 81.710 150.830 ;
        RECT 82.260 150.690 84.240 150.830 ;
        RECT 80.790 150.630 81.110 150.690 ;
        RECT 81.570 150.490 81.710 150.690 ;
        RECT 84.930 150.630 85.250 150.890 ;
        RECT 82.170 150.490 82.490 150.550 ;
        RECT 81.570 150.350 82.490 150.490 ;
        RECT 82.170 150.290 82.490 150.350 ;
        RECT 83.565 150.490 83.855 150.535 ;
        RECT 86.400 150.490 86.540 151.030 ;
        RECT 89.545 150.985 89.835 151.030 ;
        RECT 90.005 150.985 90.295 151.215 ;
        RECT 90.540 151.170 90.680 151.710 ;
        RECT 91.830 151.710 97.670 151.850 ;
        RECT 91.830 151.650 92.150 151.710 ;
        RECT 97.350 151.650 97.670 151.710 ;
        RECT 97.810 151.850 98.130 151.910 ;
        RECT 102.410 151.850 102.730 151.910 ;
        RECT 104.710 151.850 105.030 151.910 ;
        RECT 97.810 151.710 105.030 151.850 ;
        RECT 97.810 151.650 98.130 151.710 ;
        RECT 102.410 151.650 102.730 151.710 ;
        RECT 104.710 151.650 105.030 151.710 ;
        RECT 109.310 151.850 109.630 151.910 ;
        RECT 134.610 151.850 134.930 151.910 ;
        RECT 109.310 151.710 124.260 151.850 ;
        RECT 109.310 151.650 109.630 151.710 ;
        RECT 99.190 151.310 99.510 151.570 ;
        RECT 101.030 151.310 101.350 151.570 ;
        RECT 111.610 151.510 111.930 151.570 ;
        RECT 111.610 151.370 115.060 151.510 ;
        RECT 111.610 151.310 111.930 151.370 ;
        RECT 91.385 151.170 91.675 151.215 ;
        RECT 90.540 151.030 91.675 151.170 ;
        RECT 99.280 151.135 99.420 151.310 ;
        RECT 91.385 150.985 91.675 151.030 ;
        RECT 99.205 150.905 99.495 151.135 ;
        RECT 104.725 150.985 105.015 151.215 ;
        RECT 88.625 150.645 88.915 150.875 ;
        RECT 89.070 150.830 89.390 150.890 ;
        RECT 92.765 150.830 93.055 150.875 ;
        RECT 103.345 150.830 103.635 150.875 ;
        RECT 104.800 150.830 104.940 150.985 ;
        RECT 114.370 150.970 114.690 151.230 ;
        RECT 114.920 151.215 115.060 151.370 ;
        RECT 117.590 151.310 117.910 151.570 ;
        RECT 122.650 151.510 122.970 151.570 ;
        RECT 118.140 151.370 122.970 151.510 ;
        RECT 114.845 150.985 115.135 151.215 ;
        RECT 116.225 151.170 116.515 151.215 ;
        RECT 116.670 151.170 116.990 151.230 ;
        RECT 116.225 151.030 116.990 151.170 ;
        RECT 116.225 150.985 116.515 151.030 ;
        RECT 116.670 150.970 116.990 151.030 ;
        RECT 117.145 151.170 117.435 151.215 ;
        RECT 117.680 151.170 117.820 151.310 ;
        RECT 117.145 151.030 117.820 151.170 ;
        RECT 117.145 150.985 117.435 151.030 ;
        RECT 106.090 150.830 106.410 150.890 ;
        RECT 89.070 150.690 93.055 150.830 ;
        RECT 83.565 150.350 86.540 150.490 ;
        RECT 87.230 150.490 87.550 150.550 ;
        RECT 88.700 150.490 88.840 150.645 ;
        RECT 89.070 150.630 89.390 150.690 ;
        RECT 92.765 150.645 93.055 150.690 ;
        RECT 102.040 150.690 103.100 150.830 ;
        RECT 97.350 150.490 97.670 150.550 ;
        RECT 102.040 150.490 102.180 150.690 ;
        RECT 87.230 150.350 91.600 150.490 ;
        RECT 83.565 150.305 83.855 150.350 ;
        RECT 87.230 150.290 87.550 150.350 ;
        RECT 89.070 150.150 89.390 150.210 ;
        RECT 79.040 150.010 89.390 150.150 ;
        RECT 69.750 149.950 70.070 150.010 ;
        RECT 77.110 149.950 77.430 150.010 ;
        RECT 89.070 149.950 89.390 150.010 ;
        RECT 90.910 149.950 91.230 150.210 ;
        RECT 91.460 150.150 91.600 150.350 ;
        RECT 97.350 150.350 102.180 150.490 ;
        RECT 97.350 150.290 97.670 150.350 ;
        RECT 102.410 150.290 102.730 150.550 ;
        RECT 102.960 150.490 103.100 150.690 ;
        RECT 103.345 150.690 106.410 150.830 ;
        RECT 103.345 150.645 103.635 150.690 ;
        RECT 106.090 150.630 106.410 150.690 ;
        RECT 110.690 150.830 111.010 150.890 ;
        RECT 113.925 150.830 114.215 150.875 ;
        RECT 110.690 150.690 114.215 150.830 ;
        RECT 114.460 150.830 114.600 150.970 ;
        RECT 115.765 150.830 116.055 150.875 ;
        RECT 114.460 150.690 116.055 150.830 ;
        RECT 116.760 150.830 116.900 150.970 ;
        RECT 118.140 150.830 118.280 151.370 ;
        RECT 122.650 151.310 122.970 151.370 ;
        RECT 118.510 150.970 118.830 151.230 ;
        RECT 116.760 150.690 118.280 150.830 ;
        RECT 110.690 150.630 111.010 150.690 ;
        RECT 113.925 150.645 114.215 150.690 ;
        RECT 115.765 150.645 116.055 150.690 ;
        RECT 115.305 150.490 115.595 150.535 ;
        RECT 118.600 150.490 118.740 150.970 ;
        RECT 124.120 150.830 124.260 151.710 ;
        RECT 128.720 151.710 134.930 151.850 ;
        RECT 124.490 150.970 124.810 151.230 ;
        RECT 124.950 151.170 125.270 151.230 ;
        RECT 128.720 151.215 128.860 151.710 ;
        RECT 134.610 151.650 134.930 151.710 ;
        RECT 137.370 151.850 137.690 151.910 ;
        RECT 147.505 151.850 147.795 151.895 ;
        RECT 137.370 151.710 147.795 151.850 ;
        RECT 137.370 151.650 137.690 151.710 ;
        RECT 147.505 151.665 147.795 151.710 ;
        RECT 131.405 151.510 131.695 151.555 ;
        RECT 139.670 151.510 139.990 151.570 ;
        RECT 141.830 151.510 142.120 151.555 ;
        RECT 131.405 151.370 133.000 151.510 ;
        RECT 131.405 151.325 131.695 151.370 ;
        RECT 127.725 151.170 128.015 151.215 ;
        RECT 124.950 151.030 128.015 151.170 ;
        RECT 124.950 150.970 125.270 151.030 ;
        RECT 127.725 150.985 128.015 151.030 ;
        RECT 128.645 150.985 128.935 151.215 ;
        RECT 130.010 150.970 130.330 151.230 ;
        RECT 131.850 150.970 132.170 151.230 ;
        RECT 132.860 151.215 133.000 151.370 ;
        RECT 139.670 151.370 142.120 151.510 ;
        RECT 139.670 151.310 139.990 151.370 ;
        RECT 141.830 151.325 142.120 151.370 ;
        RECT 132.785 150.985 133.075 151.215 ;
        RECT 140.130 151.170 140.450 151.230 ;
        RECT 140.605 151.170 140.895 151.215 ;
        RECT 140.130 151.030 140.895 151.170 ;
        RECT 140.130 150.970 140.450 151.030 ;
        RECT 140.605 150.985 140.895 151.030 ;
        RECT 129.550 150.830 129.870 150.890 ;
        RECT 130.485 150.830 130.775 150.875 ;
        RECT 124.120 150.690 130.775 150.830 ;
        RECT 129.550 150.630 129.870 150.690 ;
        RECT 130.485 150.645 130.775 150.690 ;
        RECT 131.405 150.830 131.695 150.875 ;
        RECT 136.450 150.830 136.770 150.890 ;
        RECT 131.405 150.690 136.770 150.830 ;
        RECT 131.405 150.645 131.695 150.690 ;
        RECT 136.450 150.630 136.770 150.690 ;
        RECT 141.485 150.830 141.775 150.875 ;
        RECT 142.675 150.830 142.965 150.875 ;
        RECT 145.195 150.830 145.485 150.875 ;
        RECT 141.485 150.690 145.485 150.830 ;
        RECT 141.485 150.645 141.775 150.690 ;
        RECT 142.675 150.645 142.965 150.690 ;
        RECT 145.195 150.645 145.485 150.690 ;
        RECT 102.960 150.350 115.060 150.490 ;
        RECT 98.285 150.150 98.575 150.195 ;
        RECT 98.730 150.150 99.050 150.210 ;
        RECT 91.460 150.010 99.050 150.150 ;
        RECT 98.285 149.965 98.575 150.010 ;
        RECT 98.730 149.950 99.050 150.010 ;
        RECT 99.650 150.150 99.970 150.210 ;
        RECT 103.805 150.150 104.095 150.195 ;
        RECT 99.650 150.010 104.095 150.150 ;
        RECT 99.650 149.950 99.970 150.010 ;
        RECT 103.805 149.965 104.095 150.010 ;
        RECT 108.390 150.150 108.710 150.210 ;
        RECT 112.070 150.150 112.390 150.210 ;
        RECT 108.390 150.010 112.390 150.150 ;
        RECT 114.920 150.150 115.060 150.350 ;
        RECT 115.305 150.350 118.740 150.490 ;
        RECT 141.090 150.490 141.380 150.535 ;
        RECT 143.190 150.490 143.480 150.535 ;
        RECT 144.760 150.490 145.050 150.535 ;
        RECT 141.090 150.350 145.050 150.490 ;
        RECT 115.305 150.305 115.595 150.350 ;
        RECT 141.090 150.305 141.380 150.350 ;
        RECT 143.190 150.305 143.480 150.350 ;
        RECT 144.760 150.305 145.050 150.350 ;
        RECT 118.510 150.150 118.830 150.210 ;
        RECT 114.920 150.010 118.830 150.150 ;
        RECT 108.390 149.950 108.710 150.010 ;
        RECT 112.070 149.950 112.390 150.010 ;
        RECT 118.510 149.950 118.830 150.010 ;
        RECT 124.965 150.150 125.255 150.195 ;
        RECT 125.410 150.150 125.730 150.210 ;
        RECT 124.965 150.010 125.730 150.150 ;
        RECT 124.965 149.965 125.255 150.010 ;
        RECT 125.410 149.950 125.730 150.010 ;
        RECT 132.770 149.950 133.090 150.210 ;
        RECT 29.970 148.770 33.130 149.430 ;
        RECT 36.100 149.330 150.180 149.810 ;
        RECT 52.730 148.930 53.050 149.190 ;
        RECT 54.110 148.930 54.430 149.190 ;
        RECT 63.785 149.130 64.075 149.175 ;
        RECT 76.650 149.130 76.970 149.190 ;
        RECT 78.045 149.130 78.335 149.175 ;
        RECT 63.785 148.990 73.660 149.130 ;
        RECT 63.785 148.945 64.075 148.990 ;
        RECT 38.470 148.790 38.790 148.850 ;
        RECT 41.705 148.790 41.995 148.835 ;
        RECT 29.970 24.230 30.630 148.770 ;
        RECT 38.470 148.650 41.995 148.790 ;
        RECT 38.470 148.590 38.790 148.650 ;
        RECT 41.705 148.605 41.995 148.650 ;
        RECT 50.890 148.450 51.210 148.510 ;
        RECT 41.320 148.310 51.210 148.450 ;
        RECT 41.320 148.155 41.460 148.310 ;
        RECT 50.890 148.250 51.210 148.310 ;
        RECT 52.285 148.450 52.575 148.495 ;
        RECT 52.820 148.450 52.960 148.930 ;
        RECT 54.200 148.790 54.340 148.930 ;
        RECT 52.285 148.310 52.960 148.450 ;
        RECT 53.280 148.650 54.340 148.790 ;
        RECT 67.005 148.790 67.295 148.835 ;
        RECT 69.305 148.790 69.595 148.835 ;
        RECT 67.005 148.650 69.060 148.790 ;
        RECT 52.285 148.265 52.575 148.310 ;
        RECT 41.245 147.925 41.535 148.155 ;
        RECT 42.625 148.110 42.915 148.155 ;
        RECT 45.370 148.110 45.690 148.170 ;
        RECT 53.280 148.155 53.420 148.650 ;
        RECT 67.005 148.605 67.295 148.650 ;
        RECT 54.125 148.450 54.415 148.495 ;
        RECT 56.885 148.450 57.175 148.495 ;
        RECT 57.805 148.450 58.095 148.495 ;
        RECT 54.125 148.310 56.180 148.450 ;
        RECT 54.125 148.265 54.415 148.310 ;
        RECT 56.040 148.155 56.180 148.310 ;
        RECT 56.885 148.310 58.095 148.450 ;
        RECT 56.885 148.265 57.175 148.310 ;
        RECT 57.805 148.265 58.095 148.310 ;
        RECT 60.105 148.450 60.395 148.495 ;
        RECT 68.920 148.450 69.060 148.650 ;
        RECT 69.305 148.650 73.200 148.790 ;
        RECT 69.305 148.605 69.595 148.650 ;
        RECT 73.060 148.495 73.200 148.650 ;
        RECT 70.685 148.450 70.975 148.495 ;
        RECT 72.525 148.450 72.815 148.495 ;
        RECT 60.105 148.310 63.080 148.450 ;
        RECT 60.105 148.265 60.395 148.310 ;
        RECT 42.625 147.970 45.690 148.110 ;
        RECT 42.625 147.925 42.915 147.970 ;
        RECT 45.370 147.910 45.690 147.970 ;
        RECT 53.205 147.925 53.495 148.155 ;
        RECT 54.585 147.925 54.875 148.155 ;
        RECT 55.965 147.925 56.255 148.155 ;
        RECT 54.660 147.490 54.800 147.925 ;
        RECT 55.030 147.570 55.350 147.830 ;
        RECT 57.880 147.770 58.020 148.265 ;
        RECT 58.250 148.110 58.570 148.170 ;
        RECT 62.940 148.155 63.080 148.310 ;
        RECT 68.920 148.310 70.440 148.450 ;
        RECT 60.565 148.110 60.855 148.155 ;
        RECT 58.250 147.970 60.855 148.110 ;
        RECT 58.250 147.910 58.570 147.970 ;
        RECT 60.565 147.925 60.855 147.970 ;
        RECT 62.865 148.110 63.155 148.155 ;
        RECT 66.085 148.110 66.375 148.155 ;
        RECT 68.370 148.110 68.690 148.170 ;
        RECT 68.920 148.155 69.060 148.310 ;
        RECT 70.300 148.155 70.440 148.310 ;
        RECT 70.685 148.310 72.815 148.450 ;
        RECT 70.685 148.265 70.975 148.310 ;
        RECT 72.525 148.265 72.815 148.310 ;
        RECT 72.985 148.265 73.275 148.495 ;
        RECT 73.520 148.450 73.660 148.990 ;
        RECT 76.650 148.990 78.335 149.130 ;
        RECT 76.650 148.930 76.970 148.990 ;
        RECT 78.045 148.945 78.335 148.990 ;
        RECT 78.950 149.130 79.270 149.190 ;
        RECT 80.345 149.130 80.635 149.175 ;
        RECT 83.550 149.130 83.870 149.190 ;
        RECT 78.950 148.990 83.870 149.130 ;
        RECT 78.950 148.930 79.270 148.990 ;
        RECT 80.345 148.945 80.635 148.990 ;
        RECT 83.550 148.930 83.870 148.990 ;
        RECT 89.070 149.130 89.390 149.190 ;
        RECT 126.790 149.130 127.110 149.190 ;
        RECT 127.710 149.130 128.030 149.190 ;
        RECT 89.070 148.990 124.260 149.130 ;
        RECT 89.070 148.930 89.390 148.990 ;
        RECT 123.585 148.790 123.875 148.835 ;
        RECT 76.280 148.650 78.720 148.790 ;
        RECT 76.280 148.495 76.420 148.650 ;
        RECT 78.580 148.495 78.720 148.650 ;
        RECT 81.570 148.650 123.875 148.790 ;
        RECT 124.120 148.790 124.260 148.990 ;
        RECT 126.790 148.990 128.030 149.130 ;
        RECT 126.790 148.930 127.110 148.990 ;
        RECT 127.710 148.930 128.030 148.990 ;
        RECT 141.970 148.930 142.290 149.190 ;
        RECT 124.120 148.650 140.820 148.790 ;
        RECT 75.745 148.450 76.035 148.495 ;
        RECT 73.520 148.310 76.035 148.450 ;
        RECT 75.745 148.265 76.035 148.310 ;
        RECT 76.205 148.265 76.495 148.495 ;
        RECT 78.505 148.450 78.795 148.495 ;
        RECT 81.570 148.450 81.710 148.650 ;
        RECT 123.585 148.605 123.875 148.650 ;
        RECT 82.630 148.450 82.950 148.510 ;
        RECT 84.470 148.450 84.790 148.510 ;
        RECT 76.740 148.310 77.800 148.450 ;
        RECT 62.865 147.970 66.375 148.110 ;
        RECT 62.865 147.925 63.155 147.970 ;
        RECT 66.085 147.925 66.375 147.970 ;
        RECT 67.540 147.970 68.690 148.110 ;
        RECT 61.255 147.770 61.545 147.815 ;
        RECT 57.880 147.630 61.545 147.770 ;
        RECT 61.255 147.585 61.545 147.630 ;
        RECT 61.930 147.570 62.250 147.830 ;
        RECT 62.405 147.770 62.695 147.815 ;
        RECT 67.540 147.770 67.680 147.970 ;
        RECT 68.370 147.910 68.690 147.970 ;
        RECT 68.845 147.925 69.135 148.155 ;
        RECT 69.765 147.925 70.055 148.155 ;
        RECT 70.225 147.925 70.515 148.155 ;
        RECT 69.840 147.770 69.980 147.925 ;
        RECT 62.405 147.630 67.680 147.770 ;
        RECT 68.000 147.630 69.980 147.770 ;
        RECT 70.300 147.770 70.440 147.925 ;
        RECT 71.130 147.910 71.450 148.170 ;
        RECT 72.050 147.910 72.370 148.170 ;
        RECT 73.445 147.925 73.735 148.155 ;
        RECT 74.810 148.110 75.130 148.170 ;
        RECT 76.740 148.155 76.880 148.310 ;
        RECT 76.665 148.110 76.955 148.155 ;
        RECT 74.810 147.970 76.955 148.110 ;
        RECT 72.510 147.770 72.830 147.830 ;
        RECT 73.515 147.770 73.655 147.925 ;
        RECT 74.810 147.910 75.130 147.970 ;
        RECT 76.665 147.925 76.955 147.970 ;
        RECT 77.125 147.925 77.415 148.155 ;
        RECT 77.660 148.110 77.800 148.310 ;
        RECT 78.505 148.310 82.400 148.450 ;
        RECT 78.505 148.265 78.795 148.310 ;
        RECT 82.260 148.155 82.400 148.310 ;
        RECT 82.630 148.310 84.790 148.450 ;
        RECT 82.630 148.250 82.950 148.310 ;
        RECT 84.470 148.250 84.790 148.310 ;
        RECT 84.930 148.450 85.250 148.510 ;
        RECT 85.405 148.450 85.695 148.495 ;
        RECT 84.930 148.310 85.695 148.450 ;
        RECT 84.930 148.250 85.250 148.310 ;
        RECT 85.405 148.265 85.695 148.310 ;
        RECT 86.325 148.450 86.615 148.495 ;
        RECT 88.610 148.450 88.930 148.510 ;
        RECT 95.065 148.450 95.355 148.495 ;
        RECT 98.270 148.450 98.590 148.510 ;
        RECT 86.325 148.310 88.930 148.450 ;
        RECT 86.325 148.265 86.615 148.310 ;
        RECT 88.610 148.250 88.930 148.310 ;
        RECT 89.160 148.310 95.355 148.450 ;
        RECT 89.160 148.170 89.300 148.310 ;
        RECT 95.065 148.265 95.355 148.310 ;
        RECT 95.600 148.310 98.590 148.450 ;
        RECT 79.425 148.110 79.715 148.155 ;
        RECT 81.265 148.110 81.555 148.155 ;
        RECT 77.660 147.970 81.555 148.110 ;
        RECT 79.425 147.925 79.715 147.970 ;
        RECT 81.265 147.925 81.555 147.970 ;
        RECT 82.185 147.925 82.475 148.155 ;
        RECT 83.105 148.110 83.395 148.155 ;
        RECT 85.865 148.110 86.155 148.155 ;
        RECT 83.105 147.970 86.155 148.110 ;
        RECT 83.105 147.925 83.395 147.970 ;
        RECT 85.865 147.925 86.155 147.970 ;
        RECT 86.785 148.110 87.075 148.155 ;
        RECT 87.230 148.110 87.550 148.170 ;
        RECT 86.785 147.970 87.550 148.110 ;
        RECT 86.785 147.925 87.075 147.970 ;
        RECT 70.300 147.630 71.820 147.770 ;
        RECT 62.405 147.585 62.695 147.630 ;
        RECT 68.000 147.490 68.140 147.630 ;
        RECT 71.680 147.490 71.820 147.630 ;
        RECT 72.510 147.630 73.655 147.770 ;
        RECT 75.270 147.770 75.590 147.830 ;
        RECT 77.200 147.770 77.340 147.925 ;
        RECT 87.230 147.910 87.550 147.970 ;
        RECT 89.070 147.910 89.390 148.170 ;
        RECT 89.530 147.910 89.850 148.170 ;
        RECT 89.990 147.910 90.310 148.170 ;
        RECT 90.910 147.910 91.230 148.170 ;
        RECT 95.600 148.155 95.740 148.310 ;
        RECT 98.270 148.250 98.590 148.310 ;
        RECT 102.410 148.450 102.730 148.510 ;
        RECT 108.390 148.450 108.710 148.510 ;
        RECT 102.410 148.310 108.710 148.450 ;
        RECT 102.410 148.250 102.730 148.310 ;
        RECT 108.390 148.250 108.710 148.310 ;
        RECT 110.690 148.450 111.010 148.510 ;
        RECT 113.910 148.450 114.230 148.510 ;
        RECT 114.845 148.450 115.135 148.495 ;
        RECT 110.690 148.310 112.300 148.450 ;
        RECT 110.690 148.250 111.010 148.310 ;
        RECT 94.605 147.925 94.895 148.155 ;
        RECT 95.525 147.925 95.815 148.155 ;
        RECT 98.730 148.110 99.050 148.170 ;
        RECT 112.160 148.155 112.300 148.310 ;
        RECT 113.910 148.310 115.135 148.450 ;
        RECT 113.910 148.250 114.230 148.310 ;
        RECT 114.845 148.265 115.135 148.310 ;
        RECT 115.305 148.450 115.595 148.495 ;
        RECT 118.065 148.450 118.355 148.495 ;
        RECT 115.305 148.310 118.355 148.450 ;
        RECT 115.305 148.265 115.595 148.310 ;
        RECT 118.065 148.265 118.355 148.310 ;
        RECT 118.510 148.450 118.830 148.510 ;
        RECT 136.925 148.450 137.215 148.495 ;
        RECT 139.685 148.450 139.975 148.495 ;
        RECT 118.510 148.310 137.215 148.450 ;
        RECT 118.510 148.250 118.830 148.310 ;
        RECT 136.925 148.265 137.215 148.310 ;
        RECT 137.920 148.310 139.975 148.450 ;
        RECT 111.625 148.110 111.915 148.155 ;
        RECT 98.730 147.970 111.915 148.110 ;
        RECT 91.370 147.770 91.690 147.830 ;
        RECT 75.270 147.630 77.340 147.770 ;
        RECT 84.560 147.630 91.690 147.770 ;
        RECT 94.680 147.770 94.820 147.925 ;
        RECT 98.730 147.910 99.050 147.970 ;
        RECT 111.625 147.925 111.915 147.970 ;
        RECT 112.085 147.925 112.375 148.155 ;
        RECT 112.530 147.910 112.850 148.170 ;
        RECT 112.990 148.110 113.310 148.170 ;
        RECT 113.465 148.110 113.755 148.155 ;
        RECT 112.990 147.970 113.755 148.110 ;
        RECT 112.990 147.910 113.310 147.970 ;
        RECT 113.465 147.925 113.755 147.970 ;
        RECT 114.385 147.925 114.675 148.155 ;
        RECT 115.765 147.925 116.055 148.155 ;
        RECT 117.130 148.110 117.450 148.170 ;
        RECT 118.985 148.110 119.275 148.155 ;
        RECT 120.325 148.120 120.615 148.165 ;
        RECT 119.980 148.110 120.615 148.120 ;
        RECT 117.130 147.980 120.615 148.110 ;
        RECT 117.130 147.970 120.120 147.980 ;
        RECT 98.820 147.770 98.960 147.910 ;
        RECT 94.680 147.630 98.960 147.770 ;
        RECT 99.650 147.770 99.970 147.830 ;
        RECT 101.965 147.770 102.255 147.815 ;
        RECT 103.330 147.770 103.650 147.830 ;
        RECT 99.650 147.630 103.650 147.770 ;
        RECT 72.510 147.570 72.830 147.630 ;
        RECT 75.270 147.570 75.590 147.630 ;
        RECT 38.930 147.430 39.250 147.490 ;
        RECT 40.325 147.430 40.615 147.475 ;
        RECT 38.930 147.290 40.615 147.430 ;
        RECT 38.930 147.230 39.250 147.290 ;
        RECT 40.325 147.245 40.615 147.290 ;
        RECT 54.570 147.230 54.890 147.490 ;
        RECT 67.910 147.230 68.230 147.490 ;
        RECT 71.590 147.230 71.910 147.490 ;
        RECT 72.050 147.430 72.370 147.490 ;
        RECT 73.890 147.430 74.210 147.490 ;
        RECT 72.050 147.290 74.210 147.430 ;
        RECT 72.050 147.230 72.370 147.290 ;
        RECT 73.890 147.230 74.210 147.290 ;
        RECT 74.365 147.430 74.655 147.475 ;
        RECT 77.110 147.430 77.430 147.490 ;
        RECT 84.560 147.475 84.700 147.630 ;
        RECT 91.370 147.570 91.690 147.630 ;
        RECT 99.650 147.570 99.970 147.630 ;
        RECT 101.965 147.585 102.255 147.630 ;
        RECT 103.330 147.570 103.650 147.630 ;
        RECT 106.090 147.770 106.410 147.830 ;
        RECT 109.770 147.770 110.090 147.830 ;
        RECT 114.460 147.770 114.600 147.925 ;
        RECT 106.090 147.630 109.540 147.770 ;
        RECT 106.090 147.570 106.410 147.630 ;
        RECT 109.400 147.490 109.540 147.630 ;
        RECT 109.770 147.630 114.600 147.770 ;
        RECT 115.840 147.770 115.980 147.925 ;
        RECT 117.130 147.910 117.450 147.970 ;
        RECT 118.985 147.925 119.275 147.970 ;
        RECT 120.325 147.935 120.615 147.980 ;
        RECT 121.285 148.110 121.575 148.155 ;
        RECT 121.285 147.970 121.960 148.110 ;
        RECT 121.285 147.925 121.575 147.970 ;
        RECT 119.905 147.770 120.195 147.815 ;
        RECT 121.820 147.770 121.960 147.970 ;
        RECT 122.650 147.910 122.970 148.170 ;
        RECT 137.920 148.155 138.060 148.310 ;
        RECT 139.685 148.265 139.975 148.310 ;
        RECT 140.680 148.155 140.820 148.650 ;
        RECT 141.525 148.450 141.815 148.495 ;
        RECT 142.060 148.450 142.200 148.930 ;
        RECT 144.270 148.590 144.590 148.850 ;
        RECT 143.810 148.450 144.130 148.510 ;
        RECT 141.525 148.310 142.200 148.450 ;
        RECT 142.520 148.310 144.130 148.450 ;
        RECT 141.525 148.265 141.815 148.310 ;
        RECT 123.585 147.925 123.875 148.155 ;
        RECT 129.105 148.110 129.395 148.155 ;
        RECT 129.105 147.970 130.240 148.110 ;
        RECT 129.105 147.925 129.395 147.970 ;
        RECT 123.660 147.770 123.800 147.925 ;
        RECT 115.840 147.630 117.360 147.770 ;
        RECT 109.770 147.570 110.090 147.630 ;
        RECT 74.365 147.290 77.430 147.430 ;
        RECT 74.365 147.245 74.655 147.290 ;
        RECT 77.110 147.230 77.430 147.290 ;
        RECT 84.485 147.245 84.775 147.475 ;
        RECT 84.930 147.430 85.250 147.490 ;
        RECT 87.705 147.430 87.995 147.475 ;
        RECT 84.930 147.290 87.995 147.430 ;
        RECT 84.930 147.230 85.250 147.290 ;
        RECT 87.705 147.245 87.995 147.290 ;
        RECT 88.610 147.430 88.930 147.490 ;
        RECT 99.205 147.430 99.495 147.475 ;
        RECT 88.610 147.290 99.495 147.430 ;
        RECT 88.610 147.230 88.930 147.290 ;
        RECT 99.205 147.245 99.495 147.290 ;
        RECT 100.570 147.430 100.890 147.490 ;
        RECT 101.505 147.430 101.795 147.475 ;
        RECT 100.570 147.290 101.795 147.430 ;
        RECT 100.570 147.230 100.890 147.290 ;
        RECT 101.505 147.245 101.795 147.290 ;
        RECT 106.550 147.430 106.870 147.490 ;
        RECT 108.390 147.430 108.710 147.490 ;
        RECT 106.550 147.290 108.710 147.430 ;
        RECT 106.550 147.230 106.870 147.290 ;
        RECT 108.390 147.230 108.710 147.290 ;
        RECT 109.310 147.230 109.630 147.490 ;
        RECT 110.230 147.230 110.550 147.490 ;
        RECT 110.690 147.430 111.010 147.490 ;
        RECT 116.685 147.430 116.975 147.475 ;
        RECT 110.690 147.290 116.975 147.430 ;
        RECT 117.220 147.430 117.360 147.630 ;
        RECT 119.905 147.630 123.800 147.770 ;
        RECT 119.905 147.585 120.195 147.630 ;
        RECT 123.660 147.490 123.800 147.630 ;
        RECT 125.425 147.770 125.715 147.815 ;
        RECT 125.425 147.630 127.020 147.770 ;
        RECT 125.425 147.585 125.715 147.630 ;
        RECT 120.365 147.430 120.655 147.475 ;
        RECT 117.220 147.290 120.655 147.430 ;
        RECT 110.690 147.230 111.010 147.290 ;
        RECT 116.685 147.245 116.975 147.290 ;
        RECT 120.365 147.245 120.655 147.290 ;
        RECT 123.570 147.230 123.890 147.490 ;
        RECT 126.880 147.475 127.020 147.630 ;
        RECT 130.100 147.490 130.240 147.970 ;
        RECT 137.845 147.925 138.135 148.155 ;
        RECT 139.225 147.925 139.515 148.155 ;
        RECT 140.605 147.925 140.895 148.155 ;
        RECT 139.300 147.770 139.440 147.925 ;
        RECT 142.520 147.770 142.660 148.310 ;
        RECT 143.810 148.250 144.130 148.310 ;
        RECT 142.890 147.910 143.210 148.170 ;
        RECT 144.360 148.125 144.500 148.590 ;
        RECT 144.325 147.895 144.615 148.125 ;
        RECT 139.300 147.630 142.660 147.770 ;
        RECT 126.805 147.245 127.095 147.475 ;
        RECT 130.010 147.230 130.330 147.490 ;
        RECT 138.750 147.430 139.070 147.490 ;
        RECT 143.825 147.430 144.115 147.475 ;
        RECT 138.750 147.290 144.115 147.430 ;
        RECT 138.750 147.230 139.070 147.290 ;
        RECT 143.825 147.245 144.115 147.290 ;
        RECT 36.100 146.610 150.180 147.090 ;
        RECT 38.930 146.210 39.250 146.470 ;
        RECT 39.390 146.210 39.710 146.470 ;
        RECT 51.810 146.410 52.130 146.470 ;
        RECT 43.160 146.270 52.130 146.410 ;
        RECT 39.020 145.730 39.160 146.210 ;
        RECT 39.480 146.070 39.620 146.210 ;
        RECT 43.160 146.115 43.300 146.270 ;
        RECT 51.810 146.210 52.130 146.270 ;
        RECT 52.270 146.210 52.590 146.470 ;
        RECT 52.730 146.210 53.050 146.470 ;
        RECT 54.110 146.410 54.430 146.470 ;
        RECT 55.965 146.410 56.255 146.455 ;
        RECT 54.110 146.270 56.255 146.410 ;
        RECT 54.110 146.210 54.430 146.270 ;
        RECT 55.965 146.225 56.255 146.270 ;
        RECT 67.910 146.410 68.230 146.470 ;
        RECT 72.065 146.410 72.355 146.455 ;
        RECT 72.510 146.410 72.830 146.470 ;
        RECT 67.910 146.270 70.900 146.410 ;
        RECT 67.910 146.210 68.230 146.270 ;
        RECT 39.480 145.930 40.080 146.070 ;
        RECT 39.405 145.730 39.695 145.775 ;
        RECT 39.020 145.590 39.695 145.730 ;
        RECT 39.405 145.545 39.695 145.590 ;
        RECT 39.940 145.390 40.080 145.930 ;
        RECT 43.085 145.885 43.375 146.115 ;
        RECT 45.800 146.070 46.090 146.115 ;
        RECT 52.360 146.070 52.500 146.210 ;
        RECT 45.800 145.930 52.500 146.070 ;
        RECT 45.800 145.885 46.090 145.930 ;
        RECT 52.820 145.775 52.960 146.210 ;
        RECT 61.930 146.070 62.250 146.130 ;
        RECT 61.930 145.930 69.520 146.070 ;
        RECT 61.930 145.870 62.250 145.930 ;
        RECT 52.745 145.730 53.035 145.775 ;
        RECT 55.045 145.730 55.335 145.775 ;
        RECT 51.440 145.590 53.035 145.730 ;
        RECT 44.465 145.390 44.755 145.435 ;
        RECT 39.940 145.250 44.755 145.390 ;
        RECT 44.465 145.205 44.755 145.250 ;
        RECT 45.345 145.390 45.635 145.435 ;
        RECT 46.535 145.390 46.825 145.435 ;
        RECT 49.055 145.390 49.345 145.435 ;
        RECT 45.345 145.250 49.345 145.390 ;
        RECT 45.345 145.205 45.635 145.250 ;
        RECT 46.535 145.205 46.825 145.250 ;
        RECT 49.055 145.205 49.345 145.250 ;
        RECT 42.150 144.850 42.470 145.110 ;
        RECT 51.440 145.095 51.580 145.590 ;
        RECT 52.745 145.545 53.035 145.590 ;
        RECT 54.200 145.590 55.335 145.730 ;
        RECT 54.200 145.450 54.340 145.590 ;
        RECT 55.045 145.545 55.335 145.590 ;
        RECT 58.265 145.730 58.555 145.775 ;
        RECT 60.550 145.730 60.870 145.790 ;
        RECT 58.265 145.590 60.870 145.730 ;
        RECT 58.265 145.545 58.555 145.590 ;
        RECT 60.550 145.530 60.870 145.590 ;
        RECT 53.205 145.390 53.495 145.435 ;
        RECT 54.110 145.390 54.430 145.450 ;
        RECT 53.205 145.250 54.430 145.390 ;
        RECT 53.205 145.205 53.495 145.250 ;
        RECT 54.110 145.190 54.430 145.250 ;
        RECT 54.570 145.390 54.890 145.450 ;
        RECT 57.805 145.390 58.095 145.435 ;
        RECT 54.570 145.250 58.095 145.390 ;
        RECT 54.570 145.190 54.890 145.250 ;
        RECT 57.805 145.205 58.095 145.250 ;
        RECT 44.950 145.050 45.240 145.095 ;
        RECT 47.050 145.050 47.340 145.095 ;
        RECT 48.620 145.050 48.910 145.095 ;
        RECT 44.950 144.910 48.910 145.050 ;
        RECT 44.950 144.865 45.240 144.910 ;
        RECT 47.050 144.865 47.340 144.910 ;
        RECT 48.620 144.865 48.910 144.910 ;
        RECT 51.365 144.865 51.655 145.095 ;
        RECT 60.105 145.050 60.395 145.095 ;
        RECT 62.020 145.050 62.160 145.870 ;
        RECT 65.240 145.775 65.380 145.930 ;
        RECT 65.165 145.545 65.455 145.775 ;
        RECT 65.625 145.730 65.915 145.775 ;
        RECT 66.545 145.730 66.835 145.775 ;
        RECT 67.910 145.730 68.230 145.790 ;
        RECT 65.625 145.590 66.300 145.730 ;
        RECT 65.625 145.545 65.915 145.590 ;
        RECT 66.160 145.390 66.300 145.590 ;
        RECT 66.545 145.590 68.230 145.730 ;
        RECT 66.545 145.545 66.835 145.590 ;
        RECT 67.910 145.530 68.230 145.590 ;
        RECT 68.370 145.530 68.690 145.790 ;
        RECT 69.380 145.775 69.520 145.930 ;
        RECT 69.750 145.870 70.070 146.130 ;
        RECT 68.845 145.545 69.135 145.775 ;
        RECT 69.305 145.545 69.595 145.775 ;
        RECT 69.840 145.730 69.980 145.870 ;
        RECT 70.225 145.730 70.515 145.775 ;
        RECT 69.840 145.590 70.515 145.730 ;
        RECT 70.760 145.730 70.900 146.270 ;
        RECT 72.065 146.270 72.830 146.410 ;
        RECT 72.065 146.225 72.355 146.270 ;
        RECT 72.510 146.210 72.830 146.270 ;
        RECT 78.490 146.210 78.810 146.470 ;
        RECT 82.630 146.410 82.950 146.470 ;
        RECT 87.690 146.410 88.010 146.470 ;
        RECT 79.040 146.270 82.950 146.410 ;
        RECT 79.040 146.070 79.180 146.270 ;
        RECT 82.630 146.210 82.950 146.270 ;
        RECT 83.180 146.270 88.010 146.410 ;
        RECT 83.180 146.070 83.320 146.270 ;
        RECT 87.690 146.210 88.010 146.270 ;
        RECT 89.070 146.210 89.390 146.470 ;
        RECT 99.650 146.410 99.970 146.470 ;
        RECT 95.370 146.270 99.970 146.410 ;
        RECT 74.440 145.930 79.180 146.070 ;
        RECT 79.500 145.930 83.320 146.070 ;
        RECT 74.440 145.775 74.580 145.930 ;
        RECT 72.985 145.730 73.275 145.775 ;
        RECT 70.760 145.590 73.275 145.730 ;
        RECT 70.225 145.545 70.515 145.590 ;
        RECT 72.985 145.545 73.275 145.590 ;
        RECT 74.365 145.545 74.655 145.775 ;
        RECT 68.460 145.390 68.600 145.530 ;
        RECT 66.160 145.250 68.600 145.390 ;
        RECT 68.920 145.390 69.060 145.545 ;
        RECT 75.270 145.530 75.590 145.790 ;
        RECT 76.190 145.530 76.510 145.790 ;
        RECT 79.500 145.775 79.640 145.930 ;
        RECT 79.425 145.545 79.715 145.775 ;
        RECT 80.330 145.530 80.650 145.790 ;
        RECT 80.790 145.530 81.110 145.790 ;
        RECT 83.180 145.775 83.320 145.930 ;
        RECT 85.480 145.930 88.380 146.070 ;
        RECT 83.105 145.545 83.395 145.775 ;
        RECT 84.010 145.530 84.330 145.790 ;
        RECT 85.480 145.775 85.620 145.930 ;
        RECT 88.240 145.790 88.380 145.930 ;
        RECT 85.405 145.545 85.695 145.775 ;
        RECT 86.325 145.545 86.615 145.775 ;
        RECT 69.765 145.390 70.055 145.435 ;
        RECT 68.920 145.250 70.055 145.390 ;
        RECT 69.765 145.205 70.055 145.250 ;
        RECT 71.130 145.190 71.450 145.450 ;
        RECT 71.590 145.390 71.910 145.450 ;
        RECT 73.905 145.390 74.195 145.435 ;
        RECT 75.360 145.390 75.500 145.530 ;
        RECT 71.590 145.250 75.500 145.390 ;
        RECT 77.585 145.390 77.875 145.435 ;
        RECT 80.880 145.390 81.020 145.530 ;
        RECT 77.585 145.250 81.020 145.390 ;
        RECT 82.170 145.390 82.490 145.450 ;
        RECT 84.485 145.390 84.775 145.435 ;
        RECT 84.945 145.390 85.235 145.435 ;
        RECT 85.850 145.390 86.170 145.450 ;
        RECT 82.170 145.250 86.170 145.390 ;
        RECT 86.400 145.390 86.540 145.545 ;
        RECT 88.150 145.530 88.470 145.790 ;
        RECT 89.160 145.730 89.300 146.210 ;
        RECT 95.370 146.070 95.510 146.270 ;
        RECT 99.650 146.210 99.970 146.270 ;
        RECT 101.030 146.410 101.350 146.470 ;
        RECT 110.690 146.410 111.010 146.470 ;
        RECT 101.030 146.270 111.010 146.410 ;
        RECT 101.030 146.210 101.350 146.270 ;
        RECT 110.690 146.210 111.010 146.270 ;
        RECT 111.610 146.410 111.930 146.470 ;
        RECT 118.970 146.410 119.290 146.470 ;
        RECT 111.610 146.270 117.820 146.410 ;
        RECT 111.610 146.210 111.930 146.270 ;
        RECT 103.330 146.070 103.650 146.130 ;
        RECT 91.000 145.930 95.740 146.070 ;
        RECT 90.005 145.730 90.295 145.775 ;
        RECT 89.160 145.590 90.295 145.730 ;
        RECT 90.005 145.545 90.295 145.590 ;
        RECT 90.450 145.530 90.770 145.790 ;
        RECT 91.000 145.775 91.140 145.930 ;
        RECT 90.925 145.545 91.215 145.775 ;
        RECT 91.370 145.730 91.690 145.790 ;
        RECT 91.845 145.730 92.135 145.775 ;
        RECT 91.370 145.590 92.135 145.730 ;
        RECT 91.370 145.530 91.690 145.590 ;
        RECT 91.845 145.545 92.135 145.590 ;
        RECT 94.590 145.530 94.910 145.790 ;
        RECT 95.600 145.775 95.740 145.930 ;
        RECT 103.330 145.930 104.940 146.070 ;
        RECT 103.330 145.870 103.650 145.930 ;
        RECT 95.525 145.545 95.815 145.775 ;
        RECT 99.205 145.730 99.495 145.775 ;
        RECT 101.965 145.730 102.255 145.775 ;
        RECT 102.410 145.730 102.730 145.790 ;
        RECT 99.205 145.590 102.730 145.730 ;
        RECT 99.205 145.545 99.495 145.590 ;
        RECT 101.965 145.545 102.255 145.590 ;
        RECT 102.410 145.530 102.730 145.590 ;
        RECT 102.885 145.730 103.175 145.775 ;
        RECT 103.790 145.730 104.110 145.790 ;
        RECT 104.800 145.775 104.940 145.930 ;
        RECT 106.180 145.930 113.220 146.070 ;
        RECT 106.180 145.775 106.320 145.930 ;
        RECT 113.080 145.790 113.220 145.930 ;
        RECT 102.885 145.590 104.110 145.730 ;
        RECT 102.885 145.545 103.175 145.590 ;
        RECT 103.790 145.530 104.110 145.590 ;
        RECT 104.725 145.545 105.015 145.775 ;
        RECT 106.105 145.545 106.395 145.775 ;
        RECT 107.010 145.530 107.330 145.790 ;
        RECT 107.930 145.530 108.250 145.790 ;
        RECT 109.310 145.530 109.630 145.790 ;
        RECT 111.150 145.530 111.470 145.790 ;
        RECT 112.070 145.530 112.390 145.790 ;
        RECT 112.990 145.530 113.310 145.790 ;
        RECT 114.370 145.530 114.690 145.790 ;
        RECT 115.290 145.530 115.610 145.790 ;
        RECT 117.130 145.530 117.450 145.790 ;
        RECT 117.680 145.730 117.820 146.270 ;
        RECT 118.970 146.270 122.420 146.410 ;
        RECT 118.970 146.210 119.290 146.270 ;
        RECT 118.600 145.930 121.960 146.070 ;
        RECT 118.065 145.730 118.355 145.775 ;
        RECT 118.600 145.730 118.740 145.930 ;
        RECT 121.820 145.790 121.960 145.930 ;
        RECT 117.680 145.590 118.740 145.730 ;
        RECT 118.065 145.545 118.355 145.590 ;
        RECT 119.430 145.530 119.750 145.790 ;
        RECT 120.350 145.730 120.670 145.790 ;
        RECT 121.285 145.730 121.575 145.775 ;
        RECT 120.350 145.590 121.575 145.730 ;
        RECT 120.350 145.530 120.670 145.590 ;
        RECT 121.285 145.545 121.575 145.590 ;
        RECT 121.730 145.530 122.050 145.790 ;
        RECT 122.280 145.775 122.420 146.270 ;
        RECT 132.770 146.210 133.090 146.470 ;
        RECT 145.190 146.410 145.510 146.470 ;
        RECT 146.585 146.410 146.875 146.455 ;
        RECT 145.190 146.270 146.875 146.410 ;
        RECT 145.190 146.210 145.510 146.270 ;
        RECT 146.585 146.225 146.875 146.270 ;
        RECT 123.570 145.870 123.890 146.130 ;
        RECT 122.205 145.545 122.495 145.775 ;
        RECT 125.425 145.730 125.715 145.775 ;
        RECT 128.185 145.730 128.475 145.775 ;
        RECT 130.010 145.730 130.330 145.790 ;
        RECT 132.310 145.730 132.630 145.790 ;
        RECT 125.425 145.590 132.630 145.730 ;
        RECT 132.860 145.730 133.000 146.210 ;
        RECT 143.810 145.870 144.130 146.130 ;
        RECT 133.145 145.730 133.435 145.775 ;
        RECT 140.130 145.730 140.450 145.790 ;
        RECT 140.620 145.775 140.880 145.820 ;
        RECT 132.860 145.590 133.435 145.730 ;
        RECT 125.425 145.545 125.715 145.590 ;
        RECT 128.185 145.545 128.475 145.590 ;
        RECT 130.010 145.530 130.330 145.590 ;
        RECT 132.310 145.530 132.630 145.590 ;
        RECT 133.145 145.545 133.435 145.590 ;
        RECT 137.000 145.590 140.450 145.730 ;
        RECT 94.145 145.390 94.435 145.435 ;
        RECT 96.890 145.390 97.210 145.450 ;
        RECT 100.570 145.390 100.890 145.450 ;
        RECT 86.400 145.250 90.220 145.390 ;
        RECT 71.590 145.190 71.910 145.250 ;
        RECT 73.905 145.205 74.195 145.250 ;
        RECT 77.585 145.205 77.875 145.250 ;
        RECT 82.170 145.190 82.490 145.250 ;
        RECT 84.485 145.205 84.775 145.250 ;
        RECT 84.945 145.205 85.235 145.250 ;
        RECT 85.850 145.190 86.170 145.250 ;
        RECT 60.105 144.910 62.160 145.050 ;
        RECT 71.220 145.050 71.360 145.190 ;
        RECT 90.080 145.110 90.220 145.250 ;
        RECT 91.460 145.250 95.510 145.390 ;
        RECT 73.445 145.050 73.735 145.095 ;
        RECT 71.220 144.910 73.735 145.050 ;
        RECT 60.105 144.865 60.395 144.910 ;
        RECT 73.445 144.865 73.735 144.910 ;
        RECT 74.350 145.050 74.670 145.110 ;
        RECT 88.625 145.050 88.915 145.095 ;
        RECT 74.350 144.910 88.915 145.050 ;
        RECT 74.350 144.850 74.670 144.910 ;
        RECT 88.625 144.865 88.915 144.910 ;
        RECT 89.990 144.850 90.310 145.110 ;
        RECT 91.460 144.770 91.600 145.250 ;
        RECT 94.145 145.205 94.435 145.250 ;
        RECT 95.370 145.050 95.510 145.250 ;
        RECT 96.890 145.250 100.890 145.390 ;
        RECT 96.890 145.190 97.210 145.250 ;
        RECT 100.570 145.190 100.890 145.250 ;
        RECT 103.345 145.390 103.635 145.435 ;
        RECT 107.485 145.390 107.775 145.435 ;
        RECT 110.705 145.390 110.995 145.435 ;
        RECT 113.910 145.390 114.230 145.450 ;
        RECT 116.685 145.390 116.975 145.435 ;
        RECT 120.825 145.390 121.115 145.435 ;
        RECT 126.790 145.390 127.110 145.450 ;
        RECT 103.345 145.250 107.775 145.390 ;
        RECT 103.345 145.205 103.635 145.250 ;
        RECT 107.485 145.205 107.775 145.250 ;
        RECT 110.320 145.250 116.975 145.390 ;
        RECT 103.420 145.050 103.560 145.205 ;
        RECT 110.320 145.095 110.460 145.250 ;
        RECT 110.705 145.205 110.995 145.250 ;
        RECT 113.910 145.190 114.230 145.250 ;
        RECT 116.685 145.205 116.975 145.250 ;
        RECT 117.220 145.250 127.110 145.390 ;
        RECT 103.805 145.050 104.095 145.095 ;
        RECT 95.370 144.910 104.095 145.050 ;
        RECT 103.805 144.865 104.095 144.910 ;
        RECT 110.245 144.865 110.535 145.095 ;
        RECT 112.070 145.050 112.390 145.110 ;
        RECT 117.220 145.050 117.360 145.250 ;
        RECT 120.825 145.205 121.115 145.250 ;
        RECT 126.790 145.190 127.110 145.250 ;
        RECT 127.710 145.190 128.030 145.450 ;
        RECT 131.865 145.205 132.155 145.435 ;
        RECT 132.745 145.390 133.035 145.435 ;
        RECT 133.935 145.390 134.225 145.435 ;
        RECT 136.455 145.390 136.745 145.435 ;
        RECT 132.745 145.250 136.745 145.390 ;
        RECT 132.745 145.205 133.035 145.250 ;
        RECT 133.935 145.205 134.225 145.250 ;
        RECT 136.455 145.205 136.745 145.250 ;
        RECT 112.070 144.910 117.360 145.050 ;
        RECT 118.985 145.050 119.275 145.095 ;
        RECT 128.630 145.050 128.950 145.110 ;
        RECT 118.985 144.910 128.950 145.050 ;
        RECT 112.070 144.850 112.390 144.910 ;
        RECT 118.985 144.865 119.275 144.910 ;
        RECT 128.630 144.850 128.950 144.910 ;
        RECT 33.410 144.710 33.730 144.770 ;
        RECT 38.025 144.710 38.315 144.755 ;
        RECT 33.410 144.570 38.315 144.710 ;
        RECT 33.410 144.510 33.730 144.570 ;
        RECT 38.025 144.525 38.315 144.570 ;
        RECT 68.845 144.710 69.135 144.755 ;
        RECT 74.810 144.710 75.130 144.770 ;
        RECT 68.845 144.570 75.130 144.710 ;
        RECT 68.845 144.525 69.135 144.570 ;
        RECT 74.810 144.510 75.130 144.570 ;
        RECT 75.270 144.510 75.590 144.770 ;
        RECT 77.110 144.510 77.430 144.770 ;
        RECT 82.170 144.510 82.490 144.770 ;
        RECT 87.230 144.510 87.550 144.770 ;
        RECT 91.370 144.510 91.690 144.770 ;
        RECT 96.430 144.510 96.750 144.770 ;
        RECT 98.270 144.510 98.590 144.770 ;
        RECT 100.125 144.710 100.415 144.755 ;
        RECT 100.570 144.710 100.890 144.770 ;
        RECT 100.125 144.570 100.890 144.710 ;
        RECT 100.125 144.525 100.415 144.570 ;
        RECT 100.570 144.510 100.890 144.570 ;
        RECT 101.045 144.710 101.335 144.755 ;
        RECT 102.410 144.710 102.730 144.770 ;
        RECT 101.045 144.570 102.730 144.710 ;
        RECT 101.045 144.525 101.335 144.570 ;
        RECT 102.410 144.510 102.730 144.570 ;
        RECT 105.170 144.510 105.490 144.770 ;
        RECT 108.850 144.510 109.170 144.770 ;
        RECT 112.990 144.510 113.310 144.770 ;
        RECT 116.210 144.510 116.530 144.770 ;
        RECT 120.350 144.510 120.670 144.770 ;
        RECT 123.110 144.510 123.430 144.770 ;
        RECT 128.185 144.710 128.475 144.755 ;
        RECT 129.105 144.710 129.395 144.755 ;
        RECT 128.185 144.570 129.395 144.710 ;
        RECT 131.940 144.710 132.080 145.205 ;
        RECT 132.350 145.050 132.640 145.095 ;
        RECT 134.450 145.050 134.740 145.095 ;
        RECT 136.020 145.050 136.310 145.095 ;
        RECT 132.350 144.910 136.310 145.050 ;
        RECT 132.350 144.865 132.640 144.910 ;
        RECT 134.450 144.865 134.740 144.910 ;
        RECT 136.020 144.865 136.310 144.910 ;
        RECT 137.000 144.710 137.140 145.590 ;
        RECT 140.130 145.530 140.450 145.590 ;
        RECT 140.605 145.730 140.895 145.775 ;
        RECT 143.365 145.730 143.655 145.775 ;
        RECT 145.665 145.730 145.955 145.775 ;
        RECT 140.605 145.590 143.655 145.730 ;
        RECT 140.605 145.545 140.895 145.590 ;
        RECT 143.365 145.545 143.655 145.590 ;
        RECT 143.900 145.590 145.955 145.730 ;
        RECT 140.620 145.500 140.880 145.545 ;
        RECT 141.065 145.390 141.355 145.435 ;
        RECT 142.890 145.390 143.210 145.450 ;
        RECT 143.900 145.390 144.040 145.590 ;
        RECT 145.665 145.545 145.955 145.590 ;
        RECT 141.065 145.250 143.210 145.390 ;
        RECT 141.065 145.205 141.355 145.250 ;
        RECT 138.765 145.050 139.055 145.095 ;
        RECT 141.140 145.050 141.280 145.205 ;
        RECT 142.890 145.190 143.210 145.250 ;
        RECT 143.670 145.250 144.040 145.390 ;
        RECT 138.765 144.910 141.280 145.050 ;
        RECT 141.510 145.050 141.830 145.110 ;
        RECT 143.670 145.050 143.810 145.250 ;
        RECT 141.510 144.910 143.810 145.050 ;
        RECT 138.765 144.865 139.055 144.910 ;
        RECT 141.510 144.850 141.830 144.910 ;
        RECT 131.940 144.570 137.140 144.710 ;
        RECT 139.685 144.710 139.975 144.755 ;
        RECT 140.605 144.710 140.895 144.755 ;
        RECT 139.685 144.570 140.895 144.710 ;
        RECT 128.185 144.525 128.475 144.570 ;
        RECT 129.105 144.525 129.395 144.570 ;
        RECT 139.685 144.525 139.975 144.570 ;
        RECT 140.605 144.525 140.895 144.570 ;
        RECT 36.100 143.890 150.180 144.370 ;
        RECT 39.390 143.490 39.710 143.750 ;
        RECT 47.225 143.690 47.515 143.735 ;
        RECT 54.110 143.690 54.430 143.750 ;
        RECT 47.225 143.550 54.430 143.690 ;
        RECT 47.225 143.505 47.515 143.550 ;
        RECT 54.110 143.490 54.430 143.550 ;
        RECT 74.900 143.550 81.940 143.690 ;
        RECT 39.480 143.010 39.620 143.490 ;
        RECT 40.810 143.350 41.100 143.395 ;
        RECT 42.910 143.350 43.200 143.395 ;
        RECT 44.480 143.350 44.770 143.395 ;
        RECT 74.350 143.350 74.670 143.410 ;
        RECT 40.810 143.210 44.770 143.350 ;
        RECT 40.810 143.165 41.100 143.210 ;
        RECT 42.910 143.165 43.200 143.210 ;
        RECT 44.480 143.165 44.770 143.210 ;
        RECT 56.040 143.210 74.670 143.350 ;
        RECT 40.325 143.010 40.615 143.055 ;
        RECT 39.480 142.870 40.615 143.010 ;
        RECT 40.325 142.825 40.615 142.870 ;
        RECT 41.205 143.010 41.495 143.055 ;
        RECT 42.395 143.010 42.685 143.055 ;
        RECT 44.915 143.010 45.205 143.055 ;
        RECT 41.205 142.870 45.205 143.010 ;
        RECT 41.205 142.825 41.495 142.870 ;
        RECT 42.395 142.825 42.685 142.870 ;
        RECT 44.915 142.825 45.205 142.870 ;
        RECT 38.470 142.670 38.790 142.730 ;
        RECT 56.040 142.715 56.180 143.210 ;
        RECT 74.350 143.150 74.670 143.210 ;
        RECT 74.900 143.010 75.040 143.550 ;
        RECT 75.270 143.150 75.590 143.410 ;
        RECT 78.505 143.165 78.795 143.395 ;
        RECT 60.180 142.870 75.040 143.010 ;
        RECT 60.180 142.715 60.320 142.870 ;
        RECT 39.405 142.670 39.695 142.715 ;
        RECT 38.470 142.530 39.695 142.670 ;
        RECT 38.470 142.470 38.790 142.530 ;
        RECT 39.405 142.485 39.695 142.530 ;
        RECT 50.905 142.670 51.195 142.715 ;
        RECT 50.905 142.530 55.720 142.670 ;
        RECT 50.905 142.485 51.195 142.530 ;
        RECT 41.660 142.330 41.950 142.375 ;
        RECT 42.610 142.330 42.930 142.390 ;
        RECT 41.660 142.190 42.930 142.330 ;
        RECT 41.660 142.145 41.950 142.190 ;
        RECT 42.610 142.130 42.930 142.190 ;
        RECT 45.830 142.330 46.150 142.390 ;
        RECT 51.365 142.330 51.655 142.375 ;
        RECT 45.830 142.190 51.655 142.330 ;
        RECT 45.830 142.130 46.150 142.190 ;
        RECT 51.365 142.145 51.655 142.190 ;
        RECT 53.205 142.145 53.495 142.375 ;
        RECT 55.580 142.330 55.720 142.530 ;
        RECT 55.965 142.485 56.255 142.715 ;
        RECT 60.105 142.485 60.395 142.715 ;
        RECT 64.230 142.470 64.550 142.730 ;
        RECT 75.360 142.330 75.500 143.150 ;
        RECT 76.665 142.485 76.955 142.715 ;
        RECT 55.580 142.190 75.500 142.330 ;
        RECT 76.740 142.330 76.880 142.485 ;
        RECT 77.570 142.470 77.890 142.730 ;
        RECT 78.580 142.670 78.720 143.165 ;
        RECT 79.425 142.670 79.715 142.715 ;
        RECT 78.580 142.530 79.715 142.670 ;
        RECT 79.425 142.485 79.715 142.530 ;
        RECT 81.800 142.330 81.940 143.550 ;
        RECT 82.170 143.490 82.490 143.750 ;
        RECT 87.230 143.490 87.550 143.750 ;
        RECT 91.845 143.690 92.135 143.735 ;
        RECT 93.670 143.690 93.990 143.750 ;
        RECT 91.845 143.550 93.990 143.690 ;
        RECT 91.845 143.505 92.135 143.550 ;
        RECT 93.670 143.490 93.990 143.550 ;
        RECT 96.430 143.490 96.750 143.750 ;
        RECT 98.270 143.490 98.590 143.750 ;
        RECT 105.170 143.490 105.490 143.750 ;
        RECT 108.390 143.690 108.710 143.750 ;
        RECT 112.070 143.690 112.390 143.750 ;
        RECT 108.390 143.550 112.390 143.690 ;
        RECT 108.390 143.490 108.710 143.550 ;
        RECT 112.070 143.490 112.390 143.550 ;
        RECT 112.990 143.490 113.310 143.750 ;
        RECT 113.450 143.690 113.770 143.750 ;
        RECT 114.385 143.690 114.675 143.735 ;
        RECT 113.450 143.550 114.675 143.690 ;
        RECT 113.450 143.490 113.770 143.550 ;
        RECT 114.385 143.505 114.675 143.550 ;
        RECT 121.270 143.690 121.590 143.750 ;
        RECT 127.265 143.690 127.555 143.735 ;
        RECT 121.270 143.550 127.555 143.690 ;
        RECT 121.270 143.490 121.590 143.550 ;
        RECT 127.265 143.505 127.555 143.550 ;
        RECT 132.310 143.690 132.630 143.750 ;
        RECT 142.425 143.690 142.715 143.735 ;
        RECT 143.345 143.690 143.635 143.735 ;
        RECT 132.310 143.550 140.360 143.690 ;
        RECT 132.310 143.490 132.630 143.550 ;
        RECT 82.260 143.010 82.400 143.490 ;
        RECT 82.260 142.870 83.780 143.010 ;
        RECT 82.170 142.470 82.490 142.730 ;
        RECT 83.640 142.715 83.780 142.870 ;
        RECT 83.565 142.485 83.855 142.715 ;
        RECT 87.320 142.670 87.460 143.490 ;
        RECT 91.370 142.810 91.690 143.070 ;
        RECT 88.625 142.670 88.915 142.715 ;
        RECT 87.320 142.530 88.915 142.670 ;
        RECT 88.625 142.485 88.915 142.530 ;
        RECT 90.910 142.670 91.230 142.730 ;
        RECT 92.765 142.670 93.055 142.715 ;
        RECT 90.910 142.530 93.055 142.670 ;
        RECT 90.910 142.470 91.230 142.530 ;
        RECT 92.765 142.485 93.055 142.530 ;
        RECT 93.685 142.670 93.975 142.715 ;
        RECT 94.145 142.670 94.435 142.715 ;
        RECT 93.685 142.530 94.435 142.670 ;
        RECT 96.520 142.670 96.660 143.490 ;
        RECT 97.365 142.670 97.655 142.715 ;
        RECT 96.520 142.530 97.655 142.670 ;
        RECT 93.685 142.485 93.975 142.530 ;
        RECT 94.145 142.485 94.435 142.530 ;
        RECT 97.365 142.485 97.655 142.530 ;
        RECT 98.360 142.330 98.500 143.490 ;
        RECT 101.045 142.670 101.335 142.715 ;
        RECT 102.410 142.670 102.730 142.730 ;
        RECT 101.045 142.530 102.730 142.670 ;
        RECT 105.260 142.670 105.400 143.490 ;
        RECT 113.080 143.350 113.220 143.490 ;
        RECT 113.080 143.210 138.060 143.350 ;
        RECT 108.940 142.870 116.900 143.010 ;
        RECT 108.940 142.730 109.080 142.870 ;
        RECT 105.645 142.670 105.935 142.715 ;
        RECT 105.260 142.530 105.935 142.670 ;
        RECT 101.045 142.485 101.335 142.530 ;
        RECT 102.410 142.470 102.730 142.530 ;
        RECT 105.645 142.485 105.935 142.530 ;
        RECT 108.850 142.470 109.170 142.730 ;
        RECT 112.530 142.470 112.850 142.730 ;
        RECT 113.910 142.470 114.230 142.730 ;
        RECT 115.305 142.485 115.595 142.715 ;
        RECT 76.740 142.190 81.480 142.330 ;
        RECT 81.800 142.190 98.500 142.330 ;
        RECT 112.620 142.330 112.760 142.470 ;
        RECT 115.380 142.330 115.520 142.485 ;
        RECT 116.210 142.470 116.530 142.730 ;
        RECT 116.760 142.715 116.900 142.870 ;
        RECT 123.110 142.810 123.430 143.070 ;
        RECT 126.790 142.810 127.110 143.070 ;
        RECT 128.630 143.010 128.950 143.070 ;
        RECT 128.630 142.870 137.600 143.010 ;
        RECT 128.630 142.810 128.950 142.870 ;
        RECT 116.685 142.485 116.975 142.715 ;
        RECT 120.350 142.670 120.670 142.730 ;
        RECT 120.825 142.670 121.115 142.715 ;
        RECT 120.350 142.530 121.115 142.670 ;
        RECT 123.200 142.670 123.340 142.810 ;
        RECT 124.505 142.670 124.795 142.715 ;
        RECT 123.200 142.530 124.795 142.670 ;
        RECT 120.350 142.470 120.670 142.530 ;
        RECT 120.825 142.485 121.115 142.530 ;
        RECT 124.505 142.485 124.795 142.530 ;
        RECT 128.170 142.470 128.490 142.730 ;
        RECT 137.460 142.715 137.600 142.870 ;
        RECT 133.245 142.670 133.535 142.715 ;
        RECT 128.720 142.530 133.535 142.670 ;
        RECT 112.620 142.190 115.520 142.330 ;
        RECT 116.300 142.330 116.440 142.470 ;
        RECT 128.720 142.330 128.860 142.530 ;
        RECT 133.245 142.485 133.535 142.530 ;
        RECT 137.385 142.485 137.675 142.715 ;
        RECT 116.300 142.190 128.860 142.330 ;
        RECT 129.105 142.330 129.395 142.375 ;
        RECT 130.025 142.330 130.315 142.375 ;
        RECT 129.105 142.190 130.315 142.330 ;
        RECT 137.920 142.330 138.060 143.210 ;
        RECT 140.220 143.055 140.360 143.550 ;
        RECT 142.425 143.550 143.635 143.690 ;
        RECT 142.425 143.505 142.715 143.550 ;
        RECT 143.345 143.505 143.635 143.550 ;
        RECT 140.145 142.825 140.435 143.055 ;
        RECT 143.810 142.810 144.130 143.070 ;
        RECT 144.270 142.470 144.590 142.730 ;
        RECT 146.125 142.485 146.415 142.715 ;
        RECT 146.200 142.330 146.340 142.485 ;
        RECT 137.920 142.190 146.340 142.330 ;
        RECT 38.470 141.790 38.790 142.050 ;
        RECT 49.970 141.790 50.290 142.050 ;
        RECT 53.280 141.990 53.420 142.145 ;
        RECT 53.650 141.990 53.970 142.050 ;
        RECT 53.280 141.850 53.970 141.990 ;
        RECT 53.650 141.790 53.970 141.850 ;
        RECT 55.030 141.790 55.350 142.050 ;
        RECT 59.170 141.790 59.490 142.050 ;
        RECT 63.310 141.790 63.630 142.050 ;
        RECT 75.730 141.790 76.050 142.050 ;
        RECT 78.950 141.990 79.270 142.050 ;
        RECT 81.340 142.035 81.480 142.190 ;
        RECT 129.105 142.145 129.395 142.190 ;
        RECT 130.025 142.145 130.315 142.190 ;
        RECT 80.345 141.990 80.635 142.035 ;
        RECT 78.950 141.850 80.635 141.990 ;
        RECT 78.950 141.790 79.270 141.850 ;
        RECT 80.345 141.805 80.635 141.850 ;
        RECT 81.265 141.805 81.555 142.035 ;
        RECT 83.090 141.990 83.410 142.050 ;
        RECT 84.485 141.990 84.775 142.035 ;
        RECT 83.090 141.850 84.775 141.990 ;
        RECT 83.090 141.790 83.410 141.850 ;
        RECT 84.485 141.805 84.775 141.850 ;
        RECT 89.070 141.790 89.390 142.050 ;
        RECT 91.370 141.990 91.690 142.050 ;
        RECT 95.065 141.990 95.355 142.035 ;
        RECT 91.370 141.850 95.355 141.990 ;
        RECT 91.370 141.790 91.690 141.850 ;
        RECT 95.065 141.805 95.355 141.850 ;
        RECT 96.430 141.790 96.750 142.050 ;
        RECT 99.650 141.990 99.970 142.050 ;
        RECT 101.965 141.990 102.255 142.035 ;
        RECT 99.650 141.850 102.255 141.990 ;
        RECT 99.650 141.790 99.970 141.850 ;
        RECT 101.965 141.805 102.255 141.850 ;
        RECT 104.710 141.790 105.030 142.050 ;
        RECT 116.225 141.990 116.515 142.035 ;
        RECT 117.130 141.990 117.450 142.050 ;
        RECT 116.225 141.850 117.450 141.990 ;
        RECT 116.225 141.805 116.515 141.850 ;
        RECT 117.130 141.790 117.450 141.850 ;
        RECT 117.590 141.790 117.910 142.050 ;
        RECT 120.350 141.990 120.670 142.050 ;
        RECT 121.745 141.990 122.035 142.035 ;
        RECT 120.350 141.850 122.035 141.990 ;
        RECT 120.350 141.790 120.670 141.850 ;
        RECT 121.745 141.805 122.035 141.850 ;
        RECT 125.410 141.790 125.730 142.050 ;
        RECT 128.630 141.990 128.950 142.050 ;
        RECT 130.485 141.990 130.775 142.035 ;
        RECT 128.630 141.850 130.775 141.990 ;
        RECT 128.630 141.790 128.950 141.850 ;
        RECT 130.485 141.805 130.775 141.850 ;
        RECT 132.770 141.990 133.090 142.050 ;
        RECT 134.165 141.990 134.455 142.035 ;
        RECT 132.770 141.850 134.455 141.990 ;
        RECT 132.770 141.790 133.090 141.850 ;
        RECT 134.165 141.805 134.455 141.850 ;
        RECT 136.910 141.990 137.230 142.050 ;
        RECT 138.305 141.990 138.595 142.035 ;
        RECT 136.910 141.850 138.595 141.990 ;
        RECT 136.910 141.790 137.230 141.850 ;
        RECT 138.305 141.805 138.595 141.850 ;
        RECT 141.050 141.990 141.370 142.050 ;
        RECT 147.045 141.990 147.335 142.035 ;
        RECT 141.050 141.850 147.335 141.990 ;
        RECT 141.050 141.790 141.370 141.850 ;
        RECT 147.045 141.805 147.335 141.850 ;
        RECT 36.100 141.170 150.180 141.650 ;
        RECT 141.510 140.970 141.830 141.030 ;
        RECT 127.800 140.830 141.830 140.970 ;
        RECT 60.550 140.630 60.870 140.690 ;
        RECT 117.130 140.630 117.450 140.690 ;
        RECT 127.800 140.630 127.940 140.830 ;
        RECT 141.510 140.770 141.830 140.830 ;
        RECT 60.550 140.490 116.900 140.630 ;
        RECT 60.550 140.430 60.870 140.490 ;
        RECT 64.230 140.290 64.550 140.350 ;
        RECT 110.230 140.290 110.550 140.350 ;
        RECT 64.230 140.150 110.550 140.290 ;
        RECT 116.760 140.290 116.900 140.490 ;
        RECT 117.130 140.490 127.940 140.630 ;
        RECT 117.130 140.430 117.450 140.490 ;
        RECT 124.030 140.290 124.350 140.350 ;
        RECT 116.760 140.150 124.350 140.290 ;
        RECT 64.230 140.090 64.550 140.150 ;
        RECT 110.230 140.090 110.550 140.150 ;
        RECT 124.030 140.090 124.350 140.150 ;
        RECT 53.650 139.950 53.970 140.010 ;
        RECT 84.470 139.950 84.790 140.010 ;
        RECT 96.890 139.950 97.210 140.010 ;
        RECT 53.650 139.810 84.790 139.950 ;
        RECT 53.650 139.750 53.970 139.810 ;
        RECT 84.470 139.750 84.790 139.810 ;
        RECT 92.840 139.810 97.210 139.950 ;
        RECT 80.790 139.610 81.110 139.670 ;
        RECT 92.840 139.610 92.980 139.810 ;
        RECT 96.890 139.750 97.210 139.810 ;
        RECT 80.790 139.470 92.980 139.610 ;
        RECT 80.790 139.410 81.110 139.470 ;
        RECT 33.430 132.440 33.710 132.470 ;
        RECT 37.570 132.440 37.850 132.470 ;
        RECT 41.710 132.440 41.990 132.470 ;
        RECT 45.850 132.440 46.130 132.470 ;
        RECT 49.990 132.440 50.270 132.470 ;
        RECT 54.130 132.440 54.410 132.470 ;
        RECT 58.270 132.440 58.550 132.470 ;
        RECT 62.410 132.440 62.690 132.470 ;
        RECT 74.830 132.440 75.110 132.470 ;
        RECT 78.970 132.440 79.250 132.470 ;
        RECT 83.110 132.440 83.390 132.470 ;
        RECT 87.250 132.440 87.530 132.470 ;
        RECT 91.390 132.440 91.670 132.470 ;
        RECT 95.530 132.440 95.810 132.470 ;
        RECT 116.230 132.440 116.510 132.470 ;
        RECT 120.370 132.440 120.650 132.470 ;
        RECT 124.510 132.440 124.790 132.470 ;
        RECT 128.650 132.440 128.930 132.470 ;
        RECT 33.430 132.160 35.240 132.440 ;
        RECT 33.430 132.130 33.710 132.160 ;
        RECT 34.960 130.830 35.240 132.160 ;
        RECT 37.570 132.160 39.240 132.440 ;
        RECT 37.570 132.130 37.850 132.160 ;
        RECT 38.960 130.830 39.240 132.160 ;
        RECT 41.710 132.160 43.240 132.440 ;
        RECT 41.710 132.130 41.990 132.160 ;
        RECT 42.960 130.830 43.240 132.160 ;
        RECT 45.850 132.160 47.240 132.440 ;
        RECT 45.850 132.130 46.130 132.160 ;
        RECT 46.960 130.830 47.240 132.160 ;
        RECT 49.990 132.160 51.240 132.440 ;
        RECT 49.990 132.130 50.270 132.160 ;
        RECT 50.960 130.830 51.240 132.160 ;
        RECT 54.130 132.160 55.240 132.440 ;
        RECT 54.130 132.130 54.410 132.160 ;
        RECT 54.960 130.830 55.240 132.160 ;
        RECT 58.270 132.160 59.240 132.440 ;
        RECT 58.270 132.130 58.550 132.160 ;
        RECT 58.960 130.830 59.240 132.160 ;
        RECT 34.580 126.330 35.580 130.830 ;
        RECT 38.580 126.330 39.580 130.830 ;
        RECT 42.580 126.330 43.580 130.830 ;
        RECT 46.580 126.330 47.580 130.830 ;
        RECT 50.580 126.330 51.580 130.830 ;
        RECT 54.580 126.330 55.580 130.830 ;
        RECT 58.580 126.330 59.580 130.830 ;
        RECT 34.810 125.865 35.400 126.330 ;
        RECT 38.810 125.865 39.400 126.330 ;
        RECT 42.810 125.865 43.400 126.330 ;
        RECT 46.810 125.865 47.400 126.330 ;
        RECT 50.810 125.865 51.400 126.330 ;
        RECT 54.810 125.865 55.400 126.330 ;
        RECT 58.810 125.865 59.400 126.330 ;
        RECT 60.580 105.110 61.580 132.330 ;
        RECT 62.410 132.160 63.240 132.440 ;
        RECT 62.410 132.130 62.690 132.160 ;
        RECT 62.960 130.830 63.240 132.160 ;
        RECT 62.580 126.330 63.580 130.830 ;
        RECT 62.810 125.865 63.400 126.330 ;
        RECT 60.580 105.080 61.600 105.110 ;
        RECT 33.900 104.080 64.410 105.080 ;
        RECT 60.600 104.050 61.600 104.080 ;
        RECT 34.810 85.650 35.400 86.075 ;
        RECT 38.810 85.650 39.400 86.075 ;
        RECT 42.810 85.650 43.400 86.075 ;
        RECT 46.810 85.650 47.400 86.075 ;
        RECT 50.810 85.650 51.400 86.075 ;
        RECT 54.810 85.650 55.400 86.075 ;
        RECT 58.810 85.650 59.400 86.075 ;
        RECT 62.810 85.650 63.400 86.075 ;
        RECT 34.580 82.530 35.580 85.650 ;
        RECT 33.000 82.330 35.580 82.530 ;
        RECT 32.070 81.530 35.580 82.330 ;
        RECT 32.070 81.465 34.130 81.530 ;
        RECT 32.070 52.530 32.935 81.465 ;
        RECT 34.580 78.430 35.580 81.530 ;
        RECT 38.580 79.430 39.580 85.650 ;
        RECT 42.580 79.430 43.580 85.650 ;
        RECT 46.580 79.430 47.580 85.650 ;
        RECT 50.580 79.430 51.580 85.650 ;
        RECT 54.580 79.430 55.580 85.650 ;
        RECT 58.580 79.430 59.580 85.650 ;
        RECT 62.580 79.430 63.580 85.650 ;
        RECT 36.630 78.430 39.610 79.430 ;
        RECT 40.630 78.430 43.610 79.430 ;
        RECT 44.630 78.430 47.610 79.430 ;
        RECT 48.630 78.430 51.610 79.430 ;
        RECT 52.630 78.430 55.610 79.430 ;
        RECT 56.630 78.430 59.610 79.430 ;
        RECT 60.630 78.430 63.610 79.430 ;
        RECT 34.810 77.865 35.400 78.430 ;
        RECT 34.810 57.940 35.400 58.425 ;
        RECT 36.630 57.940 37.630 78.430 ;
        RECT 38.810 77.865 39.400 78.430 ;
        RECT 38.810 57.940 39.400 58.425 ;
        RECT 40.630 57.940 41.630 78.430 ;
        RECT 42.810 77.865 43.400 78.430 ;
        RECT 42.810 57.940 43.400 58.425 ;
        RECT 44.630 57.940 45.630 78.430 ;
        RECT 46.810 77.865 47.400 78.430 ;
        RECT 46.810 57.940 47.400 58.425 ;
        RECT 48.630 57.940 49.630 78.430 ;
        RECT 50.810 77.865 51.400 78.430 ;
        RECT 50.810 57.940 51.400 58.425 ;
        RECT 52.630 57.940 53.630 78.430 ;
        RECT 54.810 77.865 55.400 78.430 ;
        RECT 54.810 57.940 55.400 58.425 ;
        RECT 56.630 57.940 57.630 78.430 ;
        RECT 58.810 77.865 59.400 78.430 ;
        RECT 58.810 57.940 59.400 58.425 ;
        RECT 60.630 57.940 61.630 78.430 ;
        RECT 62.810 77.865 63.400 78.430 ;
        RECT 34.490 56.940 37.630 57.940 ;
        RECT 38.490 56.940 41.630 57.940 ;
        RECT 42.490 56.940 45.630 57.940 ;
        RECT 46.490 56.940 49.630 57.940 ;
        RECT 50.490 56.940 53.630 57.940 ;
        RECT 54.490 56.940 57.630 57.940 ;
        RECT 58.490 56.940 61.630 57.940 ;
        RECT 62.810 57.930 63.400 58.425 ;
        RECT 64.930 57.930 65.930 132.330 ;
        RECT 74.830 132.160 76.240 132.440 ;
        RECT 74.830 132.130 75.110 132.160 ;
        RECT 75.960 130.830 76.240 132.160 ;
        RECT 78.970 132.160 80.240 132.440 ;
        RECT 78.970 132.130 79.250 132.160 ;
        RECT 79.960 130.830 80.240 132.160 ;
        RECT 83.110 132.160 84.240 132.440 ;
        RECT 83.110 132.130 83.390 132.160 ;
        RECT 83.960 130.830 84.240 132.160 ;
        RECT 87.250 132.160 88.240 132.440 ;
        RECT 87.250 132.130 87.530 132.160 ;
        RECT 87.960 130.830 88.240 132.160 ;
        RECT 91.390 132.160 92.240 132.440 ;
        RECT 91.390 132.130 91.670 132.160 ;
        RECT 91.960 130.830 92.240 132.160 ;
        RECT 95.530 132.160 96.340 132.440 ;
        RECT 99.640 132.160 100.340 132.440 ;
        RECT 95.530 132.130 95.810 132.160 ;
        RECT 96.060 130.830 96.340 132.160 ;
        RECT 100.060 130.830 100.340 132.160 ;
        RECT 75.580 126.330 76.580 130.830 ;
        RECT 79.580 126.330 80.580 130.830 ;
        RECT 83.580 126.330 84.580 130.830 ;
        RECT 87.580 126.330 88.580 130.830 ;
        RECT 91.580 126.330 92.580 130.830 ;
        RECT 95.580 126.330 96.580 130.830 ;
        RECT 99.580 126.330 100.580 130.830 ;
        RECT 75.810 125.865 76.400 126.330 ;
        RECT 79.810 125.865 80.400 126.330 ;
        RECT 83.810 125.865 84.400 126.330 ;
        RECT 87.810 125.865 88.400 126.330 ;
        RECT 91.810 125.865 92.400 126.330 ;
        RECT 95.810 125.865 96.400 126.330 ;
        RECT 99.810 125.865 100.400 126.330 ;
        RECT 101.580 105.110 102.580 132.430 ;
        RECT 103.780 132.160 104.120 132.440 ;
        RECT 103.810 130.830 104.090 132.160 ;
        RECT 103.580 126.330 104.580 130.830 ;
        RECT 103.810 125.865 104.400 126.330 ;
        RECT 101.580 105.080 102.600 105.110 ;
        RECT 74.900 104.080 105.410 105.080 ;
        RECT 101.600 104.050 102.600 104.080 ;
        RECT 75.810 85.650 76.400 86.075 ;
        RECT 79.810 85.650 80.400 86.075 ;
        RECT 83.810 85.650 84.400 86.075 ;
        RECT 87.810 85.650 88.400 86.075 ;
        RECT 91.810 85.650 92.400 86.075 ;
        RECT 95.810 85.650 96.400 86.075 ;
        RECT 99.810 85.650 100.400 86.075 ;
        RECT 103.810 85.650 104.400 86.075 ;
        RECT 75.580 82.530 76.580 85.650 ;
        RECT 74.000 82.440 76.580 82.530 ;
        RECT 34.810 56.320 35.400 56.940 ;
        RECT 38.810 56.320 39.400 56.940 ;
        RECT 42.810 56.320 43.400 56.940 ;
        RECT 46.810 56.320 47.400 56.940 ;
        RECT 50.810 56.320 51.400 56.940 ;
        RECT 54.810 56.320 55.400 56.940 ;
        RECT 58.810 56.320 59.400 56.940 ;
        RECT 62.520 56.930 65.930 57.930 ;
        RECT 72.360 81.555 76.580 82.440 ;
        RECT 62.810 56.320 63.400 56.930 ;
        RECT 33.980 55.030 63.920 56.030 ;
        RECT 72.360 52.540 73.245 81.555 ;
        RECT 74.000 81.530 76.580 81.555 ;
        RECT 75.580 78.430 76.580 81.530 ;
        RECT 79.580 79.430 80.580 85.650 ;
        RECT 83.580 79.430 84.580 85.650 ;
        RECT 87.580 79.430 88.580 85.650 ;
        RECT 91.580 79.430 92.580 85.650 ;
        RECT 95.580 79.430 96.580 85.650 ;
        RECT 99.580 79.430 100.580 85.650 ;
        RECT 103.580 79.430 104.580 85.650 ;
        RECT 77.630 78.430 80.610 79.430 ;
        RECT 81.630 78.430 84.610 79.430 ;
        RECT 85.630 78.430 88.610 79.430 ;
        RECT 89.630 78.430 92.610 79.430 ;
        RECT 93.630 78.430 96.610 79.430 ;
        RECT 97.630 78.430 100.610 79.430 ;
        RECT 101.630 78.430 104.610 79.430 ;
        RECT 75.810 77.865 76.400 78.430 ;
        RECT 75.810 57.940 76.400 58.425 ;
        RECT 77.630 57.940 78.630 78.430 ;
        RECT 79.810 77.865 80.400 78.430 ;
        RECT 79.810 57.940 80.400 58.425 ;
        RECT 81.630 57.940 82.630 78.430 ;
        RECT 83.810 77.865 84.400 78.430 ;
        RECT 83.810 57.940 84.400 58.425 ;
        RECT 85.630 57.940 86.630 78.430 ;
        RECT 87.810 77.865 88.400 78.430 ;
        RECT 87.810 57.940 88.400 58.425 ;
        RECT 89.630 57.940 90.630 78.430 ;
        RECT 91.810 77.865 92.400 78.430 ;
        RECT 91.810 57.940 92.400 58.425 ;
        RECT 93.630 57.940 94.630 78.430 ;
        RECT 95.810 77.865 96.400 78.430 ;
        RECT 95.810 57.940 96.400 58.425 ;
        RECT 97.630 57.940 98.630 78.430 ;
        RECT 99.810 77.865 100.400 78.430 ;
        RECT 99.810 57.940 100.400 58.425 ;
        RECT 101.630 57.940 102.630 78.430 ;
        RECT 103.810 77.865 104.400 78.430 ;
        RECT 75.490 56.940 78.630 57.940 ;
        RECT 79.490 56.940 82.630 57.940 ;
        RECT 83.490 56.940 86.630 57.940 ;
        RECT 87.490 56.940 90.630 57.940 ;
        RECT 91.490 56.940 94.630 57.940 ;
        RECT 95.490 56.940 98.630 57.940 ;
        RECT 99.490 56.940 102.630 57.940 ;
        RECT 103.810 57.930 104.400 58.425 ;
        RECT 105.930 57.930 106.930 132.430 ;
        RECT 116.230 132.160 117.240 132.440 ;
        RECT 116.230 132.130 116.510 132.160 ;
        RECT 116.960 130.830 117.240 132.160 ;
        RECT 120.370 132.160 121.240 132.440 ;
        RECT 120.370 132.130 120.650 132.160 ;
        RECT 120.960 130.830 121.240 132.160 ;
        RECT 124.510 132.160 125.240 132.440 ;
        RECT 124.510 132.130 124.790 132.160 ;
        RECT 124.960 130.830 125.240 132.160 ;
        RECT 128.650 132.160 129.500 132.440 ;
        RECT 132.760 132.160 133.100 132.440 ;
        RECT 136.900 132.160 137.240 132.440 ;
        RECT 141.040 132.160 141.380 132.440 ;
        RECT 128.650 132.130 128.930 132.160 ;
        RECT 129.220 130.830 129.500 132.160 ;
        RECT 132.790 130.830 133.070 132.160 ;
        RECT 136.930 130.830 137.210 132.160 ;
        RECT 141.070 130.830 141.350 132.160 ;
        RECT 116.580 126.330 117.580 130.830 ;
        RECT 120.580 126.330 121.580 130.830 ;
        RECT 124.580 126.330 125.580 130.830 ;
        RECT 128.580 126.330 129.580 130.830 ;
        RECT 132.580 126.330 133.580 130.830 ;
        RECT 136.580 126.330 137.580 130.830 ;
        RECT 140.580 126.330 141.580 130.830 ;
        RECT 116.810 125.865 117.400 126.330 ;
        RECT 120.810 125.865 121.400 126.330 ;
        RECT 124.810 125.865 125.400 126.330 ;
        RECT 128.810 125.865 129.400 126.330 ;
        RECT 132.810 125.865 133.400 126.330 ;
        RECT 136.810 125.865 137.400 126.330 ;
        RECT 140.810 125.865 141.400 126.330 ;
        RECT 142.580 105.110 143.580 132.430 ;
        RECT 144.880 132.200 145.520 132.480 ;
        RECT 144.880 130.830 145.160 132.200 ;
        RECT 144.580 126.330 145.580 130.830 ;
        RECT 144.810 125.865 145.400 126.330 ;
        RECT 142.580 105.080 143.600 105.110 ;
        RECT 115.900 104.080 146.410 105.080 ;
        RECT 142.600 104.050 143.600 104.080 ;
        RECT 116.810 85.650 117.400 86.075 ;
        RECT 120.810 85.650 121.400 86.075 ;
        RECT 124.810 85.650 125.400 86.075 ;
        RECT 128.810 85.650 129.400 86.075 ;
        RECT 132.810 85.650 133.400 86.075 ;
        RECT 136.810 85.650 137.400 86.075 ;
        RECT 140.810 85.650 141.400 86.075 ;
        RECT 144.810 85.650 145.400 86.075 ;
        RECT 116.580 82.530 117.580 85.650 ;
        RECT 115.000 82.470 117.580 82.530 ;
        RECT 75.810 56.320 76.400 56.940 ;
        RECT 79.810 56.320 80.400 56.940 ;
        RECT 83.810 56.320 84.400 56.940 ;
        RECT 87.810 56.320 88.400 56.940 ;
        RECT 91.810 56.320 92.400 56.940 ;
        RECT 95.810 56.320 96.400 56.940 ;
        RECT 99.810 56.320 100.400 56.940 ;
        RECT 103.520 56.930 106.930 57.930 ;
        RECT 113.330 81.530 117.580 82.470 ;
        RECT 103.810 56.320 104.400 56.930 ;
        RECT 74.980 55.030 104.920 56.030 ;
        RECT 113.330 52.570 114.270 81.530 ;
        RECT 116.580 78.430 117.580 81.530 ;
        RECT 120.580 79.430 121.580 85.650 ;
        RECT 124.580 79.430 125.580 85.650 ;
        RECT 128.580 79.430 129.580 85.650 ;
        RECT 132.580 79.430 133.580 85.650 ;
        RECT 136.580 79.430 137.580 85.650 ;
        RECT 140.580 79.430 141.580 85.650 ;
        RECT 144.580 79.430 145.580 85.650 ;
        RECT 118.630 78.430 121.610 79.430 ;
        RECT 122.630 78.430 125.610 79.430 ;
        RECT 126.630 78.430 129.610 79.430 ;
        RECT 130.630 78.430 133.610 79.430 ;
        RECT 134.630 78.430 137.610 79.430 ;
        RECT 138.630 78.430 141.610 79.430 ;
        RECT 142.630 78.430 145.610 79.430 ;
        RECT 116.810 77.865 117.400 78.430 ;
        RECT 116.810 57.940 117.400 58.425 ;
        RECT 118.630 57.940 119.630 78.430 ;
        RECT 120.810 77.865 121.400 78.430 ;
        RECT 120.810 57.940 121.400 58.425 ;
        RECT 122.630 57.940 123.630 78.430 ;
        RECT 124.810 77.865 125.400 78.430 ;
        RECT 124.810 57.940 125.400 58.425 ;
        RECT 126.630 57.940 127.630 78.430 ;
        RECT 128.810 77.865 129.400 78.430 ;
        RECT 128.810 57.940 129.400 58.425 ;
        RECT 130.630 57.940 131.630 78.430 ;
        RECT 132.810 77.865 133.400 78.430 ;
        RECT 132.810 57.940 133.400 58.425 ;
        RECT 134.630 57.940 135.630 78.430 ;
        RECT 136.810 77.865 137.400 78.430 ;
        RECT 136.810 57.940 137.400 58.425 ;
        RECT 138.630 57.940 139.630 78.430 ;
        RECT 140.810 77.865 141.400 78.430 ;
        RECT 140.810 57.940 141.400 58.425 ;
        RECT 142.630 57.940 143.630 78.430 ;
        RECT 144.810 77.865 145.400 78.430 ;
        RECT 116.490 56.940 119.630 57.940 ;
        RECT 120.490 56.940 123.630 57.940 ;
        RECT 124.490 56.940 127.630 57.940 ;
        RECT 128.490 56.940 131.630 57.940 ;
        RECT 132.490 56.940 135.630 57.940 ;
        RECT 136.490 56.940 139.630 57.940 ;
        RECT 140.490 56.940 143.630 57.940 ;
        RECT 144.810 57.930 145.400 58.425 ;
        RECT 146.930 57.930 147.930 132.430 ;
        RECT 116.810 56.320 117.400 56.940 ;
        RECT 120.810 56.320 121.400 56.940 ;
        RECT 124.810 56.320 125.400 56.940 ;
        RECT 128.810 56.320 129.400 56.940 ;
        RECT 132.810 56.320 133.400 56.940 ;
        RECT 136.810 56.320 137.400 56.940 ;
        RECT 140.810 56.320 141.400 56.940 ;
        RECT 144.520 56.930 147.930 57.930 ;
        RECT 144.810 56.320 145.400 56.930 ;
        RECT 115.980 55.030 145.920 56.030 ;
        RECT 143.530 52.570 144.470 52.600 ;
        RECT 32.070 51.665 65.735 52.530 ;
        RECT 64.870 50.430 65.735 51.665 ;
        RECT 72.360 51.655 107.045 52.540 ;
        RECT 64.870 49.565 104.535 50.430 ;
        RECT 103.670 48.130 104.535 49.565 ;
        RECT 106.160 50.340 107.045 51.655 ;
        RECT 113.330 51.630 144.470 52.570 ;
        RECT 143.530 51.600 144.470 51.630 ;
        RECT 126.660 50.340 127.545 50.370 ;
        RECT 106.160 49.455 127.545 50.340 ;
        RECT 126.660 49.425 127.545 49.455 ;
        RECT 122.870 48.130 123.735 48.160 ;
        RECT 103.670 47.265 123.735 48.130 ;
        RECT 122.870 47.235 123.735 47.265 ;
        RECT 29.970 23.570 34.330 24.230 ;
        RECT 24.270 22.000 33.050 23.000 ;
        RECT 27.600 20.330 30.700 20.365 ;
        RECT 27.595 20.100 30.700 20.330 ;
        RECT 27.600 20.065 30.700 20.100 ;
        RECT 27.405 16.615 27.635 19.895 ;
        RECT 27.845 16.865 28.075 19.895 ;
        RECT 30.400 18.365 30.700 20.065 ;
        RECT 31.600 18.365 31.900 18.395 ;
        RECT 30.300 18.065 31.900 18.365 ;
        RECT 31.600 18.035 31.900 18.065 ;
        RECT 30.220 16.865 30.450 17.915 ;
        RECT 30.660 17.765 30.890 17.915 ;
        RECT 32.050 17.765 33.050 22.000 ;
        RECT 22.770 15.615 27.650 16.615 ;
        RECT 27.845 15.615 30.450 16.865 ;
        RECT 30.650 16.765 33.050 17.765 ;
        RECT 27.405 11.895 27.635 15.615 ;
        RECT 27.845 11.895 28.075 15.615 ;
        RECT 29.050 12.365 29.350 15.615 ;
        RECT 30.220 13.915 30.450 15.615 ;
        RECT 30.660 13.915 30.890 16.765 ;
        RECT 32.050 16.195 33.050 16.365 ;
        RECT 33.670 16.195 34.330 23.570 ;
        RECT 31.600 16.015 31.900 16.045 ;
        RECT 32.050 16.015 34.330 16.195 ;
        RECT 31.600 15.715 34.330 16.015 ;
        RECT 31.600 15.685 31.900 15.715 ;
        RECT 32.050 15.535 34.330 15.715 ;
        RECT 32.050 15.365 33.050 15.535 ;
        RECT 31.600 13.765 31.900 13.795 ;
        RECT 30.300 13.465 31.900 13.765 ;
        RECT 33.770 13.700 34.830 14.700 ;
        RECT 29.900 12.365 30.200 12.395 ;
        RECT 29.050 12.065 30.200 12.365 ;
        RECT 29.900 12.035 30.200 12.065 ;
        RECT 30.400 11.715 30.700 13.465 ;
        RECT 31.600 13.435 31.900 13.465 ;
        RECT 32.050 12.700 33.050 12.715 ;
        RECT 33.800 12.700 34.800 13.700 ;
        RECT 32.000 12.365 36.600 12.700 ;
        RECT 30.920 12.065 36.600 12.365 ;
        RECT 27.550 11.415 30.700 11.715 ;
        RECT 32.000 11.700 36.600 12.065 ;
        RECT 35.600 9.000 36.600 11.700 ;
        RECT 35.570 8.000 36.630 9.000 ;
      LAYER via ;
        RECT 114.400 215.570 114.660 215.830 ;
        RECT 119.460 215.570 119.720 215.830 ;
        RECT 66.100 215.230 66.360 215.490 ;
        RECT 67.020 215.230 67.280 215.490 ;
        RECT 105.660 215.230 105.920 215.490 ;
        RECT 107.040 215.230 107.300 215.490 ;
        RECT 123.600 215.230 123.860 215.490 ;
        RECT 144.760 215.230 145.020 215.490 ;
        RECT 40.170 214.720 40.430 214.980 ;
        RECT 40.490 214.720 40.750 214.980 ;
        RECT 40.810 214.720 41.070 214.980 ;
        RECT 41.130 214.720 41.390 214.980 ;
        RECT 41.450 214.720 41.710 214.980 ;
        RECT 41.770 214.720 42.030 214.980 ;
        RECT 70.170 214.720 70.430 214.980 ;
        RECT 70.490 214.720 70.750 214.980 ;
        RECT 70.810 214.720 71.070 214.980 ;
        RECT 71.130 214.720 71.390 214.980 ;
        RECT 71.450 214.720 71.710 214.980 ;
        RECT 71.770 214.720 72.030 214.980 ;
        RECT 100.170 214.720 100.430 214.980 ;
        RECT 100.490 214.720 100.750 214.980 ;
        RECT 100.810 214.720 101.070 214.980 ;
        RECT 101.130 214.720 101.390 214.980 ;
        RECT 101.450 214.720 101.710 214.980 ;
        RECT 101.770 214.720 102.030 214.980 ;
        RECT 130.170 214.720 130.430 214.980 ;
        RECT 130.490 214.720 130.750 214.980 ;
        RECT 130.810 214.720 131.070 214.980 ;
        RECT 131.130 214.720 131.390 214.980 ;
        RECT 131.450 214.720 131.710 214.980 ;
        RECT 131.770 214.720 132.030 214.980 ;
        RECT 56.440 214.210 56.700 214.470 ;
        RECT 59.200 214.210 59.460 214.470 ;
        RECT 64.260 214.210 64.520 214.470 ;
        RECT 66.560 214.210 66.820 214.470 ;
        RECT 69.780 214.210 70.040 214.470 ;
        RECT 73.920 214.210 74.180 214.470 ;
        RECT 78.980 214.210 79.240 214.470 ;
        RECT 81.280 214.210 81.540 214.470 ;
        RECT 84.960 214.210 85.220 214.470 ;
        RECT 88.640 214.210 88.900 214.470 ;
        RECT 105.660 214.210 105.920 214.470 ;
        RECT 32.470 213.070 33.130 213.730 ;
        RECT 44.480 213.190 44.740 213.450 ;
        RECT 57.820 213.190 58.080 213.450 ;
        RECT 67.020 212.850 67.280 213.110 ;
        RECT 67.940 212.850 68.200 213.110 ;
        RECT 71.620 213.530 71.880 213.790 ;
        RECT 126.360 214.210 126.620 214.470 ;
        RECT 118.540 213.870 118.800 214.130 ;
        RECT 119.920 213.870 120.180 214.130 ;
        RECT 72.540 213.190 72.800 213.450 ;
        RECT 76.220 213.190 76.480 213.450 ;
        RECT 78.060 213.190 78.320 213.450 ;
        RECT 84.040 213.190 84.300 213.450 ;
        RECT 76.680 212.850 76.940 213.110 ;
        RECT 80.820 212.850 81.080 213.110 ;
        RECT 81.740 212.850 82.000 213.110 ;
        RECT 93.240 212.850 93.500 213.110 ;
        RECT 99.680 213.190 99.940 213.450 ;
        RECT 117.160 213.530 117.420 213.790 ;
        RECT 144.760 213.870 145.020 214.130 ;
        RECT 117.620 213.190 117.880 213.450 ;
        RECT 121.760 213.190 122.020 213.450 ;
        RECT 125.440 213.190 125.700 213.450 ;
        RECT 129.120 213.190 129.380 213.450 ;
        RECT 133.720 213.190 133.980 213.450 ;
        RECT 134.180 213.190 134.440 213.450 ;
        RECT 136.480 213.190 136.740 213.450 ;
        RECT 140.160 213.190 140.420 213.450 ;
        RECT 140.620 213.190 140.880 213.450 ;
        RECT 124.520 212.850 124.780 213.110 ;
        RECT 143.840 213.190 144.100 213.450 ;
        RECT 147.520 213.190 147.780 213.450 ;
        RECT 45.860 212.510 46.120 212.770 ;
        RECT 59.200 212.510 59.460 212.770 ;
        RECT 68.860 212.510 69.120 212.770 ;
        RECT 73.000 212.510 73.260 212.770 ;
        RECT 92.780 212.510 93.040 212.770 ;
        RECT 102.440 212.510 102.700 212.770 ;
        RECT 125.900 212.510 126.160 212.770 ;
        RECT 127.740 212.510 128.000 212.770 ;
        RECT 129.580 212.510 129.840 212.770 ;
        RECT 133.260 212.510 133.520 212.770 ;
        RECT 134.180 212.510 134.440 212.770 ;
        RECT 141.080 212.510 141.340 212.770 ;
        RECT 55.170 212.000 55.430 212.260 ;
        RECT 55.490 212.000 55.750 212.260 ;
        RECT 55.810 212.000 56.070 212.260 ;
        RECT 56.130 212.000 56.390 212.260 ;
        RECT 56.450 212.000 56.710 212.260 ;
        RECT 56.770 212.000 57.030 212.260 ;
        RECT 85.170 212.000 85.430 212.260 ;
        RECT 85.490 212.000 85.750 212.260 ;
        RECT 85.810 212.000 86.070 212.260 ;
        RECT 86.130 212.000 86.390 212.260 ;
        RECT 86.450 212.000 86.710 212.260 ;
        RECT 86.770 212.000 87.030 212.260 ;
        RECT 115.170 212.000 115.430 212.260 ;
        RECT 115.490 212.000 115.750 212.260 ;
        RECT 115.810 212.000 116.070 212.260 ;
        RECT 116.130 212.000 116.390 212.260 ;
        RECT 116.450 212.000 116.710 212.260 ;
        RECT 116.770 212.000 117.030 212.260 ;
        RECT 145.170 212.000 145.430 212.260 ;
        RECT 145.490 212.000 145.750 212.260 ;
        RECT 145.810 212.000 146.070 212.260 ;
        RECT 146.130 212.000 146.390 212.260 ;
        RECT 146.450 212.000 146.710 212.260 ;
        RECT 146.770 212.000 147.030 212.260 ;
        RECT 44.480 211.490 44.740 211.750 ;
        RECT 45.400 211.490 45.660 211.750 ;
        RECT 57.820 211.490 58.080 211.750 ;
        RECT 66.560 211.490 66.820 211.750 ;
        RECT 71.620 211.490 71.880 211.750 ;
        RECT 73.000 211.490 73.260 211.750 ;
        RECT 78.060 211.490 78.320 211.750 ;
        RECT 45.860 210.810 46.120 211.070 ;
        RECT 47.700 210.810 47.960 211.070 ;
        RECT 63.800 211.150 64.060 211.410 ;
        RECT 55.060 210.810 55.320 211.070 ;
        RECT 60.120 210.810 60.380 211.070 ;
        RECT 66.100 210.810 66.360 211.070 ;
        RECT 67.020 210.810 67.280 211.070 ;
        RECT 68.860 210.810 69.120 211.070 ;
        RECT 73.460 210.810 73.720 211.070 ;
        RECT 77.140 210.810 77.400 211.070 ;
        RECT 86.800 211.490 87.060 211.750 ;
        RECT 84.500 210.810 84.760 211.070 ;
        RECT 107.040 211.490 107.300 211.750 ;
        RECT 112.100 211.490 112.360 211.750 ;
        RECT 118.080 211.490 118.340 211.750 ;
        RECT 123.600 211.490 123.860 211.750 ;
        RECT 125.440 211.490 125.700 211.750 ;
        RECT 129.580 211.490 129.840 211.750 ;
        RECT 140.620 211.490 140.880 211.750 ;
        RECT 38.500 209.790 38.760 210.050 ;
        RECT 42.640 209.790 42.900 210.050 ;
        RECT 54.600 209.790 54.860 210.050 ;
        RECT 64.260 209.790 64.520 210.050 ;
        RECT 78.980 210.470 79.240 210.730 ;
        RECT 79.900 210.470 80.160 210.730 ;
        RECT 83.580 210.130 83.840 210.390 ;
        RECT 73.920 209.790 74.180 210.050 ;
        RECT 79.900 209.790 80.160 210.050 ;
        RECT 87.260 209.790 87.520 210.050 ;
        RECT 87.720 209.790 87.980 210.050 ;
        RECT 90.020 209.790 90.280 210.050 ;
        RECT 99.680 209.790 99.940 210.050 ;
        RECT 106.120 210.810 106.380 211.070 ;
        RECT 120.380 211.150 120.640 211.410 ;
        RECT 109.340 210.470 109.600 210.730 ;
        RECT 114.860 210.470 115.120 210.730 ;
        RECT 115.780 210.810 116.040 211.070 ;
        RECT 121.300 210.810 121.560 211.070 ;
        RECT 118.540 210.470 118.800 210.730 ;
        RECT 124.520 210.810 124.780 211.070 ;
        RECT 126.360 210.810 126.620 211.070 ;
        RECT 123.140 210.470 123.400 210.730 ;
        RECT 112.560 210.130 112.820 210.390 ;
        RECT 119.000 210.130 119.260 210.390 ;
        RECT 120.840 210.130 121.100 210.390 ;
        RECT 110.260 209.790 110.520 210.050 ;
        RECT 113.940 209.790 114.200 210.050 ;
        RECT 122.680 209.790 122.940 210.050 ;
        RECT 127.280 210.470 127.540 210.730 ;
        RECT 133.260 210.810 133.520 211.070 ;
        RECT 127.740 210.130 128.000 210.390 ;
        RECT 126.360 209.790 126.620 210.050 ;
        RECT 40.170 209.280 40.430 209.540 ;
        RECT 40.490 209.280 40.750 209.540 ;
        RECT 40.810 209.280 41.070 209.540 ;
        RECT 41.130 209.280 41.390 209.540 ;
        RECT 41.450 209.280 41.710 209.540 ;
        RECT 41.770 209.280 42.030 209.540 ;
        RECT 70.170 209.280 70.430 209.540 ;
        RECT 70.490 209.280 70.750 209.540 ;
        RECT 70.810 209.280 71.070 209.540 ;
        RECT 71.130 209.280 71.390 209.540 ;
        RECT 71.450 209.280 71.710 209.540 ;
        RECT 71.770 209.280 72.030 209.540 ;
        RECT 100.170 209.280 100.430 209.540 ;
        RECT 100.490 209.280 100.750 209.540 ;
        RECT 100.810 209.280 101.070 209.540 ;
        RECT 101.130 209.280 101.390 209.540 ;
        RECT 101.450 209.280 101.710 209.540 ;
        RECT 101.770 209.280 102.030 209.540 ;
        RECT 130.170 209.280 130.430 209.540 ;
        RECT 130.490 209.280 130.750 209.540 ;
        RECT 130.810 209.280 131.070 209.540 ;
        RECT 131.130 209.280 131.390 209.540 ;
        RECT 131.450 209.280 131.710 209.540 ;
        RECT 131.770 209.280 132.030 209.540 ;
        RECT 42.640 208.770 42.900 209.030 ;
        RECT 45.400 208.770 45.660 209.030 ;
        RECT 47.700 208.770 47.960 209.030 ;
        RECT 72.540 208.770 72.800 209.030 ;
        RECT 76.220 208.770 76.480 209.030 ;
        RECT 83.580 208.770 83.840 209.030 ;
        RECT 87.720 208.770 87.980 209.030 ;
        RECT 90.020 208.770 90.280 209.030 ;
        RECT 64.720 208.430 64.980 208.690 ;
        RECT 85.880 208.430 86.140 208.690 ;
        RECT 39.420 207.750 39.680 208.010 ;
        RECT 44.020 207.750 44.280 208.010 ;
        RECT 42.180 207.410 42.440 207.670 ;
        RECT 46.780 207.750 47.040 208.010 ;
        RECT 52.760 207.750 53.020 208.010 ;
        RECT 55.060 207.750 55.320 208.010 ;
        RECT 67.480 207.750 67.740 208.010 ;
        RECT 72.080 207.750 72.340 208.010 ;
        RECT 74.380 207.750 74.640 208.010 ;
        RECT 64.260 207.410 64.520 207.670 ;
        RECT 46.320 207.070 46.580 207.330 ;
        RECT 61.040 207.070 61.300 207.330 ;
        RECT 76.220 207.750 76.480 208.010 ;
        RECT 78.980 207.750 79.240 208.010 ;
        RECT 79.900 207.750 80.160 208.010 ;
        RECT 89.100 208.430 89.360 208.690 ;
        RECT 92.780 208.430 93.040 208.690 ;
        RECT 87.260 207.750 87.520 208.010 ;
        RECT 90.480 207.750 90.740 208.010 ;
        RECT 91.400 207.750 91.660 208.010 ;
        RECT 98.300 207.750 98.560 208.010 ;
        RECT 106.120 208.770 106.380 209.030 ;
        RECT 114.400 208.770 114.660 209.030 ;
        RECT 117.620 208.770 117.880 209.030 ;
        RECT 121.300 208.770 121.560 209.030 ;
        RECT 122.680 208.770 122.940 209.030 ;
        RECT 125.440 208.770 125.700 209.030 ;
        RECT 126.360 208.770 126.620 209.030 ;
        RECT 133.720 208.770 133.980 209.030 ;
        RECT 140.620 208.770 140.880 209.030 ;
        RECT 104.280 208.430 104.540 208.690 ;
        RECT 110.260 208.090 110.520 208.350 ;
        RECT 112.100 208.090 112.360 208.350 ;
        RECT 112.560 208.090 112.820 208.350 ;
        RECT 99.220 207.750 99.480 208.010 ;
        RECT 99.680 207.750 99.940 208.010 ;
        RECT 102.440 207.750 102.700 208.010 ;
        RECT 106.580 207.750 106.840 208.010 ;
        RECT 113.940 207.750 114.200 208.010 ;
        RECT 118.540 208.090 118.800 208.350 ;
        RECT 122.680 207.750 122.940 208.010 ;
        RECT 126.820 207.750 127.080 208.010 ;
        RECT 128.200 207.750 128.460 208.010 ;
        RECT 129.120 208.090 129.380 208.350 ;
        RECT 134.180 207.750 134.440 208.010 ;
        RECT 83.120 207.070 83.380 207.330 ;
        RECT 88.180 207.070 88.440 207.330 ;
        RECT 117.160 207.070 117.420 207.330 ;
        RECT 117.620 207.070 117.880 207.330 ;
        RECT 119.920 207.070 120.180 207.330 ;
        RECT 126.820 207.070 127.080 207.330 ;
        RECT 55.170 206.560 55.430 206.820 ;
        RECT 55.490 206.560 55.750 206.820 ;
        RECT 55.810 206.560 56.070 206.820 ;
        RECT 56.130 206.560 56.390 206.820 ;
        RECT 56.450 206.560 56.710 206.820 ;
        RECT 56.770 206.560 57.030 206.820 ;
        RECT 85.170 206.560 85.430 206.820 ;
        RECT 85.490 206.560 85.750 206.820 ;
        RECT 85.810 206.560 86.070 206.820 ;
        RECT 86.130 206.560 86.390 206.820 ;
        RECT 86.450 206.560 86.710 206.820 ;
        RECT 86.770 206.560 87.030 206.820 ;
        RECT 115.170 206.560 115.430 206.820 ;
        RECT 115.490 206.560 115.750 206.820 ;
        RECT 115.810 206.560 116.070 206.820 ;
        RECT 116.130 206.560 116.390 206.820 ;
        RECT 116.450 206.560 116.710 206.820 ;
        RECT 116.770 206.560 117.030 206.820 ;
        RECT 145.170 206.560 145.430 206.820 ;
        RECT 145.490 206.560 145.750 206.820 ;
        RECT 145.810 206.560 146.070 206.820 ;
        RECT 146.130 206.560 146.390 206.820 ;
        RECT 146.450 206.560 146.710 206.820 ;
        RECT 146.770 206.560 147.030 206.820 ;
        RECT 38.960 205.710 39.220 205.970 ;
        RECT 44.480 205.710 44.740 205.970 ;
        RECT 38.500 205.370 38.760 205.630 ;
        RECT 52.760 206.050 53.020 206.310 ;
        RECT 76.220 206.050 76.480 206.310 ;
        RECT 46.320 205.710 46.580 205.970 ;
        RECT 67.940 205.710 68.200 205.970 ;
        RECT 63.800 205.370 64.060 205.630 ;
        RECT 72.080 205.710 72.340 205.970 ;
        RECT 73.920 205.710 74.180 205.970 ;
        RECT 84.500 205.710 84.760 205.970 ;
        RECT 54.140 205.030 54.400 205.290 ;
        RECT 62.420 205.030 62.680 205.290 ;
        RECT 77.140 205.370 77.400 205.630 ;
        RECT 74.380 205.030 74.640 205.290 ;
        RECT 79.900 205.030 80.160 205.290 ;
        RECT 81.280 205.030 81.540 205.290 ;
        RECT 87.260 205.370 87.520 205.630 ;
        RECT 62.880 204.690 63.140 204.950 ;
        RECT 93.700 205.710 93.960 205.970 ;
        RECT 98.760 206.050 99.020 206.310 ;
        RECT 120.840 206.050 121.100 206.310 ;
        RECT 122.220 206.050 122.480 206.310 ;
        RECT 123.600 206.050 123.860 206.310 ;
        RECT 125.440 206.050 125.700 206.310 ;
        RECT 125.900 206.050 126.160 206.310 ;
        RECT 126.820 206.050 127.080 206.310 ;
        RECT 89.100 205.370 89.360 205.630 ;
        RECT 43.560 204.350 43.820 204.610 ;
        RECT 46.780 204.350 47.040 204.610 ;
        RECT 50.460 204.350 50.720 204.610 ;
        RECT 60.120 204.350 60.380 204.610 ;
        RECT 63.800 204.350 64.060 204.610 ;
        RECT 65.640 204.350 65.900 204.610 ;
        RECT 67.940 204.350 68.200 204.610 ;
        RECT 73.460 204.350 73.720 204.610 ;
        RECT 83.120 204.350 83.380 204.610 ;
        RECT 86.800 204.350 87.060 204.610 ;
        RECT 87.720 204.350 87.980 204.610 ;
        RECT 89.100 204.690 89.360 204.950 ;
        RECT 90.940 204.690 91.200 204.950 ;
        RECT 92.320 205.030 92.580 205.290 ;
        RECT 113.020 205.030 113.280 205.290 ;
        RECT 123.140 205.710 123.400 205.970 ;
        RECT 129.120 206.050 129.380 206.310 ;
        RECT 117.620 205.370 117.880 205.630 ;
        RECT 117.160 205.030 117.420 205.290 ;
        RECT 125.900 205.370 126.160 205.630 ;
        RECT 132.340 205.370 132.600 205.630 ;
        RECT 115.320 204.690 115.580 204.950 ;
        RECT 124.980 205.030 125.240 205.290 ;
        RECT 125.440 205.030 125.700 205.290 ;
        RECT 140.620 205.710 140.880 205.970 ;
        RECT 140.160 205.370 140.420 205.630 ;
        RECT 134.640 205.030 134.900 205.290 ;
        RECT 96.920 204.350 97.180 204.610 ;
        RECT 105.660 204.350 105.920 204.610 ;
        RECT 141.080 204.690 141.340 204.950 ;
        RECT 121.300 204.350 121.560 204.610 ;
        RECT 135.560 204.350 135.820 204.610 ;
        RECT 40.170 203.840 40.430 204.100 ;
        RECT 40.490 203.840 40.750 204.100 ;
        RECT 40.810 203.840 41.070 204.100 ;
        RECT 41.130 203.840 41.390 204.100 ;
        RECT 41.450 203.840 41.710 204.100 ;
        RECT 41.770 203.840 42.030 204.100 ;
        RECT 70.170 203.840 70.430 204.100 ;
        RECT 70.490 203.840 70.750 204.100 ;
        RECT 70.810 203.840 71.070 204.100 ;
        RECT 71.130 203.840 71.390 204.100 ;
        RECT 71.450 203.840 71.710 204.100 ;
        RECT 71.770 203.840 72.030 204.100 ;
        RECT 100.170 203.840 100.430 204.100 ;
        RECT 100.490 203.840 100.750 204.100 ;
        RECT 100.810 203.840 101.070 204.100 ;
        RECT 101.130 203.840 101.390 204.100 ;
        RECT 101.450 203.840 101.710 204.100 ;
        RECT 101.770 203.840 102.030 204.100 ;
        RECT 130.170 203.840 130.430 204.100 ;
        RECT 130.490 203.840 130.750 204.100 ;
        RECT 130.810 203.840 131.070 204.100 ;
        RECT 131.130 203.840 131.390 204.100 ;
        RECT 131.450 203.840 131.710 204.100 ;
        RECT 131.770 203.840 132.030 204.100 ;
        RECT 41.720 203.330 41.980 203.590 ;
        RECT 42.180 203.330 42.440 203.590 ;
        RECT 43.560 203.330 43.820 203.590 ;
        RECT 44.480 203.330 44.740 203.590 ;
        RECT 41.260 202.650 41.520 202.910 ;
        RECT 45.400 202.990 45.660 203.250 ;
        RECT 38.960 201.970 39.220 202.230 ;
        RECT 48.160 202.990 48.420 203.250 ;
        RECT 52.760 203.330 53.020 203.590 ;
        RECT 61.040 203.330 61.300 203.590 ;
        RECT 62.880 203.330 63.140 203.590 ;
        RECT 65.640 203.330 65.900 203.590 ;
        RECT 68.400 203.330 68.660 203.590 ;
        RECT 83.580 203.330 83.840 203.590 ;
        RECT 60.120 202.650 60.380 202.910 ;
        RECT 41.720 201.630 41.980 201.890 ;
        RECT 43.100 201.630 43.360 201.890 ;
        RECT 48.160 202.310 48.420 202.570 ;
        RECT 57.360 202.310 57.620 202.570 ;
        RECT 64.720 202.310 64.980 202.570 ;
        RECT 67.020 202.990 67.280 203.250 ;
        RECT 48.160 201.630 48.420 201.890 ;
        RECT 53.220 201.630 53.480 201.890 ;
        RECT 57.820 201.630 58.080 201.890 ;
        RECT 67.480 202.310 67.740 202.570 ;
        RECT 84.040 202.990 84.300 203.250 ;
        RECT 98.300 203.330 98.560 203.590 ;
        RECT 113.020 203.330 113.280 203.590 ;
        RECT 121.300 203.330 121.560 203.590 ;
        RECT 86.800 202.650 87.060 202.910 ;
        RECT 87.720 202.650 87.980 202.910 ;
        RECT 97.840 202.990 98.100 203.250 ;
        RECT 70.700 201.970 70.960 202.230 ;
        RECT 82.660 202.310 82.920 202.570 ;
        RECT 92.780 202.650 93.040 202.910 ;
        RECT 102.440 202.650 102.700 202.910 ;
        RECT 115.320 202.990 115.580 203.250 ;
        RECT 123.600 202.650 123.860 202.910 ;
        RECT 124.980 202.650 125.240 202.910 ;
        RECT 127.280 202.650 127.540 202.910 ;
        RECT 90.020 202.310 90.280 202.570 ;
        RECT 90.940 202.310 91.200 202.570 ;
        RECT 91.400 202.310 91.660 202.570 ;
        RECT 91.860 202.310 92.120 202.570 ;
        RECT 69.780 201.630 70.040 201.890 ;
        RECT 74.380 201.630 74.640 201.890 ;
        RECT 80.820 201.630 81.080 201.890 ;
        RECT 89.560 201.970 89.820 202.230 ;
        RECT 98.760 202.310 99.020 202.570 ;
        RECT 102.900 202.310 103.160 202.570 ;
        RECT 104.740 202.310 105.000 202.570 ;
        RECT 105.200 202.310 105.460 202.570 ;
        RECT 105.660 202.310 105.920 202.570 ;
        RECT 119.460 202.310 119.720 202.570 ;
        RECT 84.500 201.630 84.760 201.890 ;
        RECT 93.240 201.630 93.500 201.890 ;
        RECT 117.620 201.970 117.880 202.230 ;
        RECT 106.580 201.630 106.840 201.890 ;
        RECT 119.920 201.630 120.180 201.890 ;
        RECT 127.280 201.630 127.540 201.890 ;
        RECT 132.340 202.310 132.600 202.570 ;
        RECT 134.640 202.310 134.900 202.570 ;
        RECT 135.560 202.310 135.820 202.570 ;
        RECT 140.160 203.330 140.420 203.590 ;
        RECT 141.080 202.650 141.340 202.910 ;
        RECT 149.820 202.650 150.080 202.910 ;
        RECT 132.800 201.970 133.060 202.230 ;
        RECT 133.260 201.970 133.520 202.230 ;
        RECT 144.300 201.970 144.560 202.230 ;
        RECT 134.180 201.630 134.440 201.890 ;
        RECT 136.940 201.630 137.200 201.890 ;
        RECT 147.520 201.630 147.780 201.890 ;
        RECT 55.170 201.120 55.430 201.380 ;
        RECT 55.490 201.120 55.750 201.380 ;
        RECT 55.810 201.120 56.070 201.380 ;
        RECT 56.130 201.120 56.390 201.380 ;
        RECT 56.450 201.120 56.710 201.380 ;
        RECT 56.770 201.120 57.030 201.380 ;
        RECT 85.170 201.120 85.430 201.380 ;
        RECT 85.490 201.120 85.750 201.380 ;
        RECT 85.810 201.120 86.070 201.380 ;
        RECT 86.130 201.120 86.390 201.380 ;
        RECT 86.450 201.120 86.710 201.380 ;
        RECT 86.770 201.120 87.030 201.380 ;
        RECT 115.170 201.120 115.430 201.380 ;
        RECT 115.490 201.120 115.750 201.380 ;
        RECT 115.810 201.120 116.070 201.380 ;
        RECT 116.130 201.120 116.390 201.380 ;
        RECT 116.450 201.120 116.710 201.380 ;
        RECT 116.770 201.120 117.030 201.380 ;
        RECT 145.170 201.120 145.430 201.380 ;
        RECT 145.490 201.120 145.750 201.380 ;
        RECT 145.810 201.120 146.070 201.380 ;
        RECT 146.130 201.120 146.390 201.380 ;
        RECT 146.450 201.120 146.710 201.380 ;
        RECT 146.770 201.120 147.030 201.380 ;
        RECT 41.720 200.610 41.980 200.870 ;
        RECT 41.260 200.270 41.520 200.530 ;
        RECT 42.640 200.270 42.900 200.530 ;
        RECT 43.100 199.930 43.360 200.190 ;
        RECT 45.400 200.270 45.660 200.530 ;
        RECT 57.360 200.610 57.620 200.870 ;
        RECT 60.120 200.610 60.380 200.870 ;
        RECT 70.700 200.610 70.960 200.870 ;
        RECT 45.860 199.930 46.120 200.190 ;
        RECT 54.600 199.930 54.860 200.190 ;
        RECT 43.560 199.590 43.820 199.850 ;
        RECT 38.960 199.250 39.220 199.510 ;
        RECT 42.180 199.250 42.440 199.510 ;
        RECT 44.940 199.250 45.200 199.510 ;
        RECT 46.320 199.590 46.580 199.850 ;
        RECT 56.440 199.930 56.700 200.190 ;
        RECT 57.820 199.930 58.080 200.190 ;
        RECT 60.120 199.930 60.380 200.190 ;
        RECT 62.880 199.930 63.140 200.190 ;
        RECT 72.540 199.930 72.800 200.190 ;
        RECT 75.760 199.930 76.020 200.190 ;
        RECT 84.500 199.930 84.760 200.190 ;
        RECT 56.900 199.590 57.160 199.850 ;
        RECT 45.400 198.910 45.660 199.170 ;
        RECT 48.160 198.910 48.420 199.170 ;
        RECT 50.920 198.910 51.180 199.170 ;
        RECT 54.140 198.910 54.400 199.170 ;
        RECT 56.440 198.910 56.700 199.170 ;
        RECT 58.740 199.250 59.000 199.510 ;
        RECT 63.340 199.250 63.600 199.510 ;
        RECT 69.780 199.590 70.040 199.850 ;
        RECT 77.140 199.590 77.400 199.850 ;
        RECT 82.200 199.590 82.460 199.850 ;
        RECT 84.040 199.590 84.300 199.850 ;
        RECT 87.720 200.270 87.980 200.530 ;
        RECT 91.400 200.610 91.660 200.870 ;
        RECT 102.440 200.610 102.700 200.870 ;
        RECT 104.740 200.610 105.000 200.870 ;
        RECT 112.100 200.610 112.360 200.870 ;
        RECT 120.380 200.610 120.640 200.870 ;
        RECT 86.800 199.590 87.060 199.850 ;
        RECT 90.940 199.590 91.200 199.850 ;
        RECT 60.580 198.910 60.840 199.170 ;
        RECT 61.500 198.910 61.760 199.170 ;
        RECT 79.900 199.250 80.160 199.510 ;
        RECT 66.560 198.910 66.820 199.170 ;
        RECT 73.000 198.910 73.260 199.170 ;
        RECT 80.360 198.910 80.620 199.170 ;
        RECT 87.720 199.250 87.980 199.510 ;
        RECT 90.480 199.250 90.740 199.510 ;
        RECT 98.300 199.930 98.560 200.190 ;
        RECT 96.460 199.590 96.720 199.850 ;
        RECT 97.380 199.590 97.640 199.850 ;
        RECT 94.160 199.250 94.420 199.510 ;
        RECT 98.760 199.250 99.020 199.510 ;
        RECT 86.340 198.910 86.600 199.170 ;
        RECT 87.260 198.910 87.520 199.170 ;
        RECT 89.560 198.910 89.820 199.170 ;
        RECT 94.620 198.910 94.880 199.170 ;
        RECT 99.680 198.910 99.940 199.170 ;
        RECT 101.980 199.930 102.240 200.190 ;
        RECT 103.820 200.270 104.080 200.530 ;
        RECT 107.040 200.270 107.300 200.530 ;
        RECT 113.020 200.270 113.280 200.530 ;
        RECT 114.400 199.930 114.660 200.190 ;
        RECT 128.660 200.270 128.920 200.530 ;
        RECT 124.980 199.930 125.240 200.190 ;
        RECT 125.440 199.930 125.700 200.190 ;
        RECT 126.820 199.930 127.080 200.190 ;
        RECT 134.640 200.270 134.900 200.530 ;
        RECT 127.280 199.590 127.540 199.850 ;
        RECT 121.300 199.250 121.560 199.510 ;
        RECT 102.440 198.910 102.700 199.170 ;
        RECT 108.880 198.910 109.140 199.170 ;
        RECT 113.020 198.910 113.280 199.170 ;
        RECT 113.940 198.910 114.200 199.170 ;
        RECT 125.900 198.910 126.160 199.170 ;
        RECT 126.360 198.910 126.620 199.170 ;
        RECT 144.760 198.910 145.020 199.170 ;
        RECT 40.170 198.400 40.430 198.660 ;
        RECT 40.490 198.400 40.750 198.660 ;
        RECT 40.810 198.400 41.070 198.660 ;
        RECT 41.130 198.400 41.390 198.660 ;
        RECT 41.450 198.400 41.710 198.660 ;
        RECT 41.770 198.400 42.030 198.660 ;
        RECT 70.170 198.400 70.430 198.660 ;
        RECT 70.490 198.400 70.750 198.660 ;
        RECT 70.810 198.400 71.070 198.660 ;
        RECT 71.130 198.400 71.390 198.660 ;
        RECT 71.450 198.400 71.710 198.660 ;
        RECT 71.770 198.400 72.030 198.660 ;
        RECT 100.170 198.400 100.430 198.660 ;
        RECT 100.490 198.400 100.750 198.660 ;
        RECT 100.810 198.400 101.070 198.660 ;
        RECT 101.130 198.400 101.390 198.660 ;
        RECT 101.450 198.400 101.710 198.660 ;
        RECT 101.770 198.400 102.030 198.660 ;
        RECT 130.170 198.400 130.430 198.660 ;
        RECT 130.490 198.400 130.750 198.660 ;
        RECT 130.810 198.400 131.070 198.660 ;
        RECT 131.130 198.400 131.390 198.660 ;
        RECT 131.450 198.400 131.710 198.660 ;
        RECT 131.770 198.400 132.030 198.660 ;
        RECT 43.560 197.890 43.820 198.150 ;
        RECT 45.860 197.890 46.120 198.150 ;
        RECT 54.600 197.550 54.860 197.810 ;
        RECT 58.740 197.890 59.000 198.150 ;
        RECT 59.200 197.890 59.460 198.150 ;
        RECT 87.720 197.890 87.980 198.150 ;
        RECT 99.680 197.890 99.940 198.150 ;
        RECT 56.900 197.550 57.160 197.810 ;
        RECT 86.800 197.550 87.060 197.810 ;
        RECT 61.960 197.210 62.220 197.470 ;
        RECT 42.180 196.870 42.440 197.130 ;
        RECT 44.940 196.870 45.200 197.130 ;
        RECT 49.540 196.870 49.800 197.130 ;
        RECT 50.920 196.870 51.180 197.130 ;
        RECT 54.600 196.870 54.860 197.130 ;
        RECT 56.900 196.870 57.160 197.130 ;
        RECT 60.580 196.870 60.840 197.130 ;
        RECT 62.880 196.870 63.140 197.130 ;
        RECT 65.640 197.210 65.900 197.470 ;
        RECT 87.720 197.210 87.980 197.470 ;
        RECT 88.180 197.210 88.440 197.470 ;
        RECT 73.000 196.870 73.260 197.130 ;
        RECT 65.640 196.530 65.900 196.790 ;
        RECT 67.480 196.530 67.740 196.790 ;
        RECT 69.320 196.530 69.580 196.790 ;
        RECT 84.500 196.530 84.760 196.790 ;
        RECT 88.640 196.870 88.900 197.130 ;
        RECT 90.940 197.550 91.200 197.810 ;
        RECT 90.480 197.210 90.740 197.470 ;
        RECT 94.160 197.550 94.420 197.810 ;
        RECT 91.860 196.870 92.120 197.130 ;
        RECT 101.980 196.870 102.240 197.130 ;
        RECT 103.820 197.890 104.080 198.150 ;
        RECT 103.820 196.870 104.080 197.130 ;
        RECT 97.840 196.530 98.100 196.790 ;
        RECT 101.520 196.530 101.780 196.790 ;
        RECT 104.740 196.530 105.000 196.790 ;
        RECT 114.400 197.890 114.660 198.150 ;
        RECT 120.380 197.890 120.640 198.150 ;
        RECT 124.980 197.890 125.240 198.150 ;
        RECT 125.900 197.890 126.160 198.150 ;
        RECT 126.820 197.890 127.080 198.150 ;
        RECT 113.940 197.210 114.200 197.470 ;
        RECT 119.000 197.210 119.260 197.470 ;
        RECT 107.960 196.870 108.220 197.130 ;
        RECT 106.580 196.530 106.840 196.790 ;
        RECT 110.260 196.870 110.520 197.130 ;
        RECT 119.460 196.870 119.720 197.130 ;
        RECT 123.140 196.870 123.400 197.130 ;
        RECT 126.360 196.870 126.620 197.130 ;
        RECT 134.640 197.210 134.900 197.470 ;
        RECT 136.480 197.210 136.740 197.470 ;
        RECT 40.800 196.190 41.060 196.450 ;
        RECT 42.640 196.190 42.900 196.450 ;
        RECT 53.220 196.190 53.480 196.450 ;
        RECT 58.740 196.190 59.000 196.450 ;
        RECT 59.200 196.190 59.460 196.450 ;
        RECT 65.180 196.190 65.440 196.450 ;
        RECT 67.020 196.190 67.280 196.450 ;
        RECT 92.780 196.190 93.040 196.450 ;
        RECT 93.700 196.190 93.960 196.450 ;
        RECT 103.360 196.190 103.620 196.450 ;
        RECT 106.120 196.190 106.380 196.450 ;
        RECT 108.420 196.190 108.680 196.450 ;
        RECT 129.120 196.870 129.380 197.130 ;
        RECT 132.800 196.870 133.060 197.130 ;
        RECT 135.100 196.870 135.360 197.130 ;
        RECT 138.780 196.870 139.040 197.130 ;
        RECT 135.560 196.530 135.820 196.790 ;
        RECT 137.860 196.530 138.120 196.790 ;
        RECT 138.320 196.190 138.580 196.450 ;
        RECT 143.840 196.190 144.100 196.450 ;
        RECT 55.170 195.680 55.430 195.940 ;
        RECT 55.490 195.680 55.750 195.940 ;
        RECT 55.810 195.680 56.070 195.940 ;
        RECT 56.130 195.680 56.390 195.940 ;
        RECT 56.450 195.680 56.710 195.940 ;
        RECT 56.770 195.680 57.030 195.940 ;
        RECT 85.170 195.680 85.430 195.940 ;
        RECT 85.490 195.680 85.750 195.940 ;
        RECT 85.810 195.680 86.070 195.940 ;
        RECT 86.130 195.680 86.390 195.940 ;
        RECT 86.450 195.680 86.710 195.940 ;
        RECT 86.770 195.680 87.030 195.940 ;
        RECT 115.170 195.680 115.430 195.940 ;
        RECT 115.490 195.680 115.750 195.940 ;
        RECT 115.810 195.680 116.070 195.940 ;
        RECT 116.130 195.680 116.390 195.940 ;
        RECT 116.450 195.680 116.710 195.940 ;
        RECT 116.770 195.680 117.030 195.940 ;
        RECT 145.170 195.680 145.430 195.940 ;
        RECT 145.490 195.680 145.750 195.940 ;
        RECT 145.810 195.680 146.070 195.940 ;
        RECT 146.130 195.680 146.390 195.940 ;
        RECT 146.450 195.680 146.710 195.940 ;
        RECT 146.770 195.680 147.030 195.940 ;
        RECT 57.820 195.170 58.080 195.430 ;
        RECT 58.740 195.170 59.000 195.430 ;
        RECT 64.260 195.170 64.520 195.430 ;
        RECT 69.320 195.170 69.580 195.430 ;
        RECT 72.540 195.170 72.800 195.430 ;
        RECT 75.760 195.170 76.020 195.430 ;
        RECT 84.500 195.170 84.760 195.430 ;
        RECT 38.500 194.490 38.760 194.750 ;
        RECT 40.800 194.490 41.060 194.750 ;
        RECT 50.000 194.490 50.260 194.750 ;
        RECT 54.140 194.490 54.400 194.750 ;
        RECT 56.900 194.490 57.160 194.750 ;
        RECT 66.560 194.830 66.820 195.090 ;
        RECT 75.300 194.830 75.560 195.090 ;
        RECT 83.120 194.830 83.380 195.090 ;
        RECT 88.640 195.170 88.900 195.430 ;
        RECT 89.560 195.170 89.820 195.430 ;
        RECT 96.000 195.170 96.260 195.430 ;
        RECT 54.600 194.150 54.860 194.410 ;
        RECT 60.120 194.490 60.380 194.750 ;
        RECT 66.100 194.490 66.360 194.750 ;
        RECT 58.280 194.150 58.540 194.410 ;
        RECT 66.560 194.150 66.820 194.410 ;
        RECT 73.920 194.150 74.180 194.410 ;
        RECT 77.600 194.490 77.860 194.750 ;
        RECT 79.440 194.490 79.700 194.750 ;
        RECT 80.360 194.490 80.620 194.750 ;
        RECT 102.440 194.830 102.700 195.090 ;
        RECT 87.720 194.490 87.980 194.750 ;
        RECT 89.100 194.150 89.360 194.410 ;
        RECT 97.380 194.490 97.640 194.750 ;
        RECT 99.220 194.490 99.480 194.750 ;
        RECT 52.760 193.810 53.020 194.070 ;
        RECT 49.540 193.470 49.800 193.730 ;
        RECT 55.060 193.810 55.320 194.070 ;
        RECT 53.680 193.470 53.940 193.730 ;
        RECT 54.600 193.470 54.860 193.730 ;
        RECT 59.200 193.810 59.460 194.070 ;
        RECT 57.360 193.470 57.620 193.730 ;
        RECT 74.380 193.470 74.640 193.730 ;
        RECT 88.640 193.810 88.900 194.070 ;
        RECT 89.560 193.810 89.820 194.070 ;
        RECT 79.440 193.470 79.700 193.730 ;
        RECT 92.780 194.150 93.040 194.410 ;
        RECT 102.900 194.490 103.160 194.750 ;
        RECT 103.820 195.170 104.080 195.430 ;
        RECT 104.740 195.170 105.000 195.430 ;
        RECT 105.660 195.170 105.920 195.430 ;
        RECT 107.960 195.170 108.220 195.430 ;
        RECT 103.820 194.490 104.080 194.750 ;
        RECT 110.260 194.830 110.520 195.090 ;
        RECT 113.940 195.170 114.200 195.430 ;
        RECT 129.120 195.170 129.380 195.430 ;
        RECT 115.320 194.830 115.580 195.090 ;
        RECT 101.520 194.150 101.780 194.410 ;
        RECT 113.940 194.490 114.200 194.750 ;
        RECT 117.160 194.490 117.420 194.750 ;
        RECT 121.300 194.490 121.560 194.750 ;
        RECT 124.520 194.830 124.780 195.090 ;
        RECT 132.800 195.170 133.060 195.430 ;
        RECT 136.020 195.170 136.280 195.430 ;
        RECT 136.480 195.170 136.740 195.430 ;
        RECT 138.320 195.170 138.580 195.430 ;
        RECT 132.340 194.830 132.600 195.090 ;
        RECT 108.880 194.150 109.140 194.410 ;
        RECT 110.260 194.150 110.520 194.410 ;
        RECT 123.140 194.150 123.400 194.410 ;
        RECT 125.440 194.490 125.700 194.750 ;
        RECT 127.280 194.490 127.540 194.750 ;
        RECT 131.880 194.150 132.140 194.410 ;
        RECT 136.480 194.490 136.740 194.750 ;
        RECT 138.780 194.490 139.040 194.750 ;
        RECT 91.400 193.810 91.660 194.070 ;
        RECT 99.680 193.810 99.940 194.070 ;
        RECT 133.720 193.810 133.980 194.070 ;
        RECT 110.720 193.470 110.980 193.730 ;
        RECT 122.220 193.470 122.480 193.730 ;
        RECT 134.640 193.470 134.900 193.730 ;
        RECT 136.940 193.470 137.200 193.730 ;
        RECT 144.760 193.470 145.020 193.730 ;
        RECT 40.170 192.960 40.430 193.220 ;
        RECT 40.490 192.960 40.750 193.220 ;
        RECT 40.810 192.960 41.070 193.220 ;
        RECT 41.130 192.960 41.390 193.220 ;
        RECT 41.450 192.960 41.710 193.220 ;
        RECT 41.770 192.960 42.030 193.220 ;
        RECT 70.170 192.960 70.430 193.220 ;
        RECT 70.490 192.960 70.750 193.220 ;
        RECT 70.810 192.960 71.070 193.220 ;
        RECT 71.130 192.960 71.390 193.220 ;
        RECT 71.450 192.960 71.710 193.220 ;
        RECT 71.770 192.960 72.030 193.220 ;
        RECT 100.170 192.960 100.430 193.220 ;
        RECT 100.490 192.960 100.750 193.220 ;
        RECT 100.810 192.960 101.070 193.220 ;
        RECT 101.130 192.960 101.390 193.220 ;
        RECT 101.450 192.960 101.710 193.220 ;
        RECT 101.770 192.960 102.030 193.220 ;
        RECT 130.170 192.960 130.430 193.220 ;
        RECT 130.490 192.960 130.750 193.220 ;
        RECT 130.810 192.960 131.070 193.220 ;
        RECT 131.130 192.960 131.390 193.220 ;
        RECT 131.450 192.960 131.710 193.220 ;
        RECT 131.770 192.960 132.030 193.220 ;
        RECT 42.180 192.450 42.440 192.710 ;
        RECT 51.840 192.450 52.100 192.710 ;
        RECT 42.180 191.770 42.440 192.030 ;
        RECT 42.640 191.430 42.900 191.690 ;
        RECT 50.920 191.430 51.180 191.690 ;
        RECT 53.680 191.430 53.940 191.690 ;
        RECT 54.140 191.430 54.400 191.690 ;
        RECT 59.660 192.450 59.920 192.710 ;
        RECT 66.560 192.450 66.820 192.710 ;
        RECT 75.300 192.450 75.560 192.710 ;
        RECT 77.600 192.450 77.860 192.710 ;
        RECT 80.820 192.450 81.080 192.710 ;
        RECT 87.720 192.450 87.980 192.710 ;
        RECT 90.020 192.450 90.280 192.710 ;
        RECT 57.360 192.110 57.620 192.370 ;
        RECT 59.200 191.770 59.460 192.030 ;
        RECT 61.040 191.770 61.300 192.030 ;
        RECT 57.360 191.430 57.620 191.690 ;
        RECT 73.920 192.110 74.180 192.370 ;
        RECT 65.640 191.770 65.900 192.030 ;
        RECT 67.480 191.770 67.740 192.030 ;
        RECT 65.180 191.430 65.440 191.690 ;
        RECT 67.940 191.430 68.200 191.690 ;
        RECT 75.760 191.430 76.020 191.690 ;
        RECT 78.060 191.770 78.320 192.030 ;
        RECT 52.300 190.750 52.560 191.010 ;
        RECT 61.960 191.090 62.220 191.350 ;
        RECT 62.420 191.090 62.680 191.350 ;
        RECT 61.040 190.750 61.300 191.010 ;
        RECT 75.760 190.750 76.020 191.010 ;
        RECT 77.600 191.430 77.860 191.690 ;
        RECT 88.640 192.110 88.900 192.370 ;
        RECT 83.120 191.770 83.380 192.030 ;
        RECT 96.460 192.450 96.720 192.710 ;
        RECT 99.220 192.450 99.480 192.710 ;
        RECT 112.560 192.450 112.820 192.710 ;
        RECT 115.320 192.450 115.580 192.710 ;
        RECT 124.520 192.450 124.780 192.710 ;
        RECT 132.340 192.450 132.600 192.710 ;
        RECT 132.800 192.450 133.060 192.710 ;
        RECT 89.100 191.430 89.360 191.690 ;
        RECT 90.480 191.430 90.740 191.690 ;
        RECT 79.440 191.090 79.700 191.350 ;
        RECT 80.360 191.090 80.620 191.350 ;
        RECT 92.320 191.430 92.580 191.690 ;
        RECT 97.380 191.770 97.640 192.030 ;
        RECT 94.160 191.430 94.420 191.690 ;
        RECT 95.540 191.430 95.800 191.690 ;
        RECT 98.300 191.430 98.560 191.690 ;
        RECT 90.020 190.750 90.280 191.010 ;
        RECT 90.480 190.750 90.740 191.010 ;
        RECT 99.220 191.430 99.480 191.690 ;
        RECT 102.900 192.110 103.160 192.370 ;
        RECT 102.440 191.770 102.700 192.030 ;
        RECT 101.980 191.430 102.240 191.690 ;
        RECT 102.900 191.430 103.160 191.690 ;
        RECT 103.820 191.430 104.080 191.690 ;
        RECT 104.280 191.430 104.540 191.690 ;
        RECT 106.120 191.430 106.380 191.690 ;
        RECT 106.580 191.430 106.840 191.690 ;
        RECT 110.260 191.770 110.520 192.030 ;
        RECT 118.540 191.770 118.800 192.030 ;
        RECT 137.860 192.450 138.120 192.710 ;
        RECT 109.800 191.430 110.060 191.690 ;
        RECT 113.940 191.430 114.200 191.690 ;
        RECT 114.400 191.430 114.660 191.690 ;
        RECT 102.440 191.090 102.700 191.350 ;
        RECT 117.160 191.430 117.420 191.690 ;
        RECT 119.000 191.430 119.260 191.690 ;
        RECT 121.300 191.430 121.560 191.690 ;
        RECT 130.040 191.430 130.300 191.690 ;
        RECT 134.640 191.770 134.900 192.030 ;
        RECT 143.840 191.770 144.100 192.030 ;
        RECT 99.220 190.750 99.480 191.010 ;
        RECT 105.660 190.750 105.920 191.010 ;
        RECT 110.260 190.750 110.520 191.010 ;
        RECT 119.460 190.750 119.720 191.010 ;
        RECT 125.900 190.750 126.160 191.010 ;
        RECT 132.340 190.750 132.600 191.010 ;
        RECT 133.260 190.750 133.520 191.010 ;
        RECT 136.940 191.430 137.200 191.690 ;
        RECT 137.400 191.430 137.660 191.690 ;
        RECT 144.760 191.430 145.020 191.690 ;
        RECT 147.520 191.770 147.780 192.030 ;
        RECT 142.460 190.750 142.720 191.010 ;
        RECT 147.980 190.750 148.240 191.010 ;
        RECT 55.170 190.240 55.430 190.500 ;
        RECT 55.490 190.240 55.750 190.500 ;
        RECT 55.810 190.240 56.070 190.500 ;
        RECT 56.130 190.240 56.390 190.500 ;
        RECT 56.450 190.240 56.710 190.500 ;
        RECT 56.770 190.240 57.030 190.500 ;
        RECT 85.170 190.240 85.430 190.500 ;
        RECT 85.490 190.240 85.750 190.500 ;
        RECT 85.810 190.240 86.070 190.500 ;
        RECT 86.130 190.240 86.390 190.500 ;
        RECT 86.450 190.240 86.710 190.500 ;
        RECT 86.770 190.240 87.030 190.500 ;
        RECT 115.170 190.240 115.430 190.500 ;
        RECT 115.490 190.240 115.750 190.500 ;
        RECT 115.810 190.240 116.070 190.500 ;
        RECT 116.130 190.240 116.390 190.500 ;
        RECT 116.450 190.240 116.710 190.500 ;
        RECT 116.770 190.240 117.030 190.500 ;
        RECT 145.170 190.240 145.430 190.500 ;
        RECT 145.490 190.240 145.750 190.500 ;
        RECT 145.810 190.240 146.070 190.500 ;
        RECT 146.130 190.240 146.390 190.500 ;
        RECT 146.450 190.240 146.710 190.500 ;
        RECT 146.770 190.240 147.030 190.500 ;
        RECT 42.180 189.730 42.440 189.990 ;
        RECT 41.720 189.050 41.980 189.310 ;
        RECT 44.020 189.730 44.280 189.990 ;
        RECT 46.780 189.390 47.040 189.650 ;
        RECT 49.540 189.390 49.800 189.650 ;
        RECT 67.020 189.730 67.280 189.990 ;
        RECT 73.920 189.730 74.180 189.990 ;
        RECT 75.760 189.730 76.020 189.990 ;
        RECT 39.420 188.710 39.680 188.970 ;
        RECT 38.960 188.030 39.220 188.290 ;
        RECT 43.560 188.030 43.820 188.290 ;
        RECT 46.320 189.050 46.580 189.310 ;
        RECT 50.000 189.050 50.260 189.310 ;
        RECT 54.600 189.050 54.860 189.310 ;
        RECT 61.040 189.390 61.300 189.650 ;
        RECT 72.540 189.050 72.800 189.310 ;
        RECT 74.840 189.050 75.100 189.310 ;
        RECT 76.680 189.050 76.940 189.310 ;
        RECT 77.600 189.390 77.860 189.650 ;
        RECT 78.520 189.050 78.780 189.310 ;
        RECT 47.240 188.370 47.500 188.630 ;
        RECT 47.700 188.370 47.960 188.630 ;
        RECT 63.340 188.370 63.600 188.630 ;
        RECT 64.260 188.370 64.520 188.630 ;
        RECT 83.120 189.050 83.380 189.310 ;
        RECT 88.640 189.730 88.900 189.990 ;
        RECT 79.900 188.710 80.160 188.970 ;
        RECT 88.180 189.050 88.440 189.310 ;
        RECT 90.480 189.730 90.740 189.990 ;
        RECT 91.860 189.730 92.120 189.990 ;
        RECT 101.980 189.730 102.240 189.990 ;
        RECT 103.820 189.730 104.080 189.990 ;
        RECT 109.800 189.730 110.060 189.990 ;
        RECT 117.160 189.730 117.420 189.990 ;
        RECT 119.000 189.730 119.260 189.990 ;
        RECT 126.820 189.730 127.080 189.990 ;
        RECT 128.660 189.730 128.920 189.990 ;
        RECT 130.040 189.730 130.300 189.990 ;
        RECT 134.180 189.730 134.440 189.990 ;
        RECT 141.080 189.730 141.340 189.990 ;
        RECT 144.300 189.730 144.560 189.990 ;
        RECT 89.560 189.050 89.820 189.310 ;
        RECT 90.020 189.050 90.280 189.310 ;
        RECT 96.460 189.390 96.720 189.650 ;
        RECT 88.640 188.710 88.900 188.970 ;
        RECT 79.440 188.370 79.700 188.630 ;
        RECT 98.300 189.050 98.560 189.310 ;
        RECT 99.220 189.050 99.480 189.310 ;
        RECT 107.040 189.390 107.300 189.650 ;
        RECT 96.920 188.710 97.180 188.970 ;
        RECT 103.360 189.050 103.620 189.310 ;
        RECT 104.740 189.050 105.000 189.310 ;
        RECT 105.660 189.050 105.920 189.310 ;
        RECT 113.480 189.050 113.740 189.310 ;
        RECT 116.700 189.050 116.960 189.310 ;
        RECT 117.620 189.050 117.880 189.310 ;
        RECT 111.180 188.710 111.440 188.970 ;
        RECT 114.400 188.710 114.660 188.970 ;
        RECT 116.240 188.710 116.500 188.970 ;
        RECT 119.920 188.710 120.180 188.970 ;
        RECT 120.840 189.050 121.100 189.310 ;
        RECT 122.220 189.050 122.480 189.310 ;
        RECT 124.980 189.050 125.240 189.310 ;
        RECT 130.040 188.710 130.300 188.970 ;
        RECT 132.340 189.050 132.600 189.310 ;
        RECT 132.800 188.710 133.060 188.970 ;
        RECT 133.720 188.710 133.980 188.970 ;
        RECT 92.320 188.370 92.580 188.630 ;
        RECT 49.080 188.030 49.340 188.290 ;
        RECT 53.680 188.030 53.940 188.290 ;
        RECT 56.900 188.030 57.160 188.290 ;
        RECT 61.040 188.030 61.300 188.290 ;
        RECT 65.640 188.030 65.900 188.290 ;
        RECT 69.780 188.030 70.040 188.290 ;
        RECT 73.000 188.030 73.260 188.290 ;
        RECT 74.840 188.030 75.100 188.290 ;
        RECT 76.680 188.030 76.940 188.290 ;
        RECT 77.600 188.030 77.860 188.290 ;
        RECT 82.200 188.030 82.460 188.290 ;
        RECT 83.120 188.030 83.380 188.290 ;
        RECT 87.720 188.030 87.980 188.290 ;
        RECT 139.240 188.370 139.500 188.630 ;
        RECT 102.900 188.030 103.160 188.290 ;
        RECT 106.580 188.030 106.840 188.290 ;
        RECT 107.040 188.030 107.300 188.290 ;
        RECT 113.940 188.030 114.200 188.290 ;
        RECT 117.160 188.030 117.420 188.290 ;
        RECT 129.580 188.030 129.840 188.290 ;
        RECT 134.640 188.030 134.900 188.290 ;
        RECT 136.480 188.030 136.740 188.290 ;
        RECT 141.540 189.050 141.800 189.310 ;
        RECT 141.080 188.710 141.340 188.970 ;
        RECT 142.000 188.710 142.260 188.970 ;
        RECT 144.300 188.710 144.560 188.970 ;
        RECT 145.680 189.050 145.940 189.310 ;
        RECT 147.060 188.030 147.320 188.290 ;
        RECT 40.170 187.520 40.430 187.780 ;
        RECT 40.490 187.520 40.750 187.780 ;
        RECT 40.810 187.520 41.070 187.780 ;
        RECT 41.130 187.520 41.390 187.780 ;
        RECT 41.450 187.520 41.710 187.780 ;
        RECT 41.770 187.520 42.030 187.780 ;
        RECT 70.170 187.520 70.430 187.780 ;
        RECT 70.490 187.520 70.750 187.780 ;
        RECT 70.810 187.520 71.070 187.780 ;
        RECT 71.130 187.520 71.390 187.780 ;
        RECT 71.450 187.520 71.710 187.780 ;
        RECT 71.770 187.520 72.030 187.780 ;
        RECT 100.170 187.520 100.430 187.780 ;
        RECT 100.490 187.520 100.750 187.780 ;
        RECT 100.810 187.520 101.070 187.780 ;
        RECT 101.130 187.520 101.390 187.780 ;
        RECT 101.450 187.520 101.710 187.780 ;
        RECT 101.770 187.520 102.030 187.780 ;
        RECT 130.170 187.520 130.430 187.780 ;
        RECT 130.490 187.520 130.750 187.780 ;
        RECT 130.810 187.520 131.070 187.780 ;
        RECT 131.130 187.520 131.390 187.780 ;
        RECT 131.450 187.520 131.710 187.780 ;
        RECT 131.770 187.520 132.030 187.780 ;
        RECT 46.320 187.010 46.580 187.270 ;
        RECT 49.540 187.010 49.800 187.270 ;
        RECT 44.940 185.990 45.200 186.250 ;
        RECT 45.400 185.990 45.660 186.250 ;
        RECT 52.760 186.330 53.020 186.590 ;
        RECT 61.040 187.010 61.300 187.270 ;
        RECT 67.940 187.010 68.200 187.270 ;
        RECT 91.400 187.010 91.660 187.270 ;
        RECT 93.240 187.010 93.500 187.270 ;
        RECT 107.040 187.010 107.300 187.270 ;
        RECT 60.580 186.670 60.840 186.930 ;
        RECT 49.080 185.990 49.340 186.250 ;
        RECT 49.540 185.990 49.800 186.250 ;
        RECT 50.920 185.990 51.180 186.250 ;
        RECT 54.140 185.990 54.400 186.250 ;
        RECT 56.900 185.990 57.160 186.250 ;
        RECT 58.280 185.990 58.540 186.250 ;
        RECT 52.760 185.650 53.020 185.910 ;
        RECT 44.480 185.310 44.740 185.570 ;
        RECT 49.080 185.310 49.340 185.570 ;
        RECT 59.660 185.990 59.920 186.250 ;
        RECT 69.780 186.330 70.040 186.590 ;
        RECT 62.880 185.990 63.140 186.250 ;
        RECT 65.640 185.990 65.900 186.250 ;
        RECT 60.120 185.650 60.380 185.910 ;
        RECT 73.920 185.990 74.180 186.250 ;
        RECT 94.160 186.330 94.420 186.590 ;
        RECT 78.060 185.990 78.320 186.250 ;
        RECT 81.740 185.990 82.000 186.250 ;
        RECT 84.500 185.990 84.760 186.250 ;
        RECT 95.540 186.330 95.800 186.590 ;
        RECT 97.840 186.330 98.100 186.590 ;
        RECT 98.760 186.330 99.020 186.590 ;
        RECT 99.220 186.330 99.480 186.590 ;
        RECT 100.600 186.330 100.860 186.590 ;
        RECT 103.360 186.330 103.620 186.590 ;
        RECT 63.340 185.650 63.600 185.910 ;
        RECT 66.100 185.650 66.360 185.910 ;
        RECT 73.000 185.650 73.260 185.910 ;
        RECT 77.600 185.650 77.860 185.910 ;
        RECT 62.880 185.310 63.140 185.570 ;
        RECT 87.260 185.650 87.520 185.910 ;
        RECT 101.980 185.990 102.240 186.250 ;
        RECT 108.420 186.670 108.680 186.930 ;
        RECT 117.160 187.010 117.420 187.270 ;
        RECT 118.540 187.010 118.800 187.270 ;
        RECT 121.760 187.010 122.020 187.270 ;
        RECT 98.760 185.650 99.020 185.910 ;
        RECT 104.280 185.650 104.540 185.910 ;
        RECT 111.180 185.990 111.440 186.250 ;
        RECT 113.020 186.330 113.280 186.590 ;
        RECT 124.980 186.670 125.240 186.930 ;
        RECT 136.480 187.010 136.740 187.270 ;
        RECT 139.240 187.010 139.500 187.270 ;
        RECT 140.160 187.010 140.420 187.270 ;
        RECT 143.840 187.010 144.100 187.270 ;
        RECT 144.300 187.010 144.560 187.270 ;
        RECT 111.640 185.650 111.900 185.910 ;
        RECT 82.200 185.310 82.460 185.570 ;
        RECT 88.180 185.310 88.440 185.570 ;
        RECT 90.020 185.310 90.280 185.570 ;
        RECT 112.560 185.310 112.820 185.570 ;
        RECT 116.700 185.990 116.960 186.250 ;
        RECT 122.680 185.990 122.940 186.250 ;
        RECT 126.360 186.330 126.620 186.590 ;
        RECT 129.120 186.330 129.380 186.590 ;
        RECT 132.800 186.670 133.060 186.930 ;
        RECT 136.020 186.670 136.280 186.930 ;
        RECT 133.720 186.330 133.980 186.590 ;
        RECT 143.380 186.670 143.640 186.930 ;
        RECT 145.680 187.010 145.940 187.270 ;
        RECT 117.620 185.650 117.880 185.910 ;
        RECT 117.160 185.310 117.420 185.570 ;
        RECT 119.460 185.310 119.720 185.570 ;
        RECT 121.760 185.310 122.020 185.570 ;
        RECT 122.220 185.310 122.480 185.570 ;
        RECT 126.820 185.650 127.080 185.910 ;
        RECT 124.060 185.310 124.320 185.570 ;
        RECT 127.280 185.310 127.540 185.570 ;
        RECT 127.740 185.310 128.000 185.570 ;
        RECT 130.960 185.650 131.220 185.910 ;
        RECT 132.800 185.820 133.060 186.080 ;
        RECT 137.400 185.990 137.660 186.250 ;
        RECT 138.780 185.990 139.040 186.250 ;
        RECT 133.260 185.310 133.520 185.570 ;
        RECT 136.940 185.310 137.200 185.570 ;
        RECT 141.540 185.990 141.800 186.250 ;
        RECT 144.300 185.990 144.560 186.250 ;
        RECT 147.520 185.990 147.780 186.250 ;
        RECT 143.840 185.650 144.100 185.910 ;
        RECT 147.060 185.650 147.320 185.910 ;
        RECT 141.540 185.310 141.800 185.570 ;
        RECT 143.380 185.310 143.640 185.570 ;
        RECT 55.170 184.800 55.430 185.060 ;
        RECT 55.490 184.800 55.750 185.060 ;
        RECT 55.810 184.800 56.070 185.060 ;
        RECT 56.130 184.800 56.390 185.060 ;
        RECT 56.450 184.800 56.710 185.060 ;
        RECT 56.770 184.800 57.030 185.060 ;
        RECT 85.170 184.800 85.430 185.060 ;
        RECT 85.490 184.800 85.750 185.060 ;
        RECT 85.810 184.800 86.070 185.060 ;
        RECT 86.130 184.800 86.390 185.060 ;
        RECT 86.450 184.800 86.710 185.060 ;
        RECT 86.770 184.800 87.030 185.060 ;
        RECT 115.170 184.800 115.430 185.060 ;
        RECT 115.490 184.800 115.750 185.060 ;
        RECT 115.810 184.800 116.070 185.060 ;
        RECT 116.130 184.800 116.390 185.060 ;
        RECT 116.450 184.800 116.710 185.060 ;
        RECT 116.770 184.800 117.030 185.060 ;
        RECT 145.170 184.800 145.430 185.060 ;
        RECT 145.490 184.800 145.750 185.060 ;
        RECT 145.810 184.800 146.070 185.060 ;
        RECT 146.130 184.800 146.390 185.060 ;
        RECT 146.450 184.800 146.710 185.060 ;
        RECT 146.770 184.800 147.030 185.060 ;
        RECT 50.920 184.290 51.180 184.550 ;
        RECT 44.020 183.610 44.280 183.870 ;
        RECT 44.480 183.610 44.740 183.870 ;
        RECT 45.400 183.610 45.660 183.870 ;
        RECT 46.320 183.610 46.580 183.870 ;
        RECT 51.380 183.950 51.640 184.210 ;
        RECT 49.540 183.610 49.800 183.870 ;
        RECT 59.660 184.290 59.920 184.550 ;
        RECT 78.060 184.290 78.320 184.550 ;
        RECT 78.980 184.290 79.240 184.550 ;
        RECT 62.420 183.950 62.680 184.210 ;
        RECT 50.000 182.930 50.260 183.190 ;
        RECT 51.380 183.270 51.640 183.530 ;
        RECT 53.680 183.610 53.940 183.870 ;
        RECT 58.280 183.610 58.540 183.870 ;
        RECT 58.740 183.610 59.000 183.870 ;
        RECT 61.040 183.610 61.300 183.870 ;
        RECT 67.480 183.610 67.740 183.870 ;
        RECT 54.600 183.270 54.860 183.530 ;
        RECT 59.660 183.270 59.920 183.530 ;
        RECT 66.560 183.270 66.820 183.530 ;
        RECT 61.500 182.930 61.760 183.190 ;
        RECT 63.800 182.930 64.060 183.190 ;
        RECT 80.360 183.610 80.620 183.870 ;
        RECT 81.740 183.950 82.000 184.210 ;
        RECT 82.200 182.930 82.460 183.190 ;
        RECT 84.960 184.290 85.220 184.550 ;
        RECT 87.260 184.290 87.520 184.550 ;
        RECT 88.180 183.610 88.440 183.870 ;
        RECT 89.560 183.610 89.820 183.870 ;
        RECT 91.400 183.270 91.660 183.530 ;
        RECT 84.500 182.930 84.760 183.190 ;
        RECT 92.320 183.610 92.580 183.870 ;
        RECT 93.240 183.610 93.500 183.870 ;
        RECT 95.080 183.950 95.340 184.210 ;
        RECT 95.540 183.610 95.800 183.870 ;
        RECT 96.920 183.610 97.180 183.870 ;
        RECT 97.380 183.610 97.640 183.870 ;
        RECT 98.300 183.950 98.560 184.210 ;
        RECT 100.600 184.290 100.860 184.550 ;
        RECT 101.980 184.290 102.240 184.550 ;
        RECT 110.720 184.290 110.980 184.550 ;
        RECT 111.180 184.290 111.440 184.550 ;
        RECT 122.220 184.290 122.480 184.550 ;
        RECT 98.760 183.610 99.020 183.870 ;
        RECT 101.520 183.610 101.780 183.870 ;
        RECT 93.700 183.270 93.960 183.530 ;
        RECT 102.900 183.610 103.160 183.870 ;
        RECT 46.780 182.590 47.040 182.850 ;
        RECT 47.240 182.590 47.500 182.850 ;
        RECT 49.080 182.590 49.340 182.850 ;
        RECT 52.300 182.590 52.560 182.850 ;
        RECT 52.760 182.590 53.020 182.850 ;
        RECT 62.880 182.590 63.140 182.850 ;
        RECT 76.680 182.590 76.940 182.850 ;
        RECT 79.900 182.590 80.160 182.850 ;
        RECT 90.480 182.590 90.740 182.850 ;
        RECT 92.320 182.590 92.580 182.850 ;
        RECT 94.620 182.590 94.880 182.850 ;
        RECT 95.080 182.590 95.340 182.850 ;
        RECT 99.220 182.590 99.480 182.850 ;
        RECT 102.900 182.930 103.160 183.190 ;
        RECT 104.740 183.610 105.000 183.870 ;
        RECT 106.580 183.270 106.840 183.530 ;
        RECT 109.800 183.610 110.060 183.870 ;
        RECT 108.420 183.270 108.680 183.530 ;
        RECT 107.960 182.930 108.220 183.190 ;
        RECT 105.660 182.590 105.920 182.850 ;
        RECT 107.500 182.590 107.760 182.850 ;
        RECT 117.160 183.950 117.420 184.210 ;
        RECT 121.300 183.950 121.560 184.210 ;
        RECT 122.680 183.950 122.940 184.210 ;
        RECT 127.280 184.290 127.540 184.550 ;
        RECT 135.560 184.290 135.820 184.550 ;
        RECT 142.000 184.290 142.260 184.550 ;
        RECT 144.300 184.290 144.560 184.550 ;
        RECT 127.740 183.950 128.000 184.210 ;
        RECT 124.980 183.610 125.240 183.870 ;
        RECT 125.900 183.610 126.160 183.870 ;
        RECT 129.120 183.610 129.380 183.870 ;
        RECT 133.720 183.950 133.980 184.210 ;
        RECT 140.620 183.950 140.880 184.210 ;
        RECT 130.040 183.610 130.300 183.870 ;
        RECT 132.340 183.610 132.600 183.870 ;
        RECT 133.260 183.610 133.520 183.870 ;
        RECT 138.320 183.610 138.580 183.870 ;
        RECT 119.460 183.270 119.720 183.530 ;
        RECT 112.100 182.590 112.360 182.850 ;
        RECT 113.020 182.590 113.280 182.850 ;
        RECT 116.700 182.590 116.960 182.850 ;
        RECT 124.060 182.930 124.320 183.190 ;
        RECT 127.280 182.930 127.540 183.190 ;
        RECT 128.660 182.930 128.920 183.190 ;
        RECT 131.880 183.270 132.140 183.530 ;
        RECT 134.180 183.270 134.440 183.530 ;
        RECT 137.860 183.270 138.120 183.530 ;
        RECT 121.760 182.590 122.020 182.850 ;
        RECT 122.220 182.590 122.480 182.850 ;
        RECT 130.040 182.590 130.300 182.850 ;
        RECT 132.800 182.590 133.060 182.850 ;
        RECT 134.640 182.590 134.900 182.850 ;
        RECT 138.320 182.590 138.580 182.850 ;
        RECT 40.170 182.080 40.430 182.340 ;
        RECT 40.490 182.080 40.750 182.340 ;
        RECT 40.810 182.080 41.070 182.340 ;
        RECT 41.130 182.080 41.390 182.340 ;
        RECT 41.450 182.080 41.710 182.340 ;
        RECT 41.770 182.080 42.030 182.340 ;
        RECT 70.170 182.080 70.430 182.340 ;
        RECT 70.490 182.080 70.750 182.340 ;
        RECT 70.810 182.080 71.070 182.340 ;
        RECT 71.130 182.080 71.390 182.340 ;
        RECT 71.450 182.080 71.710 182.340 ;
        RECT 71.770 182.080 72.030 182.340 ;
        RECT 100.170 182.080 100.430 182.340 ;
        RECT 100.490 182.080 100.750 182.340 ;
        RECT 100.810 182.080 101.070 182.340 ;
        RECT 101.130 182.080 101.390 182.340 ;
        RECT 101.450 182.080 101.710 182.340 ;
        RECT 101.770 182.080 102.030 182.340 ;
        RECT 130.170 182.080 130.430 182.340 ;
        RECT 130.490 182.080 130.750 182.340 ;
        RECT 130.810 182.080 131.070 182.340 ;
        RECT 131.130 182.080 131.390 182.340 ;
        RECT 131.450 182.080 131.710 182.340 ;
        RECT 131.770 182.080 132.030 182.340 ;
        RECT 44.940 181.570 45.200 181.830 ;
        RECT 46.320 181.570 46.580 181.830 ;
        RECT 48.620 181.570 48.880 181.830 ;
        RECT 50.460 181.570 50.720 181.830 ;
        RECT 51.840 181.570 52.100 181.830 ;
        RECT 87.720 181.570 87.980 181.830 ;
        RECT 92.320 181.570 92.580 181.830 ;
        RECT 94.620 181.570 94.880 181.830 ;
        RECT 97.840 181.570 98.100 181.830 ;
        RECT 108.420 181.570 108.680 181.830 ;
        RECT 83.120 181.230 83.380 181.490 ;
        RECT 88.640 181.230 88.900 181.490 ;
        RECT 90.940 181.230 91.200 181.490 ;
        RECT 49.540 180.890 49.800 181.150 ;
        RECT 50.000 180.550 50.260 180.810 ;
        RECT 55.060 180.890 55.320 181.150 ;
        RECT 61.040 180.890 61.300 181.150 ;
        RECT 61.500 180.890 61.760 181.150 ;
        RECT 76.680 180.890 76.940 181.150 ;
        RECT 81.740 180.890 82.000 181.150 ;
        RECT 46.780 180.210 47.040 180.470 ;
        RECT 44.480 179.870 44.740 180.130 ;
        RECT 54.140 180.210 54.400 180.470 ;
        RECT 50.000 179.870 50.260 180.130 ;
        RECT 52.300 179.870 52.560 180.130 ;
        RECT 53.680 179.870 53.940 180.130 ;
        RECT 58.740 180.550 59.000 180.810 ;
        RECT 59.200 180.550 59.460 180.810 ;
        RECT 64.720 180.550 64.980 180.810 ;
        RECT 67.020 180.550 67.280 180.810 ;
        RECT 78.980 180.550 79.240 180.810 ;
        RECT 93.240 180.890 93.500 181.150 ;
        RECT 62.880 180.210 63.140 180.470 ;
        RECT 65.640 180.210 65.900 180.470 ;
        RECT 79.900 180.210 80.160 180.470 ;
        RECT 88.640 180.210 88.900 180.470 ;
        RECT 90.020 180.550 90.280 180.810 ;
        RECT 90.940 180.550 91.200 180.810 ;
        RECT 92.780 180.550 93.040 180.810 ;
        RECT 106.580 181.230 106.840 181.490 ;
        RECT 107.500 181.230 107.760 181.490 ;
        RECT 107.960 181.230 108.220 181.490 ;
        RECT 112.560 181.570 112.820 181.830 ;
        RECT 117.160 181.570 117.420 181.830 ;
        RECT 119.460 181.570 119.720 181.830 ;
        RECT 119.920 181.570 120.180 181.830 ;
        RECT 121.300 181.570 121.560 181.830 ;
        RECT 125.440 181.570 125.700 181.830 ;
        RECT 127.740 181.570 128.000 181.830 ;
        RECT 128.660 181.570 128.920 181.830 ;
        RECT 129.580 181.570 129.840 181.830 ;
        RECT 132.340 181.570 132.600 181.830 ;
        RECT 133.720 181.570 133.980 181.830 ;
        RECT 136.940 181.570 137.200 181.830 ;
        RECT 140.160 181.570 140.420 181.830 ;
        RECT 143.380 181.570 143.640 181.830 ;
        RECT 96.000 180.890 96.260 181.150 ;
        RECT 99.220 180.890 99.480 181.150 ;
        RECT 100.140 180.890 100.400 181.150 ;
        RECT 103.820 180.890 104.080 181.150 ;
        RECT 105.660 180.890 105.920 181.150 ;
        RECT 110.260 180.890 110.520 181.150 ;
        RECT 97.840 180.210 98.100 180.470 ;
        RECT 110.720 180.550 110.980 180.810 ;
        RECT 113.480 180.550 113.740 180.810 ;
        RECT 117.620 180.890 117.880 181.150 ;
        RECT 101.980 180.210 102.240 180.470 ;
        RECT 103.360 180.210 103.620 180.470 ;
        RECT 105.660 180.210 105.920 180.470 ;
        RECT 55.060 179.870 55.320 180.130 ;
        RECT 63.340 179.870 63.600 180.130 ;
        RECT 68.400 179.870 68.660 180.130 ;
        RECT 91.860 179.870 92.120 180.130 ;
        RECT 96.000 179.870 96.260 180.130 ;
        RECT 97.380 179.870 97.640 180.130 ;
        RECT 98.760 179.870 99.020 180.130 ;
        RECT 99.220 179.870 99.480 180.130 ;
        RECT 104.280 179.870 104.540 180.130 ;
        RECT 109.800 179.870 110.060 180.130 ;
        RECT 116.240 180.550 116.500 180.810 ;
        RECT 116.700 180.550 116.960 180.810 ;
        RECT 119.920 180.550 120.180 180.810 ;
        RECT 121.760 180.550 122.020 180.810 ;
        RECT 122.680 180.550 122.940 180.810 ;
        RECT 130.040 180.550 130.300 180.810 ;
        RECT 133.260 181.230 133.520 181.490 ;
        RECT 140.620 181.230 140.880 181.490 ;
        RECT 139.700 180.890 139.960 181.150 ;
        RECT 141.540 180.890 141.800 181.150 ;
        RECT 136.020 180.550 136.280 180.810 ;
        RECT 140.160 180.550 140.420 180.810 ;
        RECT 147.980 180.890 148.240 181.150 ;
        RECT 133.260 180.210 133.520 180.470 ;
        RECT 134.640 180.210 134.900 180.470 ;
        RECT 139.240 180.210 139.500 180.470 ;
        RECT 139.700 180.210 139.960 180.470 ;
        RECT 121.300 179.870 121.560 180.130 ;
        RECT 126.820 179.870 127.080 180.130 ;
        RECT 132.340 179.870 132.600 180.130 ;
        RECT 55.170 179.360 55.430 179.620 ;
        RECT 55.490 179.360 55.750 179.620 ;
        RECT 55.810 179.360 56.070 179.620 ;
        RECT 56.130 179.360 56.390 179.620 ;
        RECT 56.450 179.360 56.710 179.620 ;
        RECT 56.770 179.360 57.030 179.620 ;
        RECT 85.170 179.360 85.430 179.620 ;
        RECT 85.490 179.360 85.750 179.620 ;
        RECT 85.810 179.360 86.070 179.620 ;
        RECT 86.130 179.360 86.390 179.620 ;
        RECT 86.450 179.360 86.710 179.620 ;
        RECT 86.770 179.360 87.030 179.620 ;
        RECT 115.170 179.360 115.430 179.620 ;
        RECT 115.490 179.360 115.750 179.620 ;
        RECT 115.810 179.360 116.070 179.620 ;
        RECT 116.130 179.360 116.390 179.620 ;
        RECT 116.450 179.360 116.710 179.620 ;
        RECT 116.770 179.360 117.030 179.620 ;
        RECT 145.170 179.360 145.430 179.620 ;
        RECT 145.490 179.360 145.750 179.620 ;
        RECT 145.810 179.360 146.070 179.620 ;
        RECT 146.130 179.360 146.390 179.620 ;
        RECT 146.450 179.360 146.710 179.620 ;
        RECT 146.770 179.360 147.030 179.620 ;
        RECT 44.480 178.850 44.740 179.110 ;
        RECT 38.960 178.170 39.220 178.430 ;
        RECT 46.780 178.170 47.040 178.430 ;
        RECT 50.460 178.850 50.720 179.110 ;
        RECT 50.920 178.850 51.180 179.110 ;
        RECT 53.680 178.850 53.940 179.110 ;
        RECT 58.280 178.850 58.540 179.110 ;
        RECT 58.740 178.850 59.000 179.110 ;
        RECT 59.200 178.850 59.460 179.110 ;
        RECT 63.340 178.850 63.600 179.110 ;
        RECT 63.800 178.850 64.060 179.110 ;
        RECT 92.780 178.850 93.040 179.110 ;
        RECT 95.540 178.850 95.800 179.110 ;
        RECT 101.980 178.850 102.240 179.110 ;
        RECT 102.440 178.850 102.700 179.110 ;
        RECT 50.000 178.510 50.260 178.770 ;
        RECT 37.580 177.830 37.840 178.090 ;
        RECT 48.620 177.830 48.880 178.090 ;
        RECT 50.920 178.170 51.180 178.430 ;
        RECT 49.080 177.490 49.340 177.750 ;
        RECT 64.260 178.510 64.520 178.770 ;
        RECT 66.560 178.510 66.820 178.770 ;
        RECT 90.940 178.510 91.200 178.770 ;
        RECT 53.220 177.490 53.480 177.750 ;
        RECT 67.480 178.170 67.740 178.430 ;
        RECT 79.900 178.170 80.160 178.430 ;
        RECT 84.500 178.170 84.760 178.430 ;
        RECT 89.100 178.170 89.360 178.430 ;
        RECT 89.560 178.170 89.820 178.430 ;
        RECT 96.000 178.510 96.260 178.770 ;
        RECT 95.080 178.170 95.340 178.430 ;
        RECT 96.920 178.170 97.180 178.430 ;
        RECT 99.680 178.170 99.940 178.430 ;
        RECT 103.360 178.170 103.620 178.430 ;
        RECT 103.820 178.170 104.080 178.430 ;
        RECT 104.280 178.170 104.540 178.430 ;
        RECT 107.500 178.850 107.760 179.110 ;
        RECT 107.960 178.850 108.220 179.110 ;
        RECT 118.540 178.850 118.800 179.110 ;
        RECT 61.500 177.830 61.760 178.090 ;
        RECT 77.600 177.830 77.860 178.090 ;
        RECT 99.220 177.830 99.480 178.090 ;
        RECT 106.580 178.170 106.840 178.430 ;
        RECT 109.800 178.170 110.060 178.430 ;
        RECT 120.840 178.510 121.100 178.770 ;
        RECT 110.720 177.830 110.980 178.090 ;
        RECT 54.140 177.150 54.400 177.410 ;
        RECT 60.120 177.150 60.380 177.410 ;
        RECT 63.340 177.150 63.600 177.410 ;
        RECT 69.320 177.150 69.580 177.410 ;
        RECT 69.780 177.150 70.040 177.410 ;
        RECT 89.100 177.490 89.360 177.750 ;
        RECT 91.400 177.490 91.660 177.750 ;
        RECT 93.240 177.150 93.500 177.410 ;
        RECT 126.820 178.170 127.080 178.430 ;
        RECT 132.340 178.170 132.600 178.430 ;
        RECT 117.160 177.830 117.420 178.090 ;
        RECT 122.220 177.830 122.480 178.090 ;
        RECT 133.260 177.830 133.520 178.090 ;
        RECT 136.020 178.170 136.280 178.430 ;
        RECT 137.400 178.170 137.660 178.430 ;
        RECT 134.640 177.830 134.900 178.090 ;
        RECT 136.940 177.830 137.200 178.090 ;
        RECT 110.720 177.150 110.980 177.410 ;
        RECT 117.160 177.150 117.420 177.410 ;
        RECT 119.000 177.150 119.260 177.410 ;
        RECT 123.140 177.150 123.400 177.410 ;
        RECT 127.280 177.150 127.540 177.410 ;
        RECT 133.260 177.150 133.520 177.410 ;
        RECT 138.780 177.150 139.040 177.410 ;
        RECT 140.160 177.150 140.420 177.410 ;
        RECT 40.170 176.640 40.430 176.900 ;
        RECT 40.490 176.640 40.750 176.900 ;
        RECT 40.810 176.640 41.070 176.900 ;
        RECT 41.130 176.640 41.390 176.900 ;
        RECT 41.450 176.640 41.710 176.900 ;
        RECT 41.770 176.640 42.030 176.900 ;
        RECT 70.170 176.640 70.430 176.900 ;
        RECT 70.490 176.640 70.750 176.900 ;
        RECT 70.810 176.640 71.070 176.900 ;
        RECT 71.130 176.640 71.390 176.900 ;
        RECT 71.450 176.640 71.710 176.900 ;
        RECT 71.770 176.640 72.030 176.900 ;
        RECT 100.170 176.640 100.430 176.900 ;
        RECT 100.490 176.640 100.750 176.900 ;
        RECT 100.810 176.640 101.070 176.900 ;
        RECT 101.130 176.640 101.390 176.900 ;
        RECT 101.450 176.640 101.710 176.900 ;
        RECT 101.770 176.640 102.030 176.900 ;
        RECT 130.170 176.640 130.430 176.900 ;
        RECT 130.490 176.640 130.750 176.900 ;
        RECT 130.810 176.640 131.070 176.900 ;
        RECT 131.130 176.640 131.390 176.900 ;
        RECT 131.450 176.640 131.710 176.900 ;
        RECT 131.770 176.640 132.030 176.900 ;
        RECT 38.960 176.130 39.220 176.390 ;
        RECT 47.700 176.130 47.960 176.390 ;
        RECT 50.000 176.130 50.260 176.390 ;
        RECT 46.320 175.450 46.580 175.710 ;
        RECT 48.160 175.450 48.420 175.710 ;
        RECT 60.580 176.130 60.840 176.390 ;
        RECT 69.320 176.130 69.580 176.390 ;
        RECT 69.780 176.130 70.040 176.390 ;
        RECT 53.680 175.790 53.940 176.050 ;
        RECT 54.140 175.790 54.400 176.050 ;
        RECT 87.720 175.790 87.980 176.050 ;
        RECT 92.780 175.790 93.040 176.050 ;
        RECT 97.380 176.130 97.640 176.390 ;
        RECT 101.060 176.130 101.320 176.390 ;
        RECT 101.980 176.130 102.240 176.390 ;
        RECT 61.500 175.450 61.760 175.710 ;
        RECT 40.340 175.110 40.600 175.370 ;
        RECT 42.640 175.110 42.900 175.370 ;
        RECT 45.400 175.110 45.660 175.370 ;
        RECT 49.540 174.770 49.800 175.030 ;
        RECT 50.920 175.110 51.180 175.370 ;
        RECT 51.840 175.110 52.100 175.370 ;
        RECT 52.300 175.110 52.560 175.370 ;
        RECT 53.680 175.110 53.940 175.370 ;
        RECT 54.600 175.110 54.860 175.370 ;
        RECT 58.280 175.110 58.540 175.370 ;
        RECT 59.200 175.110 59.460 175.370 ;
        RECT 72.540 175.450 72.800 175.710 ;
        RECT 95.540 175.450 95.800 175.710 ;
        RECT 96.000 175.450 96.260 175.710 ;
        RECT 99.220 175.450 99.480 175.710 ;
        RECT 99.680 175.450 99.940 175.710 ;
        RECT 83.120 175.110 83.380 175.370 ;
        RECT 59.660 174.770 59.920 175.030 ;
        RECT 61.040 174.770 61.300 175.030 ;
        RECT 86.800 175.110 87.060 175.370 ;
        RECT 54.600 174.430 54.860 174.690 ;
        RECT 60.580 174.430 60.840 174.690 ;
        RECT 65.640 174.430 65.900 174.690 ;
        RECT 84.500 174.770 84.760 175.030 ;
        RECT 88.180 175.110 88.440 175.370 ;
        RECT 88.640 175.110 88.900 175.370 ;
        RECT 89.100 175.110 89.360 175.370 ;
        RECT 89.560 175.110 89.820 175.370 ;
        RECT 91.860 175.110 92.120 175.370 ;
        RECT 92.320 175.110 92.580 175.370 ;
        RECT 92.780 175.110 93.040 175.370 ;
        RECT 97.380 175.110 97.640 175.370 ;
        RECT 98.300 175.110 98.560 175.370 ;
        RECT 90.020 174.430 90.280 174.690 ;
        RECT 90.940 174.430 91.200 174.690 ;
        RECT 91.400 174.430 91.660 174.690 ;
        RECT 94.160 174.430 94.420 174.690 ;
        RECT 96.000 174.770 96.260 175.030 ;
        RECT 101.060 175.110 101.320 175.370 ;
        RECT 107.040 175.790 107.300 176.050 ;
        RECT 107.500 175.790 107.760 176.050 ;
        RECT 108.880 175.790 109.140 176.050 ;
        RECT 111.640 176.130 111.900 176.390 ;
        RECT 102.440 175.450 102.700 175.710 ;
        RECT 102.900 175.450 103.160 175.710 ;
        RECT 105.660 175.450 105.920 175.710 ;
        RECT 100.600 174.770 100.860 175.030 ;
        RECT 101.520 174.770 101.780 175.030 ;
        RECT 104.280 175.110 104.540 175.370 ;
        RECT 110.720 175.450 110.980 175.710 ;
        RECT 112.560 175.450 112.820 175.710 ;
        RECT 120.380 175.790 120.640 176.050 ;
        RECT 117.160 175.450 117.420 175.710 ;
        RECT 126.820 176.130 127.080 176.390 ;
        RECT 127.280 176.130 127.540 176.390 ;
        RECT 130.040 176.130 130.300 176.390 ;
        RECT 135.100 176.130 135.360 176.390 ;
        RECT 137.400 176.130 137.660 176.390 ;
        RECT 138.780 176.130 139.040 176.390 ;
        RECT 136.020 175.790 136.280 176.050 ;
        RECT 105.660 174.770 105.920 175.030 ;
        RECT 117.620 175.110 117.880 175.370 ;
        RECT 101.980 174.430 102.240 174.690 ;
        RECT 102.440 174.430 102.700 174.690 ;
        RECT 106.580 174.430 106.840 174.690 ;
        RECT 121.760 175.110 122.020 175.370 ;
        RECT 124.060 175.110 124.320 175.370 ;
        RECT 124.980 175.110 125.240 175.370 ;
        RECT 126.820 175.110 127.080 175.370 ;
        RECT 127.740 175.110 128.000 175.370 ;
        RECT 132.340 175.110 132.600 175.370 ;
        RECT 140.160 175.110 140.420 175.370 ;
        RECT 118.540 174.430 118.800 174.690 ;
        RECT 119.460 174.430 119.720 174.690 ;
        RECT 123.140 174.430 123.400 174.690 ;
        RECT 55.170 173.920 55.430 174.180 ;
        RECT 55.490 173.920 55.750 174.180 ;
        RECT 55.810 173.920 56.070 174.180 ;
        RECT 56.130 173.920 56.390 174.180 ;
        RECT 56.450 173.920 56.710 174.180 ;
        RECT 56.770 173.920 57.030 174.180 ;
        RECT 85.170 173.920 85.430 174.180 ;
        RECT 85.490 173.920 85.750 174.180 ;
        RECT 85.810 173.920 86.070 174.180 ;
        RECT 86.130 173.920 86.390 174.180 ;
        RECT 86.450 173.920 86.710 174.180 ;
        RECT 86.770 173.920 87.030 174.180 ;
        RECT 115.170 173.920 115.430 174.180 ;
        RECT 115.490 173.920 115.750 174.180 ;
        RECT 115.810 173.920 116.070 174.180 ;
        RECT 116.130 173.920 116.390 174.180 ;
        RECT 116.450 173.920 116.710 174.180 ;
        RECT 116.770 173.920 117.030 174.180 ;
        RECT 145.170 173.920 145.430 174.180 ;
        RECT 145.490 173.920 145.750 174.180 ;
        RECT 145.810 173.920 146.070 174.180 ;
        RECT 146.130 173.920 146.390 174.180 ;
        RECT 146.450 173.920 146.710 174.180 ;
        RECT 146.770 173.920 147.030 174.180 ;
        RECT 40.340 173.410 40.600 173.670 ;
        RECT 44.020 173.410 44.280 173.670 ;
        RECT 45.400 173.410 45.660 173.670 ;
        RECT 46.320 173.070 46.580 173.330 ;
        RECT 48.160 173.070 48.420 173.330 ;
        RECT 50.920 173.410 51.180 173.670 ;
        RECT 52.300 173.410 52.560 173.670 ;
        RECT 53.680 173.410 53.940 173.670 ;
        RECT 59.660 173.410 59.920 173.670 ;
        RECT 63.800 173.410 64.060 173.670 ;
        RECT 42.180 172.390 42.440 172.650 ;
        RECT 47.700 172.730 47.960 172.990 ;
        RECT 60.580 173.070 60.840 173.330 ;
        RECT 65.180 173.410 65.440 173.670 ;
        RECT 83.120 173.410 83.380 173.670 ;
        RECT 84.500 173.410 84.760 173.670 ;
        RECT 89.100 173.410 89.360 173.670 ;
        RECT 90.020 173.410 90.280 173.670 ;
        RECT 91.860 173.410 92.120 173.670 ;
        RECT 93.700 173.410 93.960 173.670 ;
        RECT 95.080 173.410 95.340 173.670 ;
        RECT 65.640 173.070 65.900 173.330 ;
        RECT 49.540 172.390 49.800 172.650 ;
        RECT 51.380 172.730 51.640 172.990 ;
        RECT 51.840 172.730 52.100 172.990 ;
        RECT 53.220 172.730 53.480 172.990 ;
        RECT 57.360 172.730 57.620 172.990 ;
        RECT 62.880 172.730 63.140 172.990 ;
        RECT 67.020 172.730 67.280 172.990 ;
        RECT 68.400 172.730 68.660 172.990 ;
        RECT 74.840 173.070 75.100 173.330 ;
        RECT 76.220 173.070 76.480 173.330 ;
        RECT 78.520 173.070 78.780 173.330 ;
        RECT 86.800 173.070 87.060 173.330 ;
        RECT 99.220 173.410 99.480 173.670 ;
        RECT 100.600 173.410 100.860 173.670 ;
        RECT 54.600 172.390 54.860 172.650 ;
        RECT 61.500 172.390 61.760 172.650 ;
        RECT 81.280 172.730 81.540 172.990 ;
        RECT 80.360 172.390 80.620 172.650 ;
        RECT 43.100 171.710 43.360 171.970 ;
        RECT 47.700 171.710 47.960 171.970 ;
        RECT 52.300 171.710 52.560 171.970 ;
        RECT 54.140 171.710 54.400 171.970 ;
        RECT 58.740 171.710 59.000 171.970 ;
        RECT 64.720 171.710 64.980 171.970 ;
        RECT 73.460 171.710 73.720 171.970 ;
        RECT 88.640 172.730 88.900 172.990 ;
        RECT 90.020 172.730 90.280 172.990 ;
        RECT 96.460 173.070 96.720 173.330 ;
        RECT 91.400 172.730 91.660 172.990 ;
        RECT 92.780 172.730 93.040 172.990 ;
        RECT 87.720 172.050 87.980 172.310 ;
        RECT 80.360 171.710 80.620 171.970 ;
        RECT 86.340 171.710 86.600 171.970 ;
        RECT 87.260 171.710 87.520 171.970 ;
        RECT 89.560 171.710 89.820 171.970 ;
        RECT 93.700 172.390 93.960 172.650 ;
        RECT 92.780 171.710 93.040 171.970 ;
        RECT 96.920 172.390 97.180 172.650 ;
        RECT 101.980 172.730 102.240 172.990 ;
        RECT 103.360 172.730 103.620 172.990 ;
        RECT 103.820 172.730 104.080 172.990 ;
        RECT 107.040 172.730 107.300 172.990 ;
        RECT 111.640 173.070 111.900 173.330 ;
        RECT 113.940 173.070 114.200 173.330 ;
        RECT 117.160 173.410 117.420 173.670 ;
        RECT 118.540 173.410 118.800 173.670 ;
        RECT 120.380 173.410 120.640 173.670 ;
        RECT 139.700 173.410 139.960 173.670 ;
        RECT 123.140 173.070 123.400 173.330 ;
        RECT 98.760 172.050 99.020 172.310 ;
        RECT 100.600 172.050 100.860 172.310 ;
        RECT 102.900 172.050 103.160 172.310 ;
        RECT 119.460 172.390 119.720 172.650 ;
        RECT 122.680 172.730 122.940 172.990 ;
        RECT 135.100 172.730 135.360 172.990 ;
        RECT 126.820 172.390 127.080 172.650 ;
        RECT 142.460 172.730 142.720 172.990 ;
        RECT 142.920 172.730 143.180 172.990 ;
        RECT 105.660 171.710 105.920 171.970 ;
        RECT 106.580 171.710 106.840 171.970 ;
        RECT 107.960 171.710 108.220 171.970 ;
        RECT 108.880 171.710 109.140 171.970 ;
        RECT 136.940 171.710 137.200 171.970 ;
        RECT 141.540 171.710 141.800 171.970 ;
        RECT 142.000 171.710 142.260 171.970 ;
        RECT 40.170 171.200 40.430 171.460 ;
        RECT 40.490 171.200 40.750 171.460 ;
        RECT 40.810 171.200 41.070 171.460 ;
        RECT 41.130 171.200 41.390 171.460 ;
        RECT 41.450 171.200 41.710 171.460 ;
        RECT 41.770 171.200 42.030 171.460 ;
        RECT 70.170 171.200 70.430 171.460 ;
        RECT 70.490 171.200 70.750 171.460 ;
        RECT 70.810 171.200 71.070 171.460 ;
        RECT 71.130 171.200 71.390 171.460 ;
        RECT 71.450 171.200 71.710 171.460 ;
        RECT 71.770 171.200 72.030 171.460 ;
        RECT 100.170 171.200 100.430 171.460 ;
        RECT 100.490 171.200 100.750 171.460 ;
        RECT 100.810 171.200 101.070 171.460 ;
        RECT 101.130 171.200 101.390 171.460 ;
        RECT 101.450 171.200 101.710 171.460 ;
        RECT 101.770 171.200 102.030 171.460 ;
        RECT 130.170 171.200 130.430 171.460 ;
        RECT 130.490 171.200 130.750 171.460 ;
        RECT 130.810 171.200 131.070 171.460 ;
        RECT 131.130 171.200 131.390 171.460 ;
        RECT 131.450 171.200 131.710 171.460 ;
        RECT 131.770 171.200 132.030 171.460 ;
        RECT 43.100 170.690 43.360 170.950 ;
        RECT 41.720 170.350 41.980 170.610 ;
        RECT 42.180 170.010 42.440 170.270 ;
        RECT 43.100 169.670 43.360 169.930 ;
        RECT 45.400 170.690 45.660 170.950 ;
        RECT 46.320 170.690 46.580 170.950 ;
        RECT 51.380 170.690 51.640 170.950 ;
        RECT 61.040 170.690 61.300 170.950 ;
        RECT 63.340 170.690 63.600 170.950 ;
        RECT 76.220 170.690 76.480 170.950 ;
        RECT 73.460 170.350 73.720 170.610 ;
        RECT 78.520 170.350 78.780 170.610 ;
        RECT 85.880 170.690 86.140 170.950 ;
        RECT 86.340 170.690 86.600 170.950 ;
        RECT 93.700 170.690 93.960 170.950 ;
        RECT 97.380 170.690 97.640 170.950 ;
        RECT 121.300 170.690 121.560 170.950 ;
        RECT 136.940 170.690 137.200 170.950 ;
        RECT 142.460 170.690 142.720 170.950 ;
        RECT 44.480 169.670 44.740 169.930 ;
        RECT 52.300 170.010 52.560 170.270 ;
        RECT 61.040 169.670 61.300 169.930 ;
        RECT 61.960 170.010 62.220 170.270 ;
        RECT 68.860 170.010 69.120 170.270 ;
        RECT 87.720 170.010 87.980 170.270 ;
        RECT 90.940 170.350 91.200 170.610 ;
        RECT 90.480 170.010 90.740 170.270 ;
        RECT 92.780 170.010 93.040 170.270 ;
        RECT 101.980 170.350 102.240 170.610 ;
        RECT 104.280 170.350 104.540 170.610 ;
        RECT 108.420 170.350 108.680 170.610 ;
        RECT 109.800 170.010 110.060 170.270 ;
        RECT 58.280 169.330 58.540 169.590 ;
        RECT 60.580 169.330 60.840 169.590 ;
        RECT 64.260 169.670 64.520 169.930 ;
        RECT 66.100 169.670 66.360 169.930 ;
        RECT 86.340 169.670 86.600 169.930 ;
        RECT 90.940 169.670 91.200 169.930 ;
        RECT 91.400 169.670 91.660 169.930 ;
        RECT 67.020 169.330 67.280 169.590 ;
        RECT 43.100 168.990 43.360 169.250 ;
        RECT 45.400 168.990 45.660 169.250 ;
        RECT 47.240 168.990 47.500 169.250 ;
        RECT 61.960 168.990 62.220 169.250 ;
        RECT 90.020 169.330 90.280 169.590 ;
        RECT 69.320 168.990 69.580 169.250 ;
        RECT 69.780 168.990 70.040 169.250 ;
        RECT 74.840 168.990 75.100 169.250 ;
        RECT 76.220 168.990 76.480 169.250 ;
        RECT 84.500 168.990 84.760 169.250 ;
        RECT 94.160 169.330 94.420 169.590 ;
        RECT 97.380 169.330 97.640 169.590 ;
        RECT 102.440 169.670 102.700 169.930 ;
        RECT 102.900 169.670 103.160 169.930 ;
        RECT 108.420 169.670 108.680 169.930 ;
        RECT 108.880 169.670 109.140 169.930 ;
        RECT 93.240 168.990 93.500 169.250 ;
        RECT 94.620 168.990 94.880 169.250 ;
        RECT 96.000 168.990 96.260 169.250 ;
        RECT 98.300 168.990 98.560 169.250 ;
        RECT 117.620 169.670 117.880 169.930 ;
        RECT 122.680 169.670 122.940 169.930 ;
        RECT 123.140 169.670 123.400 169.930 ;
        RECT 127.280 170.010 127.540 170.270 ;
        RECT 124.980 169.670 125.240 169.930 ;
        RECT 138.320 170.010 138.580 170.270 ;
        RECT 113.020 169.330 113.280 169.590 ;
        RECT 113.940 168.990 114.200 169.250 ;
        RECT 122.220 169.330 122.480 169.590 ;
        RECT 132.340 169.670 132.600 169.930 ;
        RECT 139.700 170.010 139.960 170.270 ;
        RECT 124.060 168.990 124.320 169.250 ;
        RECT 137.860 169.330 138.120 169.590 ;
        RECT 138.320 169.330 138.580 169.590 ;
        RECT 128.660 168.990 128.920 169.250 ;
        RECT 141.080 168.990 141.340 169.250 ;
        RECT 55.170 168.480 55.430 168.740 ;
        RECT 55.490 168.480 55.750 168.740 ;
        RECT 55.810 168.480 56.070 168.740 ;
        RECT 56.130 168.480 56.390 168.740 ;
        RECT 56.450 168.480 56.710 168.740 ;
        RECT 56.770 168.480 57.030 168.740 ;
        RECT 85.170 168.480 85.430 168.740 ;
        RECT 85.490 168.480 85.750 168.740 ;
        RECT 85.810 168.480 86.070 168.740 ;
        RECT 86.130 168.480 86.390 168.740 ;
        RECT 86.450 168.480 86.710 168.740 ;
        RECT 86.770 168.480 87.030 168.740 ;
        RECT 115.170 168.480 115.430 168.740 ;
        RECT 115.490 168.480 115.750 168.740 ;
        RECT 115.810 168.480 116.070 168.740 ;
        RECT 116.130 168.480 116.390 168.740 ;
        RECT 116.450 168.480 116.710 168.740 ;
        RECT 116.770 168.480 117.030 168.740 ;
        RECT 145.170 168.480 145.430 168.740 ;
        RECT 145.490 168.480 145.750 168.740 ;
        RECT 145.810 168.480 146.070 168.740 ;
        RECT 146.130 168.480 146.390 168.740 ;
        RECT 146.450 168.480 146.710 168.740 ;
        RECT 146.770 168.480 147.030 168.740 ;
        RECT 43.100 167.970 43.360 168.230 ;
        RECT 52.300 167.970 52.560 168.230 ;
        RECT 60.580 167.970 60.840 168.230 ;
        RECT 67.020 167.970 67.280 168.230 ;
        RECT 68.400 167.970 68.660 168.230 ;
        RECT 69.320 167.970 69.580 168.230 ;
        RECT 74.380 167.970 74.640 168.230 ;
        RECT 75.300 167.970 75.560 168.230 ;
        RECT 76.220 167.970 76.480 168.230 ;
        RECT 43.560 167.630 43.820 167.890 ;
        RECT 37.580 167.290 37.840 167.550 ;
        RECT 45.400 167.290 45.660 167.550 ;
        RECT 58.280 167.290 58.540 167.550 ;
        RECT 66.560 167.630 66.820 167.890 ;
        RECT 81.740 167.970 82.000 168.230 ;
        RECT 91.400 167.970 91.660 168.230 ;
        RECT 93.700 167.970 93.960 168.230 ;
        RECT 94.620 167.970 94.880 168.230 ;
        RECT 96.000 167.970 96.260 168.230 ;
        RECT 97.380 167.970 97.640 168.230 ;
        RECT 62.880 167.290 63.140 167.550 ;
        RECT 65.640 167.290 65.900 167.550 ;
        RECT 68.860 167.290 69.120 167.550 ;
        RECT 41.720 166.950 41.980 167.210 ;
        RECT 50.000 166.950 50.260 167.210 ;
        RECT 44.480 166.270 44.740 166.530 ;
        RECT 51.840 166.270 52.100 166.530 ;
        RECT 58.740 166.950 59.000 167.210 ;
        RECT 59.660 166.950 59.920 167.210 ;
        RECT 61.960 166.950 62.220 167.210 ;
        RECT 61.500 166.610 61.760 166.870 ;
        RECT 73.000 166.950 73.260 167.210 ;
        RECT 75.300 166.950 75.560 167.210 ;
        RECT 78.520 167.290 78.780 167.550 ;
        RECT 79.900 167.290 80.160 167.550 ;
        RECT 81.280 167.290 81.540 167.550 ;
        RECT 84.040 167.290 84.300 167.550 ;
        RECT 87.720 167.290 87.980 167.550 ;
        RECT 88.180 167.290 88.440 167.550 ;
        RECT 90.940 167.630 91.200 167.890 ;
        RECT 93.240 167.630 93.500 167.890 ;
        RECT 79.440 166.950 79.700 167.210 ;
        RECT 89.100 166.610 89.360 166.870 ;
        RECT 69.320 166.270 69.580 166.530 ;
        RECT 73.000 166.270 73.260 166.530 ;
        RECT 78.520 166.270 78.780 166.530 ;
        RECT 87.260 166.270 87.520 166.530 ;
        RECT 92.320 167.290 92.580 167.550 ;
        RECT 107.960 167.970 108.220 168.230 ;
        RECT 108.420 167.970 108.680 168.230 ;
        RECT 113.020 167.970 113.280 168.230 ;
        RECT 118.540 167.970 118.800 168.230 ;
        RECT 121.300 167.970 121.560 168.230 ;
        RECT 123.140 167.970 123.400 168.230 ;
        RECT 96.920 167.290 97.180 167.550 ;
        RECT 95.080 166.950 95.340 167.210 ;
        RECT 103.360 167.630 103.620 167.890 ;
        RECT 99.220 167.290 99.480 167.550 ;
        RECT 99.680 167.290 99.940 167.550 ;
        RECT 112.100 167.630 112.360 167.890 ;
        RECT 108.420 167.290 108.680 167.550 ;
        RECT 111.180 167.290 111.440 167.550 ;
        RECT 117.620 167.290 117.880 167.550 ;
        RECT 118.540 167.290 118.800 167.550 ;
        RECT 119.460 167.630 119.720 167.890 ;
        RECT 102.900 166.950 103.160 167.210 ;
        RECT 106.580 166.950 106.840 167.210 ;
        RECT 107.960 166.950 108.220 167.210 ;
        RECT 96.000 166.270 96.260 166.530 ;
        RECT 99.220 166.270 99.480 166.530 ;
        RECT 105.660 166.270 105.920 166.530 ;
        RECT 109.340 166.270 109.600 166.530 ;
        RECT 119.460 166.610 119.720 166.870 ;
        RECT 117.620 166.270 117.880 166.530 ;
        RECT 122.680 166.950 122.940 167.210 ;
        RECT 124.060 167.290 124.320 167.550 ;
        RECT 143.840 167.970 144.100 168.230 ;
        RECT 127.280 167.290 127.540 167.550 ;
        RECT 127.740 167.290 128.000 167.550 ;
        RECT 129.120 167.290 129.380 167.550 ;
        RECT 132.340 167.290 132.600 167.550 ;
        RECT 142.460 167.290 142.720 167.550 ;
        RECT 142.920 167.290 143.180 167.550 ;
        RECT 124.520 166.950 124.780 167.210 ;
        RECT 140.160 166.610 140.420 166.870 ;
        RECT 142.000 166.610 142.260 166.870 ;
        RECT 128.660 166.270 128.920 166.530 ;
        RECT 143.840 166.270 144.100 166.530 ;
        RECT 40.170 165.760 40.430 166.020 ;
        RECT 40.490 165.760 40.750 166.020 ;
        RECT 40.810 165.760 41.070 166.020 ;
        RECT 41.130 165.760 41.390 166.020 ;
        RECT 41.450 165.760 41.710 166.020 ;
        RECT 41.770 165.760 42.030 166.020 ;
        RECT 70.170 165.760 70.430 166.020 ;
        RECT 70.490 165.760 70.750 166.020 ;
        RECT 70.810 165.760 71.070 166.020 ;
        RECT 71.130 165.760 71.390 166.020 ;
        RECT 71.450 165.760 71.710 166.020 ;
        RECT 71.770 165.760 72.030 166.020 ;
        RECT 100.170 165.760 100.430 166.020 ;
        RECT 100.490 165.760 100.750 166.020 ;
        RECT 100.810 165.760 101.070 166.020 ;
        RECT 101.130 165.760 101.390 166.020 ;
        RECT 101.450 165.760 101.710 166.020 ;
        RECT 101.770 165.760 102.030 166.020 ;
        RECT 130.170 165.760 130.430 166.020 ;
        RECT 130.490 165.760 130.750 166.020 ;
        RECT 130.810 165.760 131.070 166.020 ;
        RECT 131.130 165.760 131.390 166.020 ;
        RECT 131.450 165.760 131.710 166.020 ;
        RECT 131.770 165.760 132.030 166.020 ;
        RECT 42.180 165.250 42.440 165.510 ;
        RECT 62.880 165.250 63.140 165.510 ;
        RECT 67.940 165.250 68.200 165.510 ;
        RECT 73.000 165.250 73.260 165.510 ;
        RECT 74.840 165.250 75.100 165.510 ;
        RECT 76.220 165.250 76.480 165.510 ;
        RECT 79.900 165.250 80.160 165.510 ;
        RECT 47.240 164.910 47.500 165.170 ;
        RECT 88.640 165.250 88.900 165.510 ;
        RECT 89.100 165.250 89.360 165.510 ;
        RECT 91.860 165.250 92.120 165.510 ;
        RECT 92.320 165.250 92.580 165.510 ;
        RECT 101.980 165.250 102.240 165.510 ;
        RECT 107.500 165.250 107.760 165.510 ;
        RECT 111.180 165.250 111.440 165.510 ;
        RECT 112.100 165.250 112.360 165.510 ;
        RECT 114.400 165.250 114.660 165.510 ;
        RECT 121.300 165.250 121.560 165.510 ;
        RECT 129.120 165.250 129.380 165.510 ;
        RECT 137.860 165.250 138.120 165.510 ;
        RECT 141.080 165.250 141.340 165.510 ;
        RECT 141.540 165.250 141.800 165.510 ;
        RECT 44.940 164.570 45.200 164.830 ;
        RECT 44.480 164.230 44.740 164.490 ;
        RECT 58.740 164.570 59.000 164.830 ;
        RECT 61.500 164.570 61.760 164.830 ;
        RECT 60.580 164.230 60.840 164.490 ;
        RECT 66.560 164.570 66.820 164.830 ;
        RECT 71.620 164.570 71.880 164.830 ;
        RECT 43.100 163.550 43.360 163.810 ;
        RECT 44.940 163.550 45.200 163.810 ;
        RECT 50.920 163.550 51.180 163.810 ;
        RECT 62.420 163.550 62.680 163.810 ;
        RECT 63.800 163.550 64.060 163.810 ;
        RECT 67.480 163.550 67.740 163.810 ;
        RECT 73.000 163.550 73.260 163.810 ;
        RECT 76.680 164.230 76.940 164.490 ;
        RECT 79.440 164.230 79.700 164.490 ;
        RECT 80.360 164.230 80.620 164.490 ;
        RECT 90.020 164.910 90.280 165.170 ;
        RECT 92.780 164.910 93.040 165.170 ;
        RECT 89.100 164.230 89.360 164.490 ;
        RECT 90.480 164.230 90.740 164.490 ;
        RECT 91.860 164.570 92.120 164.830 ;
        RECT 83.120 163.890 83.380 164.150 ;
        RECT 91.400 163.890 91.660 164.150 ;
        RECT 93.240 164.230 93.500 164.490 ;
        RECT 94.160 164.230 94.420 164.490 ;
        RECT 95.540 164.230 95.800 164.490 ;
        RECT 96.000 164.230 96.260 164.490 ;
        RECT 96.460 164.230 96.720 164.490 ;
        RECT 97.380 164.230 97.640 164.490 ;
        RECT 101.520 164.230 101.780 164.490 ;
        RECT 102.440 164.230 102.700 164.490 ;
        RECT 104.280 164.230 104.540 164.490 ;
        RECT 76.220 163.550 76.480 163.810 ;
        RECT 78.520 163.550 78.780 163.810 ;
        RECT 90.940 163.550 91.200 163.810 ;
        RECT 91.860 163.550 92.120 163.810 ;
        RECT 94.160 163.550 94.420 163.810 ;
        RECT 106.120 163.890 106.380 164.150 ;
        RECT 99.220 163.550 99.480 163.810 ;
        RECT 110.260 164.570 110.520 164.830 ;
        RECT 110.720 164.570 110.980 164.830 ;
        RECT 113.020 164.570 113.280 164.830 ;
        RECT 113.480 164.570 113.740 164.830 ;
        RECT 114.400 164.570 114.660 164.830 ;
        RECT 119.460 164.570 119.720 164.830 ;
        RECT 109.340 164.230 109.600 164.490 ;
        RECT 107.500 163.890 107.760 164.150 ;
        RECT 111.640 164.230 111.900 164.490 ;
        RECT 118.540 164.230 118.800 164.490 ;
        RECT 127.740 164.910 128.000 165.170 ;
        RECT 135.100 164.910 135.360 165.170 ;
        RECT 143.840 164.570 144.100 164.830 ;
        RECT 124.520 164.230 124.780 164.490 ;
        RECT 125.440 164.230 125.700 164.490 ;
        RECT 135.100 164.230 135.360 164.490 ;
        RECT 140.160 164.230 140.420 164.490 ;
        RECT 140.620 164.230 140.880 164.490 ;
        RECT 142.460 164.230 142.720 164.490 ;
        RECT 142.920 164.230 143.180 164.490 ;
        RECT 107.960 163.550 108.220 163.810 ;
        RECT 109.340 163.550 109.600 163.810 ;
        RECT 111.640 163.550 111.900 163.810 ;
        RECT 117.620 163.550 117.880 163.810 ;
        RECT 122.680 163.550 122.940 163.810 ;
        RECT 133.260 163.890 133.520 164.150 ;
        RECT 138.780 163.890 139.040 164.150 ;
        RECT 141.080 163.550 141.340 163.810 ;
        RECT 55.170 163.040 55.430 163.300 ;
        RECT 55.490 163.040 55.750 163.300 ;
        RECT 55.810 163.040 56.070 163.300 ;
        RECT 56.130 163.040 56.390 163.300 ;
        RECT 56.450 163.040 56.710 163.300 ;
        RECT 56.770 163.040 57.030 163.300 ;
        RECT 85.170 163.040 85.430 163.300 ;
        RECT 85.490 163.040 85.750 163.300 ;
        RECT 85.810 163.040 86.070 163.300 ;
        RECT 86.130 163.040 86.390 163.300 ;
        RECT 86.450 163.040 86.710 163.300 ;
        RECT 86.770 163.040 87.030 163.300 ;
        RECT 115.170 163.040 115.430 163.300 ;
        RECT 115.490 163.040 115.750 163.300 ;
        RECT 115.810 163.040 116.070 163.300 ;
        RECT 116.130 163.040 116.390 163.300 ;
        RECT 116.450 163.040 116.710 163.300 ;
        RECT 116.770 163.040 117.030 163.300 ;
        RECT 145.170 163.040 145.430 163.300 ;
        RECT 145.490 163.040 145.750 163.300 ;
        RECT 145.810 163.040 146.070 163.300 ;
        RECT 146.130 163.040 146.390 163.300 ;
        RECT 146.450 163.040 146.710 163.300 ;
        RECT 146.770 163.040 147.030 163.300 ;
        RECT 44.940 162.530 45.200 162.790 ;
        RECT 46.780 162.530 47.040 162.790 ;
        RECT 54.140 162.530 54.400 162.790 ;
        RECT 60.580 162.530 60.840 162.790 ;
        RECT 66.560 162.530 66.820 162.790 ;
        RECT 76.680 162.530 76.940 162.790 ;
        RECT 80.360 162.530 80.620 162.790 ;
        RECT 51.840 162.190 52.100 162.450 ;
        RECT 37.580 161.850 37.840 162.110 ;
        RECT 51.380 161.850 51.640 162.110 ;
        RECT 55.060 161.850 55.320 162.110 ;
        RECT 52.300 161.510 52.560 161.770 ;
        RECT 54.140 161.510 54.400 161.770 ;
        RECT 62.880 161.510 63.140 161.770 ;
        RECT 63.800 162.190 64.060 162.450 ;
        RECT 95.080 162.530 95.340 162.790 ;
        RECT 97.380 162.530 97.640 162.790 ;
        RECT 107.040 162.530 107.300 162.790 ;
        RECT 117.620 162.530 117.880 162.790 ;
        RECT 137.400 162.530 137.660 162.790 ;
        RECT 139.240 162.530 139.500 162.790 ;
        RECT 142.920 162.530 143.180 162.790 ;
        RECT 144.760 162.530 145.020 162.790 ;
        RECT 69.320 161.850 69.580 162.110 ;
        RECT 70.700 161.850 70.960 162.110 ;
        RECT 87.260 161.850 87.520 162.110 ;
        RECT 91.860 161.850 92.120 162.110 ;
        RECT 92.780 161.850 93.040 162.110 ;
        RECT 98.760 161.850 99.020 162.110 ;
        RECT 102.900 162.190 103.160 162.450 ;
        RECT 103.360 162.190 103.620 162.450 ;
        RECT 102.440 161.850 102.700 162.110 ;
        RECT 104.280 161.850 104.540 162.110 ;
        RECT 108.880 161.850 109.140 162.110 ;
        RECT 113.020 162.190 113.280 162.450 ;
        RECT 110.260 161.850 110.520 162.110 ;
        RECT 111.180 161.850 111.440 162.110 ;
        RECT 112.100 161.850 112.360 162.110 ;
        RECT 114.400 162.190 114.660 162.450 ;
        RECT 72.080 161.510 72.340 161.770 ;
        RECT 85.880 161.510 86.140 161.770 ;
        RECT 92.320 161.510 92.580 161.770 ;
        RECT 63.800 161.170 64.060 161.430 ;
        RECT 69.320 161.170 69.580 161.430 ;
        RECT 71.620 161.170 71.880 161.430 ;
        RECT 93.240 161.170 93.500 161.430 ;
        RECT 97.380 161.510 97.640 161.770 ;
        RECT 109.800 161.510 110.060 161.770 ;
        RECT 119.460 161.850 119.720 162.110 ;
        RECT 124.520 162.190 124.780 162.450 ;
        RECT 122.680 161.850 122.940 162.110 ;
        RECT 132.340 162.190 132.600 162.450 ;
        RECT 135.560 162.190 135.820 162.450 ;
        RECT 141.540 162.190 141.800 162.450 ;
        RECT 98.760 161.170 99.020 161.430 ;
        RECT 107.500 161.170 107.760 161.430 ;
        RECT 59.200 160.830 59.460 161.090 ;
        RECT 59.660 160.830 59.920 161.090 ;
        RECT 95.080 160.830 95.340 161.090 ;
        RECT 97.840 160.830 98.100 161.090 ;
        RECT 99.680 160.830 99.940 161.090 ;
        RECT 104.280 160.830 104.540 161.090 ;
        RECT 106.120 160.830 106.380 161.090 ;
        RECT 115.320 161.170 115.580 161.430 ;
        RECT 126.820 161.510 127.080 161.770 ;
        RECT 133.260 161.850 133.520 162.110 ;
        RECT 138.320 161.850 138.580 162.110 ;
        RECT 139.700 161.850 139.960 162.110 ;
        RECT 138.780 161.510 139.040 161.770 ;
        RECT 131.420 161.170 131.680 161.430 ;
        RECT 134.180 161.170 134.440 161.430 ;
        RECT 138.320 161.170 138.580 161.430 ;
        RECT 114.400 160.830 114.660 161.090 ;
        RECT 125.440 160.830 125.700 161.090 ;
        RECT 127.740 160.830 128.000 161.090 ;
        RECT 133.260 160.830 133.520 161.090 ;
        RECT 136.940 160.830 137.200 161.090 ;
        RECT 137.400 160.830 137.660 161.090 ;
        RECT 40.170 160.320 40.430 160.580 ;
        RECT 40.490 160.320 40.750 160.580 ;
        RECT 40.810 160.320 41.070 160.580 ;
        RECT 41.130 160.320 41.390 160.580 ;
        RECT 41.450 160.320 41.710 160.580 ;
        RECT 41.770 160.320 42.030 160.580 ;
        RECT 70.170 160.320 70.430 160.580 ;
        RECT 70.490 160.320 70.750 160.580 ;
        RECT 70.810 160.320 71.070 160.580 ;
        RECT 71.130 160.320 71.390 160.580 ;
        RECT 71.450 160.320 71.710 160.580 ;
        RECT 71.770 160.320 72.030 160.580 ;
        RECT 100.170 160.320 100.430 160.580 ;
        RECT 100.490 160.320 100.750 160.580 ;
        RECT 100.810 160.320 101.070 160.580 ;
        RECT 101.130 160.320 101.390 160.580 ;
        RECT 101.450 160.320 101.710 160.580 ;
        RECT 101.770 160.320 102.030 160.580 ;
        RECT 130.170 160.320 130.430 160.580 ;
        RECT 130.490 160.320 130.750 160.580 ;
        RECT 130.810 160.320 131.070 160.580 ;
        RECT 131.130 160.320 131.390 160.580 ;
        RECT 131.450 160.320 131.710 160.580 ;
        RECT 131.770 160.320 132.030 160.580 ;
        RECT 47.240 159.810 47.500 160.070 ;
        RECT 52.300 159.810 52.560 160.070 ;
        RECT 68.400 159.810 68.660 160.070 ;
        RECT 91.400 159.810 91.660 160.070 ;
        RECT 43.100 158.790 43.360 159.050 ;
        RECT 47.240 159.130 47.500 159.390 ;
        RECT 55.060 159.130 55.320 159.390 ;
        RECT 62.880 159.470 63.140 159.730 ;
        RECT 100.600 159.470 100.860 159.730 ;
        RECT 44.480 158.790 44.740 159.050 ;
        RECT 44.940 158.790 45.200 159.050 ;
        RECT 51.380 158.790 51.640 159.050 ;
        RECT 54.140 158.790 54.400 159.050 ;
        RECT 73.000 159.130 73.260 159.390 ;
        RECT 42.640 158.110 42.900 158.370 ;
        RECT 59.200 158.790 59.460 159.050 ;
        RECT 75.760 158.790 76.020 159.050 ;
        RECT 77.600 159.130 77.860 159.390 ;
        RECT 78.520 159.130 78.780 159.390 ;
        RECT 79.900 159.130 80.160 159.390 ;
        RECT 81.280 159.130 81.540 159.390 ;
        RECT 82.660 159.130 82.920 159.390 ;
        RECT 96.000 159.130 96.260 159.390 ;
        RECT 95.540 158.790 95.800 159.050 ;
        RECT 78.520 158.450 78.780 158.710 ;
        RECT 87.720 158.450 87.980 158.710 ;
        RECT 60.120 158.110 60.380 158.370 ;
        RECT 73.460 158.110 73.720 158.370 ;
        RECT 75.300 158.110 75.560 158.370 ;
        RECT 90.480 158.110 90.740 158.370 ;
        RECT 97.380 158.790 97.640 159.050 ;
        RECT 97.840 158.790 98.100 159.050 ;
        RECT 100.140 159.130 100.400 159.390 ;
        RECT 106.120 159.810 106.380 160.070 ;
        RECT 108.880 159.810 109.140 160.070 ;
        RECT 110.260 159.470 110.520 159.730 ;
        RECT 121.760 159.810 122.020 160.070 ;
        RECT 124.520 159.810 124.780 160.070 ;
        RECT 125.900 159.810 126.160 160.070 ;
        RECT 134.180 159.810 134.440 160.070 ;
        RECT 140.160 159.810 140.420 160.070 ;
        RECT 143.380 159.810 143.640 160.070 ;
        RECT 143.840 159.810 144.100 160.070 ;
        RECT 99.220 158.790 99.480 159.050 ;
        RECT 99.680 158.790 99.940 159.050 ;
        RECT 105.660 159.130 105.920 159.390 ;
        RECT 104.280 158.790 104.540 159.050 ;
        RECT 108.880 158.450 109.140 158.710 ;
        RECT 105.660 158.110 105.920 158.370 ;
        RECT 107.500 158.110 107.760 158.370 ;
        RECT 110.260 158.790 110.520 159.050 ;
        RECT 113.020 159.130 113.280 159.390 ;
        RECT 113.480 159.130 113.740 159.390 ;
        RECT 115.320 159.130 115.580 159.390 ;
        RECT 126.820 159.130 127.080 159.390 ;
        RECT 111.180 158.790 111.440 159.050 ;
        RECT 114.400 158.790 114.660 159.050 ;
        RECT 133.720 159.470 133.980 159.730 ;
        RECT 133.260 158.790 133.520 159.050 ;
        RECT 135.100 159.130 135.360 159.390 ;
        RECT 136.480 159.470 136.740 159.730 ;
        RECT 126.360 158.450 126.620 158.710 ;
        RECT 131.420 158.450 131.680 158.710 ;
        RECT 135.560 158.790 135.820 159.050 ;
        RECT 136.480 158.790 136.740 159.050 ;
        RECT 136.940 158.790 137.200 159.050 ;
        RECT 137.400 158.790 137.660 159.050 ;
        RECT 141.080 159.470 141.340 159.730 ;
        RECT 114.860 158.110 115.120 158.370 ;
        RECT 117.160 158.110 117.420 158.370 ;
        RECT 139.240 158.110 139.500 158.370 ;
        RECT 140.620 158.790 140.880 159.050 ;
        RECT 141.540 158.790 141.800 159.050 ;
        RECT 144.760 158.790 145.020 159.050 ;
        RECT 143.380 158.450 143.640 158.710 ;
        RECT 144.300 158.450 144.560 158.710 ;
        RECT 147.520 158.790 147.780 159.050 ;
        RECT 55.170 157.600 55.430 157.860 ;
        RECT 55.490 157.600 55.750 157.860 ;
        RECT 55.810 157.600 56.070 157.860 ;
        RECT 56.130 157.600 56.390 157.860 ;
        RECT 56.450 157.600 56.710 157.860 ;
        RECT 56.770 157.600 57.030 157.860 ;
        RECT 85.170 157.600 85.430 157.860 ;
        RECT 85.490 157.600 85.750 157.860 ;
        RECT 85.810 157.600 86.070 157.860 ;
        RECT 86.130 157.600 86.390 157.860 ;
        RECT 86.450 157.600 86.710 157.860 ;
        RECT 86.770 157.600 87.030 157.860 ;
        RECT 115.170 157.600 115.430 157.860 ;
        RECT 115.490 157.600 115.750 157.860 ;
        RECT 115.810 157.600 116.070 157.860 ;
        RECT 116.130 157.600 116.390 157.860 ;
        RECT 116.450 157.600 116.710 157.860 ;
        RECT 116.770 157.600 117.030 157.860 ;
        RECT 145.170 157.600 145.430 157.860 ;
        RECT 145.490 157.600 145.750 157.860 ;
        RECT 145.810 157.600 146.070 157.860 ;
        RECT 146.130 157.600 146.390 157.860 ;
        RECT 146.450 157.600 146.710 157.860 ;
        RECT 146.770 157.600 147.030 157.860 ;
        RECT 44.940 157.090 45.200 157.350 ;
        RECT 54.140 157.090 54.400 157.350 ;
        RECT 67.940 157.090 68.200 157.350 ;
        RECT 50.460 156.750 50.720 157.010 ;
        RECT 52.300 156.750 52.560 157.010 ;
        RECT 37.580 156.410 37.840 156.670 ;
        RECT 39.420 156.410 39.680 156.670 ;
        RECT 58.280 156.410 58.540 156.670 ;
        RECT 63.800 156.410 64.060 156.670 ;
        RECT 60.120 156.070 60.380 156.330 ;
        RECT 58.740 155.730 59.000 155.990 ;
        RECT 66.560 155.730 66.820 155.990 ;
        RECT 75.760 157.090 76.020 157.350 ;
        RECT 73.460 156.750 73.720 157.010 ;
        RECT 77.600 157.090 77.860 157.350 ;
        RECT 80.820 157.090 81.080 157.350 ;
        RECT 83.580 157.090 83.840 157.350 ;
        RECT 86.340 157.090 86.600 157.350 ;
        RECT 69.780 155.730 70.040 155.990 ;
        RECT 79.900 156.410 80.160 156.670 ;
        RECT 73.920 155.730 74.180 155.990 ;
        RECT 74.840 155.730 75.100 155.990 ;
        RECT 76.680 156.070 76.940 156.330 ;
        RECT 78.520 156.070 78.780 156.330 ;
        RECT 85.420 156.750 85.680 157.010 ;
        RECT 92.320 157.090 92.580 157.350 ;
        RECT 90.480 156.750 90.740 157.010 ;
        RECT 97.840 157.090 98.100 157.350 ;
        RECT 86.340 156.410 86.600 156.670 ;
        RECT 87.720 156.410 87.980 156.670 ;
        RECT 100.600 156.750 100.860 157.010 ;
        RECT 95.080 156.410 95.340 156.670 ;
        RECT 99.220 156.410 99.480 156.670 ;
        RECT 104.280 156.750 104.540 157.010 ;
        RECT 101.520 156.410 101.780 156.670 ;
        RECT 102.900 156.410 103.160 156.670 ;
        RECT 78.980 155.730 79.240 155.990 ;
        RECT 68.400 155.390 68.660 155.650 ;
        RECT 73.000 155.390 73.260 155.650 ;
        RECT 82.200 155.730 82.460 155.990 ;
        RECT 85.880 156.070 86.140 156.330 ;
        RECT 88.640 155.730 88.900 155.990 ;
        RECT 102.440 156.070 102.700 156.330 ;
        RECT 107.960 157.090 108.220 157.350 ;
        RECT 110.260 157.090 110.520 157.350 ;
        RECT 105.660 156.410 105.920 156.670 ;
        RECT 109.800 156.410 110.060 156.670 ;
        RECT 109.340 156.070 109.600 156.330 ;
        RECT 112.100 156.410 112.360 156.670 ;
        RECT 113.480 156.410 113.740 156.670 ;
        RECT 117.160 156.750 117.420 157.010 ;
        RECT 115.320 156.410 115.580 156.670 ;
        RECT 119.460 156.410 119.720 156.670 ;
        RECT 126.360 157.090 126.620 157.350 ;
        RECT 132.800 157.090 133.060 157.350 ;
        RECT 137.400 157.090 137.660 157.350 ;
        RECT 139.240 157.090 139.500 157.350 ;
        RECT 147.520 157.090 147.780 157.350 ;
        RECT 123.140 156.410 123.400 156.670 ;
        RECT 137.860 156.750 138.120 157.010 ;
        RECT 80.820 155.390 81.080 155.650 ;
        RECT 86.340 155.390 86.600 155.650 ;
        RECT 92.320 155.390 92.580 155.650 ;
        RECT 97.380 155.390 97.640 155.650 ;
        RECT 98.760 155.390 99.020 155.650 ;
        RECT 105.660 155.390 105.920 155.650 ;
        RECT 110.720 155.730 110.980 155.990 ;
        RECT 117.620 155.730 117.880 155.990 ;
        RECT 124.980 155.730 125.240 155.990 ;
        RECT 111.180 155.390 111.440 155.650 ;
        RECT 112.100 155.390 112.360 155.650 ;
        RECT 114.400 155.390 114.660 155.650 ;
        RECT 119.920 155.390 120.180 155.650 ;
        RECT 125.900 155.390 126.160 155.650 ;
        RECT 131.420 156.410 131.680 156.670 ;
        RECT 132.340 156.410 132.600 156.670 ;
        RECT 126.820 155.730 127.080 155.990 ;
        RECT 133.260 156.070 133.520 156.330 ;
        RECT 137.400 156.410 137.660 156.670 ;
        RECT 139.700 156.410 139.960 156.670 ;
        RECT 128.660 155.390 128.920 155.650 ;
        RECT 132.800 155.390 133.060 155.650 ;
        RECT 133.720 155.390 133.980 155.650 ;
        RECT 40.170 154.880 40.430 155.140 ;
        RECT 40.490 154.880 40.750 155.140 ;
        RECT 40.810 154.880 41.070 155.140 ;
        RECT 41.130 154.880 41.390 155.140 ;
        RECT 41.450 154.880 41.710 155.140 ;
        RECT 41.770 154.880 42.030 155.140 ;
        RECT 70.170 154.880 70.430 155.140 ;
        RECT 70.490 154.880 70.750 155.140 ;
        RECT 70.810 154.880 71.070 155.140 ;
        RECT 71.130 154.880 71.390 155.140 ;
        RECT 71.450 154.880 71.710 155.140 ;
        RECT 71.770 154.880 72.030 155.140 ;
        RECT 100.170 154.880 100.430 155.140 ;
        RECT 100.490 154.880 100.750 155.140 ;
        RECT 100.810 154.880 101.070 155.140 ;
        RECT 101.130 154.880 101.390 155.140 ;
        RECT 101.450 154.880 101.710 155.140 ;
        RECT 101.770 154.880 102.030 155.140 ;
        RECT 130.170 154.880 130.430 155.140 ;
        RECT 130.490 154.880 130.750 155.140 ;
        RECT 130.810 154.880 131.070 155.140 ;
        RECT 131.130 154.880 131.390 155.140 ;
        RECT 131.450 154.880 131.710 155.140 ;
        RECT 131.770 154.880 132.030 155.140 ;
        RECT 39.420 154.370 39.680 154.630 ;
        RECT 52.760 154.370 53.020 154.630 ;
        RECT 48.620 154.030 48.880 154.290 ;
        RECT 41.260 153.350 41.520 153.610 ;
        RECT 44.940 153.350 45.200 153.610 ;
        RECT 45.860 153.350 46.120 153.610 ;
        RECT 48.620 153.350 48.880 153.610 ;
        RECT 50.460 153.350 50.720 153.610 ;
        RECT 51.380 153.350 51.640 153.610 ;
        RECT 66.560 154.370 66.820 154.630 ;
        RECT 68.400 154.370 68.660 154.630 ;
        RECT 78.520 154.030 78.780 154.290 ;
        RECT 98.300 154.370 98.560 154.630 ;
        RECT 103.360 154.370 103.620 154.630 ;
        RECT 107.040 154.370 107.300 154.630 ;
        RECT 112.100 154.370 112.360 154.630 ;
        RECT 114.400 154.370 114.660 154.630 ;
        RECT 114.860 154.370 115.120 154.630 ;
        RECT 119.920 154.370 120.180 154.630 ;
        RECT 127.740 154.370 128.000 154.630 ;
        RECT 137.860 154.370 138.120 154.630 ;
        RECT 142.000 154.370 142.260 154.630 ;
        RECT 67.480 153.690 67.740 153.950 ;
        RECT 76.220 153.690 76.480 153.950 ;
        RECT 78.980 153.690 79.240 153.950 ;
        RECT 73.000 153.350 73.260 153.610 ;
        RECT 80.820 154.030 81.080 154.290 ;
        RECT 82.200 154.030 82.460 154.290 ;
        RECT 85.880 154.030 86.140 154.290 ;
        RECT 101.520 153.690 101.780 153.950 ;
        RECT 101.980 153.690 102.240 153.950 ;
        RECT 105.660 153.690 105.920 153.950 ;
        RECT 106.120 153.690 106.380 153.950 ;
        RECT 107.500 153.690 107.760 153.950 ;
        RECT 42.180 152.670 42.440 152.930 ;
        RECT 72.540 153.010 72.800 153.270 ;
        RECT 81.740 153.350 82.000 153.610 ;
        RECT 82.200 153.350 82.460 153.610 ;
        RECT 83.580 153.350 83.840 153.610 ;
        RECT 84.500 153.350 84.760 153.610 ;
        RECT 97.840 153.350 98.100 153.610 ;
        RECT 59.200 152.670 59.460 152.930 ;
        RECT 76.680 152.670 76.940 152.930 ;
        RECT 78.520 152.670 78.780 152.930 ;
        RECT 86.340 153.010 86.600 153.270 ;
        RECT 102.440 153.350 102.700 153.610 ;
        RECT 103.360 153.350 103.620 153.610 ;
        RECT 82.200 152.670 82.460 152.930 ;
        RECT 88.640 152.670 88.900 152.930 ;
        RECT 92.320 152.670 92.580 152.930 ;
        RECT 95.080 152.670 95.340 152.930 ;
        RECT 98.760 152.670 99.020 152.930 ;
        RECT 107.500 153.010 107.760 153.270 ;
        RECT 110.720 153.350 110.980 153.610 ;
        RECT 111.180 153.350 111.440 153.610 ;
        RECT 113.480 153.690 113.740 153.950 ;
        RECT 114.860 153.690 115.120 153.950 ;
        RECT 116.240 153.350 116.500 153.610 ;
        RECT 125.900 154.030 126.160 154.290 ;
        RECT 130.500 154.030 130.760 154.290 ;
        RECT 124.980 153.690 125.240 153.950 ;
        RECT 117.160 153.010 117.420 153.270 ;
        RECT 101.060 152.670 101.320 152.930 ;
        RECT 103.820 152.670 104.080 152.930 ;
        RECT 111.180 152.670 111.440 152.930 ;
        RECT 113.020 152.670 113.280 152.930 ;
        RECT 114.400 152.670 114.660 152.930 ;
        RECT 118.540 153.350 118.800 153.610 ;
        RECT 127.280 153.350 127.540 153.610 ;
        RECT 126.820 152.670 127.080 152.930 ;
        RECT 128.660 153.350 128.920 153.610 ;
        RECT 130.040 153.350 130.300 153.610 ;
        RECT 133.720 153.010 133.980 153.270 ;
        RECT 134.640 153.010 134.900 153.270 ;
        RECT 139.700 152.670 139.960 152.930 ;
        RECT 55.170 152.160 55.430 152.420 ;
        RECT 55.490 152.160 55.750 152.420 ;
        RECT 55.810 152.160 56.070 152.420 ;
        RECT 56.130 152.160 56.390 152.420 ;
        RECT 56.450 152.160 56.710 152.420 ;
        RECT 56.770 152.160 57.030 152.420 ;
        RECT 85.170 152.160 85.430 152.420 ;
        RECT 85.490 152.160 85.750 152.420 ;
        RECT 85.810 152.160 86.070 152.420 ;
        RECT 86.130 152.160 86.390 152.420 ;
        RECT 86.450 152.160 86.710 152.420 ;
        RECT 86.770 152.160 87.030 152.420 ;
        RECT 115.170 152.160 115.430 152.420 ;
        RECT 115.490 152.160 115.750 152.420 ;
        RECT 115.810 152.160 116.070 152.420 ;
        RECT 116.130 152.160 116.390 152.420 ;
        RECT 116.450 152.160 116.710 152.420 ;
        RECT 116.770 152.160 117.030 152.420 ;
        RECT 145.170 152.160 145.430 152.420 ;
        RECT 145.490 152.160 145.750 152.420 ;
        RECT 145.810 152.160 146.070 152.420 ;
        RECT 146.130 152.160 146.390 152.420 ;
        RECT 146.450 152.160 146.710 152.420 ;
        RECT 146.770 152.160 147.030 152.420 ;
        RECT 45.860 151.650 46.120 151.910 ;
        RECT 42.180 151.310 42.440 151.570 ;
        RECT 39.420 150.970 39.680 151.230 ;
        RECT 53.680 151.650 53.940 151.910 ;
        RECT 78.060 151.650 78.320 151.910 ;
        RECT 51.380 151.310 51.640 151.570 ;
        RECT 59.200 150.970 59.460 151.230 ;
        RECT 52.760 150.630 53.020 150.890 ;
        RECT 69.780 150.630 70.040 150.890 ;
        RECT 78.520 150.290 78.780 150.550 ;
        RECT 51.840 149.950 52.100 150.210 ;
        RECT 52.300 149.950 52.560 150.210 ;
        RECT 69.780 149.950 70.040 150.210 ;
        RECT 77.140 149.950 77.400 150.210 ;
        RECT 79.440 151.310 79.700 151.570 ;
        RECT 83.120 151.650 83.380 151.910 ;
        RECT 84.500 151.650 84.760 151.910 ;
        RECT 87.260 151.650 87.520 151.910 ;
        RECT 82.660 151.310 82.920 151.570 ;
        RECT 83.580 151.310 83.840 151.570 ;
        RECT 82.200 150.970 82.460 151.230 ;
        RECT 88.640 151.310 88.900 151.570 ;
        RECT 80.820 150.630 81.080 150.890 ;
        RECT 84.960 150.630 85.220 150.890 ;
        RECT 82.200 150.290 82.460 150.550 ;
        RECT 91.860 151.650 92.120 151.910 ;
        RECT 97.380 151.650 97.640 151.910 ;
        RECT 97.840 151.650 98.100 151.910 ;
        RECT 102.440 151.650 102.700 151.910 ;
        RECT 104.740 151.650 105.000 151.910 ;
        RECT 109.340 151.650 109.600 151.910 ;
        RECT 99.220 151.310 99.480 151.570 ;
        RECT 101.060 151.310 101.320 151.570 ;
        RECT 111.640 151.310 111.900 151.570 ;
        RECT 87.260 150.290 87.520 150.550 ;
        RECT 89.100 150.630 89.360 150.890 ;
        RECT 114.400 150.970 114.660 151.230 ;
        RECT 117.620 151.310 117.880 151.570 ;
        RECT 116.700 150.970 116.960 151.230 ;
        RECT 89.100 149.950 89.360 150.210 ;
        RECT 90.940 149.950 91.200 150.210 ;
        RECT 97.380 150.290 97.640 150.550 ;
        RECT 102.440 150.290 102.700 150.550 ;
        RECT 106.120 150.630 106.380 150.890 ;
        RECT 110.720 150.630 110.980 150.890 ;
        RECT 122.680 151.310 122.940 151.570 ;
        RECT 118.540 150.970 118.800 151.230 ;
        RECT 124.520 150.970 124.780 151.230 ;
        RECT 124.980 150.970 125.240 151.230 ;
        RECT 134.640 151.650 134.900 151.910 ;
        RECT 137.400 151.650 137.660 151.910 ;
        RECT 130.040 150.970 130.300 151.230 ;
        RECT 131.880 150.970 132.140 151.230 ;
        RECT 139.700 151.310 139.960 151.570 ;
        RECT 140.160 150.970 140.420 151.230 ;
        RECT 129.580 150.630 129.840 150.890 ;
        RECT 136.480 150.630 136.740 150.890 ;
        RECT 98.760 149.950 99.020 150.210 ;
        RECT 99.680 149.950 99.940 150.210 ;
        RECT 108.420 149.950 108.680 150.210 ;
        RECT 112.100 149.950 112.360 150.210 ;
        RECT 118.540 149.950 118.800 150.210 ;
        RECT 125.440 149.950 125.700 150.210 ;
        RECT 132.800 149.950 133.060 150.210 ;
        RECT 40.170 149.440 40.430 149.700 ;
        RECT 40.490 149.440 40.750 149.700 ;
        RECT 40.810 149.440 41.070 149.700 ;
        RECT 41.130 149.440 41.390 149.700 ;
        RECT 41.450 149.440 41.710 149.700 ;
        RECT 41.770 149.440 42.030 149.700 ;
        RECT 70.170 149.440 70.430 149.700 ;
        RECT 70.490 149.440 70.750 149.700 ;
        RECT 70.810 149.440 71.070 149.700 ;
        RECT 71.130 149.440 71.390 149.700 ;
        RECT 71.450 149.440 71.710 149.700 ;
        RECT 71.770 149.440 72.030 149.700 ;
        RECT 100.170 149.440 100.430 149.700 ;
        RECT 100.490 149.440 100.750 149.700 ;
        RECT 100.810 149.440 101.070 149.700 ;
        RECT 101.130 149.440 101.390 149.700 ;
        RECT 101.450 149.440 101.710 149.700 ;
        RECT 101.770 149.440 102.030 149.700 ;
        RECT 130.170 149.440 130.430 149.700 ;
        RECT 130.490 149.440 130.750 149.700 ;
        RECT 130.810 149.440 131.070 149.700 ;
        RECT 131.130 149.440 131.390 149.700 ;
        RECT 131.450 149.440 131.710 149.700 ;
        RECT 131.770 149.440 132.030 149.700 ;
        RECT 52.760 148.930 53.020 149.190 ;
        RECT 54.140 148.930 54.400 149.190 ;
        RECT 38.500 148.590 38.760 148.850 ;
        RECT 50.920 148.250 51.180 148.510 ;
        RECT 45.400 147.910 45.660 148.170 ;
        RECT 55.060 147.570 55.320 147.830 ;
        RECT 58.280 147.910 58.540 148.170 ;
        RECT 61.960 147.570 62.220 147.830 ;
        RECT 68.400 147.910 68.660 148.170 ;
        RECT 76.680 148.930 76.940 149.190 ;
        RECT 78.980 148.930 79.240 149.190 ;
        RECT 83.580 148.930 83.840 149.190 ;
        RECT 89.100 148.930 89.360 149.190 ;
        RECT 126.820 148.930 127.080 149.190 ;
        RECT 127.740 148.930 128.000 149.190 ;
        RECT 142.000 148.930 142.260 149.190 ;
        RECT 71.160 147.910 71.420 148.170 ;
        RECT 72.080 147.910 72.340 148.170 ;
        RECT 72.540 147.570 72.800 147.830 ;
        RECT 74.840 147.910 75.100 148.170 ;
        RECT 82.660 148.250 82.920 148.510 ;
        RECT 84.500 148.250 84.760 148.510 ;
        RECT 84.960 148.250 85.220 148.510 ;
        RECT 88.640 148.250 88.900 148.510 ;
        RECT 75.300 147.570 75.560 147.830 ;
        RECT 87.260 147.910 87.520 148.170 ;
        RECT 89.100 147.910 89.360 148.170 ;
        RECT 89.560 147.910 89.820 148.170 ;
        RECT 90.020 147.910 90.280 148.170 ;
        RECT 90.940 147.910 91.200 148.170 ;
        RECT 98.300 148.250 98.560 148.510 ;
        RECT 102.440 148.250 102.700 148.510 ;
        RECT 108.420 148.250 108.680 148.510 ;
        RECT 110.720 148.250 110.980 148.510 ;
        RECT 38.960 147.230 39.220 147.490 ;
        RECT 54.600 147.230 54.860 147.490 ;
        RECT 67.940 147.230 68.200 147.490 ;
        RECT 71.620 147.230 71.880 147.490 ;
        RECT 72.080 147.230 72.340 147.490 ;
        RECT 73.920 147.230 74.180 147.490 ;
        RECT 77.140 147.230 77.400 147.490 ;
        RECT 91.400 147.570 91.660 147.830 ;
        RECT 98.760 147.910 99.020 148.170 ;
        RECT 113.940 148.250 114.200 148.510 ;
        RECT 118.540 148.250 118.800 148.510 ;
        RECT 112.560 147.910 112.820 148.170 ;
        RECT 113.020 147.910 113.280 148.170 ;
        RECT 99.680 147.570 99.940 147.830 ;
        RECT 103.360 147.570 103.620 147.830 ;
        RECT 106.120 147.570 106.380 147.830 ;
        RECT 109.800 147.570 110.060 147.830 ;
        RECT 117.160 147.910 117.420 148.170 ;
        RECT 122.680 147.910 122.940 148.170 ;
        RECT 144.300 148.590 144.560 148.850 ;
        RECT 84.960 147.230 85.220 147.490 ;
        RECT 88.640 147.230 88.900 147.490 ;
        RECT 100.600 147.230 100.860 147.490 ;
        RECT 106.580 147.230 106.840 147.490 ;
        RECT 108.420 147.230 108.680 147.490 ;
        RECT 109.340 147.230 109.600 147.490 ;
        RECT 110.260 147.230 110.520 147.490 ;
        RECT 110.720 147.230 110.980 147.490 ;
        RECT 123.600 147.230 123.860 147.490 ;
        RECT 143.840 148.250 144.100 148.510 ;
        RECT 142.920 147.910 143.180 148.170 ;
        RECT 130.040 147.230 130.300 147.490 ;
        RECT 138.780 147.230 139.040 147.490 ;
        RECT 55.170 146.720 55.430 146.980 ;
        RECT 55.490 146.720 55.750 146.980 ;
        RECT 55.810 146.720 56.070 146.980 ;
        RECT 56.130 146.720 56.390 146.980 ;
        RECT 56.450 146.720 56.710 146.980 ;
        RECT 56.770 146.720 57.030 146.980 ;
        RECT 85.170 146.720 85.430 146.980 ;
        RECT 85.490 146.720 85.750 146.980 ;
        RECT 85.810 146.720 86.070 146.980 ;
        RECT 86.130 146.720 86.390 146.980 ;
        RECT 86.450 146.720 86.710 146.980 ;
        RECT 86.770 146.720 87.030 146.980 ;
        RECT 115.170 146.720 115.430 146.980 ;
        RECT 115.490 146.720 115.750 146.980 ;
        RECT 115.810 146.720 116.070 146.980 ;
        RECT 116.130 146.720 116.390 146.980 ;
        RECT 116.450 146.720 116.710 146.980 ;
        RECT 116.770 146.720 117.030 146.980 ;
        RECT 145.170 146.720 145.430 146.980 ;
        RECT 145.490 146.720 145.750 146.980 ;
        RECT 145.810 146.720 146.070 146.980 ;
        RECT 146.130 146.720 146.390 146.980 ;
        RECT 146.450 146.720 146.710 146.980 ;
        RECT 146.770 146.720 147.030 146.980 ;
        RECT 38.960 146.210 39.220 146.470 ;
        RECT 39.420 146.210 39.680 146.470 ;
        RECT 51.840 146.210 52.100 146.470 ;
        RECT 52.300 146.210 52.560 146.470 ;
        RECT 52.760 146.210 53.020 146.470 ;
        RECT 54.140 146.210 54.400 146.470 ;
        RECT 67.940 146.210 68.200 146.470 ;
        RECT 61.960 145.870 62.220 146.130 ;
        RECT 42.180 144.850 42.440 145.110 ;
        RECT 60.580 145.530 60.840 145.790 ;
        RECT 54.140 145.190 54.400 145.450 ;
        RECT 54.600 145.190 54.860 145.450 ;
        RECT 67.940 145.530 68.200 145.790 ;
        RECT 68.400 145.530 68.660 145.790 ;
        RECT 69.780 145.870 70.040 146.130 ;
        RECT 72.540 146.210 72.800 146.470 ;
        RECT 78.520 146.210 78.780 146.470 ;
        RECT 82.660 146.210 82.920 146.470 ;
        RECT 87.720 146.210 87.980 146.470 ;
        RECT 89.100 146.210 89.360 146.470 ;
        RECT 75.300 145.530 75.560 145.790 ;
        RECT 76.220 145.530 76.480 145.790 ;
        RECT 80.360 145.530 80.620 145.790 ;
        RECT 80.820 145.530 81.080 145.790 ;
        RECT 84.040 145.530 84.300 145.790 ;
        RECT 71.160 145.190 71.420 145.450 ;
        RECT 71.620 145.190 71.880 145.450 ;
        RECT 82.200 145.190 82.460 145.450 ;
        RECT 85.880 145.190 86.140 145.450 ;
        RECT 88.180 145.530 88.440 145.790 ;
        RECT 99.680 146.210 99.940 146.470 ;
        RECT 101.060 146.210 101.320 146.470 ;
        RECT 110.720 146.210 110.980 146.470 ;
        RECT 111.640 146.210 111.900 146.470 ;
        RECT 90.480 145.530 90.740 145.790 ;
        RECT 91.400 145.530 91.660 145.790 ;
        RECT 94.620 145.530 94.880 145.790 ;
        RECT 103.360 145.870 103.620 146.130 ;
        RECT 102.440 145.530 102.700 145.790 ;
        RECT 103.820 145.530 104.080 145.790 ;
        RECT 107.040 145.530 107.300 145.790 ;
        RECT 107.960 145.530 108.220 145.790 ;
        RECT 109.340 145.530 109.600 145.790 ;
        RECT 111.180 145.530 111.440 145.790 ;
        RECT 112.100 145.530 112.360 145.790 ;
        RECT 113.020 145.530 113.280 145.790 ;
        RECT 114.400 145.530 114.660 145.790 ;
        RECT 115.320 145.530 115.580 145.790 ;
        RECT 117.160 145.530 117.420 145.790 ;
        RECT 119.000 146.210 119.260 146.470 ;
        RECT 119.460 145.530 119.720 145.790 ;
        RECT 120.380 145.530 120.640 145.790 ;
        RECT 121.760 145.530 122.020 145.790 ;
        RECT 132.800 146.210 133.060 146.470 ;
        RECT 145.220 146.210 145.480 146.470 ;
        RECT 123.600 145.870 123.860 146.130 ;
        RECT 130.040 145.530 130.300 145.790 ;
        RECT 132.340 145.530 132.600 145.790 ;
        RECT 143.840 145.870 144.100 146.130 ;
        RECT 74.380 144.850 74.640 145.110 ;
        RECT 90.020 144.850 90.280 145.110 ;
        RECT 96.920 145.190 97.180 145.450 ;
        RECT 100.600 145.190 100.860 145.450 ;
        RECT 113.940 145.190 114.200 145.450 ;
        RECT 112.100 144.850 112.360 145.110 ;
        RECT 126.820 145.190 127.080 145.450 ;
        RECT 127.740 145.190 128.000 145.450 ;
        RECT 128.660 144.850 128.920 145.110 ;
        RECT 33.440 144.510 33.700 144.770 ;
        RECT 74.840 144.510 75.100 144.770 ;
        RECT 75.300 144.510 75.560 144.770 ;
        RECT 77.140 144.510 77.400 144.770 ;
        RECT 82.200 144.510 82.460 144.770 ;
        RECT 87.260 144.510 87.520 144.770 ;
        RECT 91.400 144.510 91.660 144.770 ;
        RECT 96.460 144.510 96.720 144.770 ;
        RECT 98.300 144.510 98.560 144.770 ;
        RECT 100.600 144.510 100.860 144.770 ;
        RECT 102.440 144.510 102.700 144.770 ;
        RECT 105.200 144.510 105.460 144.770 ;
        RECT 108.880 144.510 109.140 144.770 ;
        RECT 113.020 144.510 113.280 144.770 ;
        RECT 116.240 144.510 116.500 144.770 ;
        RECT 120.380 144.510 120.640 144.770 ;
        RECT 123.140 144.510 123.400 144.770 ;
        RECT 140.160 145.530 140.420 145.790 ;
        RECT 140.620 145.530 140.880 145.790 ;
        RECT 142.920 145.190 143.180 145.450 ;
        RECT 141.540 144.850 141.800 145.110 ;
        RECT 40.170 144.000 40.430 144.260 ;
        RECT 40.490 144.000 40.750 144.260 ;
        RECT 40.810 144.000 41.070 144.260 ;
        RECT 41.130 144.000 41.390 144.260 ;
        RECT 41.450 144.000 41.710 144.260 ;
        RECT 41.770 144.000 42.030 144.260 ;
        RECT 70.170 144.000 70.430 144.260 ;
        RECT 70.490 144.000 70.750 144.260 ;
        RECT 70.810 144.000 71.070 144.260 ;
        RECT 71.130 144.000 71.390 144.260 ;
        RECT 71.450 144.000 71.710 144.260 ;
        RECT 71.770 144.000 72.030 144.260 ;
        RECT 100.170 144.000 100.430 144.260 ;
        RECT 100.490 144.000 100.750 144.260 ;
        RECT 100.810 144.000 101.070 144.260 ;
        RECT 101.130 144.000 101.390 144.260 ;
        RECT 101.450 144.000 101.710 144.260 ;
        RECT 101.770 144.000 102.030 144.260 ;
        RECT 130.170 144.000 130.430 144.260 ;
        RECT 130.490 144.000 130.750 144.260 ;
        RECT 130.810 144.000 131.070 144.260 ;
        RECT 131.130 144.000 131.390 144.260 ;
        RECT 131.450 144.000 131.710 144.260 ;
        RECT 131.770 144.000 132.030 144.260 ;
        RECT 39.420 143.490 39.680 143.750 ;
        RECT 54.140 143.490 54.400 143.750 ;
        RECT 38.500 142.470 38.760 142.730 ;
        RECT 74.380 143.150 74.640 143.410 ;
        RECT 75.300 143.150 75.560 143.410 ;
        RECT 42.640 142.130 42.900 142.390 ;
        RECT 45.860 142.130 46.120 142.390 ;
        RECT 64.260 142.470 64.520 142.730 ;
        RECT 77.600 142.470 77.860 142.730 ;
        RECT 82.200 143.490 82.460 143.750 ;
        RECT 87.260 143.490 87.520 143.750 ;
        RECT 93.700 143.490 93.960 143.750 ;
        RECT 96.460 143.490 96.720 143.750 ;
        RECT 98.300 143.490 98.560 143.750 ;
        RECT 105.200 143.490 105.460 143.750 ;
        RECT 108.420 143.490 108.680 143.750 ;
        RECT 112.100 143.490 112.360 143.750 ;
        RECT 113.020 143.490 113.280 143.750 ;
        RECT 113.480 143.490 113.740 143.750 ;
        RECT 121.300 143.490 121.560 143.750 ;
        RECT 132.340 143.490 132.600 143.750 ;
        RECT 82.200 142.470 82.460 142.730 ;
        RECT 91.400 142.810 91.660 143.070 ;
        RECT 90.940 142.470 91.200 142.730 ;
        RECT 102.440 142.470 102.700 142.730 ;
        RECT 108.880 142.470 109.140 142.730 ;
        RECT 112.560 142.470 112.820 142.730 ;
        RECT 113.940 142.470 114.200 142.730 ;
        RECT 116.240 142.470 116.500 142.730 ;
        RECT 123.140 142.810 123.400 143.070 ;
        RECT 126.820 142.810 127.080 143.070 ;
        RECT 128.660 142.810 128.920 143.070 ;
        RECT 120.380 142.470 120.640 142.730 ;
        RECT 128.200 142.470 128.460 142.730 ;
        RECT 143.840 142.810 144.100 143.070 ;
        RECT 144.300 142.470 144.560 142.730 ;
        RECT 38.500 141.790 38.760 142.050 ;
        RECT 50.000 141.790 50.260 142.050 ;
        RECT 53.680 141.790 53.940 142.050 ;
        RECT 55.060 141.790 55.320 142.050 ;
        RECT 59.200 141.790 59.460 142.050 ;
        RECT 63.340 141.790 63.600 142.050 ;
        RECT 75.760 141.790 76.020 142.050 ;
        RECT 78.980 141.790 79.240 142.050 ;
        RECT 83.120 141.790 83.380 142.050 ;
        RECT 89.100 141.790 89.360 142.050 ;
        RECT 91.400 141.790 91.660 142.050 ;
        RECT 96.460 141.790 96.720 142.050 ;
        RECT 99.680 141.790 99.940 142.050 ;
        RECT 104.740 141.790 105.000 142.050 ;
        RECT 117.160 141.790 117.420 142.050 ;
        RECT 117.620 141.790 117.880 142.050 ;
        RECT 120.380 141.790 120.640 142.050 ;
        RECT 125.440 141.790 125.700 142.050 ;
        RECT 128.660 141.790 128.920 142.050 ;
        RECT 132.800 141.790 133.060 142.050 ;
        RECT 136.940 141.790 137.200 142.050 ;
        RECT 141.080 141.790 141.340 142.050 ;
        RECT 55.170 141.280 55.430 141.540 ;
        RECT 55.490 141.280 55.750 141.540 ;
        RECT 55.810 141.280 56.070 141.540 ;
        RECT 56.130 141.280 56.390 141.540 ;
        RECT 56.450 141.280 56.710 141.540 ;
        RECT 56.770 141.280 57.030 141.540 ;
        RECT 85.170 141.280 85.430 141.540 ;
        RECT 85.490 141.280 85.750 141.540 ;
        RECT 85.810 141.280 86.070 141.540 ;
        RECT 86.130 141.280 86.390 141.540 ;
        RECT 86.450 141.280 86.710 141.540 ;
        RECT 86.770 141.280 87.030 141.540 ;
        RECT 115.170 141.280 115.430 141.540 ;
        RECT 115.490 141.280 115.750 141.540 ;
        RECT 115.810 141.280 116.070 141.540 ;
        RECT 116.130 141.280 116.390 141.540 ;
        RECT 116.450 141.280 116.710 141.540 ;
        RECT 116.770 141.280 117.030 141.540 ;
        RECT 145.170 141.280 145.430 141.540 ;
        RECT 145.490 141.280 145.750 141.540 ;
        RECT 145.810 141.280 146.070 141.540 ;
        RECT 146.130 141.280 146.390 141.540 ;
        RECT 146.450 141.280 146.710 141.540 ;
        RECT 146.770 141.280 147.030 141.540 ;
        RECT 60.580 140.430 60.840 140.690 ;
        RECT 64.260 140.090 64.520 140.350 ;
        RECT 110.260 140.090 110.520 140.350 ;
        RECT 117.160 140.430 117.420 140.690 ;
        RECT 141.540 140.770 141.800 141.030 ;
        RECT 124.060 140.090 124.320 140.350 ;
        RECT 53.680 139.750 53.940 140.010 ;
        RECT 84.500 139.750 84.760 140.010 ;
        RECT 80.820 139.410 81.080 139.670 ;
        RECT 96.920 139.750 97.180 140.010 ;
        RECT 60.580 131.300 61.580 132.300 ;
        RECT 64.930 131.300 65.930 132.300 ;
        RECT 60.600 104.080 61.600 105.080 ;
        RECT 99.670 132.160 99.950 132.440 ;
        RECT 101.580 131.400 102.580 132.400 ;
        RECT 103.810 132.160 104.090 132.440 ;
        RECT 105.930 131.400 106.930 132.400 ;
        RECT 101.600 104.080 102.600 105.080 ;
        RECT 60.600 55.030 61.600 56.030 ;
        RECT 132.790 132.160 133.070 132.440 ;
        RECT 136.930 132.160 137.210 132.440 ;
        RECT 141.070 132.160 141.350 132.440 ;
        RECT 142.580 131.400 143.580 132.400 ;
        RECT 145.210 132.200 145.490 132.480 ;
        RECT 146.930 131.400 147.930 132.400 ;
        RECT 142.600 104.080 143.600 105.080 ;
        RECT 101.600 55.030 102.600 56.030 ;
        RECT 142.600 55.030 143.600 56.030 ;
        RECT 143.530 51.630 144.470 52.570 ;
        RECT 126.660 49.455 127.545 50.340 ;
        RECT 122.870 47.265 123.735 48.130 ;
        RECT 24.300 22.000 25.300 23.000 ;
        RECT 31.600 18.065 31.900 18.365 ;
        RECT 22.800 15.615 23.800 16.615 ;
        RECT 31.600 13.465 31.900 13.765 ;
        RECT 33.800 13.700 34.800 14.700 ;
        RECT 29.900 12.065 30.200 12.365 ;
        RECT 30.950 12.065 31.250 12.365 ;
        RECT 35.600 8.000 36.600 9.000 ;
      LAYER met2 ;
        RECT 51.830 222.440 52.130 222.450 ;
        RECT 51.795 222.160 52.165 222.440 ;
        RECT 55.510 222.320 55.810 222.330 ;
        RECT 59.190 222.320 59.490 222.330 ;
        RECT 62.870 222.320 63.170 222.330 ;
        RECT 66.550 222.320 66.850 222.330 ;
        RECT 70.230 222.320 70.530 222.330 ;
        RECT 73.910 222.320 74.210 222.330 ;
        RECT 77.590 222.320 77.890 222.330 ;
        RECT 81.270 222.320 81.570 222.330 ;
        RECT 84.950 222.320 85.250 222.330 ;
        RECT 88.630 222.320 88.930 222.330 ;
        RECT 51.830 221.370 52.130 222.160 ;
        RECT 55.475 222.040 55.845 222.320 ;
        RECT 59.155 222.040 59.525 222.320 ;
        RECT 62.835 222.040 63.205 222.320 ;
        RECT 66.515 222.040 66.885 222.320 ;
        RECT 70.195 222.040 70.565 222.320 ;
        RECT 73.875 222.040 74.245 222.320 ;
        RECT 77.555 222.040 77.925 222.320 ;
        RECT 81.235 222.040 81.605 222.320 ;
        RECT 84.915 222.040 85.285 222.320 ;
        RECT 88.595 222.040 88.965 222.320 ;
        RECT 51.830 216.070 52.170 221.370 ;
        RECT 55.510 217.300 55.810 222.040 ;
        RECT 55.510 217.160 56.640 217.300 ;
        RECT 55.510 216.940 55.810 217.160 ;
        RECT 55.510 216.690 55.790 216.940 ;
        RECT 33.930 215.730 52.170 216.070 ;
        RECT 32.470 213.730 33.130 215.175 ;
        RECT 32.440 213.070 33.160 213.730 ;
        RECT 33.930 147.700 34.270 215.730 ;
        RECT 40.160 214.665 42.040 215.035 ;
        RECT 56.500 214.500 56.640 217.160 ;
        RECT 59.190 216.940 59.490 222.040 ;
        RECT 62.870 217.300 63.170 222.040 ;
        RECT 62.870 217.160 64.460 217.300 ;
        RECT 62.870 216.940 63.170 217.160 ;
        RECT 59.190 216.690 59.470 216.940 ;
        RECT 62.870 216.690 63.150 216.940 ;
        RECT 59.260 214.500 59.400 216.690 ;
        RECT 64.320 214.500 64.460 217.160 ;
        RECT 66.550 216.940 66.850 222.040 ;
        RECT 70.230 217.300 70.530 222.040 ;
        RECT 69.840 217.160 70.530 217.300 ;
        RECT 66.550 216.690 66.830 216.940 ;
        RECT 66.100 215.200 66.360 215.520 ;
        RECT 56.440 214.180 56.700 214.500 ;
        RECT 59.200 214.180 59.460 214.500 ;
        RECT 64.260 214.180 64.520 214.500 ;
        RECT 44.480 213.160 44.740 213.480 ;
        RECT 57.820 213.160 58.080 213.480 ;
        RECT 44.540 211.780 44.680 213.160 ;
        RECT 45.860 212.480 46.120 212.800 ;
        RECT 44.480 211.460 44.740 211.780 ;
        RECT 45.400 211.460 45.660 211.780 ;
        RECT 38.500 209.760 38.760 210.080 ;
        RECT 42.640 209.760 42.900 210.080 ;
        RECT 38.560 205.660 38.700 209.760 ;
        RECT 40.160 209.225 42.040 209.595 ;
        RECT 42.700 209.060 42.840 209.760 ;
        RECT 45.460 209.060 45.600 211.460 ;
        RECT 45.920 211.100 46.060 212.480 ;
        RECT 55.160 211.945 57.040 212.315 ;
        RECT 57.880 211.780 58.020 213.160 ;
        RECT 59.200 212.480 59.460 212.800 ;
        RECT 57.820 211.460 58.080 211.780 ;
        RECT 45.860 210.780 46.120 211.100 ;
        RECT 47.700 210.780 47.960 211.100 ;
        RECT 55.060 210.780 55.320 211.100 ;
        RECT 59.260 211.010 59.400 212.480 ;
        RECT 63.800 211.120 64.060 211.440 ;
        RECT 60.120 211.010 60.380 211.100 ;
        RECT 59.260 210.870 60.380 211.010 ;
        RECT 47.760 209.060 47.900 210.780 ;
        RECT 54.600 209.760 54.860 210.080 ;
        RECT 42.640 208.740 42.900 209.060 ;
        RECT 45.400 208.740 45.660 209.060 ;
        RECT 47.700 208.740 47.960 209.060 ;
        RECT 39.420 207.720 39.680 208.040 ;
        RECT 44.020 207.720 44.280 208.040 ;
        RECT 46.780 207.720 47.040 208.040 ;
        RECT 52.760 207.720 53.020 208.040 ;
        RECT 38.960 205.680 39.220 206.000 ;
        RECT 38.500 205.340 38.760 205.660 ;
        RECT 38.560 194.780 38.700 205.340 ;
        RECT 39.020 202.260 39.160 205.680 ;
        RECT 38.960 201.940 39.220 202.260 ;
        RECT 39.020 199.540 39.160 201.940 ;
        RECT 38.960 199.220 39.220 199.540 ;
        RECT 38.500 194.460 38.760 194.780 ;
        RECT 39.020 188.320 39.160 199.220 ;
        RECT 39.480 189.000 39.620 207.720 ;
        RECT 42.180 207.380 42.440 207.700 ;
        RECT 40.160 203.785 42.040 204.155 ;
        RECT 42.240 203.620 42.380 207.380 ;
        RECT 43.560 204.320 43.820 204.640 ;
        RECT 43.620 203.620 43.760 204.320 ;
        RECT 41.720 203.300 41.980 203.620 ;
        RECT 42.180 203.300 42.440 203.620 ;
        RECT 43.560 203.300 43.820 203.620 ;
        RECT 41.260 202.620 41.520 202.940 ;
        RECT 41.320 200.560 41.460 202.620 ;
        RECT 41.780 202.340 41.920 203.300 ;
        RECT 42.170 202.340 42.450 202.455 ;
        RECT 41.780 202.200 42.450 202.340 ;
        RECT 42.170 202.085 42.450 202.200 ;
        RECT 41.720 201.600 41.980 201.920 ;
        RECT 41.780 200.900 41.920 201.600 ;
        RECT 41.720 200.580 41.980 200.900 ;
        RECT 41.260 200.240 41.520 200.560 ;
        RECT 42.240 199.540 42.380 202.085 ;
        RECT 43.100 201.600 43.360 201.920 ;
        RECT 42.640 200.415 42.900 200.560 ;
        RECT 42.630 200.045 42.910 200.415 ;
        RECT 43.160 200.220 43.300 201.600 ;
        RECT 43.100 199.900 43.360 200.220 ;
        RECT 43.560 199.560 43.820 199.880 ;
        RECT 42.180 199.220 42.440 199.540 ;
        RECT 40.160 198.345 42.040 198.715 ;
        RECT 43.620 198.180 43.760 199.560 ;
        RECT 43.560 197.860 43.820 198.180 ;
        RECT 42.180 196.840 42.440 197.160 ;
        RECT 40.800 196.160 41.060 196.480 ;
        RECT 40.860 194.780 41.000 196.160 ;
        RECT 40.800 194.460 41.060 194.780 ;
        RECT 40.160 192.905 42.040 193.275 ;
        RECT 42.240 192.740 42.380 196.840 ;
        RECT 42.640 196.160 42.900 196.480 ;
        RECT 42.180 192.420 42.440 192.740 ;
        RECT 42.180 191.740 42.440 192.060 ;
        RECT 42.240 190.020 42.380 191.740 ;
        RECT 42.700 191.720 42.840 196.160 ;
        RECT 42.640 191.400 42.900 191.720 ;
        RECT 42.180 189.700 42.440 190.020 ;
        RECT 41.710 189.165 41.990 189.535 ;
        RECT 41.720 189.020 41.980 189.165 ;
        RECT 39.420 188.680 39.680 189.000 ;
        RECT 38.960 188.000 39.220 188.320 ;
        RECT 40.160 187.465 42.040 187.835 ;
        RECT 40.160 182.025 42.040 182.395 ;
        RECT 38.960 178.140 39.220 178.460 ;
        RECT 37.580 177.800 37.840 178.120 ;
        RECT 37.640 167.580 37.780 177.800 ;
        RECT 39.020 176.420 39.160 178.140 ;
        RECT 40.160 176.585 42.040 176.955 ;
        RECT 38.960 176.100 39.220 176.420 ;
        RECT 40.340 175.080 40.600 175.400 ;
        RECT 40.400 173.700 40.540 175.080 ;
        RECT 40.340 173.380 40.600 173.700 ;
        RECT 42.240 172.680 42.380 189.700 ;
        RECT 42.700 175.400 42.840 191.400 ;
        RECT 44.080 190.020 44.220 207.720 ;
        RECT 46.320 207.040 46.580 207.360 ;
        RECT 46.380 206.000 46.520 207.040 ;
        RECT 44.480 205.680 44.740 206.000 ;
        RECT 46.320 205.680 46.580 206.000 ;
        RECT 44.540 203.620 44.680 205.680 ;
        RECT 46.840 204.640 46.980 207.720 ;
        RECT 52.820 206.340 52.960 207.720 ;
        RECT 52.760 206.020 53.020 206.340 ;
        RECT 46.780 204.320 47.040 204.640 ;
        RECT 50.460 204.320 50.720 204.640 ;
        RECT 44.480 203.300 44.740 203.620 ;
        RECT 45.400 203.190 45.660 203.280 ;
        RECT 45.400 203.050 46.520 203.190 ;
        RECT 45.400 202.960 45.660 203.050 ;
        RECT 45.400 200.240 45.660 200.560 ;
        RECT 44.940 199.220 45.200 199.540 ;
        RECT 45.000 197.160 45.140 199.220 ;
        RECT 45.460 199.200 45.600 200.240 ;
        RECT 45.850 200.045 46.130 200.415 ;
        RECT 45.860 199.900 46.120 200.045 ;
        RECT 45.400 198.880 45.660 199.200 ;
        RECT 45.920 198.180 46.060 199.900 ;
        RECT 46.380 199.880 46.520 203.050 ;
        RECT 48.160 202.960 48.420 203.280 ;
        RECT 48.220 202.600 48.360 202.960 ;
        RECT 48.160 202.455 48.420 202.600 ;
        RECT 48.150 202.085 48.430 202.455 ;
        RECT 48.160 201.600 48.420 201.920 ;
        RECT 46.320 199.560 46.580 199.880 ;
        RECT 48.220 199.200 48.360 201.600 ;
        RECT 48.160 198.880 48.420 199.200 ;
        RECT 45.860 197.860 46.120 198.180 ;
        RECT 46.310 197.580 46.590 197.695 ;
        RECT 45.920 197.440 46.590 197.580 ;
        RECT 44.940 196.840 45.200 197.160 ;
        RECT 44.020 189.700 44.280 190.020 ;
        RECT 43.560 188.000 43.820 188.320 ;
        RECT 42.640 175.080 42.900 175.400 ;
        RECT 42.180 172.360 42.440 172.680 ;
        RECT 40.160 171.145 42.040 171.515 ;
        RECT 41.720 170.320 41.980 170.640 ;
        RECT 37.580 167.260 37.840 167.580 ;
        RECT 37.640 162.140 37.780 167.260 ;
        RECT 41.780 167.240 41.920 170.320 ;
        RECT 42.240 170.300 42.380 172.360 ;
        RECT 43.100 171.680 43.360 172.000 ;
        RECT 43.160 170.980 43.300 171.680 ;
        RECT 43.100 170.660 43.360 170.980 ;
        RECT 42.180 169.980 42.440 170.300 ;
        RECT 41.720 166.920 41.980 167.240 ;
        RECT 40.160 165.705 42.040 166.075 ;
        RECT 42.240 165.540 42.380 169.980 ;
        RECT 43.100 169.640 43.360 169.960 ;
        RECT 43.160 169.280 43.300 169.640 ;
        RECT 43.100 168.960 43.360 169.280 ;
        RECT 43.160 168.260 43.300 168.960 ;
        RECT 43.100 167.940 43.360 168.260 ;
        RECT 43.620 167.920 43.760 188.000 ;
        RECT 44.940 185.960 45.200 186.280 ;
        RECT 45.400 185.960 45.660 186.280 ;
        RECT 44.480 185.280 44.740 185.600 ;
        RECT 44.540 183.900 44.680 185.280 ;
        RECT 44.020 183.580 44.280 183.900 ;
        RECT 44.480 183.580 44.740 183.900 ;
        RECT 44.080 182.055 44.220 183.580 ;
        RECT 44.010 181.685 44.290 182.055 ;
        RECT 45.000 181.860 45.140 185.960 ;
        RECT 45.460 183.900 45.600 185.960 ;
        RECT 45.400 183.580 45.660 183.900 ;
        RECT 44.080 173.700 44.220 181.685 ;
        RECT 44.940 181.540 45.200 181.860 ;
        RECT 44.480 179.840 44.740 180.160 ;
        RECT 44.540 179.140 44.680 179.840 ;
        RECT 44.480 178.820 44.740 179.140 ;
        RECT 45.400 175.080 45.660 175.400 ;
        RECT 45.460 173.700 45.600 175.080 ;
        RECT 44.020 173.380 44.280 173.700 ;
        RECT 45.400 173.380 45.660 173.700 ;
        RECT 45.400 170.890 45.660 170.980 ;
        RECT 45.000 170.750 45.660 170.890 ;
        RECT 44.480 169.870 44.740 169.960 ;
        RECT 45.000 169.870 45.140 170.750 ;
        RECT 45.400 170.660 45.660 170.750 ;
        RECT 44.480 169.730 45.140 169.870 ;
        RECT 44.480 169.640 44.740 169.730 ;
        RECT 45.400 168.960 45.660 169.280 ;
        RECT 43.560 167.600 43.820 167.920 ;
        RECT 45.460 167.580 45.600 168.960 ;
        RECT 45.400 167.260 45.660 167.580 ;
        RECT 45.920 166.980 46.060 197.440 ;
        RECT 46.310 197.325 46.590 197.440 ;
        RECT 48.220 196.335 48.360 198.880 ;
        RECT 50.520 197.695 50.660 204.320 ;
        RECT 52.820 203.620 52.960 206.020 ;
        RECT 54.140 205.000 54.400 205.320 ;
        RECT 52.760 203.300 53.020 203.620 ;
        RECT 53.220 201.600 53.480 201.920 ;
        RECT 50.920 198.880 51.180 199.200 ;
        RECT 50.450 197.325 50.730 197.695 ;
        RECT 50.980 197.160 51.120 198.880 ;
        RECT 49.540 196.840 49.800 197.160 ;
        RECT 50.920 196.840 51.180 197.160 ;
        RECT 48.150 195.965 48.430 196.335 ;
        RECT 49.600 193.760 49.740 196.840 ;
        RECT 50.000 194.460 50.260 194.780 ;
        RECT 49.540 193.440 49.800 193.760 ;
        RECT 46.770 191.205 47.050 191.575 ;
        RECT 46.840 189.680 46.980 191.205 ;
        RECT 46.780 189.360 47.040 189.680 ;
        RECT 49.540 189.360 49.800 189.680 ;
        RECT 46.320 189.020 46.580 189.340 ;
        RECT 46.380 187.300 46.520 189.020 ;
        RECT 47.240 188.340 47.500 188.660 ;
        RECT 47.700 188.340 47.960 188.660 ;
        RECT 46.320 186.980 46.580 187.300 ;
        RECT 46.320 183.580 46.580 183.900 ;
        RECT 46.380 181.860 46.520 183.580 ;
        RECT 47.300 182.880 47.440 188.340 ;
        RECT 46.780 182.560 47.040 182.880 ;
        RECT 47.240 182.560 47.500 182.880 ;
        RECT 46.320 181.540 46.580 181.860 ;
        RECT 46.380 175.740 46.520 181.540 ;
        RECT 46.840 180.500 46.980 182.560 ;
        RECT 46.780 180.180 47.040 180.500 ;
        RECT 46.780 178.140 47.040 178.460 ;
        RECT 46.320 175.420 46.580 175.740 ;
        RECT 46.320 173.040 46.580 173.360 ;
        RECT 46.380 170.980 46.520 173.040 ;
        RECT 46.320 170.660 46.580 170.980 ;
        RECT 45.460 166.840 46.060 166.980 ;
        RECT 44.480 166.240 44.740 166.560 ;
        RECT 42.180 165.220 42.440 165.540 ;
        RECT 44.540 164.940 44.680 166.240 ;
        RECT 44.540 164.860 45.140 164.940 ;
        RECT 44.540 164.800 45.200 164.860 ;
        RECT 44.940 164.540 45.200 164.800 ;
        RECT 44.480 164.200 44.740 164.520 ;
        RECT 43.100 163.520 43.360 163.840 ;
        RECT 37.580 161.820 37.840 162.140 ;
        RECT 37.640 156.700 37.780 161.820 ;
        RECT 40.160 160.265 42.040 160.635 ;
        RECT 43.160 159.080 43.300 163.520 ;
        RECT 44.540 159.080 44.680 164.200 ;
        RECT 44.940 163.520 45.200 163.840 ;
        RECT 45.000 162.820 45.140 163.520 ;
        RECT 44.940 162.500 45.200 162.820 ;
        RECT 43.100 158.760 43.360 159.080 ;
        RECT 44.480 158.760 44.740 159.080 ;
        RECT 44.940 158.760 45.200 159.080 ;
        RECT 42.640 158.080 42.900 158.400 ;
        RECT 37.580 156.380 37.840 156.700 ;
        RECT 39.420 156.380 39.680 156.700 ;
        RECT 37.640 152.560 37.780 156.380 ;
        RECT 39.480 154.660 39.620 156.380 ;
        RECT 40.160 154.825 42.040 155.195 ;
        RECT 39.420 154.340 39.680 154.660 ;
        RECT 41.260 153.495 41.520 153.640 ;
        RECT 41.250 153.125 41.530 153.495 ;
        RECT 42.180 152.640 42.440 152.960 ;
        RECT 37.640 152.420 39.620 152.560 ;
        RECT 39.480 151.260 39.620 152.420 ;
        RECT 42.240 151.600 42.380 152.640 ;
        RECT 42.180 151.280 42.440 151.600 ;
        RECT 39.420 150.940 39.680 151.260 ;
        RECT 38.500 148.560 38.760 148.880 ;
        RECT 31.400 146.700 34.600 147.700 ;
        RECT 31.400 85.600 32.400 146.700 ;
        RECT 33.440 144.480 33.700 144.800 ;
        RECT 33.500 140.690 33.640 144.480 ;
        RECT 38.560 142.760 38.700 148.560 ;
        RECT 38.960 147.200 39.220 147.520 ;
        RECT 39.020 146.500 39.160 147.200 ;
        RECT 39.480 146.500 39.620 150.940 ;
        RECT 40.160 149.385 42.040 149.755 ;
        RECT 38.960 146.180 39.220 146.500 ;
        RECT 39.420 146.180 39.680 146.500 ;
        RECT 39.480 143.780 39.620 146.180 ;
        RECT 42.180 144.820 42.440 145.140 ;
        RECT 40.160 143.945 42.040 144.315 ;
        RECT 39.420 143.460 39.680 143.780 ;
        RECT 38.500 142.440 38.760 142.760 ;
        RECT 38.500 141.760 38.760 142.080 ;
        RECT 42.240 141.820 42.380 144.820 ;
        RECT 42.700 142.420 42.840 158.080 ;
        RECT 45.000 157.380 45.140 158.760 ;
        RECT 44.940 157.060 45.200 157.380 ;
        RECT 45.000 153.640 45.140 157.060 ;
        RECT 44.940 153.320 45.200 153.640 ;
        RECT 45.460 148.200 45.600 166.840 ;
        RECT 46.840 162.820 46.980 178.140 ;
        RECT 47.760 176.420 47.900 188.340 ;
        RECT 49.080 188.000 49.340 188.320 ;
        RECT 49.140 186.280 49.280 188.000 ;
        RECT 49.600 187.300 49.740 189.360 ;
        RECT 50.060 189.340 50.200 194.460 ;
        RECT 50.980 191.720 51.120 196.840 ;
        RECT 53.280 196.480 53.420 201.600 ;
        RECT 54.200 199.620 54.340 205.000 ;
        RECT 54.660 200.220 54.800 209.760 ;
        RECT 55.120 208.040 55.260 210.780 ;
        RECT 55.060 207.720 55.320 208.040 ;
        RECT 55.160 206.505 57.040 206.875 ;
        RECT 57.360 202.280 57.620 202.600 ;
        RECT 55.160 201.065 57.040 201.435 ;
        RECT 57.420 200.900 57.560 202.280 ;
        RECT 57.820 201.600 58.080 201.920 ;
        RECT 57.360 200.860 57.620 200.900 ;
        RECT 56.500 200.720 57.620 200.860 ;
        RECT 56.500 200.220 56.640 200.720 ;
        RECT 57.360 200.580 57.620 200.720 ;
        RECT 57.880 200.220 58.020 201.600 ;
        RECT 54.600 199.900 54.860 200.220 ;
        RECT 56.440 199.900 56.700 200.220 ;
        RECT 57.820 199.900 58.080 200.220 ;
        RECT 54.200 199.480 54.800 199.620 ;
        RECT 54.140 198.880 54.400 199.200 ;
        RECT 53.220 196.160 53.480 196.480 ;
        RECT 52.760 193.780 53.020 194.100 ;
        RECT 51.840 192.420 52.100 192.740 ;
        RECT 50.920 191.400 51.180 191.720 ;
        RECT 50.000 189.020 50.260 189.340 ;
        RECT 49.540 186.980 49.800 187.300 ;
        RECT 49.080 185.960 49.340 186.280 ;
        RECT 49.540 185.960 49.800 186.280 ;
        RECT 49.080 185.280 49.340 185.600 ;
        RECT 49.140 183.300 49.280 185.280 ;
        RECT 49.600 183.900 49.740 185.960 ;
        RECT 49.540 183.580 49.800 183.900 ;
        RECT 49.140 183.160 49.740 183.300 ;
        RECT 50.060 183.220 50.200 189.020 ;
        RECT 50.920 185.960 51.180 186.280 ;
        RECT 50.980 184.580 51.120 185.960 ;
        RECT 50.920 184.260 51.180 184.580 ;
        RECT 51.380 183.980 51.640 184.240 ;
        RECT 50.980 183.920 51.640 183.980 ;
        RECT 50.980 183.840 51.580 183.920 ;
        RECT 50.980 183.300 51.120 183.840 ;
        RECT 49.080 182.560 49.340 182.880 ;
        RECT 48.610 181.685 48.890 182.055 ;
        RECT 48.620 181.540 48.880 181.685 ;
        RECT 48.620 177.800 48.880 178.120 ;
        RECT 47.700 176.100 47.960 176.420 ;
        RECT 47.690 175.565 47.970 175.935 ;
        RECT 47.760 173.020 47.900 175.565 ;
        RECT 48.160 175.420 48.420 175.740 ;
        RECT 48.220 173.360 48.360 175.420 ;
        RECT 48.160 173.040 48.420 173.360 ;
        RECT 47.700 172.700 47.960 173.020 ;
        RECT 47.760 172.000 47.900 172.700 ;
        RECT 47.700 171.680 47.960 172.000 ;
        RECT 47.240 168.960 47.500 169.280 ;
        RECT 47.300 165.200 47.440 168.960 ;
        RECT 47.240 164.880 47.500 165.200 ;
        RECT 46.780 162.500 47.040 162.820 ;
        RECT 46.840 159.330 46.980 162.500 ;
        RECT 47.300 160.100 47.440 164.880 ;
        RECT 47.240 159.780 47.500 160.100 ;
        RECT 47.240 159.330 47.500 159.420 ;
        RECT 46.840 159.190 47.500 159.330 ;
        RECT 47.240 159.100 47.500 159.190 ;
        RECT 48.680 154.320 48.820 177.800 ;
        RECT 49.140 177.780 49.280 182.560 ;
        RECT 49.600 181.180 49.740 183.160 ;
        RECT 50.000 182.900 50.260 183.220 ;
        RECT 50.520 183.160 51.120 183.300 ;
        RECT 51.380 183.240 51.640 183.560 ;
        RECT 50.520 182.620 50.660 183.160 ;
        RECT 50.060 182.480 50.660 182.620 ;
        RECT 49.540 180.860 49.800 181.180 ;
        RECT 50.060 180.840 50.200 182.480 ;
        RECT 50.460 181.540 50.720 181.860 ;
        RECT 51.440 181.770 51.580 183.240 ;
        RECT 51.900 181.860 52.040 192.420 ;
        RECT 52.300 190.720 52.560 191.040 ;
        RECT 52.360 186.815 52.500 190.720 ;
        RECT 52.290 186.445 52.570 186.815 ;
        RECT 52.820 186.620 52.960 193.780 ;
        RECT 52.760 186.300 53.020 186.620 ;
        RECT 52.760 185.620 53.020 185.940 ;
        RECT 52.820 182.880 52.960 185.620 ;
        RECT 53.280 183.810 53.420 196.160 ;
        RECT 54.200 194.780 54.340 198.880 ;
        RECT 54.660 197.840 54.800 199.480 ;
        RECT 56.500 199.200 56.640 199.900 ;
        RECT 56.900 199.790 57.160 199.880 ;
        RECT 56.900 199.650 57.560 199.790 ;
        RECT 56.900 199.560 57.160 199.650 ;
        RECT 56.440 198.880 56.700 199.200 ;
        RECT 54.600 197.520 54.860 197.840 ;
        RECT 56.900 197.520 57.160 197.840 ;
        RECT 56.960 197.160 57.100 197.520 ;
        RECT 54.600 196.840 54.860 197.160 ;
        RECT 56.900 196.840 57.160 197.160 ;
        RECT 54.140 194.460 54.400 194.780 ;
        RECT 54.660 194.440 54.800 196.840 ;
        RECT 55.160 195.625 57.040 195.995 ;
        RECT 56.900 194.460 57.160 194.780 ;
        RECT 54.600 194.120 54.860 194.440 ;
        RECT 55.050 193.925 55.330 194.295 ;
        RECT 55.060 193.780 55.320 193.925 ;
        RECT 53.680 193.440 53.940 193.760 ;
        RECT 54.600 193.440 54.860 193.760 ;
        RECT 53.740 191.720 53.880 193.440 ;
        RECT 53.680 191.400 53.940 191.720 ;
        RECT 54.140 191.400 54.400 191.720 ;
        RECT 53.670 188.485 53.950 188.855 ;
        RECT 53.740 188.320 53.880 188.485 ;
        RECT 53.680 188.000 53.940 188.320 ;
        RECT 54.200 187.060 54.340 191.400 ;
        RECT 54.660 189.340 54.800 193.440 ;
        RECT 56.960 191.630 57.100 194.460 ;
        RECT 57.420 193.760 57.560 199.650 ;
        RECT 57.880 195.460 58.020 199.900 ;
        RECT 58.740 199.220 59.000 199.540 ;
        RECT 58.800 198.180 58.940 199.220 ;
        RECT 59.260 198.180 59.400 210.870 ;
        RECT 60.120 210.780 60.380 210.870 ;
        RECT 61.040 207.040 61.300 207.360 ;
        RECT 60.120 204.320 60.380 204.640 ;
        RECT 60.180 202.940 60.320 204.320 ;
        RECT 61.100 203.620 61.240 207.040 ;
        RECT 63.860 205.660 64.000 211.120 ;
        RECT 66.160 211.100 66.300 215.200 ;
        RECT 66.620 214.500 66.760 216.690 ;
        RECT 67.020 215.200 67.280 215.520 ;
        RECT 66.560 214.180 66.820 214.500 ;
        RECT 67.080 213.900 67.220 215.200 ;
        RECT 69.840 214.500 69.980 217.160 ;
        RECT 70.230 216.940 70.530 217.160 ;
        RECT 73.910 216.940 74.210 222.040 ;
        RECT 77.590 217.300 77.890 222.040 ;
        RECT 77.590 217.160 79.180 217.300 ;
        RECT 77.590 216.940 77.890 217.160 ;
        RECT 70.230 216.690 70.510 216.940 ;
        RECT 73.910 216.690 74.190 216.940 ;
        RECT 77.590 216.690 77.870 216.940 ;
        RECT 70.160 214.665 72.040 215.035 ;
        RECT 73.980 214.500 74.120 216.690 ;
        RECT 79.040 214.500 79.180 217.160 ;
        RECT 81.270 216.940 81.570 222.040 ;
        RECT 84.950 216.940 85.250 222.040 ;
        RECT 88.630 216.940 88.930 222.040 ;
        RECT 121.750 221.320 122.050 221.330 ;
        RECT 125.430 221.320 125.730 221.330 ;
        RECT 129.110 221.320 129.410 221.330 ;
        RECT 132.790 221.320 133.090 221.330 ;
        RECT 136.470 221.320 136.770 221.330 ;
        RECT 140.150 221.320 140.450 221.330 ;
        RECT 143.830 221.320 144.130 221.330 ;
        RECT 147.510 221.320 147.810 221.330 ;
        RECT 121.715 221.040 122.085 221.320 ;
        RECT 125.395 221.040 125.765 221.320 ;
        RECT 129.075 221.040 129.445 221.320 ;
        RECT 132.755 221.040 133.125 221.320 ;
        RECT 136.435 221.040 136.805 221.320 ;
        RECT 140.115 221.040 140.485 221.320 ;
        RECT 143.795 221.040 144.165 221.320 ;
        RECT 147.475 221.040 147.845 221.320 ;
        RECT 121.750 216.940 122.050 221.040 ;
        RECT 125.430 216.940 125.730 221.040 ;
        RECT 129.110 216.940 129.410 221.040 ;
        RECT 132.790 217.300 133.090 221.040 ;
        RECT 132.790 217.160 134.380 217.300 ;
        RECT 132.790 216.940 133.090 217.160 ;
        RECT 81.270 216.690 81.550 216.940 ;
        RECT 84.950 216.690 85.230 216.940 ;
        RECT 88.630 216.690 88.910 216.940 ;
        RECT 121.750 216.690 122.030 216.940 ;
        RECT 125.430 216.690 125.710 216.940 ;
        RECT 129.110 216.690 129.390 216.940 ;
        RECT 132.790 216.690 133.070 216.940 ;
        RECT 81.340 214.500 81.480 216.690 ;
        RECT 85.020 214.500 85.160 216.690 ;
        RECT 88.700 214.500 88.840 216.690 ;
        RECT 114.400 215.540 114.660 215.860 ;
        RECT 119.460 215.540 119.720 215.860 ;
        RECT 105.660 215.200 105.920 215.520 ;
        RECT 107.040 215.200 107.300 215.520 ;
        RECT 100.160 214.665 102.040 215.035 ;
        RECT 105.720 214.500 105.860 215.200 ;
        RECT 69.780 214.180 70.040 214.500 ;
        RECT 73.920 214.180 74.180 214.500 ;
        RECT 78.980 214.180 79.240 214.500 ;
        RECT 81.280 214.180 81.540 214.500 ;
        RECT 84.960 214.180 85.220 214.500 ;
        RECT 88.640 214.180 88.900 214.500 ;
        RECT 105.660 214.180 105.920 214.500 ;
        RECT 66.620 213.760 67.220 213.900 ;
        RECT 66.620 211.780 66.760 213.760 ;
        RECT 71.620 213.500 71.880 213.820 ;
        RECT 67.020 212.820 67.280 213.140 ;
        RECT 67.940 212.820 68.200 213.140 ;
        RECT 66.560 211.460 66.820 211.780 ;
        RECT 66.100 210.780 66.360 211.100 ;
        RECT 64.260 209.760 64.520 210.080 ;
        RECT 64.320 207.700 64.460 209.760 ;
        RECT 64.720 208.400 64.980 208.720 ;
        RECT 64.260 207.380 64.520 207.700 ;
        RECT 63.800 205.340 64.060 205.660 ;
        RECT 62.420 205.000 62.680 205.320 ;
        RECT 61.040 203.300 61.300 203.620 ;
        RECT 60.120 202.850 60.380 202.940 ;
        RECT 59.720 202.710 60.380 202.850 ;
        RECT 58.740 197.860 59.000 198.180 ;
        RECT 59.200 197.860 59.460 198.180 ;
        RECT 59.190 196.900 59.470 197.015 ;
        RECT 58.340 196.760 59.470 196.900 ;
        RECT 57.820 195.140 58.080 195.460 ;
        RECT 57.810 194.605 58.090 194.975 ;
        RECT 57.360 193.440 57.620 193.760 ;
        RECT 57.420 192.400 57.560 193.440 ;
        RECT 57.360 192.080 57.620 192.400 ;
        RECT 57.360 191.630 57.620 191.720 ;
        RECT 56.960 191.490 57.620 191.630 ;
        RECT 57.360 191.400 57.620 191.490 ;
        RECT 55.160 190.185 57.040 190.555 ;
        RECT 54.600 189.020 54.860 189.340 ;
        RECT 56.900 188.000 57.160 188.320 ;
        RECT 54.200 186.920 54.800 187.060 ;
        RECT 54.140 185.960 54.400 186.280 ;
        RECT 53.680 183.810 53.940 183.900 ;
        RECT 53.280 183.670 53.940 183.810 ;
        RECT 53.680 183.580 53.940 183.670 ;
        RECT 52.300 182.560 52.560 182.880 ;
        RECT 52.760 182.560 53.020 182.880 ;
        RECT 50.980 181.630 51.580 181.770 ;
        RECT 50.000 180.520 50.260 180.840 ;
        RECT 50.000 179.840 50.260 180.160 ;
        RECT 50.060 178.800 50.200 179.840 ;
        RECT 50.520 179.140 50.660 181.540 ;
        RECT 50.980 179.140 51.120 181.630 ;
        RECT 51.840 181.540 52.100 181.860 ;
        RECT 52.360 181.260 52.500 182.560 ;
        RECT 51.440 181.120 52.500 181.260 ;
        RECT 50.460 178.820 50.720 179.140 ;
        RECT 50.920 178.820 51.180 179.140 ;
        RECT 50.000 178.480 50.260 178.800 ;
        RECT 49.080 177.460 49.340 177.780 ;
        RECT 50.060 176.420 50.200 178.480 ;
        RECT 50.910 178.285 51.190 178.655 ;
        RECT 50.920 178.140 51.180 178.285 ;
        RECT 50.000 176.100 50.260 176.420 ;
        RECT 50.920 175.080 51.180 175.400 ;
        RECT 49.540 174.740 49.800 175.060 ;
        RECT 49.600 172.680 49.740 174.740 ;
        RECT 50.980 173.700 51.120 175.080 ;
        RECT 50.920 173.380 51.180 173.700 ;
        RECT 51.440 173.020 51.580 181.120 ;
        RECT 52.300 180.070 52.560 180.160 ;
        RECT 51.900 179.930 52.560 180.070 ;
        RECT 51.900 175.400 52.040 179.930 ;
        RECT 52.300 179.840 52.560 179.930 ;
        RECT 51.840 175.080 52.100 175.400 ;
        RECT 52.300 175.080 52.560 175.400 ;
        RECT 52.360 173.700 52.500 175.080 ;
        RECT 52.300 173.380 52.560 173.700 ;
        RECT 51.380 172.700 51.640 173.020 ;
        RECT 51.840 172.700 52.100 173.020 ;
        RECT 49.540 172.590 49.800 172.680 ;
        RECT 49.540 172.450 50.200 172.590 ;
        RECT 49.540 172.360 49.800 172.450 ;
        RECT 50.060 167.240 50.200 172.450 ;
        RECT 51.440 170.980 51.580 172.700 ;
        RECT 51.380 170.660 51.640 170.980 ;
        RECT 50.000 166.920 50.260 167.240 ;
        RECT 51.900 166.560 52.040 172.700 ;
        RECT 52.300 171.680 52.560 172.000 ;
        RECT 52.360 170.300 52.500 171.680 ;
        RECT 52.300 169.980 52.560 170.300 ;
        RECT 52.360 168.260 52.500 169.980 ;
        RECT 52.300 167.940 52.560 168.260 ;
        RECT 51.840 166.240 52.100 166.560 ;
        RECT 50.920 163.520 51.180 163.840 ;
        RECT 50.460 156.720 50.720 157.040 ;
        RECT 48.620 154.000 48.880 154.320 ;
        RECT 48.680 153.640 48.820 154.000 ;
        RECT 50.520 153.640 50.660 156.720 ;
        RECT 45.860 153.320 46.120 153.640 ;
        RECT 48.620 153.320 48.880 153.640 ;
        RECT 50.460 153.320 50.720 153.640 ;
        RECT 45.920 151.940 46.060 153.320 ;
        RECT 45.860 151.620 46.120 151.940 ;
        RECT 50.980 148.540 51.120 163.520 ;
        RECT 51.900 162.480 52.040 166.240 ;
        RECT 51.840 162.160 52.100 162.480 ;
        RECT 51.380 161.820 51.640 162.140 ;
        RECT 51.440 159.080 51.580 161.820 ;
        RECT 52.300 161.480 52.560 161.800 ;
        RECT 52.360 160.100 52.500 161.480 ;
        RECT 52.300 159.780 52.560 160.100 ;
        RECT 51.380 158.760 51.640 159.080 ;
        RECT 51.440 153.640 51.580 158.760 ;
        RECT 52.360 157.040 52.500 159.780 ;
        RECT 52.300 156.720 52.560 157.040 ;
        RECT 52.820 154.660 52.960 182.560 ;
        RECT 54.200 180.500 54.340 185.960 ;
        RECT 54.660 183.560 54.800 186.920 ;
        RECT 56.960 186.280 57.100 188.000 ;
        RECT 56.900 185.960 57.160 186.280 ;
        RECT 55.160 184.745 57.040 185.115 ;
        RECT 54.600 183.240 54.860 183.560 ;
        RECT 55.060 180.860 55.320 181.180 ;
        RECT 54.140 180.180 54.400 180.500 ;
        RECT 55.120 180.160 55.260 180.860 ;
        RECT 53.680 179.840 53.940 180.160 ;
        RECT 55.060 180.070 55.320 180.160 ;
        RECT 54.660 179.930 55.320 180.070 ;
        RECT 53.740 179.140 53.880 179.840 ;
        RECT 53.680 178.820 53.940 179.140 ;
        RECT 53.220 177.460 53.480 177.780 ;
        RECT 53.280 173.020 53.420 177.460 ;
        RECT 54.140 177.120 54.400 177.440 ;
        RECT 54.200 176.080 54.340 177.120 ;
        RECT 53.680 175.935 53.940 176.080 ;
        RECT 53.670 175.565 53.950 175.935 ;
        RECT 54.140 175.760 54.400 176.080 ;
        RECT 54.660 175.400 54.800 179.930 ;
        RECT 55.060 179.840 55.320 179.930 ;
        RECT 55.160 179.305 57.040 179.675 ;
        RECT 53.680 175.080 53.940 175.400 ;
        RECT 54.600 175.080 54.860 175.400 ;
        RECT 53.740 173.700 53.880 175.080 ;
        RECT 54.600 174.460 54.860 174.720 ;
        RECT 54.200 174.400 54.860 174.460 ;
        RECT 54.200 174.320 54.800 174.400 ;
        RECT 53.680 173.380 53.940 173.700 ;
        RECT 53.220 172.700 53.480 173.020 ;
        RECT 54.200 172.000 54.340 174.320 ;
        RECT 55.160 173.865 57.040 174.235 ;
        RECT 57.420 173.020 57.560 191.400 ;
        RECT 57.880 186.190 58.020 194.605 ;
        RECT 58.340 194.440 58.480 196.760 ;
        RECT 59.190 196.645 59.470 196.760 ;
        RECT 58.740 196.160 59.000 196.480 ;
        RECT 59.200 196.160 59.460 196.480 ;
        RECT 58.800 195.460 58.940 196.160 ;
        RECT 58.740 195.140 59.000 195.460 ;
        RECT 58.280 194.120 58.540 194.440 ;
        RECT 59.260 194.100 59.400 196.160 ;
        RECT 59.720 194.690 59.860 202.710 ;
        RECT 60.120 202.620 60.380 202.710 ;
        RECT 60.120 200.580 60.380 200.900 ;
        RECT 60.180 200.220 60.320 200.580 ;
        RECT 60.120 199.900 60.380 200.220 ;
        RECT 60.580 199.110 60.840 199.200 ;
        RECT 60.180 198.970 60.840 199.110 ;
        RECT 60.180 195.655 60.320 198.970 ;
        RECT 60.580 198.880 60.840 198.970 ;
        RECT 60.580 196.840 60.840 197.160 ;
        RECT 60.110 195.285 60.390 195.655 ;
        RECT 60.120 194.690 60.380 194.780 ;
        RECT 59.720 194.550 60.380 194.690 ;
        RECT 59.200 193.780 59.460 194.100 ;
        RECT 59.260 192.060 59.400 193.780 ;
        RECT 59.720 192.740 59.860 194.550 ;
        RECT 60.120 194.460 60.380 194.550 ;
        RECT 59.660 192.420 59.920 192.740 ;
        RECT 59.200 191.740 59.460 192.060 ;
        RECT 60.640 186.960 60.780 196.840 ;
        RECT 61.100 192.060 61.240 203.300 ;
        RECT 61.500 198.880 61.760 199.200 ;
        RECT 61.560 197.580 61.700 198.880 ;
        RECT 61.560 197.500 62.160 197.580 ;
        RECT 61.560 197.440 62.220 197.500 ;
        RECT 61.960 197.180 62.220 197.440 ;
        RECT 61.040 191.740 61.300 192.060 ;
        RECT 62.480 191.970 62.620 205.000 ;
        RECT 62.880 204.660 63.140 204.980 ;
        RECT 62.940 203.620 63.080 204.660 ;
        RECT 63.800 204.320 64.060 204.640 ;
        RECT 62.880 203.300 63.140 203.620 ;
        RECT 62.880 199.900 63.140 200.220 ;
        RECT 62.940 197.160 63.080 199.900 ;
        RECT 63.340 199.220 63.600 199.540 ;
        RECT 62.880 196.840 63.140 197.160 ;
        RECT 62.020 191.830 62.620 191.970 ;
        RECT 62.020 191.380 62.160 191.830 ;
        RECT 61.960 191.060 62.220 191.380 ;
        RECT 62.420 191.060 62.680 191.380 ;
        RECT 61.040 190.720 61.300 191.040 ;
        RECT 61.100 189.680 61.240 190.720 ;
        RECT 61.040 189.360 61.300 189.680 ;
        RECT 61.040 188.000 61.300 188.320 ;
        RECT 61.100 187.300 61.240 188.000 ;
        RECT 61.040 186.980 61.300 187.300 ;
        RECT 60.580 186.640 60.840 186.960 ;
        RECT 62.480 186.700 62.620 191.060 ;
        RECT 63.400 189.250 63.540 199.220 ;
        RECT 62.020 186.560 62.620 186.700 ;
        RECT 62.940 189.110 63.540 189.250 ;
        RECT 58.280 186.190 58.540 186.280 ;
        RECT 57.880 186.050 59.400 186.190 ;
        RECT 58.280 185.960 58.540 186.050 ;
        RECT 58.280 183.580 58.540 183.900 ;
        RECT 58.740 183.580 59.000 183.900 ;
        RECT 58.340 179.140 58.480 183.580 ;
        RECT 58.800 180.840 58.940 183.580 ;
        RECT 59.260 180.840 59.400 186.050 ;
        RECT 59.660 185.960 59.920 186.280 ;
        RECT 59.720 184.580 59.860 185.960 ;
        RECT 60.120 185.620 60.380 185.940 ;
        RECT 59.660 184.260 59.920 184.580 ;
        RECT 60.180 183.980 60.320 185.620 ;
        RECT 59.720 183.840 60.320 183.980 ;
        RECT 59.720 183.560 59.860 183.840 ;
        RECT 61.040 183.580 61.300 183.900 ;
        RECT 59.660 183.240 59.920 183.560 ;
        RECT 58.740 180.520 59.000 180.840 ;
        RECT 59.200 180.520 59.460 180.840 ;
        RECT 58.800 179.140 58.940 180.520 ;
        RECT 58.280 178.820 58.540 179.140 ;
        RECT 58.740 178.820 59.000 179.140 ;
        RECT 59.200 178.820 59.460 179.140 ;
        RECT 59.260 175.400 59.400 178.820 ;
        RECT 58.280 175.080 58.540 175.400 ;
        RECT 59.200 175.080 59.460 175.400 ;
        RECT 57.360 172.700 57.620 173.020 ;
        RECT 54.600 172.360 54.860 172.680 ;
        RECT 54.140 171.680 54.400 172.000 ;
        RECT 54.200 162.820 54.340 171.680 ;
        RECT 54.140 162.500 54.400 162.820 ;
        RECT 54.140 161.480 54.400 161.800 ;
        RECT 54.200 159.080 54.340 161.480 ;
        RECT 54.140 158.760 54.400 159.080 ;
        RECT 54.200 157.380 54.340 158.760 ;
        RECT 54.140 157.060 54.400 157.380 ;
        RECT 52.760 154.340 53.020 154.660 ;
        RECT 51.380 153.320 51.640 153.640 ;
        RECT 51.440 151.600 51.580 153.320 ;
        RECT 54.660 152.560 54.800 172.360 ;
        RECT 58.340 169.620 58.480 175.080 ;
        RECT 59.720 175.060 59.860 183.240 ;
        RECT 61.100 181.180 61.240 183.580 ;
        RECT 61.500 182.900 61.760 183.220 ;
        RECT 61.560 181.180 61.700 182.900 ;
        RECT 61.040 180.860 61.300 181.180 ;
        RECT 61.500 180.860 61.760 181.180 ;
        RECT 61.560 178.120 61.700 180.860 ;
        RECT 61.500 177.800 61.760 178.120 ;
        RECT 60.120 177.120 60.380 177.440 ;
        RECT 60.180 176.330 60.320 177.120 ;
        RECT 60.580 176.330 60.840 176.420 ;
        RECT 60.180 176.190 60.840 176.330 ;
        RECT 60.580 176.100 60.840 176.190 ;
        RECT 61.030 175.565 61.310 175.935 ;
        RECT 61.560 175.740 61.700 177.800 ;
        RECT 61.100 175.060 61.240 175.565 ;
        RECT 61.500 175.420 61.760 175.740 ;
        RECT 59.660 174.740 59.920 175.060 ;
        RECT 61.040 174.740 61.300 175.060 ;
        RECT 60.580 174.400 60.840 174.720 ;
        RECT 59.660 173.380 59.920 173.700 ;
        RECT 58.740 171.680 59.000 172.000 ;
        RECT 58.280 169.300 58.540 169.620 ;
        RECT 55.160 168.425 57.040 168.795 ;
        RECT 58.280 167.260 58.540 167.580 ;
        RECT 55.160 162.985 57.040 163.355 ;
        RECT 55.060 161.820 55.320 162.140 ;
        RECT 55.120 159.420 55.260 161.820 ;
        RECT 55.060 159.100 55.320 159.420 ;
        RECT 55.160 157.545 57.040 157.915 ;
        RECT 58.340 156.700 58.480 167.260 ;
        RECT 58.800 167.240 58.940 171.680 ;
        RECT 59.720 167.240 59.860 173.380 ;
        RECT 60.640 173.360 60.780 174.400 ;
        RECT 60.580 173.040 60.840 173.360 ;
        RECT 60.640 169.620 60.780 173.040 ;
        RECT 61.560 172.680 61.700 175.420 ;
        RECT 61.500 172.360 61.760 172.680 ;
        RECT 61.040 170.660 61.300 170.980 ;
        RECT 61.100 169.960 61.240 170.660 ;
        RECT 62.020 170.300 62.160 186.560 ;
        RECT 62.940 186.280 63.080 189.110 ;
        RECT 63.340 188.340 63.600 188.660 ;
        RECT 62.880 185.960 63.140 186.280 ;
        RECT 63.400 185.940 63.540 188.340 ;
        RECT 63.340 185.620 63.600 185.940 ;
        RECT 62.880 185.280 63.140 185.600 ;
        RECT 62.420 183.920 62.680 184.240 ;
        RECT 61.960 169.980 62.220 170.300 ;
        RECT 61.040 169.640 61.300 169.960 ;
        RECT 60.580 169.300 60.840 169.620 ;
        RECT 61.960 168.960 62.220 169.280 ;
        RECT 60.580 167.940 60.840 168.260 ;
        RECT 58.740 166.920 59.000 167.240 ;
        RECT 59.660 166.920 59.920 167.240 ;
        RECT 58.800 164.860 58.940 166.920 ;
        RECT 58.740 164.540 59.000 164.860 ;
        RECT 59.720 161.120 59.860 166.920 ;
        RECT 60.640 164.520 60.780 167.940 ;
        RECT 62.020 167.240 62.160 168.960 ;
        RECT 61.960 166.920 62.220 167.240 ;
        RECT 61.500 166.580 61.760 166.900 ;
        RECT 61.560 164.860 61.700 166.580 ;
        RECT 61.500 164.540 61.760 164.860 ;
        RECT 60.580 164.200 60.840 164.520 ;
        RECT 60.640 162.820 60.780 164.200 ;
        RECT 62.480 163.840 62.620 183.920 ;
        RECT 62.940 182.880 63.080 185.280 ;
        RECT 63.860 183.220 64.000 204.320 ;
        RECT 64.780 202.600 64.920 208.400 ;
        RECT 65.640 204.320 65.900 204.640 ;
        RECT 65.700 203.620 65.840 204.320 ;
        RECT 65.640 203.300 65.900 203.620 ;
        RECT 64.720 202.280 64.980 202.600 ;
        RECT 64.260 195.140 64.520 195.460 ;
        RECT 64.320 188.660 64.460 195.140 ;
        RECT 64.260 188.340 64.520 188.660 ;
        RECT 63.800 182.900 64.060 183.220 ;
        RECT 62.880 182.560 63.140 182.880 ;
        RECT 62.940 180.500 63.080 182.560 ;
        RECT 64.780 180.840 64.920 202.280 ;
        RECT 66.620 200.860 66.760 211.460 ;
        RECT 67.080 211.100 67.220 212.820 ;
        RECT 67.020 210.780 67.280 211.100 ;
        RECT 67.080 203.280 67.220 210.780 ;
        RECT 67.480 207.720 67.740 208.040 ;
        RECT 67.020 202.960 67.280 203.280 ;
        RECT 67.540 202.600 67.680 207.720 ;
        RECT 68.000 206.000 68.140 212.820 ;
        RECT 68.860 212.480 69.120 212.800 ;
        RECT 68.920 211.100 69.060 212.480 ;
        RECT 71.680 211.780 71.820 213.500 ;
        RECT 72.540 213.160 72.800 213.480 ;
        RECT 76.220 213.160 76.480 213.480 ;
        RECT 78.060 213.160 78.320 213.480 ;
        RECT 84.040 213.160 84.300 213.480 ;
        RECT 99.680 213.160 99.940 213.480 ;
        RECT 71.620 211.460 71.880 211.780 ;
        RECT 68.860 210.780 69.120 211.100 ;
        RECT 70.160 209.225 72.040 209.595 ;
        RECT 72.600 209.060 72.740 213.160 ;
        RECT 73.000 212.480 73.260 212.800 ;
        RECT 73.060 211.780 73.200 212.480 ;
        RECT 73.000 211.460 73.260 211.780 ;
        RECT 73.460 210.780 73.720 211.100 ;
        RECT 72.540 208.740 72.800 209.060 ;
        RECT 72.080 207.720 72.340 208.040 ;
        RECT 72.140 206.000 72.280 207.720 ;
        RECT 67.940 205.910 68.200 206.000 ;
        RECT 67.940 205.770 68.600 205.910 ;
        RECT 67.940 205.680 68.200 205.770 ;
        RECT 67.940 204.320 68.200 204.640 ;
        RECT 67.480 202.280 67.740 202.600 ;
        RECT 66.160 200.720 66.760 200.860 ;
        RECT 65.640 197.180 65.900 197.500 ;
        RECT 65.700 196.820 65.840 197.180 ;
        RECT 65.640 196.500 65.900 196.820 ;
        RECT 65.180 196.160 65.440 196.480 ;
        RECT 65.240 191.720 65.380 196.160 ;
        RECT 65.700 192.060 65.840 196.500 ;
        RECT 66.160 194.780 66.300 200.720 ;
        RECT 66.560 198.880 66.820 199.200 ;
        RECT 66.620 195.120 66.760 198.880 ;
        RECT 68.000 197.580 68.140 204.320 ;
        RECT 68.460 203.620 68.600 205.770 ;
        RECT 72.080 205.680 72.340 206.000 ;
        RECT 73.520 205.060 73.660 210.780 ;
        RECT 73.920 209.760 74.180 210.080 ;
        RECT 73.980 206.000 74.120 209.760 ;
        RECT 76.280 209.060 76.420 213.160 ;
        RECT 76.680 212.820 76.940 213.140 ;
        RECT 76.220 208.740 76.480 209.060 ;
        RECT 74.380 207.720 74.640 208.040 ;
        RECT 76.220 207.720 76.480 208.040 ;
        RECT 73.920 205.680 74.180 206.000 ;
        RECT 74.440 205.320 74.580 207.720 ;
        RECT 76.280 206.340 76.420 207.720 ;
        RECT 76.220 206.020 76.480 206.340 ;
        RECT 73.910 205.060 74.190 205.175 ;
        RECT 73.520 204.920 74.190 205.060 ;
        RECT 74.380 205.000 74.640 205.320 ;
        RECT 73.520 204.640 73.660 204.920 ;
        RECT 73.910 204.805 74.190 204.920 ;
        RECT 73.460 204.320 73.720 204.640 ;
        RECT 70.160 203.785 72.040 204.155 ;
        RECT 68.400 203.300 68.660 203.620 ;
        RECT 70.700 201.940 70.960 202.260 ;
        RECT 69.780 201.600 70.040 201.920 ;
        RECT 69.840 199.880 69.980 201.600 ;
        RECT 70.760 200.900 70.900 201.940 ;
        RECT 74.440 201.920 74.580 205.000 ;
        RECT 74.380 201.600 74.640 201.920 ;
        RECT 70.700 200.580 70.960 200.900 ;
        RECT 76.740 200.860 76.880 212.820 ;
        RECT 78.120 211.780 78.260 213.160 ;
        RECT 80.820 212.820 81.080 213.140 ;
        RECT 81.740 212.820 82.000 213.140 ;
        RECT 78.060 211.460 78.320 211.780 ;
        RECT 77.140 210.780 77.400 211.100 ;
        RECT 77.200 205.660 77.340 210.780 ;
        RECT 78.980 210.440 79.240 210.760 ;
        RECT 79.900 210.440 80.160 210.760 ;
        RECT 79.040 208.040 79.180 210.440 ;
        RECT 79.960 210.080 80.100 210.440 ;
        RECT 79.900 209.760 80.160 210.080 ;
        RECT 79.960 208.040 80.100 209.760 ;
        RECT 78.980 207.720 79.240 208.040 ;
        RECT 79.900 207.720 80.160 208.040 ;
        RECT 77.140 205.340 77.400 205.660 ;
        RECT 76.740 200.720 77.340 200.860 ;
        RECT 72.540 199.900 72.800 200.220 ;
        RECT 75.760 199.900 76.020 200.220 ;
        RECT 69.780 199.560 70.040 199.880 ;
        RECT 67.080 197.440 68.140 197.580 ;
        RECT 67.080 196.480 67.220 197.440 ;
        RECT 67.470 196.645 67.750 197.015 ;
        RECT 67.480 196.500 67.740 196.645 ;
        RECT 69.320 196.500 69.580 196.820 ;
        RECT 67.020 196.160 67.280 196.480 ;
        RECT 66.560 194.800 66.820 195.120 ;
        RECT 66.100 194.460 66.360 194.780 ;
        RECT 65.640 191.740 65.900 192.060 ;
        RECT 65.180 191.400 65.440 191.720 ;
        RECT 65.640 188.000 65.900 188.320 ;
        RECT 65.700 186.280 65.840 188.000 ;
        RECT 65.640 185.960 65.900 186.280 ;
        RECT 64.720 180.520 64.980 180.840 ;
        RECT 65.700 180.500 65.840 185.960 ;
        RECT 66.160 185.940 66.300 194.460 ;
        RECT 66.560 194.120 66.820 194.440 ;
        RECT 66.620 192.740 66.760 194.120 ;
        RECT 66.560 192.420 66.820 192.740 ;
        RECT 66.100 185.620 66.360 185.940 ;
        RECT 62.880 180.180 63.140 180.500 ;
        RECT 65.640 180.180 65.900 180.500 ;
        RECT 62.940 173.020 63.080 180.180 ;
        RECT 63.340 179.840 63.600 180.160 ;
        RECT 63.400 179.140 63.540 179.840 ;
        RECT 63.340 178.820 63.600 179.140 ;
        RECT 63.800 178.820 64.060 179.140 ;
        RECT 63.340 177.350 63.600 177.440 ;
        RECT 63.860 177.350 64.000 178.820 ;
        RECT 64.260 178.710 64.520 178.800 ;
        RECT 65.700 178.710 65.840 180.180 ;
        RECT 64.260 178.570 65.840 178.710 ;
        RECT 64.260 178.480 64.520 178.570 ;
        RECT 63.340 177.210 64.000 177.350 ;
        RECT 63.340 177.120 63.600 177.210 ;
        RECT 63.860 173.700 64.000 177.210 ;
        RECT 65.640 174.400 65.900 174.720 ;
        RECT 63.800 173.380 64.060 173.700 ;
        RECT 65.180 173.610 65.440 173.700 ;
        RECT 64.780 173.470 65.440 173.610 ;
        RECT 62.880 172.700 63.140 173.020 ;
        RECT 63.340 170.890 63.600 170.980 ;
        RECT 63.860 170.890 64.000 173.380 ;
        RECT 64.780 172.000 64.920 173.470 ;
        RECT 65.180 173.380 65.440 173.470 ;
        RECT 65.700 173.360 65.840 174.400 ;
        RECT 65.640 173.040 65.900 173.360 ;
        RECT 64.720 171.680 64.980 172.000 ;
        RECT 63.340 170.750 64.000 170.890 ;
        RECT 63.340 170.660 63.600 170.750 ;
        RECT 63.860 169.870 64.000 170.750 ;
        RECT 64.260 169.870 64.520 169.960 ;
        RECT 63.860 169.730 64.520 169.870 ;
        RECT 64.260 169.640 64.520 169.730 ;
        RECT 65.700 167.580 65.840 173.040 ;
        RECT 66.160 169.960 66.300 185.620 ;
        RECT 66.620 183.560 66.760 192.420 ;
        RECT 67.080 190.020 67.220 196.160 ;
        RECT 69.380 195.460 69.520 196.500 ;
        RECT 69.320 195.140 69.580 195.460 ;
        RECT 69.380 194.295 69.520 195.140 ;
        RECT 69.310 193.925 69.590 194.295 ;
        RECT 67.480 191.740 67.740 192.060 ;
        RECT 67.020 189.700 67.280 190.020 ;
        RECT 67.540 187.210 67.680 191.740 ;
        RECT 67.940 191.400 68.200 191.720 ;
        RECT 68.000 190.895 68.140 191.400 ;
        RECT 67.930 190.525 68.210 190.895 ;
        RECT 69.840 188.320 69.980 199.560 ;
        RECT 70.160 198.345 72.040 198.715 ;
        RECT 72.600 195.460 72.740 199.900 ;
        RECT 73.000 198.880 73.260 199.200 ;
        RECT 73.060 197.160 73.200 198.880 ;
        RECT 73.000 196.840 73.260 197.160 ;
        RECT 75.820 195.460 75.960 199.900 ;
        RECT 77.200 199.880 77.340 200.720 ;
        RECT 77.140 199.560 77.400 199.880 ;
        RECT 72.540 195.140 72.800 195.460 ;
        RECT 75.760 195.140 76.020 195.460 ;
        RECT 75.300 194.800 75.560 195.120 ;
        RECT 73.920 194.120 74.180 194.440 ;
        RECT 70.160 192.905 72.040 193.275 ;
        RECT 73.980 192.400 74.120 194.120 ;
        RECT 74.380 193.440 74.640 193.760 ;
        RECT 73.920 192.080 74.180 192.400 ;
        RECT 74.440 192.255 74.580 193.440 ;
        RECT 75.360 192.740 75.500 194.800 ;
        RECT 75.300 192.420 75.560 192.740 ;
        RECT 73.980 190.020 74.120 192.080 ;
        RECT 74.370 191.885 74.650 192.255 ;
        RECT 73.920 189.700 74.180 190.020 ;
        RECT 72.540 189.020 72.800 189.340 ;
        RECT 69.780 188.000 70.040 188.320 ;
        RECT 67.940 187.210 68.200 187.300 ;
        RECT 67.540 187.070 68.200 187.210 ;
        RECT 67.940 186.980 68.200 187.070 ;
        RECT 69.840 186.620 69.980 188.000 ;
        RECT 70.160 187.465 72.040 187.835 ;
        RECT 69.780 186.300 70.040 186.620 ;
        RECT 67.480 183.580 67.740 183.900 ;
        RECT 66.560 183.240 66.820 183.560 ;
        RECT 66.620 178.800 66.760 183.240 ;
        RECT 67.020 180.520 67.280 180.840 ;
        RECT 66.560 178.480 66.820 178.800 ;
        RECT 67.080 173.020 67.220 180.520 ;
        RECT 67.540 178.460 67.680 183.580 ;
        RECT 70.160 182.025 72.040 182.395 ;
        RECT 68.400 179.840 68.660 180.160 ;
        RECT 67.480 178.140 67.740 178.460 ;
        RECT 68.460 173.020 68.600 179.840 ;
        RECT 69.320 177.120 69.580 177.440 ;
        RECT 69.780 177.120 70.040 177.440 ;
        RECT 69.380 176.420 69.520 177.120 ;
        RECT 69.840 176.420 69.980 177.120 ;
        RECT 70.160 176.585 72.040 176.955 ;
        RECT 69.320 176.100 69.580 176.420 ;
        RECT 69.780 176.100 70.040 176.420 ;
        RECT 72.600 175.740 72.740 189.020 ;
        RECT 74.440 188.740 74.580 191.885 ;
        RECT 75.760 191.630 76.020 191.720 ;
        RECT 75.760 191.490 76.880 191.630 ;
        RECT 75.760 191.400 76.020 191.490 ;
        RECT 75.760 190.720 76.020 191.040 ;
        RECT 75.820 190.020 75.960 190.720 ;
        RECT 75.760 189.700 76.020 190.020 ;
        RECT 76.740 189.340 76.880 191.490 ;
        RECT 74.840 189.250 75.100 189.340 ;
        RECT 74.840 189.110 76.420 189.250 ;
        RECT 74.840 189.020 75.100 189.110 ;
        RECT 74.440 188.600 75.960 188.740 ;
        RECT 73.000 188.000 73.260 188.320 ;
        RECT 74.840 188.000 75.100 188.320 ;
        RECT 73.060 185.940 73.200 188.000 ;
        RECT 73.920 186.190 74.180 186.280 ;
        RECT 74.900 186.190 75.040 188.000 ;
        RECT 73.920 186.050 75.040 186.190 ;
        RECT 73.920 185.960 74.180 186.050 ;
        RECT 73.000 185.620 73.260 185.940 ;
        RECT 73.060 181.260 73.200 185.620 ;
        RECT 73.060 181.120 73.660 181.260 ;
        RECT 72.540 175.420 72.800 175.740 ;
        RECT 67.020 172.700 67.280 173.020 ;
        RECT 68.400 172.700 68.660 173.020 ;
        RECT 73.520 172.000 73.660 181.120 ;
        RECT 74.840 173.270 75.100 173.360 ;
        RECT 74.840 173.130 75.500 173.270 ;
        RECT 74.840 173.040 75.100 173.130 ;
        RECT 73.460 171.680 73.720 172.000 ;
        RECT 70.160 171.145 72.040 171.515 ;
        RECT 73.520 170.640 73.660 171.680 ;
        RECT 73.460 170.320 73.720 170.640 ;
        RECT 68.860 169.980 69.120 170.300 ;
        RECT 66.100 169.640 66.360 169.960 ;
        RECT 67.020 169.300 67.280 169.620 ;
        RECT 67.080 168.260 67.220 169.300 ;
        RECT 67.020 167.940 67.280 168.260 ;
        RECT 68.400 167.940 68.660 168.260 ;
        RECT 66.560 167.600 66.820 167.920 ;
        RECT 62.880 167.260 63.140 167.580 ;
        RECT 65.640 167.260 65.900 167.580 ;
        RECT 62.940 165.540 63.080 167.260 ;
        RECT 62.880 165.220 63.140 165.540 ;
        RECT 66.620 164.860 66.760 167.600 ;
        RECT 67.940 165.220 68.200 165.540 ;
        RECT 66.560 164.540 66.820 164.860 ;
        RECT 62.420 163.520 62.680 163.840 ;
        RECT 63.800 163.520 64.060 163.840 ;
        RECT 60.580 162.500 60.840 162.820 ;
        RECT 63.860 162.480 64.000 163.520 ;
        RECT 66.620 162.820 66.760 164.540 ;
        RECT 67.480 163.520 67.740 163.840 ;
        RECT 66.560 162.500 66.820 162.820 ;
        RECT 63.800 162.160 64.060 162.480 ;
        RECT 62.880 161.480 63.140 161.800 ;
        RECT 59.200 160.800 59.460 161.120 ;
        RECT 59.660 160.800 59.920 161.120 ;
        RECT 59.260 159.080 59.400 160.800 ;
        RECT 62.940 159.760 63.080 161.480 ;
        RECT 63.790 161.285 64.070 161.655 ;
        RECT 63.800 161.140 64.060 161.285 ;
        RECT 62.880 159.440 63.140 159.760 ;
        RECT 59.200 158.760 59.460 159.080 ;
        RECT 60.120 158.080 60.380 158.400 ;
        RECT 58.280 156.380 58.540 156.700 ;
        RECT 60.180 156.360 60.320 158.080 ;
        RECT 63.860 156.700 64.000 161.140 ;
        RECT 63.800 156.380 64.060 156.700 ;
        RECT 66.550 156.525 66.830 156.895 ;
        RECT 60.120 156.040 60.380 156.360 ;
        RECT 66.620 156.020 66.760 156.525 ;
        RECT 58.740 155.700 59.000 156.020 ;
        RECT 66.560 155.700 66.820 156.020 ;
        RECT 58.800 152.560 58.940 155.700 ;
        RECT 66.620 154.660 66.760 155.700 ;
        RECT 66.560 154.340 66.820 154.660 ;
        RECT 67.540 153.980 67.680 163.520 ;
        RECT 68.000 157.380 68.140 165.220 ;
        RECT 68.460 160.100 68.600 167.940 ;
        RECT 68.920 167.580 69.060 169.980 ;
        RECT 69.320 168.960 69.580 169.280 ;
        RECT 69.780 168.960 70.040 169.280 ;
        RECT 74.840 168.960 75.100 169.280 ;
        RECT 69.380 168.260 69.520 168.960 ;
        RECT 69.320 167.940 69.580 168.260 ;
        RECT 68.860 167.260 69.120 167.580 ;
        RECT 69.320 166.240 69.580 166.560 ;
        RECT 69.380 162.140 69.520 166.240 ;
        RECT 69.840 165.055 69.980 168.960 ;
        RECT 74.380 167.940 74.640 168.260 ;
        RECT 73.000 167.150 73.260 167.240 ;
        RECT 72.600 167.010 73.260 167.150 ;
        RECT 74.440 167.095 74.580 167.940 ;
        RECT 70.160 165.705 72.040 166.075 ;
        RECT 69.770 164.685 70.050 165.055 ;
        RECT 71.620 164.540 71.880 164.860 ;
        RECT 69.320 161.820 69.580 162.140 ;
        RECT 70.700 161.820 70.960 162.140 ;
        RECT 69.320 161.370 69.580 161.460 ;
        RECT 70.760 161.370 70.900 161.820 ;
        RECT 71.680 161.460 71.820 164.540 ;
        RECT 72.080 161.655 72.340 161.800 ;
        RECT 69.320 161.230 70.900 161.370 ;
        RECT 69.320 161.140 69.580 161.230 ;
        RECT 71.620 161.140 71.880 161.460 ;
        RECT 72.070 161.285 72.350 161.655 ;
        RECT 70.160 160.265 72.040 160.635 ;
        RECT 68.400 159.780 68.660 160.100 ;
        RECT 67.940 157.060 68.200 157.380 ;
        RECT 68.460 156.215 68.600 159.780 ;
        RECT 68.390 155.845 68.670 156.215 ;
        RECT 69.780 155.700 70.040 156.020 ;
        RECT 68.400 155.360 68.660 155.680 ;
        RECT 68.460 154.660 68.600 155.360 ;
        RECT 68.400 154.340 68.660 154.660 ;
        RECT 67.480 153.660 67.740 153.980 ;
        RECT 59.200 152.640 59.460 152.960 ;
        RECT 54.200 152.420 54.800 152.560 ;
        RECT 53.680 151.620 53.940 151.940 ;
        RECT 51.380 151.280 51.640 151.600 ;
        RECT 53.740 151.455 53.880 151.620 ;
        RECT 53.670 151.085 53.950 151.455 ;
        RECT 52.760 150.600 53.020 150.920 ;
        RECT 51.840 149.920 52.100 150.240 ;
        RECT 52.300 149.920 52.560 150.240 ;
        RECT 50.920 148.220 51.180 148.540 ;
        RECT 45.400 147.880 45.660 148.200 ;
        RECT 51.900 146.500 52.040 149.920 ;
        RECT 52.360 146.500 52.500 149.920 ;
        RECT 52.820 149.220 52.960 150.600 ;
        RECT 54.200 149.220 54.340 152.420 ;
        RECT 55.160 152.105 57.040 152.475 ;
        RECT 58.340 152.420 58.940 152.560 ;
        RECT 52.760 148.900 53.020 149.220 ;
        RECT 54.140 148.900 54.400 149.220 ;
        RECT 52.820 146.500 52.960 148.900 ;
        RECT 54.200 146.500 54.340 148.900 ;
        RECT 58.340 148.200 58.480 152.420 ;
        RECT 59.260 151.260 59.400 152.640 ;
        RECT 59.200 150.940 59.460 151.260 ;
        RECT 69.840 150.920 69.980 155.700 ;
        RECT 70.160 154.825 72.040 155.195 ;
        RECT 72.600 153.495 72.740 167.010 ;
        RECT 73.000 166.920 73.260 167.010 ;
        RECT 74.370 166.980 74.650 167.095 ;
        RECT 73.980 166.840 74.650 166.980 ;
        RECT 73.000 166.240 73.260 166.560 ;
        RECT 73.060 165.540 73.200 166.240 ;
        RECT 73.000 165.220 73.260 165.540 ;
        RECT 73.000 163.520 73.260 163.840 ;
        RECT 73.060 159.420 73.200 163.520 ;
        RECT 73.000 159.100 73.260 159.420 ;
        RECT 73.460 158.080 73.720 158.400 ;
        RECT 73.520 157.575 73.660 158.080 ;
        RECT 73.450 157.205 73.730 157.575 ;
        RECT 73.520 157.040 73.660 157.205 ;
        RECT 73.460 156.720 73.720 157.040 ;
        RECT 73.980 156.020 74.120 166.840 ;
        RECT 74.370 166.725 74.650 166.840 ;
        RECT 74.900 165.540 75.040 168.960 ;
        RECT 75.360 168.260 75.500 173.130 ;
        RECT 75.820 170.890 75.960 188.600 ;
        RECT 76.280 173.360 76.420 189.110 ;
        RECT 76.680 189.020 76.940 189.340 ;
        RECT 76.740 188.320 76.880 189.020 ;
        RECT 76.680 188.000 76.940 188.320 ;
        RECT 76.680 182.560 76.940 182.880 ;
        RECT 76.740 181.180 76.880 182.560 ;
        RECT 76.680 180.860 76.940 181.180 ;
        RECT 76.220 173.040 76.480 173.360 ;
        RECT 76.220 170.890 76.480 170.980 ;
        RECT 75.820 170.750 76.480 170.890 ;
        RECT 76.220 170.660 76.480 170.750 ;
        RECT 76.220 168.960 76.480 169.280 ;
        RECT 76.280 168.260 76.420 168.960 ;
        RECT 75.300 167.940 75.560 168.260 ;
        RECT 76.220 167.940 76.480 168.260 ;
        RECT 75.300 166.920 75.560 167.240 ;
        RECT 74.840 165.220 75.100 165.540 ;
        RECT 74.370 161.965 74.650 162.335 ;
        RECT 73.920 155.700 74.180 156.020 ;
        RECT 73.000 155.360 73.260 155.680 ;
        RECT 73.060 153.640 73.200 155.360 ;
        RECT 72.530 153.125 72.810 153.495 ;
        RECT 73.000 153.320 73.260 153.640 ;
        RECT 72.540 152.980 72.800 153.125 ;
        RECT 69.780 150.600 70.040 150.920 ;
        RECT 69.780 149.920 70.040 150.240 ;
        RECT 55.050 147.685 55.330 148.055 ;
        RECT 58.280 147.880 58.540 148.200 ;
        RECT 68.400 147.880 68.660 148.200 ;
        RECT 55.060 147.540 55.320 147.685 ;
        RECT 61.960 147.540 62.220 147.860 ;
        RECT 54.600 147.200 54.860 147.520 ;
        RECT 51.840 146.180 52.100 146.500 ;
        RECT 52.300 146.180 52.560 146.500 ;
        RECT 52.760 146.180 53.020 146.500 ;
        RECT 54.140 146.180 54.400 146.500 ;
        RECT 54.660 145.480 54.800 147.200 ;
        RECT 55.160 146.665 57.040 147.035 ;
        RECT 62.020 146.160 62.160 147.540 ;
        RECT 67.940 147.200 68.200 147.520 ;
        RECT 68.000 146.500 68.140 147.200 ;
        RECT 67.940 146.180 68.200 146.500 ;
        RECT 61.960 145.840 62.220 146.160 ;
        RECT 68.000 145.820 68.140 146.180 ;
        RECT 68.460 145.900 68.600 147.880 ;
        RECT 69.840 146.160 69.980 149.920 ;
        RECT 70.160 149.385 72.040 149.755 ;
        RECT 71.150 148.365 71.430 148.735 ;
        RECT 71.220 148.200 71.360 148.365 ;
        RECT 71.160 147.880 71.420 148.200 ;
        RECT 72.080 147.880 72.340 148.200 ;
        RECT 69.780 145.900 70.040 146.160 ;
        RECT 68.460 145.840 70.040 145.900 ;
        RECT 68.460 145.820 69.980 145.840 ;
        RECT 60.580 145.500 60.840 145.820 ;
        RECT 67.940 145.500 68.200 145.820 ;
        RECT 68.400 145.760 69.980 145.820 ;
        RECT 68.400 145.500 68.660 145.760 ;
        RECT 54.140 145.160 54.400 145.480 ;
        RECT 54.600 145.160 54.860 145.480 ;
        RECT 54.200 143.780 54.340 145.160 ;
        RECT 54.140 143.460 54.400 143.780 ;
        RECT 42.640 142.100 42.900 142.420 ;
        RECT 45.860 142.100 46.120 142.420 ;
        RECT 38.560 141.140 38.700 141.760 ;
        RECT 37.640 141.000 38.700 141.140 ;
        RECT 41.780 141.680 42.380 141.820 ;
        RECT 37.640 140.690 37.780 141.000 ;
        RECT 41.780 140.690 41.920 141.680 ;
        RECT 45.920 140.690 46.060 142.100 ;
        RECT 50.000 141.760 50.260 142.080 ;
        RECT 53.680 141.760 53.940 142.080 ;
        RECT 55.060 141.990 55.320 142.080 ;
        RECT 59.200 141.990 59.460 142.080 ;
        RECT 54.200 141.850 55.320 141.990 ;
        RECT 50.060 140.690 50.200 141.760 ;
        RECT 33.430 132.440 33.710 140.690 ;
        RECT 37.570 132.440 37.850 140.690 ;
        RECT 41.710 132.440 41.990 140.690 ;
        RECT 45.850 132.440 46.130 140.690 ;
        RECT 49.990 132.440 50.270 140.690 ;
        RECT 53.740 140.040 53.880 141.760 ;
        RECT 54.200 140.690 54.340 141.850 ;
        RECT 55.060 141.760 55.320 141.850 ;
        RECT 58.340 141.850 59.460 141.990 ;
        RECT 55.160 141.225 57.040 141.595 ;
        RECT 58.340 140.690 58.480 141.850 ;
        RECT 59.200 141.760 59.460 141.850 ;
        RECT 60.640 140.720 60.780 145.500 ;
        RECT 71.220 145.480 71.360 147.880 ;
        RECT 72.140 147.520 72.280 147.880 ;
        RECT 72.540 147.540 72.800 147.860 ;
        RECT 71.620 147.200 71.880 147.520 ;
        RECT 72.080 147.200 72.340 147.520 ;
        RECT 71.680 145.480 71.820 147.200 ;
        RECT 72.600 146.500 72.740 147.540 ;
        RECT 73.920 147.430 74.180 147.520 ;
        RECT 74.440 147.430 74.580 161.965 ;
        RECT 75.360 158.400 75.500 166.920 ;
        RECT 76.220 165.220 76.480 165.540 ;
        RECT 76.280 163.840 76.420 165.220 ;
        RECT 76.680 164.200 76.940 164.520 ;
        RECT 76.220 163.520 76.480 163.840 ;
        RECT 76.740 162.820 76.880 164.200 ;
        RECT 76.680 162.500 76.940 162.820 ;
        RECT 75.760 158.760 76.020 159.080 ;
        RECT 75.300 158.080 75.560 158.400 ;
        RECT 75.360 156.950 75.500 158.080 ;
        RECT 75.820 157.380 75.960 158.760 ;
        RECT 75.760 157.060 76.020 157.380 ;
        RECT 74.900 156.810 75.500 156.950 ;
        RECT 74.900 156.020 75.040 156.810 ;
        RECT 76.680 156.040 76.940 156.360 ;
        RECT 74.840 155.700 75.100 156.020 ;
        RECT 76.220 153.660 76.480 153.980 ;
        RECT 76.280 149.415 76.420 153.660 ;
        RECT 76.740 152.960 76.880 156.040 ;
        RECT 76.680 152.640 76.940 152.960 ;
        RECT 76.210 149.045 76.490 149.415 ;
        RECT 76.740 149.220 76.880 152.640 ;
        RECT 77.200 152.560 77.340 199.560 ;
        RECT 77.600 194.460 77.860 194.780 ;
        RECT 77.660 192.740 77.800 194.460 ;
        RECT 77.600 192.420 77.860 192.740 ;
        RECT 78.060 191.740 78.320 192.060 ;
        RECT 77.600 191.400 77.860 191.720 ;
        RECT 77.660 189.680 77.800 191.400 ;
        RECT 77.600 189.360 77.860 189.680 ;
        RECT 78.120 189.250 78.260 191.740 ;
        RECT 78.520 189.250 78.780 189.340 ;
        RECT 78.120 189.110 78.780 189.250 ;
        RECT 78.520 189.020 78.780 189.110 ;
        RECT 77.600 188.000 77.860 188.320 ;
        RECT 77.660 185.940 77.800 188.000 ;
        RECT 78.580 187.495 78.720 189.020 ;
        RECT 78.510 187.125 78.790 187.495 ;
        RECT 78.060 185.960 78.320 186.280 ;
        RECT 77.600 185.620 77.860 185.940 ;
        RECT 78.120 184.580 78.260 185.960 ;
        RECT 79.040 184.580 79.180 207.720 ;
        RECT 79.900 205.000 80.160 205.320 ;
        RECT 79.960 199.540 80.100 205.000 ;
        RECT 80.880 203.135 81.020 212.820 ;
        RECT 81.280 205.000 81.540 205.320 ;
        RECT 80.810 202.765 81.090 203.135 ;
        RECT 80.820 201.600 81.080 201.920 ;
        RECT 79.900 199.220 80.160 199.540 ;
        RECT 80.360 198.880 80.620 199.200 ;
        RECT 80.420 194.780 80.560 198.880 ;
        RECT 79.440 194.460 79.700 194.780 ;
        RECT 80.360 194.460 80.620 194.780 ;
        RECT 79.500 193.760 79.640 194.460 ;
        RECT 79.440 193.440 79.700 193.760 ;
        RECT 79.500 191.380 79.640 193.440 ;
        RECT 80.880 192.740 81.020 201.600 ;
        RECT 80.820 192.420 81.080 192.740 ;
        RECT 79.440 191.060 79.700 191.380 ;
        RECT 80.360 191.060 80.620 191.380 ;
        RECT 79.500 188.660 79.640 191.060 ;
        RECT 80.420 190.895 80.560 191.060 ;
        RECT 80.350 190.525 80.630 190.895 ;
        RECT 79.900 188.680 80.160 189.000 ;
        RECT 79.440 188.340 79.700 188.660 ;
        RECT 78.060 184.260 78.320 184.580 ;
        RECT 78.980 184.260 79.240 184.580 ;
        RECT 79.960 182.880 80.100 188.680 ;
        RECT 80.360 183.580 80.620 183.900 ;
        RECT 79.900 182.560 80.160 182.880 ;
        RECT 78.980 180.520 79.240 180.840 ;
        RECT 79.040 178.655 79.180 180.520 ;
        RECT 79.900 180.410 80.160 180.500 ;
        RECT 80.420 180.410 80.560 183.580 ;
        RECT 79.900 180.270 80.560 180.410 ;
        RECT 80.810 180.325 81.090 180.695 ;
        RECT 79.900 180.180 80.160 180.270 ;
        RECT 78.970 178.285 79.250 178.655 ;
        RECT 79.960 178.460 80.100 180.180 ;
        RECT 79.900 178.140 80.160 178.460 ;
        RECT 77.600 177.800 77.860 178.120 ;
        RECT 77.660 159.420 77.800 177.800 ;
        RECT 80.880 177.180 81.020 180.325 ;
        RECT 80.420 177.040 81.020 177.180 ;
        RECT 78.520 173.040 78.780 173.360 ;
        RECT 78.580 170.640 78.720 173.040 ;
        RECT 80.420 172.680 80.560 177.040 ;
        RECT 81.340 176.330 81.480 205.000 ;
        RECT 81.800 202.455 81.940 212.820 ;
        RECT 83.580 210.100 83.840 210.420 ;
        RECT 83.640 209.060 83.780 210.100 ;
        RECT 83.580 208.740 83.840 209.060 ;
        RECT 84.100 208.460 84.240 213.160 ;
        RECT 93.240 212.820 93.500 213.140 ;
        RECT 92.780 212.480 93.040 212.800 ;
        RECT 85.160 211.945 87.040 212.315 ;
        RECT 86.800 211.460 87.060 211.780 ;
        RECT 84.500 210.780 84.760 211.100 ;
        RECT 83.640 208.320 84.240 208.460 ;
        RECT 83.120 207.040 83.380 207.360 ;
        RECT 83.180 204.640 83.320 207.040 ;
        RECT 83.120 204.320 83.380 204.640 ;
        RECT 81.730 202.085 82.010 202.455 ;
        RECT 82.660 202.280 82.920 202.600 ;
        RECT 81.800 186.280 81.940 202.085 ;
        RECT 82.200 199.560 82.460 199.880 ;
        RECT 82.260 199.055 82.400 199.560 ;
        RECT 82.190 198.685 82.470 199.055 ;
        RECT 82.260 188.320 82.400 198.685 ;
        RECT 82.200 188.000 82.460 188.320 ;
        RECT 81.740 185.960 82.000 186.280 ;
        RECT 82.200 185.280 82.460 185.600 ;
        RECT 81.740 183.920 82.000 184.240 ;
        RECT 81.800 181.180 81.940 183.920 ;
        RECT 82.260 183.220 82.400 185.280 ;
        RECT 82.200 182.900 82.460 183.220 ;
        RECT 82.720 182.735 82.860 202.280 ;
        RECT 83.180 195.120 83.320 204.320 ;
        RECT 83.640 203.620 83.780 208.320 ;
        RECT 84.560 206.000 84.700 210.780 ;
        RECT 85.880 208.400 86.140 208.720 ;
        RECT 85.940 207.895 86.080 208.400 ;
        RECT 85.870 207.525 86.150 207.895 ;
        RECT 86.860 207.270 87.000 211.460 ;
        RECT 87.260 209.760 87.520 210.080 ;
        RECT 87.720 209.760 87.980 210.080 ;
        RECT 90.020 209.760 90.280 210.080 ;
        RECT 87.320 208.040 87.460 209.760 ;
        RECT 87.780 209.060 87.920 209.760 ;
        RECT 90.080 209.060 90.220 209.760 ;
        RECT 87.720 208.740 87.980 209.060 ;
        RECT 90.020 208.740 90.280 209.060 ;
        RECT 92.840 208.720 92.980 212.480 ;
        RECT 89.100 208.400 89.360 208.720 ;
        RECT 92.780 208.400 93.040 208.720 ;
        RECT 87.260 207.720 87.520 208.040 ;
        RECT 86.860 207.130 87.460 207.270 ;
        RECT 85.160 206.505 87.040 206.875 ;
        RECT 84.500 205.680 84.760 206.000 ;
        RECT 87.320 205.660 87.460 207.130 ;
        RECT 88.180 207.040 88.440 207.360 ;
        RECT 87.260 205.340 87.520 205.660 ;
        RECT 86.800 204.320 87.060 204.640 ;
        RECT 87.720 204.320 87.980 204.640 ;
        RECT 83.580 203.300 83.840 203.620 ;
        RECT 83.120 194.800 83.380 195.120 ;
        RECT 83.180 192.060 83.320 194.800 ;
        RECT 83.120 191.740 83.380 192.060 ;
        RECT 83.180 189.340 83.320 191.740 ;
        RECT 83.120 189.020 83.380 189.340 ;
        RECT 83.120 188.000 83.380 188.320 ;
        RECT 82.650 182.365 82.930 182.735 ;
        RECT 83.180 181.940 83.320 188.000 ;
        RECT 82.260 181.800 83.320 181.940 ;
        RECT 81.740 180.860 82.000 181.180 ;
        RECT 80.880 176.190 81.480 176.330 ;
        RECT 80.360 172.590 80.620 172.680 ;
        RECT 79.960 172.450 80.620 172.590 ;
        RECT 78.520 170.320 78.780 170.640 ;
        RECT 79.960 167.580 80.100 172.450 ;
        RECT 80.360 172.360 80.620 172.450 ;
        RECT 80.360 171.680 80.620 172.000 ;
        RECT 78.520 167.260 78.780 167.580 ;
        RECT 79.900 167.260 80.160 167.580 ;
        RECT 78.580 166.560 78.720 167.260 ;
        RECT 79.440 166.920 79.700 167.240 ;
        RECT 78.520 166.240 78.780 166.560 ;
        RECT 79.500 164.520 79.640 166.920 ;
        RECT 79.960 165.540 80.100 167.260 ;
        RECT 79.900 165.220 80.160 165.540 ;
        RECT 80.420 164.520 80.560 171.680 ;
        RECT 79.440 164.200 79.700 164.520 ;
        RECT 80.360 164.200 80.620 164.520 ;
        RECT 78.520 163.520 78.780 163.840 ;
        RECT 78.580 159.420 78.720 163.520 ;
        RECT 80.420 162.820 80.560 164.200 ;
        RECT 80.360 162.500 80.620 162.820 ;
        RECT 77.600 159.100 77.860 159.420 ;
        RECT 78.520 159.100 78.780 159.420 ;
        RECT 79.900 159.100 80.160 159.420 ;
        RECT 77.660 157.380 77.800 159.100 ;
        RECT 78.520 158.420 78.780 158.740 ;
        RECT 77.600 157.060 77.860 157.380 ;
        RECT 78.580 156.360 78.720 158.420 ;
        RECT 78.970 157.205 79.250 157.575 ;
        RECT 78.520 156.040 78.780 156.360 ;
        RECT 78.580 154.320 78.720 156.040 ;
        RECT 79.040 156.020 79.180 157.205 ;
        RECT 79.960 156.700 80.100 159.100 ;
        RECT 80.880 157.380 81.020 176.190 ;
        RECT 81.270 175.565 81.550 175.935 ;
        RECT 81.340 173.020 81.480 175.565 ;
        RECT 81.280 172.700 81.540 173.020 ;
        RECT 81.730 172.165 82.010 172.535 ;
        RECT 81.270 169.445 81.550 169.815 ;
        RECT 81.340 167.580 81.480 169.445 ;
        RECT 81.800 168.260 81.940 172.165 ;
        RECT 81.740 167.940 82.000 168.260 ;
        RECT 81.280 167.260 81.540 167.580 ;
        RECT 81.280 159.100 81.540 159.420 ;
        RECT 81.340 158.255 81.480 159.100 ;
        RECT 81.270 157.885 81.550 158.255 ;
        RECT 80.820 157.060 81.080 157.380 ;
        RECT 82.260 156.780 82.400 181.800 ;
        RECT 82.650 181.005 82.930 181.375 ;
        RECT 83.120 181.200 83.380 181.520 ;
        RECT 82.720 159.420 82.860 181.005 ;
        RECT 83.180 175.400 83.320 181.200 ;
        RECT 83.120 175.080 83.380 175.400 ;
        RECT 83.120 173.380 83.380 173.700 ;
        RECT 83.180 164.180 83.320 173.380 ;
        RECT 83.640 165.735 83.780 203.300 ;
        RECT 84.040 202.960 84.300 203.280 ;
        RECT 84.100 200.415 84.240 202.960 ;
        RECT 86.860 202.940 87.000 204.320 ;
        RECT 87.780 202.940 87.920 204.320 ;
        RECT 86.800 202.620 87.060 202.940 ;
        RECT 87.720 202.620 87.980 202.940 ;
        RECT 84.500 201.600 84.760 201.920 ;
        RECT 84.030 200.045 84.310 200.415 ;
        RECT 84.560 200.220 84.700 201.600 ;
        RECT 85.160 201.065 87.040 201.435 ;
        RECT 87.720 200.470 87.980 200.560 ;
        RECT 88.240 200.470 88.380 207.040 ;
        RECT 89.160 205.660 89.300 208.400 ;
        RECT 90.480 207.950 90.740 208.040 ;
        RECT 91.400 207.950 91.660 208.040 ;
        RECT 90.480 207.810 91.660 207.950 ;
        RECT 90.480 207.720 90.740 207.810 ;
        RECT 91.400 207.720 91.660 207.810 ;
        RECT 89.100 205.340 89.360 205.660 ;
        RECT 92.320 205.175 92.580 205.320 ;
        RECT 89.100 204.660 89.360 204.980 ;
        RECT 90.940 204.660 91.200 204.980 ;
        RECT 92.310 204.805 92.590 205.175 ;
        RECT 89.160 202.455 89.300 204.660 ;
        RECT 91.000 202.600 91.140 204.660 ;
        RECT 92.780 202.620 93.040 202.940 ;
        RECT 89.090 202.085 89.370 202.455 ;
        RECT 90.020 202.280 90.280 202.600 ;
        RECT 90.940 202.280 91.200 202.600 ;
        RECT 91.400 202.280 91.660 202.600 ;
        RECT 91.860 202.280 92.120 202.600 ;
        RECT 89.560 201.940 89.820 202.260 ;
        RECT 89.090 201.405 89.370 201.775 ;
        RECT 87.720 200.330 88.380 200.470 ;
        RECT 87.720 200.240 87.980 200.330 ;
        RECT 84.500 199.900 84.760 200.220 ;
        RECT 84.040 199.560 84.300 199.880 ;
        RECT 84.100 167.580 84.240 199.560 ;
        RECT 86.330 199.365 86.610 199.735 ;
        RECT 86.800 199.560 87.060 199.880 ;
        RECT 86.400 199.200 86.540 199.365 ;
        RECT 86.340 198.880 86.600 199.200 ;
        RECT 86.860 197.840 87.000 199.560 ;
        RECT 87.720 199.220 87.980 199.540 ;
        RECT 87.260 198.880 87.520 199.200 ;
        RECT 86.800 197.520 87.060 197.840 ;
        RECT 87.320 197.410 87.460 198.880 ;
        RECT 87.780 198.180 87.920 199.220 ;
        RECT 87.720 197.860 87.980 198.180 ;
        RECT 89.160 198.090 89.300 201.405 ;
        RECT 89.620 199.200 89.760 201.940 ;
        RECT 89.560 198.880 89.820 199.200 ;
        RECT 88.240 197.950 89.300 198.090 ;
        RECT 88.240 197.500 88.380 197.950 ;
        RECT 87.720 197.410 87.980 197.500 ;
        RECT 87.320 197.270 87.980 197.410 ;
        RECT 87.720 197.180 87.980 197.270 ;
        RECT 88.180 197.180 88.440 197.500 ;
        RECT 84.500 196.500 84.760 196.820 ;
        RECT 84.560 195.460 84.700 196.500 ;
        RECT 85.160 195.625 87.040 195.995 ;
        RECT 84.500 195.140 84.760 195.460 ;
        RECT 87.720 194.460 87.980 194.780 ;
        RECT 87.780 192.740 87.920 194.460 ;
        RECT 87.720 192.420 87.980 192.740 ;
        RECT 85.160 190.185 87.040 190.555 ;
        RECT 88.240 189.930 88.380 197.180 ;
        RECT 88.640 197.070 88.900 197.160 ;
        RECT 88.640 196.930 89.300 197.070 ;
        RECT 88.640 196.840 88.900 196.930 ;
        RECT 89.160 196.220 89.300 196.930 ;
        RECT 88.700 196.080 89.300 196.220 ;
        RECT 88.700 195.460 88.840 196.080 ;
        RECT 88.640 195.140 88.900 195.460 ;
        RECT 89.090 195.285 89.370 195.655 ;
        RECT 89.160 194.440 89.300 195.285 ;
        RECT 89.560 195.140 89.820 195.460 ;
        RECT 89.100 194.120 89.360 194.440 ;
        RECT 89.620 194.100 89.760 195.140 ;
        RECT 88.640 193.780 88.900 194.100 ;
        RECT 89.560 193.780 89.820 194.100 ;
        RECT 88.700 192.400 88.840 193.780 ;
        RECT 90.080 192.740 90.220 202.280 ;
        RECT 91.460 200.900 91.600 202.280 ;
        RECT 91.400 200.580 91.660 200.900 ;
        RECT 90.930 200.045 91.210 200.415 ;
        RECT 91.000 199.880 91.140 200.045 ;
        RECT 90.940 199.560 91.200 199.880 ;
        RECT 90.480 199.220 90.740 199.540 ;
        RECT 90.540 197.500 90.680 199.220 ;
        RECT 91.000 197.840 91.140 199.560 ;
        RECT 91.390 198.940 91.670 199.055 ;
        RECT 91.920 198.940 92.060 202.280 ;
        RECT 91.390 198.800 92.060 198.940 ;
        RECT 91.390 198.685 91.670 198.800 ;
        RECT 90.940 197.520 91.200 197.840 ;
        RECT 90.480 197.180 90.740 197.500 ;
        RECT 90.540 194.010 90.680 197.180 ;
        RECT 91.860 196.840 92.120 197.160 ;
        RECT 91.400 194.010 91.660 194.100 ;
        RECT 90.540 193.870 91.660 194.010 ;
        RECT 91.400 193.780 91.660 193.870 ;
        RECT 90.020 192.420 90.280 192.740 ;
        RECT 88.640 192.080 88.900 192.400 ;
        RECT 88.700 190.020 88.840 192.080 ;
        RECT 89.100 191.400 89.360 191.720 ;
        RECT 90.480 191.630 90.740 191.720 ;
        RECT 90.480 191.490 91.140 191.630 ;
        RECT 90.480 191.400 90.740 191.490 ;
        RECT 86.860 189.790 88.380 189.930 ;
        RECT 84.500 185.960 84.760 186.280 ;
        RECT 86.860 186.135 87.000 189.790 ;
        RECT 88.640 189.700 88.900 190.020 ;
        RECT 88.180 189.020 88.440 189.340 ;
        RECT 87.720 188.000 87.980 188.320 ;
        RECT 84.560 184.490 84.700 185.960 ;
        RECT 86.790 185.765 87.070 186.135 ;
        RECT 87.260 185.620 87.520 185.940 ;
        RECT 85.160 184.745 87.040 185.115 ;
        RECT 87.320 184.580 87.460 185.620 ;
        RECT 84.960 184.490 85.220 184.580 ;
        RECT 84.560 184.350 85.220 184.490 ;
        RECT 84.960 184.260 85.220 184.350 ;
        RECT 87.260 184.260 87.520 184.580 ;
        RECT 84.490 183.045 84.770 183.415 ;
        RECT 84.500 182.900 84.760 183.045 ;
        RECT 85.020 180.070 85.160 184.260 ;
        RECT 87.780 181.860 87.920 188.000 ;
        RECT 88.240 185.600 88.380 189.020 ;
        RECT 88.640 188.680 88.900 189.000 ;
        RECT 88.180 185.280 88.440 185.600 ;
        RECT 88.240 183.900 88.380 185.280 ;
        RECT 88.180 183.580 88.440 183.900 ;
        RECT 87.720 181.540 87.980 181.860 ;
        RECT 84.560 179.930 85.160 180.070 ;
        RECT 84.560 178.460 84.700 179.930 ;
        RECT 85.160 179.305 87.040 179.675 ;
        RECT 84.500 178.140 84.760 178.460 ;
        RECT 84.490 176.245 84.770 176.615 ;
        RECT 84.560 175.060 84.700 176.245 ;
        RECT 87.720 175.760 87.980 176.080 ;
        RECT 86.800 175.310 87.060 175.400 ;
        RECT 86.800 175.170 87.460 175.310 ;
        RECT 86.800 175.080 87.060 175.170 ;
        RECT 84.500 174.740 84.760 175.060 ;
        RECT 84.560 173.700 84.700 174.740 ;
        RECT 85.160 173.865 87.040 174.235 ;
        RECT 84.500 173.380 84.760 173.700 ;
        RECT 86.800 173.270 87.060 173.360 ;
        RECT 87.320 173.270 87.460 175.170 ;
        RECT 86.800 173.130 87.460 173.270 ;
        RECT 86.800 173.040 87.060 173.130 ;
        RECT 87.780 172.340 87.920 175.760 ;
        RECT 88.240 175.400 88.380 183.580 ;
        RECT 88.700 181.520 88.840 188.680 ;
        RECT 88.640 181.200 88.900 181.520 ;
        RECT 88.640 180.180 88.900 180.500 ;
        RECT 88.700 175.400 88.840 180.180 ;
        RECT 89.160 178.460 89.300 191.400 ;
        RECT 90.020 190.720 90.280 191.040 ;
        RECT 90.480 190.720 90.740 191.040 ;
        RECT 90.080 189.340 90.220 190.720 ;
        RECT 90.540 190.020 90.680 190.720 ;
        RECT 90.480 189.700 90.740 190.020 ;
        RECT 89.560 189.020 89.820 189.340 ;
        RECT 90.020 189.020 90.280 189.340 ;
        RECT 89.620 183.900 89.760 189.020 ;
        RECT 90.020 185.280 90.280 185.600 ;
        RECT 89.560 183.580 89.820 183.900 ;
        RECT 90.080 180.840 90.220 185.280 ;
        RECT 90.480 182.560 90.740 182.880 ;
        RECT 90.020 180.520 90.280 180.840 ;
        RECT 89.100 178.140 89.360 178.460 ;
        RECT 89.560 178.140 89.820 178.460 ;
        RECT 89.100 177.460 89.360 177.780 ;
        RECT 89.160 175.400 89.300 177.460 ;
        RECT 89.620 175.400 89.760 178.140 ;
        RECT 88.180 175.080 88.440 175.400 ;
        RECT 88.640 175.080 88.900 175.400 ;
        RECT 89.100 175.080 89.360 175.400 ;
        RECT 89.560 175.080 89.820 175.400 ;
        RECT 87.720 172.020 87.980 172.340 ;
        RECT 85.870 171.485 86.150 171.855 ;
        RECT 86.340 171.680 86.600 172.000 ;
        RECT 87.260 171.680 87.520 172.000 ;
        RECT 85.940 170.980 86.080 171.485 ;
        RECT 86.400 170.980 86.540 171.680 ;
        RECT 85.880 170.660 86.140 170.980 ;
        RECT 86.340 170.660 86.600 170.980 ;
        RECT 86.400 169.960 86.540 170.660 ;
        RECT 86.340 169.640 86.600 169.960 ;
        RECT 84.500 168.960 84.760 169.280 ;
        RECT 84.040 167.260 84.300 167.580 ;
        RECT 83.570 165.365 83.850 165.735 ;
        RECT 83.120 163.860 83.380 164.180 ;
        RECT 84.560 159.500 84.700 168.960 ;
        RECT 85.160 168.425 87.040 168.795 ;
        RECT 87.320 166.980 87.460 171.680 ;
        RECT 87.710 170.125 87.990 170.495 ;
        RECT 87.720 169.980 87.980 170.125 ;
        RECT 87.710 168.765 87.990 169.135 ;
        RECT 87.780 167.580 87.920 168.765 ;
        RECT 88.240 167.580 88.380 175.080 ;
        RECT 89.100 173.610 89.360 173.700 ;
        RECT 89.620 173.610 89.760 175.080 ;
        RECT 90.080 174.720 90.220 180.520 ;
        RECT 90.020 174.400 90.280 174.720 ;
        RECT 89.100 173.470 89.760 173.610 ;
        RECT 89.100 173.380 89.360 173.470 ;
        RECT 90.020 173.380 90.280 173.700 ;
        RECT 88.640 172.700 88.900 173.020 ;
        RECT 87.720 167.260 87.980 167.580 ;
        RECT 88.180 167.260 88.440 167.580 ;
        RECT 87.320 166.840 88.380 166.980 ;
        RECT 87.260 166.240 87.520 166.560 ;
        RECT 85.160 162.985 87.040 163.355 ;
        RECT 87.320 162.140 87.460 166.240 ;
        RECT 87.260 161.820 87.520 162.140 ;
        RECT 85.880 161.655 86.140 161.800 ;
        RECT 85.870 161.285 86.150 161.655 ;
        RECT 82.660 159.100 82.920 159.420 ;
        RECT 84.100 159.360 84.700 159.500 ;
        RECT 83.570 157.205 83.850 157.575 ;
        RECT 83.580 157.060 83.840 157.205 ;
        RECT 79.900 156.380 80.160 156.700 ;
        RECT 81.340 156.640 82.400 156.780 ;
        RECT 78.980 155.700 79.240 156.020 ;
        RECT 78.520 154.230 78.780 154.320 ;
        RECT 78.120 154.090 78.780 154.230 ;
        RECT 77.200 152.420 77.800 152.560 ;
        RECT 77.140 150.095 77.400 150.240 ;
        RECT 77.130 149.725 77.410 150.095 ;
        RECT 76.680 148.900 76.940 149.220 ;
        RECT 74.840 147.880 75.100 148.200 ;
        RECT 73.920 147.290 74.580 147.430 ;
        RECT 73.920 147.200 74.180 147.290 ;
        RECT 72.540 146.180 72.800 146.500 ;
        RECT 71.160 145.160 71.420 145.480 ;
        RECT 71.620 145.160 71.880 145.480 ;
        RECT 74.380 144.820 74.640 145.140 ;
        RECT 70.160 143.945 72.040 144.315 ;
        RECT 74.440 143.440 74.580 144.820 ;
        RECT 74.900 144.800 75.040 147.880 ;
        RECT 75.300 147.540 75.560 147.860 ;
        RECT 75.360 145.820 75.500 147.540 ;
        RECT 77.140 147.200 77.400 147.520 ;
        RECT 75.300 145.500 75.560 145.820 ;
        RECT 76.210 145.645 76.490 146.015 ;
        RECT 76.220 145.500 76.480 145.645 ;
        RECT 77.200 144.800 77.340 147.200 ;
        RECT 74.840 144.480 75.100 144.800 ;
        RECT 75.300 144.480 75.560 144.800 ;
        RECT 77.140 144.480 77.400 144.800 ;
        RECT 75.360 143.440 75.500 144.480 ;
        RECT 74.380 143.120 74.640 143.440 ;
        RECT 75.300 143.120 75.560 143.440 ;
        RECT 77.660 142.760 77.800 152.420 ;
        RECT 78.120 151.940 78.260 154.090 ;
        RECT 78.520 154.000 78.780 154.090 ;
        RECT 79.040 153.980 79.180 155.700 ;
        RECT 80.820 155.360 81.080 155.680 ;
        RECT 81.340 155.535 81.480 156.640 ;
        RECT 84.100 156.270 84.240 159.360 ;
        RECT 85.160 157.545 87.040 157.915 ;
        RECT 86.340 157.060 86.600 157.380 ;
        RECT 85.420 156.720 85.680 157.040 ;
        RECT 84.100 156.130 85.160 156.270 ;
        RECT 82.200 155.700 82.460 156.020 ;
        RECT 80.880 154.855 81.020 155.360 ;
        RECT 81.270 155.165 81.550 155.535 ;
        RECT 80.810 154.485 81.090 154.855 ;
        RECT 82.260 154.320 82.400 155.700 ;
        RECT 83.110 154.740 83.390 154.855 ;
        RECT 85.020 154.740 85.160 156.130 ;
        RECT 85.480 154.855 85.620 156.720 ;
        RECT 86.400 156.700 86.540 157.060 ;
        RECT 86.340 156.380 86.600 156.700 ;
        RECT 85.880 156.040 86.140 156.360 ;
        RECT 83.110 154.600 83.780 154.740 ;
        RECT 83.110 154.485 83.390 154.600 ;
        RECT 80.820 154.060 81.080 154.320 ;
        RECT 81.730 154.060 82.010 154.175 ;
        RECT 80.820 154.000 82.010 154.060 ;
        RECT 82.200 154.000 82.460 154.320 ;
        RECT 83.640 154.060 83.780 154.600 ;
        RECT 78.980 153.660 79.240 153.980 ;
        RECT 80.880 153.920 82.010 154.000 ;
        RECT 81.730 153.805 82.010 153.920 ;
        RECT 82.260 153.640 82.400 154.000 ;
        RECT 83.180 153.920 83.780 154.060 ;
        RECT 84.100 154.600 85.160 154.740 ;
        RECT 81.740 153.550 82.000 153.640 ;
        RECT 81.340 153.410 82.000 153.550 ;
        RECT 78.520 152.640 78.780 152.960 ;
        RECT 79.890 152.700 80.170 152.815 ;
        RECT 81.340 152.700 81.480 153.410 ;
        RECT 81.740 153.320 82.000 153.410 ;
        RECT 82.200 153.380 82.460 153.640 ;
        RECT 82.200 153.320 82.860 153.380 ;
        RECT 82.260 153.240 82.860 153.320 ;
        RECT 82.200 152.815 82.460 152.960 ;
        RECT 78.060 151.620 78.320 151.940 ;
        RECT 78.580 151.510 78.720 152.640 ;
        RECT 79.890 152.560 81.480 152.700 ;
        RECT 79.890 152.445 80.170 152.560 ;
        RECT 82.190 152.445 82.470 152.815 ;
        RECT 80.810 151.765 81.090 152.135 ;
        RECT 82.190 151.765 82.470 152.135 ;
        RECT 79.440 151.510 79.700 151.600 ;
        RECT 78.580 151.370 79.700 151.510 ;
        RECT 79.440 151.280 79.700 151.370 ;
        RECT 80.880 150.920 81.020 151.765 ;
        RECT 82.260 151.260 82.400 151.765 ;
        RECT 82.720 151.600 82.860 153.240 ;
        RECT 83.180 151.940 83.320 153.920 ;
        RECT 83.580 153.320 83.840 153.640 ;
        RECT 83.640 152.135 83.780 153.320 ;
        RECT 83.120 151.620 83.380 151.940 ;
        RECT 83.570 151.765 83.850 152.135 ;
        RECT 82.660 151.280 82.920 151.600 ;
        RECT 83.580 151.280 83.840 151.600 ;
        RECT 82.200 150.940 82.460 151.260 ;
        RECT 78.520 150.260 78.780 150.580 ;
        RECT 80.350 150.405 80.630 150.775 ;
        RECT 80.820 150.600 81.080 150.920 ;
        RECT 78.580 146.500 78.720 150.260 ;
        RECT 78.980 148.900 79.240 149.220 ;
        RECT 79.040 148.735 79.180 148.900 ;
        RECT 78.970 148.365 79.250 148.735 ;
        RECT 78.520 146.180 78.780 146.500 ;
        RECT 80.420 145.820 80.560 150.405 ;
        RECT 82.200 150.260 82.460 150.580 ;
        RECT 80.810 147.005 81.090 147.375 ;
        RECT 80.880 145.820 81.020 147.005 ;
        RECT 80.360 145.500 80.620 145.820 ;
        RECT 80.820 145.500 81.080 145.820 ;
        RECT 64.260 142.440 64.520 142.760 ;
        RECT 77.600 142.440 77.860 142.760 ;
        RECT 63.340 141.990 63.600 142.080 ;
        RECT 62.480 141.850 63.600 141.990 ;
        RECT 53.680 139.720 53.940 140.040 ;
        RECT 54.130 132.440 54.410 140.690 ;
        RECT 58.270 132.440 58.550 140.690 ;
        RECT 60.580 140.400 60.840 140.720 ;
        RECT 62.480 140.690 62.620 141.850 ;
        RECT 63.340 141.760 63.600 141.850 ;
        RECT 33.400 132.160 33.740 132.440 ;
        RECT 37.540 132.160 37.880 132.440 ;
        RECT 41.680 132.160 42.020 132.440 ;
        RECT 45.820 132.160 46.160 132.440 ;
        RECT 49.960 132.160 50.300 132.440 ;
        RECT 54.100 132.160 54.440 132.440 ;
        RECT 58.240 132.160 58.580 132.440 ;
        RECT 60.580 132.300 61.580 134.445 ;
        RECT 62.410 132.440 62.690 140.690 ;
        RECT 64.320 140.380 64.460 142.440 ;
        RECT 75.760 141.990 76.020 142.080 ;
        RECT 74.900 141.850 76.020 141.990 ;
        RECT 74.900 140.690 75.040 141.850 ;
        RECT 75.760 141.760 76.020 141.850 ;
        RECT 78.980 141.760 79.240 142.080 ;
        RECT 79.040 140.690 79.180 141.760 ;
        RECT 64.260 140.060 64.520 140.380 ;
        RECT 60.550 131.300 61.610 132.300 ;
        RECT 62.380 132.160 62.720 132.440 ;
        RECT 64.930 132.300 65.930 134.445 ;
        RECT 74.830 132.440 75.110 140.690 ;
        RECT 78.970 132.440 79.250 140.690 ;
        RECT 80.880 139.700 81.020 145.500 ;
        RECT 82.260 145.480 82.400 150.260 ;
        RECT 83.640 149.220 83.780 151.280 ;
        RECT 83.580 148.900 83.840 149.220 ;
        RECT 82.660 148.220 82.920 148.540 ;
        RECT 82.720 146.500 82.860 148.220 ;
        RECT 82.660 146.180 82.920 146.500 ;
        RECT 84.100 145.820 84.240 154.600 ;
        RECT 85.410 154.485 85.690 154.855 ;
        RECT 85.940 154.320 86.080 156.040 ;
        RECT 86.340 155.360 86.600 155.680 ;
        RECT 85.880 154.000 86.140 154.320 ;
        RECT 84.500 153.320 84.760 153.640 ;
        RECT 84.560 151.940 84.700 153.320 ;
        RECT 86.400 153.300 86.540 155.360 ;
        RECT 86.340 152.980 86.600 153.300 ;
        RECT 85.160 152.105 87.040 152.475 ;
        RECT 87.320 151.940 87.460 161.820 ;
        RECT 87.720 158.420 87.980 158.740 ;
        RECT 87.780 156.700 87.920 158.420 ;
        RECT 87.720 156.380 87.980 156.700 ;
        RECT 84.500 151.620 84.760 151.940 ;
        RECT 87.260 151.620 87.520 151.940 ;
        RECT 84.560 148.540 84.700 151.620 ;
        RECT 84.960 150.600 85.220 150.920 ;
        RECT 85.020 148.540 85.160 150.600 ;
        RECT 87.260 150.260 87.520 150.580 ;
        RECT 84.500 148.220 84.760 148.540 ;
        RECT 84.960 148.220 85.220 148.540 ;
        RECT 87.320 148.200 87.460 150.260 ;
        RECT 87.710 148.365 87.990 148.735 ;
        RECT 84.560 147.800 85.160 147.940 ;
        RECT 87.260 147.880 87.520 148.200 ;
        RECT 84.040 145.500 84.300 145.820 ;
        RECT 82.200 145.160 82.460 145.480 ;
        RECT 82.200 144.480 82.460 144.800 ;
        RECT 82.260 143.780 82.400 144.480 ;
        RECT 82.200 143.460 82.460 143.780 ;
        RECT 82.190 142.925 82.470 143.295 ;
        RECT 82.260 142.760 82.400 142.925 ;
        RECT 82.200 142.440 82.460 142.760 ;
        RECT 83.120 141.760 83.380 142.080 ;
        RECT 83.180 140.690 83.320 141.760 ;
        RECT 80.820 139.380 81.080 139.700 ;
        RECT 83.110 132.440 83.390 140.690 ;
        RECT 84.560 140.040 84.700 147.800 ;
        RECT 85.020 147.520 85.160 147.800 ;
        RECT 84.960 147.200 85.220 147.520 ;
        RECT 85.160 146.665 87.040 147.035 ;
        RECT 87.780 146.500 87.920 148.365 ;
        RECT 87.720 146.180 87.980 146.500 ;
        RECT 88.240 145.820 88.380 166.840 ;
        RECT 88.700 165.540 88.840 172.700 ;
        RECT 89.160 166.900 89.300 173.380 ;
        RECT 90.080 173.020 90.220 173.380 ;
        RECT 90.020 172.700 90.280 173.020 ;
        RECT 89.560 171.680 89.820 172.000 ;
        RECT 89.100 166.580 89.360 166.900 ;
        RECT 88.640 165.220 88.900 165.540 ;
        RECT 89.100 165.220 89.360 165.540 ;
        RECT 89.160 164.520 89.300 165.220 ;
        RECT 88.630 164.005 88.910 164.375 ;
        RECT 89.100 164.200 89.360 164.520 ;
        RECT 88.700 156.020 88.840 164.005 ;
        RECT 88.640 155.700 88.900 156.020 ;
        RECT 88.630 155.165 88.910 155.535 ;
        RECT 88.700 154.060 88.840 155.165 ;
        RECT 88.700 153.920 89.300 154.060 ;
        RECT 88.640 152.640 88.900 152.960 ;
        RECT 88.700 151.600 88.840 152.640 ;
        RECT 88.640 151.280 88.900 151.600 ;
        RECT 89.160 150.920 89.300 153.920 ;
        RECT 89.100 150.830 89.360 150.920 ;
        RECT 88.700 150.690 89.360 150.830 ;
        RECT 88.700 148.540 88.840 150.690 ;
        RECT 89.100 150.600 89.360 150.690 ;
        RECT 89.100 149.920 89.360 150.240 ;
        RECT 89.160 149.220 89.300 149.920 ;
        RECT 89.100 148.900 89.360 149.220 ;
        RECT 88.640 148.220 88.900 148.540 ;
        RECT 89.620 148.200 89.760 171.680 ;
        RECT 90.540 170.300 90.680 182.560 ;
        RECT 91.000 181.520 91.140 191.490 ;
        RECT 91.390 189.845 91.670 190.215 ;
        RECT 91.920 190.020 92.060 196.840 ;
        RECT 92.840 196.480 92.980 202.620 ;
        RECT 93.300 201.920 93.440 212.820 ;
        RECT 99.740 210.080 99.880 213.160 ;
        RECT 102.440 212.480 102.700 212.800 ;
        RECT 99.680 209.760 99.940 210.080 ;
        RECT 99.740 208.040 99.880 209.760 ;
        RECT 100.160 209.225 102.040 209.595 ;
        RECT 102.500 208.575 102.640 212.480 ;
        RECT 107.100 211.780 107.240 215.200 ;
        RECT 107.040 211.460 107.300 211.780 ;
        RECT 112.100 211.460 112.360 211.780 ;
        RECT 106.120 210.780 106.380 211.100 ;
        RECT 106.180 209.060 106.320 210.780 ;
        RECT 109.340 210.440 109.600 210.760 ;
        RECT 106.120 208.740 106.380 209.060 ;
        RECT 102.430 208.205 102.710 208.575 ;
        RECT 104.280 208.400 104.540 208.720 ;
        RECT 102.500 208.040 102.640 208.205 ;
        RECT 98.300 207.720 98.560 208.040 ;
        RECT 99.220 207.720 99.480 208.040 ;
        RECT 99.680 207.720 99.940 208.040 ;
        RECT 102.440 207.720 102.700 208.040 ;
        RECT 93.700 205.680 93.960 206.000 ;
        RECT 93.240 201.600 93.500 201.920 ;
        RECT 93.760 196.480 93.900 205.680 ;
        RECT 96.920 204.320 97.180 204.640 ;
        RECT 96.460 199.560 96.720 199.880 ;
        RECT 94.160 199.220 94.420 199.540 ;
        RECT 94.220 197.840 94.360 199.220 ;
        RECT 94.620 198.880 94.880 199.200 ;
        RECT 94.160 197.520 94.420 197.840 ;
        RECT 92.780 196.160 93.040 196.480 ;
        RECT 93.700 196.160 93.960 196.480 ;
        RECT 92.780 194.120 93.040 194.440 ;
        RECT 92.320 191.400 92.580 191.720 ;
        RECT 91.460 187.300 91.600 189.845 ;
        RECT 91.860 189.700 92.120 190.020 ;
        RECT 92.380 188.660 92.520 191.400 ;
        RECT 92.320 188.340 92.580 188.660 ;
        RECT 91.400 186.980 91.660 187.300 ;
        RECT 92.310 183.725 92.590 184.095 ;
        RECT 92.320 183.580 92.580 183.725 ;
        RECT 91.400 183.240 91.660 183.560 ;
        RECT 90.940 181.200 91.200 181.520 ;
        RECT 90.940 180.520 91.200 180.840 ;
        RECT 91.000 178.800 91.140 180.520 ;
        RECT 90.940 178.480 91.200 178.800 ;
        RECT 91.460 177.780 91.600 183.240 ;
        RECT 92.320 182.560 92.580 182.880 ;
        RECT 92.380 181.860 92.520 182.560 ;
        RECT 92.320 181.540 92.580 181.860 ;
        RECT 92.840 181.260 92.980 194.120 ;
        RECT 94.160 191.400 94.420 191.720 ;
        RECT 93.240 186.980 93.500 187.300 ;
        RECT 93.300 183.900 93.440 186.980 ;
        RECT 94.220 186.620 94.360 191.400 ;
        RECT 94.680 190.895 94.820 198.880 ;
        RECT 96.000 195.140 96.260 195.460 ;
        RECT 95.540 191.400 95.800 191.720 ;
        RECT 94.610 190.525 94.890 190.895 ;
        RECT 95.600 186.620 95.740 191.400 ;
        RECT 94.160 186.300 94.420 186.620 ;
        RECT 95.540 186.300 95.800 186.620 ;
        RECT 93.240 183.580 93.500 183.900 ;
        RECT 92.380 181.120 92.980 181.260 ;
        RECT 93.300 181.180 93.440 183.580 ;
        RECT 93.700 183.240 93.960 183.560 ;
        RECT 91.860 179.840 92.120 180.160 ;
        RECT 91.400 177.460 91.660 177.780 ;
        RECT 91.920 175.400 92.060 179.840 ;
        RECT 92.380 175.400 92.520 181.120 ;
        RECT 93.240 180.860 93.500 181.180 ;
        RECT 92.780 180.520 93.040 180.840 ;
        RECT 92.840 179.140 92.980 180.520 ;
        RECT 92.780 178.820 93.040 179.140 ;
        RECT 93.240 177.120 93.500 177.440 ;
        RECT 92.780 175.760 93.040 176.080 ;
        RECT 92.840 175.400 92.980 175.760 ;
        RECT 91.860 175.080 92.120 175.400 ;
        RECT 92.320 175.255 92.580 175.400 ;
        RECT 92.310 174.885 92.590 175.255 ;
        RECT 92.780 175.080 93.040 175.400 ;
        RECT 90.940 174.400 91.200 174.720 ;
        RECT 91.400 174.400 91.660 174.720 ;
        RECT 91.000 173.895 91.140 174.400 ;
        RECT 90.930 173.525 91.210 173.895 ;
        RECT 90.930 172.845 91.210 173.215 ;
        RECT 91.460 173.020 91.600 174.400 ;
        RECT 91.860 173.380 92.120 173.700 ;
        RECT 91.000 170.640 91.140 172.845 ;
        RECT 91.400 172.700 91.660 173.020 ;
        RECT 90.940 170.320 91.200 170.640 ;
        RECT 90.480 169.980 90.740 170.300 ;
        RECT 90.940 169.640 91.200 169.960 ;
        RECT 91.400 169.640 91.660 169.960 ;
        RECT 90.020 169.300 90.280 169.620 ;
        RECT 90.080 168.455 90.220 169.300 ;
        RECT 90.010 168.085 90.290 168.455 ;
        RECT 91.000 167.920 91.140 169.640 ;
        RECT 91.460 168.260 91.600 169.640 ;
        RECT 91.400 167.940 91.660 168.260 ;
        RECT 90.940 167.600 91.200 167.920 ;
        RECT 91.920 165.540 92.060 173.380 ;
        RECT 92.380 167.580 92.520 174.885 ;
        RECT 92.770 173.525 93.050 173.895 ;
        RECT 92.840 173.020 92.980 173.525 ;
        RECT 92.780 172.700 93.040 173.020 ;
        RECT 92.780 171.680 93.040 172.000 ;
        RECT 92.840 170.300 92.980 171.680 ;
        RECT 92.780 169.980 93.040 170.300 ;
        RECT 92.840 167.830 92.980 169.980 ;
        RECT 93.300 169.870 93.440 177.120 ;
        RECT 93.760 173.700 93.900 183.240 ;
        RECT 94.220 176.615 94.360 186.300 ;
        RECT 95.070 185.085 95.350 185.455 ;
        RECT 95.140 184.240 95.280 185.085 ;
        RECT 95.080 183.920 95.340 184.240 ;
        RECT 95.600 183.900 95.740 186.300 ;
        RECT 95.540 183.580 95.800 183.900 ;
        RECT 94.680 183.160 95.740 183.300 ;
        RECT 94.680 182.880 94.820 183.160 ;
        RECT 94.620 182.560 94.880 182.880 ;
        RECT 95.080 182.560 95.340 182.880 ;
        RECT 94.620 181.540 94.880 181.860 ;
        RECT 94.150 176.245 94.430 176.615 ;
        RECT 94.680 175.140 94.820 181.540 ;
        RECT 95.140 178.460 95.280 182.560 ;
        RECT 95.600 180.015 95.740 183.160 ;
        RECT 96.060 181.180 96.200 195.140 ;
        RECT 96.520 192.740 96.660 199.560 ;
        RECT 96.460 192.420 96.720 192.740 ;
        RECT 96.460 189.360 96.720 189.680 ;
        RECT 96.000 180.860 96.260 181.180 ;
        RECT 95.530 179.645 95.810 180.015 ;
        RECT 96.000 179.840 96.260 180.160 ;
        RECT 96.060 179.335 96.200 179.840 ;
        RECT 95.540 178.820 95.800 179.140 ;
        RECT 95.990 178.965 96.270 179.335 ;
        RECT 95.080 178.140 95.340 178.460 ;
        RECT 95.600 175.740 95.740 178.820 ;
        RECT 96.060 178.800 96.200 178.965 ;
        RECT 96.000 178.480 96.260 178.800 ;
        RECT 96.060 175.740 96.200 178.480 ;
        RECT 95.540 175.420 95.800 175.740 ;
        RECT 96.000 175.420 96.260 175.740 ;
        RECT 94.680 175.000 95.740 175.140 ;
        RECT 94.160 174.400 94.420 174.720 ;
        RECT 94.220 173.895 94.360 174.400 ;
        RECT 93.700 173.380 93.960 173.700 ;
        RECT 94.150 173.525 94.430 173.895 ;
        RECT 95.080 173.380 95.340 173.700 ;
        RECT 93.700 172.360 93.960 172.680 ;
        RECT 93.760 170.980 93.900 172.360 ;
        RECT 94.150 171.485 94.430 171.855 ;
        RECT 93.700 170.660 93.960 170.980 ;
        RECT 93.300 169.730 93.900 169.870 ;
        RECT 93.240 168.960 93.500 169.280 ;
        RECT 93.760 169.020 93.900 169.730 ;
        RECT 94.220 169.620 94.360 171.485 ;
        RECT 94.160 169.300 94.420 169.620 ;
        RECT 93.300 168.455 93.440 168.960 ;
        RECT 93.760 168.880 94.360 169.020 ;
        RECT 94.620 168.960 94.880 169.280 ;
        RECT 93.230 168.085 93.510 168.455 ;
        RECT 93.700 167.940 93.960 168.260 ;
        RECT 93.240 167.830 93.500 167.920 ;
        RECT 92.840 167.690 93.500 167.830 ;
        RECT 93.240 167.600 93.500 167.690 ;
        RECT 92.320 167.260 92.580 167.580 ;
        RECT 91.860 165.220 92.120 165.540 ;
        RECT 92.320 165.220 92.580 165.540 ;
        RECT 90.020 164.880 90.280 165.200 ;
        RECT 92.380 164.940 92.520 165.220 ;
        RECT 90.080 163.695 90.220 164.880 ;
        RECT 91.920 164.860 92.520 164.940 ;
        RECT 92.780 164.880 93.040 165.200 ;
        RECT 91.860 164.800 92.520 164.860 ;
        RECT 91.860 164.540 92.120 164.800 ;
        RECT 90.480 164.200 90.740 164.520 ;
        RECT 90.010 163.325 90.290 163.695 ;
        RECT 90.540 158.400 90.680 164.200 ;
        RECT 91.400 163.860 91.660 164.180 ;
        RECT 90.940 163.520 91.200 163.840 ;
        RECT 90.480 158.080 90.740 158.400 ;
        RECT 90.540 157.040 90.680 158.080 ;
        RECT 90.480 156.720 90.740 157.040 ;
        RECT 91.000 152.560 91.140 163.520 ;
        RECT 91.460 160.100 91.600 163.860 ;
        RECT 91.860 163.520 92.120 163.840 ;
        RECT 91.920 162.140 92.060 163.520 ;
        RECT 92.840 162.140 92.980 164.880 ;
        RECT 93.300 164.520 93.440 167.600 ;
        RECT 93.240 164.200 93.500 164.520 ;
        RECT 91.860 161.820 92.120 162.140 ;
        RECT 92.780 161.820 93.040 162.140 ;
        RECT 92.320 161.480 92.580 161.800 ;
        RECT 91.400 159.780 91.660 160.100 ;
        RECT 92.380 157.380 92.520 161.480 ;
        RECT 93.300 161.460 93.440 164.200 ;
        RECT 93.240 161.140 93.500 161.460 ;
        RECT 92.320 157.060 92.580 157.380 ;
        RECT 92.320 155.360 92.580 155.680 ;
        RECT 92.380 154.175 92.520 155.360 ;
        RECT 92.310 153.805 92.590 154.175 ;
        RECT 92.320 152.640 92.580 152.960 ;
        RECT 90.540 152.420 91.140 152.560 ;
        RECT 90.010 150.405 90.290 150.775 ;
        RECT 90.080 148.200 90.220 150.405 ;
        RECT 89.100 147.880 89.360 148.200 ;
        RECT 89.560 147.880 89.820 148.200 ;
        RECT 90.020 147.880 90.280 148.200 ;
        RECT 88.640 147.200 88.900 147.520 ;
        RECT 88.180 145.500 88.440 145.820 ;
        RECT 85.880 145.390 86.140 145.480 ;
        RECT 85.880 145.250 87.000 145.390 ;
        RECT 85.880 145.160 86.140 145.250 ;
        RECT 86.860 145.220 87.000 145.250 ;
        RECT 88.700 145.220 88.840 147.200 ;
        RECT 89.160 146.500 89.300 147.880 ;
        RECT 89.100 146.180 89.360 146.500 ;
        RECT 86.860 145.080 88.840 145.220 ;
        RECT 90.080 145.140 90.220 147.880 ;
        RECT 90.540 145.820 90.680 152.420 ;
        RECT 91.860 151.620 92.120 151.940 ;
        RECT 90.940 149.920 91.200 150.240 ;
        RECT 91.920 150.095 92.060 151.620 ;
        RECT 91.000 148.200 91.140 149.920 ;
        RECT 91.850 149.725 92.130 150.095 ;
        RECT 92.380 149.415 92.520 152.640 ;
        RECT 92.310 149.045 92.590 149.415 ;
        RECT 90.940 147.880 91.200 148.200 ;
        RECT 91.400 147.540 91.660 147.860 ;
        RECT 90.480 145.500 90.740 145.820 ;
        RECT 90.930 145.645 91.210 146.015 ;
        RECT 91.460 145.820 91.600 147.540 ;
        RECT 90.020 144.820 90.280 145.140 ;
        RECT 87.260 144.480 87.520 144.800 ;
        RECT 87.320 143.780 87.460 144.480 ;
        RECT 87.260 143.460 87.520 143.780 ;
        RECT 91.000 142.760 91.140 145.645 ;
        RECT 91.400 145.500 91.660 145.820 ;
        RECT 91.400 144.480 91.660 144.800 ;
        RECT 91.460 143.100 91.600 144.480 ;
        RECT 93.760 143.780 93.900 167.940 ;
        RECT 94.220 164.520 94.360 168.880 ;
        RECT 94.680 168.260 94.820 168.960 ;
        RECT 94.620 167.940 94.880 168.260 ;
        RECT 95.140 167.660 95.280 173.380 ;
        RECT 94.680 167.520 95.280 167.660 ;
        RECT 94.160 164.200 94.420 164.520 ;
        RECT 94.160 163.520 94.420 163.840 ;
        RECT 94.220 152.560 94.360 163.520 ;
        RECT 94.680 152.870 94.820 167.520 ;
        RECT 95.080 166.920 95.340 167.240 ;
        RECT 95.140 162.820 95.280 166.920 ;
        RECT 95.600 164.520 95.740 175.000 ;
        RECT 96.000 174.740 96.260 175.060 ;
        RECT 96.060 173.215 96.200 174.740 ;
        RECT 96.520 173.360 96.660 189.360 ;
        RECT 96.980 189.000 97.120 204.320 ;
        RECT 98.360 203.620 98.500 207.720 ;
        RECT 98.760 206.020 99.020 206.340 ;
        RECT 98.300 203.300 98.560 203.620 ;
        RECT 97.840 203.135 98.100 203.280 ;
        RECT 97.830 202.765 98.110 203.135 ;
        RECT 98.820 202.600 98.960 206.020 ;
        RECT 98.760 202.280 99.020 202.600 ;
        RECT 98.300 199.900 98.560 200.220 ;
        RECT 97.380 199.620 97.640 199.880 ;
        RECT 97.380 199.560 98.040 199.620 ;
        RECT 97.440 199.480 98.040 199.560 ;
        RECT 97.900 196.820 98.040 199.480 ;
        RECT 98.360 197.695 98.500 199.900 ;
        RECT 98.760 199.220 99.020 199.540 ;
        RECT 98.290 197.325 98.570 197.695 ;
        RECT 97.840 196.500 98.100 196.820 ;
        RECT 97.380 194.460 97.640 194.780 ;
        RECT 97.440 192.060 97.580 194.460 ;
        RECT 97.380 191.740 97.640 192.060 ;
        RECT 96.920 188.680 97.180 189.000 ;
        RECT 97.900 187.060 98.040 196.500 ;
        RECT 98.300 191.400 98.560 191.720 ;
        RECT 98.360 189.340 98.500 191.400 ;
        RECT 98.300 189.020 98.560 189.340 ;
        RECT 96.980 186.920 98.040 187.060 ;
        RECT 96.980 185.455 97.120 186.920 ;
        RECT 97.840 186.300 98.100 186.620 ;
        RECT 96.910 185.085 97.190 185.455 ;
        RECT 96.920 183.580 97.180 183.900 ;
        RECT 97.380 183.580 97.640 183.900 ;
        RECT 96.980 179.050 97.120 183.580 ;
        RECT 97.440 180.160 97.580 183.580 ;
        RECT 97.900 181.860 98.040 186.300 ;
        RECT 98.360 184.240 98.500 189.020 ;
        RECT 98.820 186.620 98.960 199.220 ;
        RECT 99.280 194.780 99.420 207.720 ;
        RECT 100.160 203.785 102.040 204.155 ;
        RECT 102.440 202.620 102.700 202.940 ;
        RECT 101.970 201.405 102.250 201.775 ;
        RECT 102.040 200.220 102.180 201.405 ;
        RECT 102.500 200.900 102.640 202.620 ;
        RECT 102.900 202.280 103.160 202.600 ;
        RECT 102.440 200.580 102.700 200.900 ;
        RECT 101.980 199.900 102.240 200.220 ;
        RECT 99.680 198.880 99.940 199.200 ;
        RECT 102.440 198.880 102.700 199.200 ;
        RECT 99.740 198.180 99.880 198.880 ;
        RECT 100.160 198.345 102.040 198.715 ;
        RECT 99.680 197.860 99.940 198.180 ;
        RECT 101.980 196.900 102.240 197.160 ;
        RECT 102.500 196.900 102.640 198.880 ;
        RECT 101.980 196.840 102.640 196.900 ;
        RECT 101.520 196.500 101.780 196.820 ;
        RECT 102.040 196.760 102.640 196.840 ;
        RECT 99.220 194.460 99.480 194.780 ;
        RECT 101.580 194.440 101.720 196.500 ;
        RECT 102.960 195.655 103.100 202.280 ;
        RECT 103.820 200.240 104.080 200.560 ;
        RECT 103.880 198.180 104.020 200.240 ;
        RECT 103.820 197.860 104.080 198.180 ;
        RECT 103.820 196.840 104.080 197.160 ;
        RECT 103.360 196.160 103.620 196.480 ;
        RECT 102.890 195.285 103.170 195.655 ;
        RECT 102.440 194.800 102.700 195.120 ;
        RECT 101.520 194.120 101.780 194.440 ;
        RECT 102.500 194.295 102.640 194.800 ;
        RECT 102.900 194.460 103.160 194.780 ;
        RECT 103.420 194.690 103.560 196.160 ;
        RECT 103.880 195.460 104.020 196.840 ;
        RECT 103.820 195.140 104.080 195.460 ;
        RECT 103.820 194.690 104.080 194.780 ;
        RECT 103.420 194.550 104.080 194.690 ;
        RECT 103.820 194.460 104.080 194.550 ;
        RECT 99.680 193.780 99.940 194.100 ;
        RECT 102.430 193.925 102.710 194.295 ;
        RECT 99.220 192.420 99.480 192.740 ;
        RECT 99.280 191.720 99.420 192.420 ;
        RECT 99.220 191.400 99.480 191.720 ;
        RECT 99.220 190.720 99.480 191.040 ;
        RECT 99.280 190.215 99.420 190.720 ;
        RECT 99.210 189.845 99.490 190.215 ;
        RECT 99.220 189.020 99.480 189.340 ;
        RECT 99.280 186.620 99.420 189.020 ;
        RECT 98.760 186.300 99.020 186.620 ;
        RECT 99.220 186.300 99.480 186.620 ;
        RECT 98.760 185.620 99.020 185.940 ;
        RECT 98.300 183.920 98.560 184.240 ;
        RECT 98.820 183.900 98.960 185.620 ;
        RECT 98.760 183.580 99.020 183.900 ;
        RECT 99.220 182.560 99.480 182.880 ;
        RECT 97.840 181.540 98.100 181.860 ;
        RECT 99.280 181.180 99.420 182.560 ;
        RECT 99.220 180.860 99.480 181.180 ;
        RECT 97.840 180.180 98.100 180.500 ;
        RECT 97.380 179.840 97.640 180.160 ;
        RECT 96.980 178.910 97.580 179.050 ;
        RECT 96.920 178.140 97.180 178.460 ;
        RECT 95.990 172.845 96.270 173.215 ;
        RECT 96.460 173.040 96.720 173.360 ;
        RECT 96.980 172.680 97.120 178.140 ;
        RECT 97.440 176.420 97.580 178.910 ;
        RECT 97.380 176.100 97.640 176.420 ;
        RECT 97.380 175.080 97.640 175.400 ;
        RECT 96.920 172.360 97.180 172.680 ;
        RECT 96.000 168.960 96.260 169.280 ;
        RECT 96.060 168.260 96.200 168.960 ;
        RECT 96.000 167.940 96.260 168.260 ;
        RECT 96.980 167.580 97.120 172.360 ;
        RECT 97.440 170.980 97.580 175.080 ;
        RECT 97.380 170.660 97.640 170.980 ;
        RECT 97.380 169.300 97.640 169.620 ;
        RECT 97.440 168.260 97.580 169.300 ;
        RECT 97.380 167.940 97.640 168.260 ;
        RECT 96.920 167.260 97.180 167.580 ;
        RECT 97.370 166.725 97.650 167.095 ;
        RECT 96.000 166.240 96.260 166.560 ;
        RECT 96.060 164.520 96.200 166.240 ;
        RECT 97.440 164.940 97.580 166.725 ;
        RECT 96.520 164.800 97.580 164.940 ;
        RECT 96.520 164.520 96.660 164.800 ;
        RECT 95.540 164.200 95.800 164.520 ;
        RECT 96.000 164.200 96.260 164.520 ;
        RECT 96.460 164.200 96.720 164.520 ;
        RECT 97.380 164.200 97.640 164.520 ;
        RECT 95.080 162.500 95.340 162.820 ;
        RECT 95.080 160.800 95.340 161.120 ;
        RECT 95.140 156.700 95.280 160.800 ;
        RECT 95.600 159.080 95.740 164.200 ;
        RECT 96.060 159.420 96.200 164.200 ;
        RECT 97.440 162.820 97.580 164.200 ;
        RECT 97.380 162.500 97.640 162.820 ;
        RECT 97.380 161.480 97.640 161.800 ;
        RECT 96.000 159.100 96.260 159.420 ;
        RECT 97.440 159.080 97.580 161.480 ;
        RECT 97.900 161.120 98.040 180.180 ;
        RECT 98.760 179.840 99.020 180.160 ;
        RECT 99.220 179.840 99.480 180.160 ;
        RECT 98.820 175.990 98.960 179.840 ;
        RECT 99.280 178.120 99.420 179.840 ;
        RECT 99.740 178.460 99.880 193.780 ;
        RECT 100.160 192.905 102.040 193.275 ;
        RECT 102.500 192.060 102.640 193.925 ;
        RECT 102.960 192.400 103.100 194.460 ;
        RECT 102.900 192.080 103.160 192.400 ;
        RECT 102.440 191.740 102.700 192.060 ;
        RECT 104.340 191.720 104.480 208.400 ;
        RECT 106.580 207.895 106.840 208.040 ;
        RECT 106.570 207.525 106.850 207.895 ;
        RECT 105.660 204.320 105.920 204.640 ;
        RECT 105.720 202.600 105.860 204.320 ;
        RECT 104.740 202.280 105.000 202.600 ;
        RECT 105.200 202.280 105.460 202.600 ;
        RECT 105.660 202.280 105.920 202.600 ;
        RECT 104.800 200.900 104.940 202.280 ;
        RECT 104.740 200.580 105.000 200.900 ;
        RECT 104.740 196.500 105.000 196.820 ;
        RECT 104.800 195.460 104.940 196.500 ;
        RECT 104.740 195.140 105.000 195.460 ;
        RECT 101.980 191.400 102.240 191.720 ;
        RECT 102.900 191.400 103.160 191.720 ;
        RECT 103.820 191.400 104.080 191.720 ;
        RECT 104.280 191.400 104.540 191.720 ;
        RECT 102.040 190.020 102.180 191.400 ;
        RECT 102.440 191.060 102.700 191.380 ;
        RECT 101.980 189.700 102.240 190.020 ;
        RECT 100.160 187.465 102.040 187.835 ;
        RECT 102.500 187.060 102.640 191.060 ;
        RECT 102.960 188.320 103.100 191.400 ;
        RECT 103.880 190.020 104.020 191.400 ;
        RECT 103.820 189.700 104.080 190.020 ;
        RECT 103.360 189.020 103.620 189.340 ;
        RECT 102.900 188.000 103.160 188.320 ;
        RECT 100.200 186.920 102.640 187.060 ;
        RECT 100.200 184.775 100.340 186.920 ;
        RECT 102.960 186.700 103.100 188.000 ;
        RECT 100.600 186.300 100.860 186.620 ;
        RECT 102.500 186.560 103.100 186.700 ;
        RECT 103.420 186.620 103.560 189.020 ;
        RECT 104.340 187.380 104.480 191.400 ;
        RECT 104.800 189.340 104.940 195.140 ;
        RECT 104.740 189.020 105.000 189.340 ;
        RECT 104.340 187.240 104.940 187.380 ;
        RECT 100.130 184.405 100.410 184.775 ;
        RECT 100.660 184.580 100.800 186.300 ;
        RECT 101.980 185.960 102.240 186.280 ;
        RECT 102.040 184.580 102.180 185.960 ;
        RECT 100.600 184.260 100.860 184.580 ;
        RECT 101.980 184.260 102.240 184.580 ;
        RECT 101.510 183.725 101.790 184.095 ;
        RECT 101.520 183.580 101.780 183.725 ;
        RECT 101.580 182.790 101.720 183.580 ;
        RECT 102.500 183.130 102.640 186.560 ;
        RECT 103.360 186.300 103.620 186.620 ;
        RECT 103.420 183.980 103.560 186.300 ;
        RECT 104.280 185.620 104.540 185.940 ;
        RECT 102.960 183.900 103.560 183.980 ;
        RECT 102.900 183.840 103.560 183.900 ;
        RECT 102.900 183.580 103.160 183.840 ;
        RECT 102.900 183.130 103.160 183.220 ;
        RECT 102.500 182.990 103.160 183.130 ;
        RECT 102.900 182.900 103.160 182.990 ;
        RECT 101.580 182.650 102.640 182.790 ;
        RECT 100.160 182.025 102.040 182.395 ;
        RECT 100.140 180.860 100.400 181.180 ;
        RECT 99.680 178.140 99.940 178.460 ;
        RECT 99.220 177.800 99.480 178.120 ;
        RECT 100.200 177.860 100.340 180.860 ;
        RECT 101.980 180.410 102.240 180.500 ;
        RECT 101.580 180.270 102.240 180.410 ;
        RECT 101.580 178.030 101.720 180.270 ;
        RECT 101.980 180.180 102.240 180.270 ;
        RECT 102.500 179.140 102.640 182.650 ;
        RECT 101.980 178.820 102.240 179.140 ;
        RECT 102.440 178.820 102.700 179.140 ;
        RECT 102.040 178.655 102.180 178.820 ;
        RECT 101.970 178.285 102.250 178.655 ;
        RECT 101.580 177.890 102.640 178.030 ;
        RECT 98.360 175.850 98.960 175.990 ;
        RECT 99.740 177.720 100.340 177.860 ;
        RECT 98.360 175.400 98.500 175.850 ;
        RECT 99.740 175.740 99.880 177.720 ;
        RECT 100.160 176.585 102.040 176.955 ;
        RECT 101.060 176.100 101.320 176.420 ;
        RECT 101.980 176.100 102.240 176.420 ;
        RECT 99.220 175.420 99.480 175.740 ;
        RECT 99.680 175.420 99.940 175.740 ;
        RECT 98.300 175.080 98.560 175.400 ;
        RECT 99.280 173.700 99.420 175.420 ;
        RECT 101.120 175.400 101.260 176.100 ;
        RECT 101.060 175.080 101.320 175.400 ;
        RECT 100.600 174.740 100.860 175.060 ;
        RECT 100.660 173.700 100.800 174.740 ;
        RECT 99.220 173.380 99.480 173.700 ;
        RECT 100.600 173.380 100.860 173.700 ;
        RECT 98.760 172.020 99.020 172.340 ;
        RECT 98.300 168.960 98.560 169.280 ;
        RECT 98.360 163.015 98.500 168.960 ;
        RECT 98.290 162.645 98.570 163.015 ;
        RECT 98.820 162.140 98.960 172.020 ;
        RECT 99.280 167.580 99.420 173.380 ;
        RECT 100.600 172.250 100.860 172.340 ;
        RECT 101.120 172.250 101.260 175.080 ;
        RECT 101.520 174.740 101.780 175.060 ;
        RECT 101.580 172.930 101.720 174.740 ;
        RECT 102.040 174.720 102.180 176.100 ;
        RECT 102.500 175.740 102.640 177.890 ;
        RECT 102.960 175.740 103.100 182.900 ;
        RECT 103.420 180.500 103.560 183.840 ;
        RECT 103.820 180.860 104.080 181.180 ;
        RECT 103.360 180.180 103.620 180.500 ;
        RECT 103.350 178.965 103.630 179.335 ;
        RECT 103.420 178.460 103.560 178.965 ;
        RECT 103.880 178.460 104.020 180.860 ;
        RECT 104.340 180.160 104.480 185.620 ;
        RECT 104.800 183.900 104.940 187.240 ;
        RECT 104.740 183.580 105.000 183.900 ;
        RECT 104.280 179.840 104.540 180.160 ;
        RECT 104.340 178.460 104.480 179.840 ;
        RECT 103.360 178.140 103.620 178.460 ;
        RECT 103.820 178.140 104.080 178.460 ;
        RECT 104.280 178.140 104.540 178.460 ;
        RECT 104.340 177.860 104.480 178.140 ;
        RECT 103.880 177.720 104.480 177.860 ;
        RECT 103.880 177.690 104.020 177.720 ;
        RECT 103.420 177.550 104.020 177.690 ;
        RECT 102.440 175.420 102.700 175.740 ;
        RECT 102.900 175.420 103.160 175.740 ;
        RECT 101.980 174.400 102.240 174.720 ;
        RECT 102.440 174.400 102.700 174.720 ;
        RECT 101.980 172.930 102.240 173.020 ;
        RECT 101.580 172.790 102.240 172.930 ;
        RECT 101.580 172.535 101.720 172.790 ;
        RECT 101.980 172.700 102.240 172.790 ;
        RECT 100.600 172.110 101.260 172.250 ;
        RECT 101.510 172.165 101.790 172.535 ;
        RECT 100.600 172.020 100.860 172.110 ;
        RECT 100.160 171.145 102.040 171.515 ;
        RECT 101.980 170.320 102.240 170.640 ;
        RECT 102.040 169.190 102.180 170.320 ;
        RECT 102.500 169.960 102.640 174.400 ;
        RECT 103.420 173.020 103.560 177.550 ;
        RECT 104.270 176.500 104.550 176.615 ;
        RECT 103.880 176.360 104.550 176.500 ;
        RECT 103.880 173.020 104.020 176.360 ;
        RECT 104.270 176.245 104.550 176.360 ;
        RECT 104.280 175.255 104.540 175.400 ;
        RECT 104.270 174.885 104.550 175.255 ;
        RECT 103.360 172.700 103.620 173.020 ;
        RECT 103.820 172.700 104.080 173.020 ;
        RECT 102.900 172.020 103.160 172.340 ;
        RECT 102.960 171.175 103.100 172.020 ;
        RECT 102.890 170.805 103.170 171.175 ;
        RECT 102.960 169.960 103.100 170.805 ;
        RECT 103.880 170.495 104.020 172.700 ;
        RECT 103.810 170.125 104.090 170.495 ;
        RECT 104.280 170.320 104.540 170.640 ;
        RECT 102.440 169.640 102.700 169.960 ;
        RECT 102.900 169.640 103.160 169.960 ;
        RECT 102.040 169.050 102.640 169.190 ;
        RECT 99.220 167.260 99.480 167.580 ;
        RECT 99.680 167.260 99.940 167.580 ;
        RECT 99.740 167.095 99.880 167.260 ;
        RECT 99.670 166.725 99.950 167.095 ;
        RECT 99.220 166.240 99.480 166.560 ;
        RECT 99.280 164.375 99.420 166.240 ;
        RECT 100.160 165.705 102.040 166.075 ;
        RECT 101.980 165.220 102.240 165.540 ;
        RECT 99.210 164.005 99.490 164.375 ;
        RECT 101.520 164.200 101.780 164.520 ;
        RECT 99.220 163.520 99.480 163.840 ;
        RECT 101.580 163.695 101.720 164.200 ;
        RECT 98.760 162.050 99.020 162.140 ;
        RECT 98.360 161.910 99.020 162.050 ;
        RECT 97.840 160.800 98.100 161.120 ;
        RECT 95.540 158.760 95.800 159.080 ;
        RECT 97.380 158.935 97.640 159.080 ;
        RECT 97.370 158.565 97.650 158.935 ;
        RECT 97.840 158.760 98.100 159.080 ;
        RECT 95.080 156.380 95.340 156.700 ;
        RECT 95.140 153.495 95.280 156.380 ;
        RECT 97.440 155.680 97.580 158.565 ;
        RECT 97.900 157.380 98.040 158.760 ;
        RECT 97.840 157.060 98.100 157.380 ;
        RECT 97.380 155.360 97.640 155.680 ;
        RECT 98.360 154.660 98.500 161.910 ;
        RECT 98.760 161.820 99.020 161.910 ;
        RECT 98.760 161.140 99.020 161.460 ;
        RECT 98.820 155.680 98.960 161.140 ;
        RECT 99.280 159.080 99.420 163.520 ;
        RECT 101.510 163.325 101.790 163.695 ;
        RECT 102.040 162.050 102.180 165.220 ;
        RECT 102.500 164.520 102.640 169.050 ;
        RECT 103.360 167.600 103.620 167.920 ;
        RECT 102.900 166.920 103.160 167.240 ;
        RECT 102.440 164.200 102.700 164.520 ;
        RECT 102.960 162.480 103.100 166.920 ;
        RECT 103.420 162.480 103.560 167.600 ;
        RECT 104.340 164.520 104.480 170.320 ;
        RECT 104.280 164.200 104.540 164.520 ;
        RECT 102.900 162.160 103.160 162.480 ;
        RECT 103.360 162.160 103.620 162.480 ;
        RECT 102.440 162.050 102.700 162.140 ;
        RECT 104.280 162.050 104.540 162.140 ;
        RECT 102.040 161.910 102.700 162.050 ;
        RECT 102.440 161.820 102.700 161.910 ;
        RECT 103.880 161.910 104.540 162.050 ;
        RECT 99.680 160.800 99.940 161.120 ;
        RECT 99.740 159.080 99.880 160.800 ;
        RECT 100.160 160.265 102.040 160.635 ;
        RECT 102.500 160.010 102.640 161.820 ;
        RECT 101.120 159.870 102.640 160.010 ;
        RECT 100.600 159.615 100.860 159.760 ;
        RECT 100.140 159.100 100.400 159.420 ;
        RECT 100.590 159.245 100.870 159.615 ;
        RECT 99.220 158.760 99.480 159.080 ;
        RECT 99.680 158.760 99.940 159.080 ;
        RECT 99.280 156.700 99.420 158.760 ;
        RECT 99.220 156.380 99.480 156.700 ;
        RECT 98.760 155.360 99.020 155.680 ;
        RECT 100.200 155.590 100.340 159.100 ;
        RECT 100.600 156.950 100.860 157.040 ;
        RECT 101.120 156.950 101.260 159.870 ;
        RECT 103.880 159.670 104.020 161.910 ;
        RECT 104.280 161.820 104.540 161.910 ;
        RECT 104.280 160.800 104.540 161.120 ;
        RECT 100.600 156.810 101.260 156.950 ;
        RECT 101.580 159.530 104.020 159.670 ;
        RECT 100.600 156.720 100.860 156.810 ;
        RECT 101.580 156.700 101.720 159.530 ;
        RECT 104.340 159.080 104.480 160.800 ;
        RECT 104.280 158.760 104.540 159.080 ;
        RECT 104.340 157.040 104.480 158.760 ;
        RECT 104.280 156.720 104.540 157.040 ;
        RECT 101.520 156.380 101.780 156.700 ;
        RECT 102.900 156.380 103.160 156.700 ;
        RECT 102.440 156.040 102.700 156.360 ;
        RECT 99.740 155.450 100.340 155.590 ;
        RECT 98.300 154.570 98.560 154.660 ;
        RECT 98.300 154.430 99.420 154.570 ;
        RECT 98.300 154.340 98.560 154.430 ;
        RECT 95.070 153.125 95.350 153.495 ;
        RECT 97.840 153.320 98.100 153.640 ;
        RECT 95.080 152.870 95.340 152.960 ;
        RECT 94.680 152.730 95.340 152.870 ;
        RECT 95.080 152.640 95.340 152.730 ;
        RECT 94.220 152.420 94.820 152.560 ;
        RECT 94.680 145.820 94.820 152.420 ;
        RECT 97.900 151.940 98.040 153.320 ;
        RECT 98.760 152.640 99.020 152.960 ;
        RECT 97.380 151.620 97.640 151.940 ;
        RECT 97.840 151.620 98.100 151.940 ;
        RECT 98.290 151.765 98.570 152.135 ;
        RECT 97.440 150.580 97.580 151.620 ;
        RECT 97.380 150.260 97.640 150.580 ;
        RECT 98.360 148.540 98.500 151.765 ;
        RECT 98.820 150.830 98.960 152.640 ;
        RECT 99.280 151.600 99.420 154.430 ;
        RECT 99.740 153.890 99.880 155.450 ;
        RECT 100.160 154.825 102.040 155.195 ;
        RECT 101.520 153.890 101.780 153.980 ;
        RECT 99.740 153.750 101.780 153.890 ;
        RECT 101.520 153.660 101.780 153.750 ;
        RECT 101.980 153.660 102.240 153.980 ;
        RECT 101.060 152.870 101.320 152.960 ;
        RECT 102.040 152.870 102.180 153.660 ;
        RECT 102.500 153.640 102.640 156.040 ;
        RECT 102.440 153.320 102.700 153.640 ;
        RECT 102.960 152.870 103.100 156.380 ;
        RECT 103.360 154.340 103.620 154.660 ;
        RECT 103.420 153.640 103.560 154.340 ;
        RECT 103.360 153.320 103.620 153.640 ;
        RECT 101.060 152.730 103.100 152.870 ;
        RECT 101.060 152.640 101.320 152.730 ;
        RECT 103.820 152.640 104.080 152.960 ;
        RECT 101.050 151.765 101.330 152.135 ;
        RECT 101.120 151.600 101.260 151.765 ;
        RECT 102.440 151.620 102.700 151.940 ;
        RECT 99.220 151.280 99.480 151.600 ;
        RECT 101.060 151.280 101.320 151.600 ;
        RECT 98.820 150.690 99.880 150.830 ;
        RECT 99.740 150.240 99.880 150.690 ;
        RECT 102.500 150.580 102.640 151.620 ;
        RECT 102.440 150.260 102.700 150.580 ;
        RECT 98.760 149.920 99.020 150.240 ;
        RECT 99.680 149.920 99.940 150.240 ;
        RECT 98.300 148.220 98.560 148.540 ;
        RECT 98.820 148.200 98.960 149.920 ;
        RECT 98.760 147.880 99.020 148.200 ;
        RECT 99.740 147.860 99.880 149.920 ;
        RECT 100.160 149.385 102.040 149.755 ;
        RECT 102.440 148.220 102.700 148.540 ;
        RECT 99.680 147.540 99.940 147.860 ;
        RECT 100.600 147.200 100.860 147.520 ;
        RECT 99.680 146.410 99.940 146.500 ;
        RECT 100.130 146.410 100.410 146.695 ;
        RECT 99.680 146.325 100.410 146.410 ;
        RECT 99.680 146.270 100.340 146.325 ;
        RECT 99.680 146.180 99.940 146.270 ;
        RECT 94.620 145.500 94.880 145.820 ;
        RECT 100.660 145.480 100.800 147.200 ;
        RECT 101.060 146.180 101.320 146.500 ;
        RECT 96.920 145.160 97.180 145.480 ;
        RECT 100.600 145.160 100.860 145.480 ;
        RECT 96.460 144.480 96.720 144.800 ;
        RECT 96.520 143.780 96.660 144.480 ;
        RECT 93.700 143.460 93.960 143.780 ;
        RECT 96.460 143.460 96.720 143.780 ;
        RECT 91.400 142.780 91.660 143.100 ;
        RECT 90.940 142.440 91.200 142.760 ;
        RECT 89.100 141.760 89.360 142.080 ;
        RECT 91.400 141.760 91.660 142.080 ;
        RECT 96.460 141.760 96.720 142.080 ;
        RECT 85.160 141.225 87.040 141.595 ;
        RECT 87.320 141.000 87.920 141.140 ;
        RECT 87.320 140.690 87.460 141.000 ;
        RECT 84.500 139.720 84.760 140.040 ;
        RECT 87.250 132.440 87.530 140.690 ;
        RECT 87.780 140.460 87.920 141.000 ;
        RECT 89.160 140.460 89.300 141.760 ;
        RECT 91.460 140.690 91.600 141.760 ;
        RECT 96.520 141.140 96.660 141.760 ;
        RECT 95.600 141.000 96.660 141.140 ;
        RECT 95.600 140.690 95.740 141.000 ;
        RECT 87.780 140.320 89.300 140.460 ;
        RECT 91.390 132.440 91.670 140.690 ;
        RECT 95.530 132.440 95.810 140.690 ;
        RECT 96.980 140.040 97.120 145.160 ;
        RECT 98.300 144.480 98.560 144.800 ;
        RECT 100.600 144.710 100.860 144.800 ;
        RECT 101.120 144.710 101.260 146.180 ;
        RECT 102.500 145.820 102.640 148.220 ;
        RECT 103.360 147.540 103.620 147.860 ;
        RECT 103.420 146.160 103.560 147.540 ;
        RECT 103.360 145.840 103.620 146.160 ;
        RECT 103.880 145.820 104.020 152.640 ;
        RECT 104.800 151.940 104.940 183.580 ;
        RECT 105.260 152.560 105.400 202.280 ;
        RECT 106.580 201.775 106.840 201.920 ;
        RECT 106.570 201.405 106.850 201.775 ;
        RECT 107.040 200.240 107.300 200.560 ;
        RECT 106.580 196.500 106.840 196.820 ;
        RECT 106.120 196.160 106.380 196.480 ;
        RECT 105.660 195.140 105.920 195.460 ;
        RECT 105.720 191.040 105.860 195.140 ;
        RECT 106.180 191.720 106.320 196.160 ;
        RECT 106.640 195.655 106.780 196.500 ;
        RECT 106.570 195.285 106.850 195.655 ;
        RECT 106.120 191.400 106.380 191.720 ;
        RECT 106.580 191.400 106.840 191.720 ;
        RECT 105.660 190.720 105.920 191.040 ;
        RECT 105.720 189.340 105.860 190.720 ;
        RECT 106.110 190.525 106.390 190.895 ;
        RECT 105.660 189.020 105.920 189.340 ;
        RECT 105.660 182.560 105.920 182.880 ;
        RECT 105.720 181.180 105.860 182.560 ;
        RECT 105.660 180.860 105.920 181.180 ;
        RECT 105.660 180.180 105.920 180.500 ;
        RECT 105.720 175.740 105.860 180.180 ;
        RECT 105.660 175.420 105.920 175.740 ;
        RECT 105.660 174.740 105.920 175.060 ;
        RECT 105.720 172.000 105.860 174.740 ;
        RECT 105.660 171.680 105.920 172.000 ;
        RECT 105.660 166.240 105.920 166.560 ;
        RECT 105.720 159.420 105.860 166.240 ;
        RECT 106.180 164.770 106.320 190.525 ;
        RECT 106.640 188.320 106.780 191.400 ;
        RECT 107.100 190.215 107.240 200.240 ;
        RECT 108.880 198.880 109.140 199.200 ;
        RECT 107.960 196.840 108.220 197.160 ;
        RECT 108.020 195.460 108.160 196.840 ;
        RECT 108.420 196.160 108.680 196.480 ;
        RECT 107.960 195.140 108.220 195.460 ;
        RECT 107.030 189.845 107.310 190.215 ;
        RECT 107.100 189.680 107.240 189.845 ;
        RECT 107.040 189.360 107.300 189.680 ;
        RECT 106.580 188.000 106.840 188.320 ;
        RECT 107.040 188.000 107.300 188.320 ;
        RECT 107.100 187.300 107.240 188.000 ;
        RECT 107.040 186.980 107.300 187.300 ;
        RECT 108.480 186.960 108.620 196.160 ;
        RECT 108.940 194.440 109.080 198.880 ;
        RECT 108.880 194.120 109.140 194.440 ;
        RECT 108.420 186.640 108.680 186.960 ;
        RECT 106.570 183.725 106.850 184.095 ;
        RECT 106.640 183.560 106.780 183.725 ;
        RECT 108.480 183.560 108.620 186.640 ;
        RECT 106.580 183.240 106.840 183.560 ;
        RECT 108.420 183.240 108.680 183.560 ;
        RECT 106.640 181.520 106.780 183.240 ;
        RECT 107.960 182.900 108.220 183.220 ;
        RECT 107.500 182.560 107.760 182.880 ;
        RECT 107.560 181.520 107.700 182.560 ;
        RECT 108.020 181.520 108.160 182.900 ;
        RECT 108.480 182.735 108.620 183.240 ;
        RECT 108.410 182.365 108.690 182.735 ;
        RECT 108.420 181.540 108.680 181.860 ;
        RECT 106.580 181.200 106.840 181.520 ;
        RECT 107.500 181.200 107.760 181.520 ;
        RECT 107.960 181.200 108.220 181.520 ;
        RECT 107.560 179.140 107.700 181.200 ;
        RECT 107.500 178.820 107.760 179.140 ;
        RECT 107.960 178.820 108.220 179.140 ;
        RECT 106.580 178.370 106.840 178.460 ;
        RECT 106.580 178.230 107.700 178.370 ;
        RECT 106.580 178.140 106.840 178.230 ;
        RECT 107.560 176.615 107.700 178.230 ;
        RECT 107.490 176.245 107.770 176.615 ;
        RECT 107.040 175.760 107.300 176.080 ;
        RECT 107.500 175.760 107.760 176.080 ;
        RECT 106.580 174.400 106.840 174.720 ;
        RECT 106.640 172.420 106.780 174.400 ;
        RECT 107.100 173.020 107.240 175.760 ;
        RECT 107.040 172.700 107.300 173.020 ;
        RECT 106.640 172.280 107.240 172.420 ;
        RECT 106.580 171.680 106.840 172.000 ;
        RECT 106.640 167.240 106.780 171.680 ;
        RECT 107.100 169.135 107.240 172.280 ;
        RECT 107.030 168.765 107.310 169.135 ;
        RECT 107.030 167.405 107.310 167.775 ;
        RECT 106.580 166.920 106.840 167.240 ;
        RECT 106.180 164.630 106.780 164.770 ;
        RECT 106.120 163.860 106.380 164.180 ;
        RECT 106.180 161.120 106.320 163.860 ;
        RECT 106.120 160.800 106.380 161.120 ;
        RECT 106.180 160.100 106.320 160.800 ;
        RECT 106.120 159.780 106.380 160.100 ;
        RECT 105.660 159.100 105.920 159.420 ;
        RECT 105.660 158.080 105.920 158.400 ;
        RECT 105.720 156.700 105.860 158.080 ;
        RECT 105.660 156.380 105.920 156.700 ;
        RECT 105.660 155.360 105.920 155.680 ;
        RECT 105.720 153.980 105.860 155.360 ;
        RECT 106.640 154.175 106.780 164.630 ;
        RECT 107.100 162.820 107.240 167.405 ;
        RECT 107.560 165.540 107.700 175.760 ;
        RECT 108.020 172.000 108.160 178.820 ;
        RECT 107.960 171.680 108.220 172.000 ;
        RECT 108.480 170.640 108.620 181.540 ;
        RECT 108.940 176.080 109.080 194.120 ;
        RECT 108.880 175.760 109.140 176.080 ;
        RECT 108.880 171.680 109.140 172.000 ;
        RECT 108.420 170.320 108.680 170.640 ;
        RECT 108.940 169.960 109.080 171.680 ;
        RECT 108.420 169.640 108.680 169.960 ;
        RECT 108.880 169.640 109.140 169.960 ;
        RECT 108.480 168.260 108.620 169.640 ;
        RECT 107.960 167.940 108.220 168.260 ;
        RECT 108.420 167.940 108.680 168.260 ;
        RECT 108.020 167.240 108.160 167.940 ;
        RECT 108.480 167.580 108.620 167.940 ;
        RECT 108.420 167.260 108.680 167.580 ;
        RECT 107.960 166.920 108.220 167.240 ;
        RECT 109.400 166.980 109.540 210.440 ;
        RECT 110.260 209.760 110.520 210.080 ;
        RECT 110.320 208.380 110.460 209.760 ;
        RECT 112.160 208.380 112.300 211.460 ;
        RECT 112.550 210.245 112.830 210.615 ;
        RECT 112.560 210.100 112.820 210.245 ;
        RECT 113.940 209.760 114.200 210.080 ;
        RECT 110.260 208.060 110.520 208.380 ;
        RECT 112.100 208.060 112.360 208.380 ;
        RECT 112.560 208.060 112.820 208.380 ;
        RECT 110.320 197.160 110.460 208.060 ;
        RECT 112.160 200.900 112.300 208.060 ;
        RECT 112.620 207.215 112.760 208.060 ;
        RECT 114.000 208.040 114.140 209.760 ;
        RECT 114.460 209.060 114.600 215.540 ;
        RECT 118.540 213.840 118.800 214.160 ;
        RECT 117.160 213.500 117.420 213.820 ;
        RECT 115.160 211.945 117.040 212.315 ;
        RECT 117.220 211.180 117.360 213.500 ;
        RECT 117.620 213.160 117.880 213.480 ;
        RECT 114.920 211.040 117.360 211.180 ;
        RECT 114.920 210.760 115.060 211.040 ;
        RECT 115.780 210.780 116.040 211.040 ;
        RECT 114.860 210.440 115.120 210.760 ;
        RECT 117.680 209.060 117.820 213.160 ;
        RECT 118.080 211.460 118.340 211.780 ;
        RECT 114.400 208.740 114.660 209.060 ;
        RECT 117.620 208.740 117.880 209.060 ;
        RECT 113.940 207.720 114.200 208.040 ;
        RECT 112.550 206.845 112.830 207.215 ;
        RECT 117.160 207.040 117.420 207.360 ;
        RECT 117.620 207.040 117.880 207.360 ;
        RECT 115.160 206.505 117.040 206.875 ;
        RECT 117.220 205.320 117.360 207.040 ;
        RECT 117.680 205.660 117.820 207.040 ;
        RECT 117.620 205.340 117.880 205.660 ;
        RECT 113.020 205.000 113.280 205.320 ;
        RECT 117.160 205.000 117.420 205.320 ;
        RECT 113.080 203.620 113.220 205.000 ;
        RECT 115.320 204.660 115.580 204.980 ;
        RECT 113.020 203.300 113.280 203.620 ;
        RECT 115.380 203.280 115.520 204.660 ;
        RECT 115.320 202.960 115.580 203.280 ;
        RECT 117.680 202.260 117.820 205.340 ;
        RECT 117.620 201.940 117.880 202.260 ;
        RECT 112.100 200.580 112.360 200.900 ;
        RECT 112.550 200.725 112.830 201.095 ;
        RECT 115.160 201.065 117.040 201.435 ;
        RECT 110.260 196.840 110.520 197.160 ;
        RECT 110.320 195.120 110.460 196.840 ;
        RECT 110.260 195.030 110.520 195.120 ;
        RECT 109.860 194.890 110.520 195.030 ;
        RECT 109.860 191.720 110.000 194.890 ;
        RECT 110.260 194.800 110.520 194.890 ;
        RECT 110.260 194.120 110.520 194.440 ;
        RECT 110.320 192.060 110.460 194.120 ;
        RECT 110.720 193.440 110.980 193.760 ;
        RECT 110.260 191.740 110.520 192.060 ;
        RECT 109.800 191.400 110.060 191.720 ;
        RECT 110.260 190.720 110.520 191.040 ;
        RECT 109.800 189.700 110.060 190.020 ;
        RECT 109.860 183.900 110.000 189.700 ;
        RECT 110.320 184.095 110.460 190.720 ;
        RECT 110.780 188.910 110.920 193.440 ;
        RECT 112.620 192.740 112.760 200.725 ;
        RECT 113.020 200.240 113.280 200.560 ;
        RECT 113.080 199.200 113.220 200.240 ;
        RECT 114.400 199.900 114.660 200.220 ;
        RECT 113.020 198.880 113.280 199.200 ;
        RECT 113.940 198.880 114.200 199.200 ;
        RECT 113.470 197.325 113.750 197.695 ;
        RECT 114.000 197.500 114.140 198.880 ;
        RECT 114.460 198.180 114.600 199.900 ;
        RECT 114.400 197.860 114.660 198.180 ;
        RECT 112.560 192.420 112.820 192.740 ;
        RECT 113.540 189.340 113.680 197.325 ;
        RECT 113.940 197.180 114.200 197.500 ;
        RECT 117.150 197.325 117.430 197.695 ;
        RECT 114.000 195.460 114.140 197.180 ;
        RECT 115.160 195.625 117.040 195.995 ;
        RECT 113.940 195.140 114.200 195.460 ;
        RECT 114.000 194.780 114.140 195.140 ;
        RECT 115.320 194.800 115.580 195.120 ;
        RECT 113.940 194.460 114.200 194.780 ;
        RECT 115.380 192.740 115.520 194.800 ;
        RECT 117.220 194.780 117.360 197.325 ;
        RECT 117.160 194.460 117.420 194.780 ;
        RECT 115.320 192.420 115.580 192.740 ;
        RECT 113.940 191.400 114.200 191.720 ;
        RECT 114.400 191.400 114.660 191.720 ;
        RECT 117.160 191.400 117.420 191.720 ;
        RECT 113.480 189.020 113.740 189.340 ;
        RECT 111.180 188.910 111.440 189.000 ;
        RECT 110.780 188.770 111.440 188.910 ;
        RECT 111.180 188.680 111.440 188.770 ;
        RECT 111.240 186.280 111.380 188.680 ;
        RECT 114.000 188.320 114.140 191.400 ;
        RECT 114.460 189.000 114.600 191.400 ;
        RECT 115.160 190.185 117.040 190.555 ;
        RECT 117.220 190.020 117.360 191.400 ;
        RECT 117.610 191.205 117.890 191.575 ;
        RECT 117.160 189.700 117.420 190.020 ;
        RECT 117.680 189.340 117.820 191.205 ;
        RECT 116.700 189.020 116.960 189.340 ;
        RECT 117.620 189.020 117.880 189.340 ;
        RECT 114.400 188.680 114.660 189.000 ;
        RECT 116.240 188.680 116.500 189.000 ;
        RECT 113.940 188.000 114.200 188.320 ;
        RECT 113.020 186.300 113.280 186.620 ;
        RECT 111.180 185.960 111.440 186.280 ;
        RECT 111.240 184.580 111.380 185.960 ;
        RECT 111.640 185.620 111.900 185.940 ;
        RECT 110.720 184.260 110.980 184.580 ;
        RECT 111.180 184.260 111.440 184.580 ;
        RECT 109.800 183.580 110.060 183.900 ;
        RECT 110.250 183.725 110.530 184.095 ;
        RECT 110.320 181.180 110.460 183.725 ;
        RECT 110.780 181.375 110.920 184.260 ;
        RECT 110.260 180.860 110.520 181.180 ;
        RECT 110.710 181.005 110.990 181.375 ;
        RECT 110.720 180.520 110.980 180.840 ;
        RECT 109.800 179.840 110.060 180.160 ;
        RECT 109.860 178.460 110.000 179.840 ;
        RECT 109.800 178.370 110.060 178.460 ;
        RECT 109.800 178.230 110.460 178.370 ;
        RECT 109.800 178.140 110.060 178.230 ;
        RECT 109.790 174.885 110.070 175.255 ;
        RECT 109.860 170.300 110.000 174.885 ;
        RECT 109.800 169.980 110.060 170.300 ;
        RECT 108.480 166.840 109.540 166.980 ;
        RECT 107.500 165.220 107.760 165.540 ;
        RECT 107.500 163.860 107.760 164.180 ;
        RECT 107.040 162.500 107.300 162.820 ;
        RECT 107.560 161.460 107.700 163.860 ;
        RECT 107.960 163.520 108.220 163.840 ;
        RECT 107.500 161.140 107.760 161.460 ;
        RECT 107.500 158.080 107.760 158.400 ;
        RECT 107.040 154.340 107.300 154.660 ;
        RECT 105.660 153.660 105.920 153.980 ;
        RECT 106.120 153.890 106.380 153.980 ;
        RECT 106.570 153.890 106.850 154.175 ;
        RECT 106.120 153.805 106.850 153.890 ;
        RECT 106.120 153.750 106.780 153.805 ;
        RECT 106.120 153.660 106.380 153.750 ;
        RECT 105.260 152.420 106.780 152.560 ;
        RECT 104.740 151.620 105.000 151.940 ;
        RECT 106.120 150.600 106.380 150.920 ;
        RECT 106.180 147.860 106.320 150.600 ;
        RECT 106.120 147.540 106.380 147.860 ;
        RECT 106.640 147.520 106.780 152.420 ;
        RECT 106.580 147.200 106.840 147.520 ;
        RECT 107.100 145.820 107.240 154.340 ;
        RECT 107.560 153.980 107.700 158.080 ;
        RECT 108.020 157.380 108.160 163.520 ;
        RECT 107.960 157.060 108.220 157.380 ;
        RECT 107.500 153.660 107.760 153.980 ;
        RECT 107.490 153.125 107.770 153.495 ;
        RECT 107.500 152.980 107.760 153.125 ;
        RECT 108.480 150.240 108.620 166.840 ;
        RECT 109.340 166.240 109.600 166.560 ;
        RECT 109.400 164.520 109.540 166.240 ;
        RECT 110.320 164.860 110.460 178.230 ;
        RECT 110.780 178.120 110.920 180.520 ;
        RECT 110.720 177.800 110.980 178.120 ;
        RECT 110.720 177.120 110.980 177.440 ;
        RECT 110.780 175.740 110.920 177.120 ;
        RECT 110.720 175.420 110.980 175.740 ;
        RECT 111.240 167.580 111.380 184.260 ;
        RECT 111.700 180.015 111.840 185.620 ;
        RECT 112.560 185.280 112.820 185.600 ;
        RECT 112.100 182.560 112.360 182.880 ;
        RECT 111.630 179.645 111.910 180.015 ;
        RECT 111.700 176.420 111.840 179.645 ;
        RECT 111.640 176.100 111.900 176.420 ;
        RECT 111.640 173.040 111.900 173.360 ;
        RECT 111.180 167.260 111.440 167.580 ;
        RECT 111.180 165.220 111.440 165.540 ;
        RECT 110.260 164.540 110.520 164.860 ;
        RECT 110.710 164.685 110.990 165.055 ;
        RECT 110.720 164.540 110.980 164.685 ;
        RECT 109.340 164.430 109.600 164.520 ;
        RECT 109.340 164.290 110.000 164.430 ;
        RECT 109.340 164.200 109.600 164.290 ;
        RECT 109.340 163.520 109.600 163.840 ;
        RECT 108.880 161.820 109.140 162.140 ;
        RECT 108.940 160.100 109.080 161.820 ;
        RECT 109.400 160.180 109.540 163.520 ;
        RECT 109.860 161.800 110.000 164.290 ;
        RECT 110.320 162.140 110.460 164.540 ;
        RECT 110.260 161.820 110.520 162.140 ;
        RECT 109.800 161.480 110.060 161.800 ;
        RECT 108.880 159.780 109.140 160.100 ;
        RECT 109.400 160.040 110.000 160.180 ;
        RECT 108.880 158.420 109.140 158.740 ;
        RECT 108.420 149.920 108.680 150.240 ;
        RECT 107.950 149.045 108.230 149.415 ;
        RECT 108.020 145.820 108.160 149.045 ;
        RECT 108.480 148.540 108.620 149.920 ;
        RECT 108.420 148.220 108.680 148.540 ;
        RECT 108.940 147.940 109.080 158.420 ;
        RECT 109.860 156.700 110.000 160.040 ;
        RECT 110.320 159.760 110.460 161.820 ;
        RECT 110.780 161.655 110.920 164.540 ;
        RECT 111.240 162.140 111.380 165.220 ;
        RECT 111.700 164.520 111.840 173.040 ;
        RECT 112.160 167.920 112.300 182.560 ;
        RECT 112.620 181.860 112.760 185.280 ;
        RECT 113.080 182.880 113.220 186.300 ;
        RECT 113.020 182.560 113.280 182.880 ;
        RECT 112.560 181.540 112.820 181.860 ;
        RECT 112.620 175.740 112.760 181.540 ;
        RECT 113.080 180.070 113.220 182.560 ;
        RECT 113.470 182.365 113.750 182.735 ;
        RECT 113.540 180.840 113.680 182.365 ;
        RECT 113.480 180.520 113.740 180.840 ;
        RECT 113.080 179.930 113.680 180.070 ;
        RECT 112.560 175.420 112.820 175.740 ;
        RECT 113.010 170.805 113.290 171.175 ;
        RECT 113.080 169.620 113.220 170.805 ;
        RECT 113.020 169.300 113.280 169.620 ;
        RECT 113.080 168.260 113.220 169.300 ;
        RECT 113.020 167.940 113.280 168.260 ;
        RECT 112.100 167.600 112.360 167.920 ;
        RECT 112.160 165.540 112.300 167.600 ;
        RECT 113.010 166.045 113.290 166.415 ;
        RECT 112.100 165.220 112.360 165.540 ;
        RECT 113.080 164.860 113.220 166.045 ;
        RECT 113.540 164.860 113.680 179.930 ;
        RECT 114.000 173.360 114.140 188.000 ;
        RECT 116.300 187.060 116.440 188.680 ;
        RECT 114.460 186.920 116.440 187.060 ;
        RECT 114.460 184.490 114.600 186.920 ;
        RECT 116.760 186.280 116.900 189.020 ;
        RECT 117.160 188.000 117.420 188.320 ;
        RECT 117.220 187.300 117.360 188.000 ;
        RECT 117.160 186.980 117.420 187.300 ;
        RECT 116.700 186.135 116.960 186.280 ;
        RECT 116.690 185.765 116.970 186.135 ;
        RECT 117.620 185.620 117.880 185.940 ;
        RECT 117.160 185.280 117.420 185.600 ;
        RECT 115.160 184.745 117.040 185.115 ;
        RECT 114.460 184.350 115.060 184.490 ;
        RECT 114.920 180.070 115.060 184.350 ;
        RECT 117.220 184.240 117.360 185.280 ;
        RECT 117.160 183.920 117.420 184.240 ;
        RECT 116.700 182.560 116.960 182.880 ;
        RECT 116.760 180.840 116.900 182.560 ;
        RECT 117.160 181.540 117.420 181.860 ;
        RECT 116.240 180.695 116.500 180.840 ;
        RECT 116.230 180.325 116.510 180.695 ;
        RECT 116.700 180.520 116.960 180.840 ;
        RECT 117.220 180.580 117.360 181.540 ;
        RECT 117.680 181.180 117.820 185.620 ;
        RECT 117.620 180.860 117.880 181.180 ;
        RECT 117.220 180.440 117.820 180.580 ;
        RECT 114.920 179.930 117.360 180.070 ;
        RECT 115.160 179.305 117.040 179.675 ;
        RECT 117.220 178.120 117.360 179.930 ;
        RECT 117.160 177.800 117.420 178.120 ;
        RECT 117.160 177.120 117.420 177.440 ;
        RECT 117.220 175.740 117.360 177.120 ;
        RECT 117.160 175.420 117.420 175.740 ;
        RECT 114.390 173.525 114.670 173.895 ;
        RECT 115.160 173.865 117.040 174.235 ;
        RECT 117.220 173.700 117.360 175.420 ;
        RECT 117.680 175.400 117.820 180.440 ;
        RECT 117.620 175.080 117.880 175.400 ;
        RECT 113.940 173.040 114.200 173.360 ;
        RECT 113.940 168.960 114.200 169.280 ;
        RECT 113.020 164.540 113.280 164.860 ;
        RECT 113.480 164.540 113.740 164.860 ;
        RECT 111.640 164.200 111.900 164.520 ;
        RECT 111.640 163.750 111.900 163.840 ;
        RECT 111.640 163.610 112.760 163.750 ;
        RECT 111.640 163.520 111.900 163.610 ;
        RECT 111.180 162.050 111.440 162.140 ;
        RECT 111.180 161.910 111.840 162.050 ;
        RECT 111.180 161.820 111.440 161.910 ;
        RECT 110.710 161.285 110.990 161.655 ;
        RECT 110.260 159.440 110.520 159.760 ;
        RECT 110.260 158.760 110.520 159.080 ;
        RECT 111.180 158.990 111.440 159.080 ;
        RECT 111.700 158.990 111.840 161.910 ;
        RECT 112.100 161.820 112.360 162.140 ;
        RECT 111.180 158.850 111.840 158.990 ;
        RECT 111.180 158.760 111.440 158.850 ;
        RECT 110.320 157.380 110.460 158.760 ;
        RECT 110.260 157.060 110.520 157.380 ;
        RECT 112.160 156.700 112.300 161.820 ;
        RECT 109.800 156.380 110.060 156.700 ;
        RECT 112.100 156.380 112.360 156.700 ;
        RECT 109.340 156.040 109.600 156.360 ;
        RECT 109.400 151.940 109.540 156.040 ;
        RECT 110.720 155.700 110.980 156.020 ;
        RECT 110.780 153.640 110.920 155.700 ;
        RECT 111.180 155.535 111.440 155.680 ;
        RECT 111.170 155.165 111.450 155.535 ;
        RECT 112.100 155.360 112.360 155.680 ;
        RECT 111.240 153.640 111.380 155.165 ;
        RECT 112.160 154.660 112.300 155.360 ;
        RECT 112.100 154.340 112.360 154.660 ;
        RECT 112.090 153.805 112.370 154.175 ;
        RECT 110.720 153.320 110.980 153.640 ;
        RECT 111.180 153.550 111.440 153.640 ;
        RECT 111.180 153.410 111.840 153.550 ;
        RECT 111.180 153.320 111.440 153.410 ;
        RECT 111.180 152.640 111.440 152.960 ;
        RECT 109.340 151.620 109.600 151.940 ;
        RECT 110.720 150.600 110.980 150.920 ;
        RECT 110.780 148.540 110.920 150.600 ;
        RECT 110.720 148.220 110.980 148.540 ;
        RECT 108.940 147.860 110.000 147.940 ;
        RECT 108.940 147.800 110.060 147.860 ;
        RECT 109.800 147.540 110.060 147.800 ;
        RECT 108.420 147.200 108.680 147.520 ;
        RECT 109.340 147.200 109.600 147.520 ;
        RECT 110.260 147.200 110.520 147.520 ;
        RECT 110.720 147.200 110.980 147.520 ;
        RECT 102.440 145.500 102.700 145.820 ;
        RECT 103.820 145.500 104.080 145.820 ;
        RECT 107.040 145.500 107.300 145.820 ;
        RECT 107.960 145.500 108.220 145.820 ;
        RECT 100.600 144.570 101.260 144.710 ;
        RECT 100.600 144.480 100.860 144.570 ;
        RECT 102.440 144.480 102.700 144.800 ;
        RECT 105.200 144.480 105.460 144.800 ;
        RECT 98.360 143.780 98.500 144.480 ;
        RECT 100.160 143.945 102.040 144.315 ;
        RECT 98.300 143.460 98.560 143.780 ;
        RECT 102.500 142.760 102.640 144.480 ;
        RECT 105.260 143.780 105.400 144.480 ;
        RECT 108.480 143.780 108.620 147.200 ;
        RECT 109.400 145.820 109.540 147.200 ;
        RECT 109.340 145.500 109.600 145.820 ;
        RECT 108.880 144.480 109.140 144.800 ;
        RECT 105.200 143.460 105.460 143.780 ;
        RECT 108.420 143.460 108.680 143.780 ;
        RECT 108.940 142.760 109.080 144.480 ;
        RECT 102.440 142.440 102.700 142.760 ;
        RECT 108.880 142.440 109.140 142.760 ;
        RECT 99.680 141.760 99.940 142.080 ;
        RECT 104.740 141.760 105.000 142.080 ;
        RECT 99.740 140.690 99.880 141.760 ;
        RECT 104.800 141.140 104.940 141.760 ;
        RECT 103.880 141.000 104.940 141.140 ;
        RECT 103.880 140.690 104.020 141.000 ;
        RECT 96.920 139.720 97.180 140.040 ;
        RECT 64.900 131.300 65.960 132.300 ;
        RECT 74.800 132.160 75.140 132.440 ;
        RECT 78.940 132.160 79.280 132.440 ;
        RECT 83.080 132.160 83.420 132.440 ;
        RECT 87.220 132.160 87.560 132.440 ;
        RECT 91.360 132.160 91.700 132.440 ;
        RECT 95.500 132.160 95.840 132.440 ;
        RECT 99.670 132.130 99.950 140.690 ;
        RECT 101.580 132.400 102.580 134.445 ;
        RECT 101.550 131.400 102.610 132.400 ;
        RECT 103.810 132.130 104.090 140.690 ;
        RECT 110.320 140.380 110.460 147.200 ;
        RECT 110.780 146.500 110.920 147.200 ;
        RECT 110.720 146.180 110.980 146.500 ;
        RECT 111.240 145.820 111.380 152.640 ;
        RECT 111.700 151.600 111.840 153.410 ;
        RECT 111.640 151.280 111.900 151.600 ;
        RECT 112.160 150.660 112.300 153.805 ;
        RECT 111.700 150.520 112.300 150.660 ;
        RECT 111.700 149.415 111.840 150.520 ;
        RECT 112.100 149.920 112.360 150.240 ;
        RECT 111.630 149.045 111.910 149.415 ;
        RECT 111.630 146.325 111.910 146.695 ;
        RECT 111.640 146.180 111.900 146.325 ;
        RECT 112.160 145.820 112.300 149.920 ;
        RECT 112.620 148.200 112.760 163.610 ;
        RECT 113.020 162.160 113.280 162.480 ;
        RECT 113.080 159.420 113.220 162.160 ;
        RECT 113.470 161.285 113.750 161.655 ;
        RECT 113.540 159.420 113.680 161.285 ;
        RECT 113.020 159.100 113.280 159.420 ;
        RECT 113.480 159.100 113.740 159.420 ;
        RECT 113.480 156.380 113.740 156.700 ;
        RECT 113.540 153.980 113.680 156.380 ;
        RECT 113.480 153.660 113.740 153.980 ;
        RECT 113.020 152.700 113.280 152.960 ;
        RECT 113.020 152.640 113.680 152.700 ;
        RECT 113.080 152.560 113.680 152.640 ;
        RECT 113.010 149.725 113.290 150.095 ;
        RECT 113.080 148.200 113.220 149.725 ;
        RECT 112.560 147.880 112.820 148.200 ;
        RECT 113.020 147.880 113.280 148.200 ;
        RECT 113.080 145.820 113.220 147.880 ;
        RECT 111.180 145.500 111.440 145.820 ;
        RECT 112.100 145.500 112.360 145.820 ;
        RECT 113.020 145.500 113.280 145.820 ;
        RECT 113.080 145.220 113.220 145.500 ;
        RECT 112.100 144.820 112.360 145.140 ;
        RECT 112.620 145.080 113.220 145.220 ;
        RECT 112.160 143.780 112.300 144.820 ;
        RECT 112.100 143.460 112.360 143.780 ;
        RECT 112.620 142.760 112.760 145.080 ;
        RECT 113.020 144.480 113.280 144.800 ;
        RECT 113.080 143.780 113.220 144.480 ;
        RECT 113.540 143.780 113.680 152.560 ;
        RECT 114.000 150.660 114.140 168.960 ;
        RECT 114.460 165.540 114.600 173.525 ;
        RECT 117.160 173.380 117.420 173.700 ;
        RECT 117.680 169.960 117.820 175.080 ;
        RECT 117.620 169.640 117.880 169.960 ;
        RECT 115.160 168.425 117.040 168.795 ;
        RECT 117.620 167.260 117.880 167.580 ;
        RECT 117.680 166.560 117.820 167.260 ;
        RECT 117.620 166.240 117.880 166.560 ;
        RECT 118.140 166.415 118.280 211.460 ;
        RECT 118.600 210.760 118.740 213.840 ;
        RECT 118.540 210.440 118.800 210.760 ;
        RECT 118.600 208.380 118.740 210.440 ;
        RECT 118.990 210.245 119.270 210.615 ;
        RECT 119.000 210.100 119.260 210.245 ;
        RECT 118.540 208.060 118.800 208.380 ;
        RECT 119.520 202.600 119.660 215.540 ;
        RECT 119.920 213.840 120.180 214.160 ;
        RECT 119.980 207.360 120.120 213.840 ;
        RECT 121.820 213.480 121.960 216.690 ;
        RECT 123.600 215.200 123.860 215.520 ;
        RECT 121.760 213.160 122.020 213.480 ;
        RECT 123.660 211.780 123.800 215.200 ;
        RECT 125.500 213.480 125.640 216.690 ;
        RECT 126.360 214.180 126.620 214.500 ;
        RECT 125.440 213.160 125.700 213.480 ;
        RECT 124.520 212.820 124.780 213.140 ;
        RECT 123.600 211.460 123.860 211.780 ;
        RECT 120.380 211.120 120.640 211.440 ;
        RECT 119.920 207.040 120.180 207.360 ;
        RECT 119.460 202.280 119.720 202.600 ;
        RECT 119.000 197.180 119.260 197.500 ;
        RECT 119.060 192.255 119.200 197.180 ;
        RECT 119.520 197.160 119.660 202.280 ;
        RECT 119.920 201.600 120.180 201.920 ;
        RECT 119.460 196.840 119.720 197.160 ;
        RECT 118.990 192.140 119.270 192.255 ;
        RECT 118.540 191.740 118.800 192.060 ;
        RECT 118.990 192.000 119.660 192.140 ;
        RECT 118.990 191.885 119.270 192.000 ;
        RECT 118.600 187.300 118.740 191.740 ;
        RECT 119.000 191.400 119.260 191.720 ;
        RECT 119.060 190.020 119.200 191.400 ;
        RECT 119.520 191.040 119.660 192.000 ;
        RECT 119.460 190.720 119.720 191.040 ;
        RECT 119.000 189.700 119.260 190.020 ;
        RECT 119.980 189.420 120.120 201.600 ;
        RECT 120.440 200.900 120.580 211.120 ;
        RECT 121.300 210.780 121.560 211.100 ;
        RECT 123.130 210.925 123.410 211.295 ;
        RECT 124.580 211.100 124.720 212.820 ;
        RECT 125.900 212.480 126.160 212.800 ;
        RECT 125.440 211.460 125.700 211.780 ;
        RECT 120.840 210.100 121.100 210.420 ;
        RECT 120.900 206.340 121.040 210.100 ;
        RECT 121.360 209.060 121.500 210.780 ;
        RECT 123.200 210.760 123.340 210.925 ;
        RECT 124.520 210.780 124.780 211.100 ;
        RECT 123.140 210.440 123.400 210.760 ;
        RECT 122.680 209.760 122.940 210.080 ;
        RECT 122.740 209.060 122.880 209.760 ;
        RECT 125.500 209.060 125.640 211.460 ;
        RECT 121.300 208.740 121.560 209.060 ;
        RECT 122.680 208.970 122.940 209.060 ;
        RECT 122.280 208.830 122.940 208.970 ;
        RECT 122.280 206.340 122.420 208.830 ;
        RECT 122.680 208.740 122.940 208.830 ;
        RECT 125.440 208.740 125.700 209.060 ;
        RECT 122.680 207.720 122.940 208.040 ;
        RECT 120.840 206.020 121.100 206.340 ;
        RECT 122.220 206.020 122.480 206.340 ;
        RECT 121.300 204.320 121.560 204.640 ;
        RECT 121.360 203.620 121.500 204.320 ;
        RECT 121.300 203.300 121.560 203.620 ;
        RECT 120.380 200.580 120.640 200.900 ;
        RECT 120.370 199.365 120.650 199.735 ;
        RECT 120.440 198.180 120.580 199.365 ;
        RECT 121.300 199.220 121.560 199.540 ;
        RECT 120.380 197.860 120.640 198.180 ;
        RECT 120.440 189.930 120.580 197.860 ;
        RECT 121.360 194.780 121.500 199.220 ;
        RECT 121.300 194.460 121.560 194.780 ;
        RECT 121.360 191.720 121.500 194.460 ;
        RECT 122.220 193.440 122.480 193.760 ;
        RECT 121.300 191.400 121.560 191.720 ;
        RECT 120.440 189.790 121.960 189.930 ;
        RECT 119.980 189.280 120.580 189.420 ;
        RECT 119.920 188.680 120.180 189.000 ;
        RECT 118.540 186.980 118.800 187.300 ;
        RECT 118.600 179.140 118.740 186.980 ;
        RECT 119.460 185.280 119.720 185.600 ;
        RECT 119.520 183.560 119.660 185.280 ;
        RECT 119.460 183.240 119.720 183.560 ;
        RECT 119.450 181.685 119.730 182.055 ;
        RECT 119.980 181.860 120.120 188.680 ;
        RECT 119.460 181.540 119.720 181.685 ;
        RECT 119.920 181.540 120.180 181.860 ;
        RECT 119.910 181.005 120.190 181.375 ;
        RECT 119.980 180.840 120.120 181.005 ;
        RECT 119.920 180.520 120.180 180.840 ;
        RECT 118.540 178.820 118.800 179.140 ;
        RECT 119.000 177.120 119.260 177.440 ;
        RECT 118.540 174.400 118.800 174.720 ;
        RECT 118.600 173.700 118.740 174.400 ;
        RECT 118.540 173.380 118.800 173.700 ;
        RECT 118.540 167.940 118.800 168.260 ;
        RECT 118.600 167.580 118.740 167.940 ;
        RECT 118.540 167.260 118.800 167.580 ;
        RECT 118.070 166.045 118.350 166.415 ;
        RECT 114.400 165.220 114.660 165.540 ;
        RECT 114.400 164.540 114.660 164.860 ;
        RECT 114.460 162.480 114.600 164.540 ;
        RECT 118.070 164.005 118.350 164.375 ;
        RECT 118.540 164.200 118.800 164.520 ;
        RECT 117.620 163.520 117.880 163.840 ;
        RECT 115.160 162.985 117.040 163.355 ;
        RECT 117.680 162.820 117.820 163.520 ;
        RECT 117.620 162.500 117.880 162.820 ;
        RECT 114.400 162.160 114.660 162.480 ;
        RECT 115.320 161.140 115.580 161.460 ;
        RECT 114.400 160.800 114.660 161.120 ;
        RECT 114.460 159.080 114.600 160.800 ;
        RECT 115.380 159.420 115.520 161.140 ;
        RECT 115.320 159.100 115.580 159.420 ;
        RECT 114.400 158.760 114.660 159.080 ;
        RECT 114.860 158.310 115.120 158.400 ;
        RECT 114.460 158.170 115.120 158.310 ;
        RECT 114.460 156.100 114.600 158.170 ;
        RECT 114.860 158.080 115.120 158.170 ;
        RECT 117.160 158.080 117.420 158.400 ;
        RECT 115.160 157.545 117.040 157.915 ;
        RECT 117.220 157.040 117.360 158.080 ;
        RECT 117.160 156.720 117.420 157.040 ;
        RECT 115.320 156.380 115.580 156.700 ;
        RECT 114.460 155.960 115.060 156.100 ;
        RECT 114.400 155.360 114.660 155.680 ;
        RECT 114.460 154.660 114.600 155.360 ;
        RECT 114.920 154.660 115.060 155.960 ;
        RECT 115.380 155.535 115.520 156.380 ;
        RECT 116.230 155.845 116.510 156.215 ;
        RECT 115.310 155.165 115.590 155.535 ;
        RECT 114.400 154.340 114.660 154.660 ;
        RECT 114.860 154.340 115.120 154.660 ;
        RECT 114.390 153.890 114.670 154.175 ;
        RECT 114.860 153.890 115.120 153.980 ;
        RECT 114.390 153.805 115.120 153.890 ;
        RECT 114.460 153.750 115.120 153.805 ;
        RECT 114.860 153.660 115.120 153.750 ;
        RECT 116.300 153.640 116.440 155.845 ;
        RECT 117.620 155.700 117.880 156.020 ;
        RECT 116.240 153.320 116.500 153.640 ;
        RECT 117.160 152.980 117.420 153.300 ;
        RECT 114.400 152.640 114.660 152.960 ;
        RECT 114.460 151.260 114.600 152.640 ;
        RECT 115.160 152.105 117.040 152.475 ;
        RECT 114.400 150.940 114.660 151.260 ;
        RECT 116.700 151.170 116.960 151.260 ;
        RECT 117.220 151.170 117.360 152.980 ;
        RECT 117.680 151.600 117.820 155.700 ;
        RECT 117.620 151.280 117.880 151.600 ;
        RECT 116.700 151.030 117.360 151.170 ;
        RECT 116.700 150.940 116.960 151.030 ;
        RECT 114.000 150.520 114.600 150.660 ;
        RECT 113.930 149.045 114.210 149.415 ;
        RECT 114.000 148.540 114.140 149.045 ;
        RECT 113.940 148.220 114.200 148.540 ;
        RECT 114.460 145.820 114.600 150.520 ;
        RECT 117.220 148.200 117.360 151.030 ;
        RECT 117.160 147.880 117.420 148.200 ;
        RECT 115.160 146.665 117.040 147.035 ;
        RECT 114.400 145.500 114.660 145.820 ;
        RECT 115.310 145.645 115.590 146.015 ;
        RECT 117.160 145.730 117.420 145.820 ;
        RECT 118.140 145.730 118.280 164.005 ;
        RECT 118.600 162.335 118.740 164.200 ;
        RECT 118.530 161.965 118.810 162.335 ;
        RECT 118.540 153.320 118.800 153.640 ;
        RECT 118.600 151.260 118.740 153.320 ;
        RECT 118.540 150.940 118.800 151.260 ;
        RECT 118.540 149.920 118.800 150.240 ;
        RECT 118.600 148.540 118.740 149.920 ;
        RECT 119.060 148.735 119.200 177.120 ;
        RECT 120.440 176.500 120.580 189.280 ;
        RECT 120.840 189.020 121.100 189.340 ;
        RECT 120.900 178.800 121.040 189.020 ;
        RECT 121.820 187.300 121.960 189.790 ;
        RECT 122.280 189.340 122.420 193.440 ;
        RECT 122.220 189.020 122.480 189.340 ;
        RECT 121.760 186.980 122.020 187.300 ;
        RECT 121.820 185.600 121.960 186.980 ;
        RECT 122.280 186.700 122.420 189.020 ;
        RECT 122.740 187.060 122.880 207.720 ;
        RECT 125.960 206.340 126.100 212.480 ;
        RECT 126.420 211.100 126.560 214.180 ;
        RECT 129.180 213.480 129.320 216.690 ;
        RECT 130.160 214.665 132.040 215.035 ;
        RECT 134.240 213.480 134.380 217.160 ;
        RECT 136.470 216.940 136.770 221.040 ;
        RECT 140.150 216.940 140.450 221.040 ;
        RECT 143.830 216.940 144.130 221.040 ;
        RECT 147.510 216.940 147.810 221.040 ;
        RECT 136.470 216.690 136.750 216.940 ;
        RECT 140.150 216.690 140.430 216.940 ;
        RECT 143.830 216.690 144.110 216.940 ;
        RECT 147.510 216.690 147.790 216.940 ;
        RECT 136.540 213.480 136.680 216.690 ;
        RECT 140.220 213.480 140.360 216.690 ;
        RECT 143.900 213.480 144.040 216.690 ;
        RECT 144.760 215.200 145.020 215.520 ;
        RECT 144.820 214.160 144.960 215.200 ;
        RECT 144.760 213.840 145.020 214.160 ;
        RECT 147.580 213.480 147.720 216.690 ;
        RECT 129.120 213.160 129.380 213.480 ;
        RECT 133.720 213.160 133.980 213.480 ;
        RECT 134.180 213.160 134.440 213.480 ;
        RECT 136.480 213.160 136.740 213.480 ;
        RECT 140.160 213.160 140.420 213.480 ;
        RECT 140.620 213.160 140.880 213.480 ;
        RECT 143.840 213.160 144.100 213.480 ;
        RECT 147.520 213.160 147.780 213.480 ;
        RECT 127.740 212.480 128.000 212.800 ;
        RECT 129.580 212.480 129.840 212.800 ;
        RECT 133.260 212.480 133.520 212.800 ;
        RECT 127.800 211.295 127.940 212.480 ;
        RECT 129.640 211.780 129.780 212.480 ;
        RECT 129.580 211.460 129.840 211.780 ;
        RECT 126.360 210.780 126.620 211.100 ;
        RECT 127.730 210.925 128.010 211.295 ;
        RECT 133.320 211.100 133.460 212.480 ;
        RECT 126.420 210.500 126.560 210.780 ;
        RECT 126.420 210.360 127.020 210.500 ;
        RECT 127.280 210.440 127.540 210.760 ;
        RECT 126.360 209.760 126.620 210.080 ;
        RECT 126.420 209.060 126.560 209.760 ;
        RECT 126.360 208.740 126.620 209.060 ;
        RECT 126.420 208.575 126.560 208.740 ;
        RECT 126.350 208.205 126.630 208.575 ;
        RECT 126.880 208.040 127.020 210.360 ;
        RECT 126.350 207.780 126.630 207.895 ;
        RECT 126.820 207.780 127.080 208.040 ;
        RECT 126.350 207.720 127.080 207.780 ;
        RECT 126.350 207.640 127.020 207.720 ;
        RECT 126.350 207.525 126.630 207.640 ;
        RECT 126.820 207.040 127.080 207.360 ;
        RECT 126.880 206.340 127.020 207.040 ;
        RECT 123.600 206.020 123.860 206.340 ;
        RECT 125.440 206.020 125.700 206.340 ;
        RECT 125.900 206.020 126.160 206.340 ;
        RECT 126.820 206.020 127.080 206.340 ;
        RECT 123.140 205.680 123.400 206.000 ;
        RECT 123.200 200.860 123.340 205.680 ;
        RECT 123.660 202.940 123.800 206.020 ;
        RECT 125.500 205.320 125.640 206.020 ;
        RECT 125.960 205.660 126.100 206.020 ;
        RECT 125.900 205.340 126.160 205.660 ;
        RECT 124.980 205.000 125.240 205.320 ;
        RECT 125.440 205.000 125.700 205.320 ;
        RECT 125.040 202.940 125.180 205.000 ;
        RECT 127.340 202.940 127.480 210.440 ;
        RECT 127.800 210.420 127.940 210.925 ;
        RECT 133.260 210.780 133.520 211.100 ;
        RECT 127.740 210.100 128.000 210.420 ;
        RECT 130.160 209.225 132.040 209.595 ;
        RECT 133.780 209.060 133.920 213.160 ;
        RECT 134.180 212.480 134.440 212.800 ;
        RECT 133.720 208.740 133.980 209.060 ;
        RECT 129.120 208.060 129.380 208.380 ;
        RECT 133.710 208.205 133.990 208.575 ;
        RECT 128.200 207.720 128.460 208.040 ;
        RECT 127.730 205.740 128.010 205.855 ;
        RECT 128.260 205.740 128.400 207.720 ;
        RECT 129.180 206.340 129.320 208.060 ;
        RECT 129.120 206.020 129.380 206.340 ;
        RECT 127.730 205.600 128.400 205.740 ;
        RECT 127.730 205.485 128.010 205.600 ;
        RECT 132.340 205.340 132.600 205.660 ;
        RECT 130.160 203.785 132.040 204.155 ;
        RECT 123.600 202.620 123.860 202.940 ;
        RECT 124.980 202.620 125.240 202.940 ;
        RECT 127.280 202.620 127.540 202.940 ;
        RECT 132.400 202.600 132.540 205.340 ;
        RECT 132.340 202.280 132.600 202.600 ;
        RECT 132.800 201.940 133.060 202.260 ;
        RECT 133.260 201.940 133.520 202.260 ;
        RECT 127.280 201.600 127.540 201.920 ;
        RECT 127.340 200.860 127.480 201.600 ;
        RECT 123.200 200.720 123.800 200.860 ;
        RECT 127.340 200.720 128.400 200.860 ;
        RECT 123.140 196.840 123.400 197.160 ;
        RECT 123.200 194.440 123.340 196.840 ;
        RECT 123.140 194.295 123.400 194.440 ;
        RECT 123.130 193.925 123.410 194.295 ;
        RECT 122.740 186.920 123.340 187.060 ;
        RECT 122.280 186.560 122.880 186.700 ;
        RECT 122.740 186.280 122.880 186.560 ;
        RECT 122.210 185.765 122.490 186.135 ;
        RECT 122.680 185.960 122.940 186.280 ;
        RECT 122.280 185.600 122.420 185.765 ;
        RECT 121.760 185.280 122.020 185.600 ;
        RECT 122.220 185.280 122.480 185.600 ;
        RECT 122.280 184.580 122.420 185.280 ;
        RECT 122.220 184.260 122.480 184.580 ;
        RECT 121.300 183.920 121.560 184.240 ;
        RECT 122.680 183.920 122.940 184.240 ;
        RECT 121.360 181.860 121.500 183.920 ;
        RECT 121.760 182.560 122.020 182.880 ;
        RECT 122.220 182.560 122.480 182.880 ;
        RECT 121.300 181.540 121.560 181.860 ;
        RECT 121.820 180.840 121.960 182.560 ;
        RECT 122.280 182.055 122.420 182.560 ;
        RECT 122.210 181.685 122.490 182.055 ;
        RECT 122.210 181.005 122.490 181.375 ;
        RECT 121.760 180.520 122.020 180.840 ;
        RECT 121.300 179.840 121.560 180.160 ;
        RECT 120.840 178.655 121.100 178.800 ;
        RECT 120.830 178.285 121.110 178.655 ;
        RECT 120.440 176.360 121.040 176.500 ;
        RECT 120.380 175.935 120.640 176.080 ;
        RECT 120.370 175.565 120.650 175.935 ;
        RECT 119.460 174.400 119.720 174.720 ;
        RECT 119.520 172.680 119.660 174.400 ;
        RECT 120.380 173.380 120.640 173.700 ;
        RECT 119.910 172.845 120.190 173.215 ;
        RECT 119.460 172.360 119.720 172.680 ;
        RECT 119.460 167.600 119.720 167.920 ;
        RECT 119.520 166.900 119.660 167.600 ;
        RECT 119.460 166.580 119.720 166.900 ;
        RECT 119.520 164.860 119.660 166.580 ;
        RECT 119.460 164.540 119.720 164.860 ;
        RECT 119.460 161.820 119.720 162.140 ;
        RECT 119.520 156.700 119.660 161.820 ;
        RECT 119.460 156.380 119.720 156.700 ;
        RECT 119.980 156.100 120.120 172.845 ;
        RECT 119.520 155.960 120.120 156.100 ;
        RECT 118.540 148.220 118.800 148.540 ;
        RECT 118.990 148.365 119.270 148.735 ;
        RECT 119.060 146.500 119.200 148.365 ;
        RECT 119.000 146.180 119.260 146.500 ;
        RECT 119.520 145.820 119.660 155.960 ;
        RECT 119.920 155.360 120.180 155.680 ;
        RECT 119.980 154.660 120.120 155.360 ;
        RECT 119.920 154.340 120.180 154.660 ;
        RECT 120.440 145.820 120.580 173.380 ;
        RECT 120.900 150.095 121.040 176.360 ;
        RECT 121.360 170.980 121.500 179.840 ;
        RECT 122.280 178.120 122.420 181.005 ;
        RECT 122.740 180.840 122.880 183.920 ;
        RECT 122.680 180.520 122.940 180.840 ;
        RECT 122.220 177.800 122.480 178.120 ;
        RECT 121.760 175.255 122.020 175.400 ;
        RECT 121.750 174.885 122.030 175.255 ;
        RECT 121.300 170.660 121.560 170.980 ;
        RECT 121.360 168.260 121.500 170.660 ;
        RECT 121.300 167.940 121.560 168.260 ;
        RECT 121.300 165.220 121.560 165.540 ;
        RECT 120.830 149.725 121.110 150.095 ;
        RECT 115.320 145.500 115.580 145.645 ;
        RECT 117.160 145.590 118.280 145.730 ;
        RECT 117.160 145.500 117.420 145.590 ;
        RECT 119.460 145.500 119.720 145.820 ;
        RECT 120.380 145.500 120.640 145.820 ;
        RECT 113.940 145.160 114.200 145.480 ;
        RECT 113.020 143.460 113.280 143.780 ;
        RECT 113.480 143.460 113.740 143.780 ;
        RECT 114.000 142.760 114.140 145.160 ;
        RECT 116.240 144.480 116.500 144.800 ;
        RECT 120.380 144.480 120.640 144.800 ;
        RECT 116.300 142.760 116.440 144.480 ;
        RECT 120.440 142.760 120.580 144.480 ;
        RECT 121.360 143.780 121.500 165.220 ;
        RECT 121.820 160.100 121.960 174.885 ;
        RECT 122.740 173.020 122.880 180.520 ;
        RECT 123.200 177.440 123.340 186.920 ;
        RECT 123.140 177.120 123.400 177.440 ;
        RECT 123.140 174.400 123.400 174.720 ;
        RECT 123.200 173.360 123.340 174.400 ;
        RECT 123.140 173.040 123.400 173.360 ;
        RECT 122.680 172.700 122.940 173.020 ;
        RECT 122.740 169.960 122.880 172.700 ;
        RECT 122.680 169.640 122.940 169.960 ;
        RECT 123.140 169.640 123.400 169.960 ;
        RECT 122.220 169.300 122.480 169.620 ;
        RECT 122.280 163.750 122.420 169.300 ;
        RECT 122.740 167.240 122.880 169.640 ;
        RECT 123.200 168.260 123.340 169.640 ;
        RECT 123.140 167.940 123.400 168.260 ;
        RECT 122.680 166.920 122.940 167.240 ;
        RECT 122.680 163.750 122.940 163.840 ;
        RECT 122.280 163.610 122.940 163.750 ;
        RECT 122.680 163.520 122.940 163.610 ;
        RECT 122.740 162.140 122.880 163.520 ;
        RECT 122.680 161.820 122.940 162.140 ;
        RECT 121.760 159.780 122.020 160.100 ;
        RECT 123.140 156.380 123.400 156.700 ;
        RECT 123.200 156.215 123.340 156.380 ;
        RECT 123.130 155.845 123.410 156.215 ;
        RECT 122.680 151.280 122.940 151.600 ;
        RECT 122.740 148.200 122.880 151.280 ;
        RECT 122.680 147.880 122.940 148.200 ;
        RECT 123.660 147.940 123.800 200.720 ;
        RECT 124.970 200.045 125.250 200.415 ;
        RECT 124.980 199.900 125.240 200.045 ;
        RECT 125.440 199.900 125.700 200.220 ;
        RECT 126.820 199.900 127.080 200.220 ;
        RECT 125.040 198.180 125.180 199.900 ;
        RECT 124.980 197.860 125.240 198.180 ;
        RECT 124.520 194.800 124.780 195.120 ;
        RECT 124.580 192.740 124.720 194.800 ;
        RECT 125.500 194.780 125.640 199.900 ;
        RECT 125.900 198.880 126.160 199.200 ;
        RECT 126.360 198.880 126.620 199.200 ;
        RECT 125.960 198.180 126.100 198.880 ;
        RECT 125.900 197.860 126.160 198.180 ;
        RECT 126.420 197.160 126.560 198.880 ;
        RECT 126.880 198.180 127.020 199.900 ;
        RECT 127.280 199.560 127.540 199.880 ;
        RECT 126.820 197.860 127.080 198.180 ;
        RECT 126.360 196.840 126.620 197.160 ;
        RECT 125.440 194.460 125.700 194.780 ;
        RECT 124.520 192.420 124.780 192.740 ;
        RECT 124.060 185.280 124.320 185.600 ;
        RECT 124.120 183.220 124.260 185.280 ;
        RECT 124.060 182.900 124.320 183.220 ;
        RECT 124.580 179.220 124.720 192.420 ;
        RECT 124.980 189.020 125.240 189.340 ;
        RECT 125.040 186.960 125.180 189.020 ;
        RECT 124.980 186.640 125.240 186.960 ;
        RECT 125.040 183.900 125.180 186.640 ;
        RECT 124.980 183.580 125.240 183.900 ;
        RECT 125.500 181.860 125.640 194.460 ;
        RECT 125.900 190.720 126.160 191.040 ;
        RECT 125.960 186.020 126.100 190.720 ;
        RECT 126.420 186.620 126.560 196.840 ;
        RECT 127.340 194.780 127.480 199.560 ;
        RECT 127.280 194.460 127.540 194.780 ;
        RECT 126.820 189.700 127.080 190.020 ;
        RECT 126.360 186.300 126.620 186.620 ;
        RECT 125.960 185.880 126.560 186.020 ;
        RECT 126.880 185.940 127.020 189.700 ;
        RECT 125.900 183.580 126.160 183.900 ;
        RECT 125.440 181.540 125.700 181.860 ;
        RECT 124.120 179.080 124.720 179.220 ;
        RECT 124.120 175.400 124.260 179.080 ;
        RECT 124.970 177.605 125.250 177.975 ;
        RECT 125.040 175.400 125.180 177.605 ;
        RECT 124.060 175.080 124.320 175.400 ;
        RECT 124.980 175.080 125.240 175.400 ;
        RECT 124.120 169.280 124.260 175.080 ;
        RECT 125.040 169.960 125.180 175.080 ;
        RECT 125.960 171.910 126.100 183.580 ;
        RECT 126.420 182.620 126.560 185.880 ;
        RECT 126.820 185.620 127.080 185.940 ;
        RECT 127.280 185.280 127.540 185.600 ;
        RECT 127.740 185.280 128.000 185.600 ;
        RECT 127.340 184.580 127.480 185.280 ;
        RECT 127.280 184.260 127.540 184.580 ;
        RECT 127.800 184.240 127.940 185.280 ;
        RECT 127.740 183.920 128.000 184.240 ;
        RECT 127.280 182.900 127.540 183.220 ;
        RECT 127.340 182.620 127.480 182.900 ;
        RECT 126.420 182.480 127.480 182.620 ;
        RECT 127.340 180.695 127.480 182.480 ;
        RECT 127.740 181.540 128.000 181.860 ;
        RECT 127.270 180.325 127.550 180.695 ;
        RECT 126.820 179.840 127.080 180.160 ;
        RECT 126.880 178.460 127.020 179.840 ;
        RECT 126.820 178.140 127.080 178.460 ;
        RECT 126.880 176.420 127.020 178.140 ;
        RECT 127.280 177.120 127.540 177.440 ;
        RECT 127.340 176.420 127.480 177.120 ;
        RECT 126.820 176.100 127.080 176.420 ;
        RECT 127.280 176.100 127.540 176.420 ;
        RECT 127.800 175.400 127.940 181.540 ;
        RECT 126.820 175.080 127.080 175.400 ;
        RECT 127.740 175.080 128.000 175.400 ;
        RECT 126.880 172.680 127.020 175.080 ;
        RECT 126.820 172.360 127.080 172.680 ;
        RECT 125.960 171.770 127.020 171.910 ;
        RECT 124.980 169.640 125.240 169.960 ;
        RECT 124.060 168.960 124.320 169.280 ;
        RECT 124.120 167.580 124.260 168.960 ;
        RECT 124.060 167.260 124.320 167.580 ;
        RECT 124.520 166.920 124.780 167.240 ;
        RECT 124.580 164.520 124.720 166.920 ;
        RECT 124.520 164.200 124.780 164.520 ;
        RECT 125.440 164.200 125.700 164.520 ;
        RECT 124.520 162.160 124.780 162.480 ;
        RECT 124.580 160.100 124.720 162.160 ;
        RECT 125.500 161.120 125.640 164.200 ;
        RECT 126.880 161.800 127.020 171.770 ;
        RECT 127.280 169.980 127.540 170.300 ;
        RECT 127.340 167.580 127.480 169.980 ;
        RECT 127.280 167.260 127.540 167.580 ;
        RECT 127.740 167.260 128.000 167.580 ;
        RECT 127.800 165.200 127.940 167.260 ;
        RECT 127.740 164.880 128.000 165.200 ;
        RECT 126.820 161.480 127.080 161.800 ;
        RECT 125.440 160.800 125.700 161.120 ;
        RECT 124.520 159.780 124.780 160.100 ;
        RECT 124.980 155.700 125.240 156.020 ;
        RECT 125.040 153.980 125.180 155.700 ;
        RECT 124.980 153.660 125.240 153.980 ;
        RECT 124.510 151.765 124.790 152.135 ;
        RECT 124.580 151.260 124.720 151.765 ;
        RECT 125.040 151.260 125.180 153.660 ;
        RECT 124.520 150.940 124.780 151.260 ;
        RECT 124.980 150.940 125.240 151.260 ;
        RECT 124.580 148.110 124.720 150.940 ;
        RECT 125.500 150.240 125.640 160.800 ;
        RECT 125.900 159.780 126.160 160.100 ;
        RECT 125.960 159.615 126.100 159.780 ;
        RECT 125.890 159.245 126.170 159.615 ;
        RECT 126.880 159.420 127.020 161.480 ;
        RECT 127.740 160.800 128.000 161.120 ;
        RECT 126.820 159.100 127.080 159.420 ;
        RECT 125.890 158.565 126.170 158.935 ;
        RECT 125.960 155.680 126.100 158.565 ;
        RECT 126.360 158.420 126.620 158.740 ;
        RECT 126.420 157.380 126.560 158.420 ;
        RECT 126.360 157.290 126.620 157.380 ;
        RECT 126.360 157.150 127.480 157.290 ;
        RECT 126.360 157.060 126.620 157.150 ;
        RECT 126.350 155.930 126.630 156.215 ;
        RECT 126.820 155.930 127.080 156.020 ;
        RECT 126.350 155.845 127.080 155.930 ;
        RECT 126.420 155.790 127.080 155.845 ;
        RECT 126.820 155.700 127.080 155.790 ;
        RECT 125.900 155.360 126.160 155.680 ;
        RECT 125.960 154.320 126.100 155.360 ;
        RECT 125.900 154.000 126.160 154.320 ;
        RECT 127.340 153.640 127.480 157.150 ;
        RECT 127.800 156.895 127.940 160.800 ;
        RECT 127.730 156.525 128.010 156.895 ;
        RECT 127.800 154.660 127.940 156.525 ;
        RECT 127.740 154.340 128.000 154.660 ;
        RECT 127.280 153.320 127.540 153.640 ;
        RECT 126.820 152.640 127.080 152.960 ;
        RECT 125.440 149.920 125.700 150.240 ;
        RECT 123.200 147.800 123.800 147.940 ;
        RECT 124.120 147.970 124.720 148.110 ;
        RECT 125.500 148.055 125.640 149.920 ;
        RECT 126.880 149.220 127.020 152.640 ;
        RECT 128.260 151.850 128.400 200.720 ;
        RECT 128.660 200.240 128.920 200.560 ;
        RECT 128.720 190.020 128.860 200.240 ;
        RECT 130.160 198.345 132.040 198.715 ;
        RECT 132.860 197.160 133.000 201.940 ;
        RECT 129.120 196.840 129.380 197.160 ;
        RECT 132.800 196.840 133.060 197.160 ;
        RECT 129.180 195.460 129.320 196.840 ;
        RECT 129.120 195.140 129.380 195.460 ;
        RECT 132.800 195.140 133.060 195.460 ;
        RECT 132.340 194.800 132.600 195.120 ;
        RECT 131.880 194.295 132.140 194.440 ;
        RECT 131.870 193.925 132.150 194.295 ;
        RECT 130.160 192.905 132.040 193.275 ;
        RECT 132.400 192.740 132.540 194.800 ;
        RECT 132.860 192.740 133.000 195.140 ;
        RECT 133.320 193.500 133.460 201.940 ;
        RECT 133.780 194.100 133.920 208.205 ;
        RECT 134.240 208.040 134.380 212.480 ;
        RECT 140.680 211.780 140.820 213.160 ;
        RECT 141.080 212.480 141.340 212.800 ;
        RECT 140.620 211.460 140.880 211.780 ;
        RECT 140.680 209.060 140.820 211.460 ;
        RECT 140.620 208.740 140.880 209.060 ;
        RECT 134.180 207.720 134.440 208.040 ;
        RECT 134.240 201.920 134.380 207.720 ;
        RECT 140.620 205.680 140.880 206.000 ;
        RECT 140.160 205.340 140.420 205.660 ;
        RECT 134.640 205.000 134.900 205.320 ;
        RECT 134.700 202.600 134.840 205.000 ;
        RECT 135.560 204.320 135.820 204.640 ;
        RECT 135.620 202.600 135.760 204.320 ;
        RECT 140.220 203.620 140.360 205.340 ;
        RECT 140.680 203.700 140.820 205.680 ;
        RECT 141.140 204.980 141.280 212.480 ;
        RECT 145.160 211.945 147.040 212.315 ;
        RECT 145.160 206.505 147.040 206.875 ;
        RECT 141.080 204.660 141.340 204.980 ;
        RECT 140.160 203.300 140.420 203.620 ;
        RECT 140.680 203.560 141.740 203.700 ;
        RECT 141.080 202.620 141.340 202.940 ;
        RECT 134.640 202.280 134.900 202.600 ;
        RECT 135.560 202.280 135.820 202.600 ;
        RECT 134.180 201.600 134.440 201.920 ;
        RECT 134.700 200.560 134.840 202.280 ;
        RECT 136.940 201.600 137.200 201.920 ;
        RECT 134.640 200.240 134.900 200.560 ;
        RECT 134.700 197.500 134.840 200.240 ;
        RECT 134.640 197.180 134.900 197.500 ;
        RECT 136.480 197.180 136.740 197.500 ;
        RECT 135.100 196.840 135.360 197.160 ;
        RECT 133.720 193.780 133.980 194.100 ;
        RECT 133.320 193.360 134.380 193.500 ;
        RECT 134.640 193.440 134.900 193.760 ;
        RECT 132.340 192.420 132.600 192.740 ;
        RECT 132.800 192.420 133.060 192.740 ;
        RECT 130.040 191.630 130.300 191.720 ;
        RECT 129.640 191.490 130.300 191.630 ;
        RECT 128.660 189.700 128.920 190.020 ;
        RECT 128.650 189.420 128.930 189.535 ;
        RECT 129.640 189.420 129.780 191.490 ;
        RECT 130.040 191.400 130.300 191.490 ;
        RECT 132.860 191.460 133.000 192.420 ;
        RECT 132.860 191.320 133.920 191.460 ;
        RECT 132.340 190.720 132.600 191.040 ;
        RECT 133.260 190.720 133.520 191.040 ;
        RECT 130.040 189.700 130.300 190.020 ;
        RECT 128.650 189.280 129.780 189.420 ;
        RECT 128.650 189.165 128.930 189.280 ;
        RECT 129.180 186.620 129.320 189.280 ;
        RECT 130.100 189.000 130.240 189.700 ;
        RECT 132.400 189.340 132.540 190.720 ;
        RECT 132.340 189.020 132.600 189.340 ;
        RECT 130.040 188.855 130.300 189.000 ;
        RECT 130.030 188.485 130.310 188.855 ;
        RECT 129.580 188.000 129.840 188.320 ;
        RECT 132.400 188.060 132.540 189.020 ;
        RECT 132.800 188.680 133.060 189.000 ;
        RECT 132.860 188.175 133.000 188.680 ;
        RECT 129.640 187.210 129.780 188.000 ;
        RECT 132.400 187.920 132.585 188.060 ;
        RECT 130.160 187.465 132.040 187.835 ;
        RECT 132.445 187.380 132.585 187.920 ;
        RECT 132.790 187.805 133.070 188.175 ;
        RECT 133.320 187.380 133.460 190.720 ;
        RECT 133.780 189.000 133.920 191.320 ;
        RECT 134.240 190.020 134.380 193.360 ;
        RECT 134.700 192.060 134.840 193.440 ;
        RECT 134.640 191.740 134.900 192.060 ;
        RECT 134.180 189.700 134.440 190.020 ;
        RECT 133.720 188.910 133.980 189.000 ;
        RECT 133.720 188.770 134.380 188.910 ;
        RECT 133.720 188.680 133.980 188.770 ;
        RECT 132.400 187.240 132.585 187.380 ;
        RECT 132.860 187.240 133.460 187.380 ;
        RECT 129.640 187.070 130.700 187.210 ;
        RECT 129.120 186.300 129.380 186.620 ;
        RECT 130.030 186.445 130.310 186.815 ;
        RECT 130.100 183.900 130.240 186.445 ;
        RECT 130.560 184.775 130.700 187.070 ;
        RECT 130.960 185.620 131.220 185.940 ;
        RECT 130.490 184.405 130.770 184.775 ;
        RECT 129.120 183.580 129.380 183.900 ;
        RECT 130.040 183.580 130.300 183.900 ;
        RECT 129.180 183.300 129.320 183.580 ;
        RECT 131.020 183.300 131.160 185.620 ;
        RECT 131.870 183.725 132.150 184.095 ;
        RECT 132.400 183.900 132.540 187.240 ;
        RECT 132.860 186.960 133.000 187.240 ;
        RECT 132.800 186.640 133.060 186.960 ;
        RECT 133.250 186.700 133.530 186.815 ;
        RECT 132.860 186.110 133.000 186.640 ;
        RECT 133.250 186.620 133.920 186.700 ;
        RECT 133.250 186.560 133.980 186.620 ;
        RECT 133.250 186.445 133.530 186.560 ;
        RECT 133.720 186.300 133.980 186.560 ;
        RECT 132.800 185.790 133.060 186.110 ;
        RECT 133.260 185.280 133.520 185.600 ;
        RECT 133.320 183.900 133.460 185.280 ;
        RECT 133.720 183.920 133.980 184.240 ;
        RECT 131.940 183.560 132.080 183.725 ;
        RECT 132.340 183.580 132.600 183.900 ;
        RECT 133.260 183.580 133.520 183.900 ;
        RECT 128.660 182.900 128.920 183.220 ;
        RECT 129.180 183.160 131.160 183.300 ;
        RECT 131.880 183.240 132.140 183.560 ;
        RECT 128.720 181.860 128.860 182.900 ;
        RECT 130.040 182.790 130.300 182.880 ;
        RECT 129.640 182.650 130.300 182.790 ;
        RECT 129.640 181.860 129.780 182.650 ;
        RECT 130.040 182.560 130.300 182.650 ;
        RECT 130.160 182.025 132.040 182.395 ;
        RECT 132.400 181.860 132.540 183.580 ;
        RECT 132.800 182.560 133.060 182.880 ;
        RECT 128.660 181.540 128.920 181.860 ;
        RECT 129.580 181.540 129.840 181.860 ;
        RECT 132.340 181.540 132.600 181.860 ;
        RECT 130.040 180.520 130.300 180.840 ;
        RECT 130.100 177.350 130.240 180.520 ;
        RECT 132.340 179.840 132.600 180.160 ;
        RECT 132.400 178.460 132.540 179.840 ;
        RECT 132.340 178.140 132.600 178.460 ;
        RECT 129.640 177.210 130.240 177.350 ;
        RECT 129.640 176.330 129.780 177.210 ;
        RECT 130.160 176.585 132.040 176.955 ;
        RECT 130.040 176.330 130.300 176.420 ;
        RECT 129.640 176.190 130.300 176.330 ;
        RECT 130.040 176.100 130.300 176.190 ;
        RECT 132.340 175.080 132.600 175.400 ;
        RECT 130.160 171.145 132.040 171.515 ;
        RECT 132.400 169.960 132.540 175.080 ;
        RECT 132.340 169.640 132.600 169.960 ;
        RECT 128.660 168.960 128.920 169.280 ;
        RECT 128.720 166.560 128.860 168.960 ;
        RECT 132.400 167.580 132.540 169.640 ;
        RECT 129.120 167.260 129.380 167.580 ;
        RECT 132.340 167.260 132.600 167.580 ;
        RECT 128.660 166.240 128.920 166.560 ;
        RECT 129.180 165.540 129.320 167.260 ;
        RECT 130.160 165.705 132.040 166.075 ;
        RECT 129.120 165.220 129.380 165.540 ;
        RECT 132.340 162.160 132.600 162.480 ;
        RECT 131.410 161.285 131.690 161.655 ;
        RECT 131.420 161.140 131.680 161.285 ;
        RECT 130.160 160.265 132.040 160.635 ;
        RECT 131.420 158.420 131.680 158.740 ;
        RECT 131.480 156.700 131.620 158.420 ;
        RECT 132.400 156.700 132.540 162.160 ;
        RECT 132.860 157.380 133.000 182.560 ;
        RECT 133.320 181.520 133.460 183.580 ;
        RECT 133.780 181.860 133.920 183.920 ;
        RECT 134.240 183.560 134.380 188.770 ;
        RECT 134.640 188.000 134.900 188.320 ;
        RECT 134.700 186.815 134.840 188.000 ;
        RECT 134.630 186.445 134.910 186.815 ;
        RECT 134.180 183.240 134.440 183.560 ;
        RECT 134.640 182.790 134.900 182.880 ;
        RECT 134.240 182.650 134.900 182.790 ;
        RECT 133.720 181.540 133.980 181.860 ;
        RECT 133.260 181.200 133.520 181.520 ;
        RECT 134.240 180.580 134.380 182.650 ;
        RECT 134.640 182.560 134.900 182.650 ;
        RECT 133.320 180.500 134.380 180.580 ;
        RECT 133.260 180.440 134.380 180.500 ;
        RECT 133.260 180.180 133.520 180.440 ;
        RECT 134.640 180.180 134.900 180.500 ;
        RECT 134.700 180.015 134.840 180.180 ;
        RECT 133.250 179.645 133.530 180.015 ;
        RECT 134.630 179.645 134.910 180.015 ;
        RECT 133.320 178.120 133.460 179.645 ;
        RECT 135.160 178.540 135.300 196.840 ;
        RECT 135.560 196.500 135.820 196.820 ;
        RECT 135.620 184.580 135.760 196.500 ;
        RECT 136.540 195.460 136.680 197.180 ;
        RECT 137.000 197.015 137.140 201.600 ;
        RECT 136.930 196.900 137.210 197.015 ;
        RECT 136.930 196.760 137.600 196.900 ;
        RECT 138.780 196.840 139.040 197.160 ;
        RECT 136.930 196.645 137.210 196.760 ;
        RECT 136.020 195.140 136.280 195.460 ;
        RECT 136.480 195.140 136.740 195.460 ;
        RECT 136.080 186.960 136.220 195.140 ;
        RECT 136.480 194.460 136.740 194.780 ;
        RECT 136.540 194.295 136.680 194.460 ;
        RECT 136.470 193.925 136.750 194.295 ;
        RECT 136.940 193.440 137.200 193.760 ;
        RECT 137.000 191.720 137.140 193.440 ;
        RECT 137.460 191.720 137.600 196.760 ;
        RECT 137.860 196.500 138.120 196.820 ;
        RECT 137.920 192.740 138.060 196.500 ;
        RECT 138.320 196.160 138.580 196.480 ;
        RECT 138.380 195.460 138.520 196.160 ;
        RECT 138.320 195.140 138.580 195.460 ;
        RECT 138.840 194.780 138.980 196.840 ;
        RECT 138.780 194.460 139.040 194.780 ;
        RECT 137.860 192.420 138.120 192.740 ;
        RECT 136.940 191.400 137.200 191.720 ;
        RECT 137.400 191.400 137.660 191.720 ;
        RECT 141.140 190.020 141.280 202.620 ;
        RECT 141.080 189.700 141.340 190.020 ;
        RECT 141.600 189.340 141.740 203.560 ;
        RECT 149.810 202.765 150.090 203.135 ;
        RECT 149.820 202.620 150.080 202.765 ;
        RECT 144.300 201.940 144.560 202.260 ;
        RECT 143.840 196.160 144.100 196.480 ;
        RECT 143.900 192.060 144.040 196.160 ;
        RECT 143.840 191.740 144.100 192.060 ;
        RECT 142.460 190.720 142.720 191.040 ;
        RECT 141.540 189.020 141.800 189.340 ;
        RECT 141.080 188.680 141.340 189.000 ;
        RECT 142.000 188.680 142.260 189.000 ;
        RECT 139.240 188.340 139.500 188.660 ;
        RECT 136.480 188.000 136.740 188.320 ;
        RECT 136.540 187.300 136.680 188.000 ;
        RECT 138.310 187.805 138.590 188.175 ;
        RECT 136.480 186.980 136.740 187.300 ;
        RECT 136.020 186.640 136.280 186.960 ;
        RECT 135.560 184.260 135.820 184.580 ;
        RECT 133.780 178.400 135.300 178.540 ;
        RECT 133.260 177.800 133.520 178.120 ;
        RECT 133.260 177.120 133.520 177.440 ;
        RECT 133.320 169.815 133.460 177.120 ;
        RECT 133.250 169.445 133.530 169.815 ;
        RECT 133.260 163.860 133.520 164.180 ;
        RECT 133.320 162.140 133.460 163.860 ;
        RECT 133.260 161.820 133.520 162.140 ;
        RECT 133.260 160.800 133.520 161.120 ;
        RECT 133.320 159.080 133.460 160.800 ;
        RECT 133.780 159.760 133.920 178.400 ;
        RECT 134.640 177.800 134.900 178.120 ;
        RECT 134.180 161.140 134.440 161.460 ;
        RECT 134.240 160.100 134.380 161.140 ;
        RECT 134.180 159.780 134.440 160.100 ;
        RECT 133.720 159.440 133.980 159.760 ;
        RECT 133.260 158.760 133.520 159.080 ;
        RECT 132.800 157.060 133.060 157.380 ;
        RECT 131.420 156.380 131.680 156.700 ;
        RECT 132.340 156.380 132.600 156.700 ;
        RECT 133.250 156.525 133.530 156.895 ;
        RECT 133.320 156.360 133.460 156.525 ;
        RECT 133.260 156.040 133.520 156.360 ;
        RECT 128.660 155.360 128.920 155.680 ;
        RECT 132.800 155.360 133.060 155.680 ;
        RECT 133.720 155.360 133.980 155.680 ;
        RECT 128.720 153.640 128.860 155.360 ;
        RECT 130.160 154.825 132.040 155.195 ;
        RECT 130.500 154.000 130.760 154.320 ;
        RECT 128.660 153.320 128.920 153.640 ;
        RECT 130.040 153.320 130.300 153.640 ;
        RECT 130.100 152.560 130.240 153.320 ;
        RECT 127.800 151.710 128.400 151.850 ;
        RECT 129.640 152.420 130.240 152.560 ;
        RECT 127.800 150.775 127.940 151.710 ;
        RECT 129.640 150.920 129.780 152.420 ;
        RECT 130.560 151.850 130.700 154.000 ;
        RECT 131.870 153.380 132.150 153.495 ;
        RECT 132.860 153.380 133.000 155.360 ;
        RECT 131.870 153.240 133.000 153.380 ;
        RECT 133.780 153.300 133.920 155.360 ;
        RECT 134.700 153.300 134.840 177.800 ;
        RECT 135.100 176.100 135.360 176.420 ;
        RECT 135.160 173.020 135.300 176.100 ;
        RECT 135.100 172.700 135.360 173.020 ;
        RECT 135.100 164.880 135.360 165.200 ;
        RECT 135.160 164.520 135.300 164.880 ;
        RECT 135.100 164.200 135.360 164.520 ;
        RECT 135.160 159.420 135.300 164.200 ;
        RECT 135.620 162.480 135.760 184.260 ;
        RECT 136.020 180.520 136.280 180.840 ;
        RECT 136.080 178.460 136.220 180.520 ;
        RECT 136.020 178.140 136.280 178.460 ;
        RECT 136.080 176.080 136.220 178.140 ;
        RECT 136.020 175.760 136.280 176.080 ;
        RECT 135.560 162.160 135.820 162.480 ;
        RECT 135.100 159.100 135.360 159.420 ;
        RECT 135.620 159.080 135.760 162.160 ;
        RECT 136.540 159.760 136.680 186.980 ;
        RECT 137.400 185.960 137.660 186.280 ;
        RECT 136.940 185.280 137.200 185.600 ;
        RECT 137.000 181.860 137.140 185.280 ;
        RECT 137.460 183.415 137.600 185.960 ;
        RECT 138.380 183.900 138.520 187.805 ;
        RECT 139.300 187.300 139.440 188.340 ;
        RECT 139.240 186.980 139.500 187.300 ;
        RECT 140.160 186.980 140.420 187.300 ;
        RECT 139.690 186.445 139.970 186.815 ;
        RECT 138.780 186.135 139.040 186.280 ;
        RECT 138.770 185.765 139.050 186.135 ;
        RECT 138.320 183.580 138.580 183.900 ;
        RECT 137.390 183.045 137.670 183.415 ;
        RECT 137.860 183.240 138.120 183.560 ;
        RECT 136.940 181.540 137.200 181.860 ;
        RECT 136.930 180.325 137.210 180.695 ;
        RECT 137.000 178.120 137.140 180.325 ;
        RECT 137.400 178.140 137.660 178.460 ;
        RECT 136.940 177.800 137.200 178.120 ;
        RECT 137.460 176.420 137.600 178.140 ;
        RECT 137.400 176.100 137.660 176.420 ;
        RECT 136.940 171.680 137.200 172.000 ;
        RECT 137.000 170.980 137.140 171.680 ;
        RECT 136.940 170.660 137.200 170.980 ;
        RECT 137.000 161.120 137.140 170.660 ;
        RECT 137.920 170.210 138.060 183.240 ;
        RECT 138.320 182.560 138.580 182.880 ;
        RECT 138.380 170.300 138.520 182.560 ;
        RECT 139.760 181.180 139.900 186.445 ;
        RECT 140.220 184.095 140.360 186.980 ;
        RECT 140.150 183.725 140.430 184.095 ;
        RECT 140.620 183.920 140.880 184.240 ;
        RECT 140.220 181.860 140.360 183.725 ;
        RECT 140.160 181.540 140.420 181.860 ;
        RECT 140.680 181.520 140.820 183.920 ;
        RECT 140.620 181.200 140.880 181.520 ;
        RECT 139.700 180.860 139.960 181.180 ;
        RECT 140.160 180.520 140.420 180.840 ;
        RECT 139.240 180.180 139.500 180.500 ;
        RECT 139.700 180.180 139.960 180.500 ;
        RECT 138.780 177.120 139.040 177.440 ;
        RECT 138.840 176.420 138.980 177.120 ;
        RECT 138.780 176.100 139.040 176.420 ;
        RECT 137.460 170.070 138.060 170.210 ;
        RECT 137.460 162.820 137.600 170.070 ;
        RECT 138.320 169.980 138.580 170.300 ;
        RECT 137.860 169.300 138.120 169.620 ;
        RECT 138.320 169.300 138.580 169.620 ;
        RECT 137.920 165.540 138.060 169.300 ;
        RECT 137.860 165.220 138.120 165.540 ;
        RECT 137.400 162.500 137.660 162.820 ;
        RECT 138.380 162.140 138.520 169.300 ;
        RECT 138.780 163.860 139.040 164.180 ;
        RECT 138.320 161.820 138.580 162.140 ;
        RECT 138.380 161.460 138.520 161.820 ;
        RECT 138.840 161.800 138.980 163.860 ;
        RECT 139.300 162.820 139.440 180.180 ;
        RECT 139.760 180.015 139.900 180.180 ;
        RECT 139.690 179.645 139.970 180.015 ;
        RECT 139.760 173.700 139.900 179.645 ;
        RECT 140.220 177.440 140.360 180.520 ;
        RECT 140.160 177.120 140.420 177.440 ;
        RECT 140.220 175.400 140.360 177.120 ;
        RECT 140.160 175.080 140.420 175.400 ;
        RECT 139.700 173.380 139.960 173.700 ;
        RECT 139.700 169.980 139.960 170.300 ;
        RECT 139.240 162.500 139.500 162.820 ;
        RECT 139.760 162.140 139.900 169.980 ;
        RECT 140.150 166.725 140.430 167.095 ;
        RECT 140.160 166.580 140.420 166.725 ;
        RECT 140.680 164.520 140.820 181.200 ;
        RECT 141.140 169.280 141.280 188.680 ;
        RECT 141.530 186.445 141.810 186.815 ;
        RECT 141.600 186.280 141.740 186.445 ;
        RECT 141.540 185.960 141.800 186.280 ;
        RECT 141.540 185.280 141.800 185.600 ;
        RECT 141.600 181.375 141.740 185.280 ;
        RECT 142.060 184.580 142.200 188.680 ;
        RECT 142.000 184.260 142.260 184.580 ;
        RECT 141.530 181.005 141.810 181.375 ;
        RECT 141.540 180.860 141.800 181.005 ;
        RECT 142.520 173.020 142.660 190.720 ;
        RECT 143.900 187.300 144.040 191.740 ;
        RECT 144.360 190.020 144.500 201.940 ;
        RECT 147.520 201.600 147.780 201.920 ;
        RECT 145.160 201.065 147.040 201.435 ;
        RECT 144.760 198.880 145.020 199.200 ;
        RECT 144.820 193.760 144.960 198.880 ;
        RECT 145.160 195.625 147.040 195.995 ;
        RECT 144.760 193.440 145.020 193.760 ;
        RECT 144.820 191.720 144.960 193.440 ;
        RECT 147.580 192.060 147.720 201.600 ;
        RECT 147.520 191.740 147.780 192.060 ;
        RECT 144.760 191.400 145.020 191.720 ;
        RECT 144.300 189.700 144.560 190.020 ;
        RECT 144.300 188.680 144.560 189.000 ;
        RECT 144.360 187.300 144.500 188.680 ;
        RECT 143.840 186.980 144.100 187.300 ;
        RECT 144.300 186.980 144.560 187.300 ;
        RECT 143.380 186.700 143.640 186.960 ;
        RECT 144.820 186.700 144.960 191.400 ;
        RECT 145.160 190.185 147.040 190.555 ;
        RECT 145.680 189.020 145.940 189.340 ;
        RECT 145.740 187.300 145.880 189.020 ;
        RECT 147.060 188.000 147.320 188.320 ;
        RECT 145.680 186.980 145.940 187.300 ;
        RECT 143.380 186.640 144.960 186.700 ;
        RECT 143.440 186.560 144.960 186.640 ;
        RECT 143.830 185.765 144.110 186.135 ;
        RECT 144.300 185.960 144.560 186.280 ;
        RECT 143.840 185.620 144.100 185.765 ;
        RECT 143.380 185.280 143.640 185.600 ;
        RECT 143.440 181.860 143.580 185.280 ;
        RECT 143.380 181.540 143.640 181.860 ;
        RECT 142.460 172.700 142.720 173.020 ;
        RECT 142.920 172.700 143.180 173.020 ;
        RECT 141.540 171.680 141.800 172.000 ;
        RECT 142.000 171.680 142.260 172.000 ;
        RECT 141.080 168.960 141.340 169.280 ;
        RECT 141.600 165.540 141.740 171.680 ;
        RECT 142.060 166.900 142.200 171.680 ;
        RECT 142.460 170.890 142.720 170.980 ;
        RECT 142.980 170.890 143.120 172.700 ;
        RECT 142.460 170.750 143.120 170.890 ;
        RECT 142.460 170.660 142.720 170.750 ;
        RECT 142.520 167.580 142.660 170.660 ;
        RECT 143.900 168.260 144.040 185.620 ;
        RECT 144.360 184.580 144.500 185.960 ;
        RECT 147.120 185.940 147.260 188.000 ;
        RECT 147.580 186.280 147.720 191.740 ;
        RECT 147.980 190.720 148.240 191.040 ;
        RECT 147.520 185.960 147.780 186.280 ;
        RECT 147.060 185.620 147.320 185.940 ;
        RECT 145.160 184.745 147.040 185.115 ;
        RECT 144.300 184.260 144.560 184.580 ;
        RECT 148.040 181.180 148.180 190.720 ;
        RECT 147.980 180.860 148.240 181.180 ;
        RECT 145.160 179.305 147.040 179.675 ;
        RECT 145.160 173.865 147.040 174.235 ;
        RECT 145.160 168.425 147.040 168.795 ;
        RECT 143.840 167.940 144.100 168.260 ;
        RECT 142.460 167.260 142.720 167.580 ;
        RECT 142.920 167.260 143.180 167.580 ;
        RECT 142.000 166.580 142.260 166.900 ;
        RECT 141.080 165.220 141.340 165.540 ;
        RECT 141.540 165.220 141.800 165.540 ;
        RECT 140.160 164.200 140.420 164.520 ;
        RECT 140.620 164.200 140.880 164.520 ;
        RECT 139.700 161.820 139.960 162.140 ;
        RECT 138.780 161.480 139.040 161.800 ;
        RECT 138.320 161.140 138.580 161.460 ;
        RECT 136.940 160.800 137.200 161.120 ;
        RECT 137.400 160.800 137.660 161.120 ;
        RECT 136.480 159.440 136.740 159.760 ;
        RECT 137.460 159.670 137.600 160.800 ;
        RECT 137.000 159.530 137.600 159.670 ;
        RECT 137.000 159.080 137.140 159.530 ;
        RECT 135.560 158.760 135.820 159.080 ;
        RECT 136.480 158.760 136.740 159.080 ;
        RECT 136.940 158.760 137.200 159.080 ;
        RECT 137.400 158.760 137.660 159.080 ;
        RECT 131.870 153.125 132.150 153.240 ;
        RECT 130.100 151.710 130.700 151.850 ;
        RECT 130.100 151.260 130.240 151.710 ;
        RECT 131.940 151.260 132.080 153.125 ;
        RECT 133.720 152.980 133.980 153.300 ;
        RECT 134.640 152.980 134.900 153.300 ;
        RECT 134.700 151.940 134.840 152.980 ;
        RECT 134.640 151.620 134.900 151.940 ;
        RECT 130.040 150.940 130.300 151.260 ;
        RECT 131.880 150.940 132.140 151.260 ;
        RECT 136.540 150.920 136.680 158.760 ;
        RECT 137.460 157.380 137.600 158.760 ;
        RECT 137.400 157.060 137.660 157.380 ;
        RECT 137.860 156.720 138.120 157.040 ;
        RECT 137.400 156.380 137.660 156.700 ;
        RECT 137.460 151.940 137.600 156.380 ;
        RECT 137.920 154.660 138.060 156.720 ;
        RECT 137.860 154.340 138.120 154.660 ;
        RECT 137.400 151.620 137.660 151.940 ;
        RECT 127.730 150.660 128.010 150.775 ;
        RECT 127.730 150.520 128.400 150.660 ;
        RECT 129.580 150.600 129.840 150.920 ;
        RECT 136.480 150.600 136.740 150.920 ;
        RECT 127.730 150.405 128.010 150.520 ;
        RECT 126.820 148.900 127.080 149.220 ;
        RECT 127.740 148.900 128.000 149.220 ;
        RECT 121.760 145.730 122.020 145.820 ;
        RECT 123.200 145.730 123.340 147.800 ;
        RECT 123.600 147.200 123.860 147.520 ;
        RECT 123.660 146.160 123.800 147.200 ;
        RECT 123.600 145.840 123.860 146.160 ;
        RECT 121.760 145.590 123.340 145.730 ;
        RECT 121.760 145.500 122.020 145.590 ;
        RECT 123.140 144.480 123.400 144.800 ;
        RECT 121.300 143.460 121.560 143.780 ;
        RECT 123.200 143.100 123.340 144.480 ;
        RECT 123.140 142.780 123.400 143.100 ;
        RECT 112.560 142.440 112.820 142.760 ;
        RECT 113.940 142.440 114.200 142.760 ;
        RECT 116.240 142.440 116.500 142.760 ;
        RECT 120.380 142.440 120.640 142.760 ;
        RECT 117.160 141.760 117.420 142.080 ;
        RECT 117.620 141.760 117.880 142.080 ;
        RECT 120.380 141.760 120.640 142.080 ;
        RECT 115.160 141.225 117.040 141.595 ;
        RECT 116.300 140.830 116.900 140.970 ;
        RECT 116.300 140.690 116.440 140.830 ;
        RECT 110.260 140.060 110.520 140.380 ;
        RECT 105.930 132.400 106.930 134.445 ;
        RECT 116.230 132.440 116.510 140.690 ;
        RECT 116.760 139.780 116.900 140.830 ;
        RECT 117.220 140.720 117.360 141.760 ;
        RECT 117.160 140.400 117.420 140.720 ;
        RECT 117.680 139.780 117.820 141.760 ;
        RECT 120.440 140.690 120.580 141.760 ;
        RECT 116.760 139.640 117.820 139.780 ;
        RECT 120.370 132.440 120.650 140.690 ;
        RECT 124.120 140.380 124.260 147.970 ;
        RECT 125.430 147.685 125.710 148.055 ;
        RECT 127.800 145.480 127.940 148.900 ;
        RECT 126.820 145.160 127.080 145.480 ;
        RECT 127.740 145.160 128.000 145.480 ;
        RECT 126.880 143.100 127.020 145.160 ;
        RECT 126.820 142.780 127.080 143.100 ;
        RECT 128.260 142.760 128.400 150.520 ;
        RECT 132.800 149.920 133.060 150.240 ;
        RECT 130.160 149.385 132.040 149.755 ;
        RECT 130.040 147.200 130.300 147.520 ;
        RECT 130.100 145.820 130.240 147.200 ;
        RECT 132.860 146.500 133.000 149.920 ;
        RECT 138.840 147.520 138.980 161.480 ;
        RECT 139.240 158.080 139.500 158.400 ;
        RECT 139.300 157.380 139.440 158.080 ;
        RECT 139.240 157.060 139.500 157.380 ;
        RECT 139.760 156.700 139.900 161.820 ;
        RECT 140.220 160.100 140.360 164.200 ;
        RECT 141.140 163.840 141.280 165.220 ;
        RECT 142.520 164.520 142.660 167.260 ;
        RECT 142.980 164.520 143.120 167.260 ;
        RECT 143.840 166.240 144.100 166.560 ;
        RECT 143.900 164.860 144.040 166.240 ;
        RECT 143.840 164.540 144.100 164.860 ;
        RECT 142.460 164.200 142.720 164.520 ;
        RECT 142.920 164.200 143.180 164.520 ;
        RECT 141.080 163.520 141.340 163.840 ;
        RECT 140.610 161.285 140.890 161.655 ;
        RECT 140.160 159.780 140.420 160.100 ;
        RECT 140.680 159.080 140.820 161.285 ;
        RECT 141.140 159.760 141.280 163.520 ;
        RECT 142.980 162.820 143.120 164.200 ;
        RECT 142.920 162.500 143.180 162.820 ;
        RECT 141.540 162.160 141.800 162.480 ;
        RECT 141.080 159.440 141.340 159.760 ;
        RECT 141.600 159.080 141.740 162.160 ;
        RECT 143.900 160.100 144.040 164.540 ;
        RECT 145.160 162.985 147.040 163.355 ;
        RECT 144.760 162.500 145.020 162.820 ;
        RECT 143.380 159.780 143.640 160.100 ;
        RECT 143.840 159.780 144.100 160.100 ;
        RECT 140.620 158.760 140.880 159.080 ;
        RECT 141.540 158.760 141.800 159.080 ;
        RECT 141.070 156.780 141.350 156.895 ;
        RECT 141.600 156.780 141.740 158.760 ;
        RECT 143.440 158.740 143.580 159.780 ;
        RECT 144.820 159.080 144.960 162.500 ;
        RECT 144.760 158.760 145.020 159.080 ;
        RECT 147.520 158.760 147.780 159.080 ;
        RECT 143.380 158.420 143.640 158.740 ;
        RECT 144.300 158.420 144.560 158.740 ;
        RECT 139.700 156.610 139.960 156.700 ;
        RECT 141.070 156.640 141.740 156.780 ;
        RECT 139.700 156.470 140.360 156.610 ;
        RECT 141.070 156.525 141.350 156.640 ;
        RECT 139.700 156.380 139.960 156.470 ;
        RECT 139.700 152.640 139.960 152.960 ;
        RECT 139.760 151.600 139.900 152.640 ;
        RECT 139.700 151.280 139.960 151.600 ;
        RECT 140.220 151.260 140.360 156.470 ;
        RECT 142.000 154.340 142.260 154.660 ;
        RECT 140.160 150.940 140.420 151.260 ;
        RECT 140.610 151.085 140.890 151.455 ;
        RECT 138.780 147.200 139.040 147.520 ;
        RECT 132.800 146.180 133.060 146.500 ;
        RECT 140.220 145.820 140.360 150.940 ;
        RECT 140.680 145.820 140.820 151.085 ;
        RECT 142.060 149.220 142.200 154.340 ;
        RECT 142.000 148.900 142.260 149.220 ;
        RECT 144.360 148.880 144.500 158.420 ;
        RECT 145.160 157.545 147.040 157.915 ;
        RECT 147.580 157.380 147.720 158.760 ;
        RECT 147.520 157.060 147.780 157.380 ;
        RECT 145.160 152.105 147.040 152.475 ;
        RECT 144.300 148.560 144.560 148.880 ;
        RECT 143.840 148.220 144.100 148.540 ;
        RECT 142.920 147.880 143.180 148.200 ;
        RECT 130.040 145.500 130.300 145.820 ;
        RECT 132.340 145.500 132.600 145.820 ;
        RECT 140.160 145.500 140.420 145.820 ;
        RECT 140.620 145.500 140.880 145.820 ;
        RECT 128.660 144.820 128.920 145.140 ;
        RECT 128.720 143.100 128.860 144.820 ;
        RECT 130.160 143.945 132.040 144.315 ;
        RECT 132.400 143.780 132.540 145.500 ;
        RECT 142.980 145.480 143.120 147.880 ;
        RECT 143.900 146.160 144.040 148.220 ;
        RECT 143.840 145.840 144.100 146.160 ;
        RECT 142.920 145.160 143.180 145.480 ;
        RECT 141.540 144.820 141.800 145.140 ;
        RECT 132.340 143.460 132.600 143.780 ;
        RECT 128.660 142.780 128.920 143.100 ;
        RECT 128.200 142.440 128.460 142.760 ;
        RECT 125.440 141.760 125.700 142.080 ;
        RECT 128.660 141.760 128.920 142.080 ;
        RECT 132.800 141.760 133.060 142.080 ;
        RECT 136.940 141.760 137.200 142.080 ;
        RECT 141.080 141.760 141.340 142.080 ;
        RECT 125.500 141.140 125.640 141.760 ;
        RECT 124.580 141.000 125.640 141.140 ;
        RECT 124.580 140.690 124.720 141.000 ;
        RECT 128.720 140.690 128.860 141.760 ;
        RECT 132.860 140.690 133.000 141.760 ;
        RECT 137.000 140.690 137.140 141.760 ;
        RECT 141.140 140.690 141.280 141.760 ;
        RECT 141.600 141.060 141.740 144.820 ;
        RECT 143.900 143.100 144.040 145.840 ;
        RECT 143.840 142.780 144.100 143.100 ;
        RECT 144.360 142.760 144.500 148.560 ;
        RECT 145.160 146.665 147.040 147.035 ;
        RECT 145.220 146.180 145.480 146.500 ;
        RECT 144.300 142.440 144.560 142.760 ;
        RECT 145.280 142.500 145.420 146.180 ;
        RECT 144.820 142.360 145.420 142.500 ;
        RECT 141.540 140.740 141.800 141.060 ;
        RECT 144.820 140.970 144.960 142.360 ;
        RECT 145.160 141.225 147.040 141.595 ;
        RECT 144.820 140.830 145.420 140.970 ;
        RECT 145.280 140.690 145.420 140.830 ;
        RECT 124.060 140.060 124.320 140.380 ;
        RECT 124.510 132.440 124.790 140.690 ;
        RECT 128.650 132.440 128.930 140.690 ;
        RECT 105.900 131.400 106.960 132.400 ;
        RECT 116.200 132.160 116.540 132.440 ;
        RECT 120.340 132.160 120.680 132.440 ;
        RECT 124.480 132.160 124.820 132.440 ;
        RECT 128.620 132.160 128.960 132.440 ;
        RECT 132.790 132.130 133.070 140.690 ;
        RECT 136.930 132.130 137.210 140.690 ;
        RECT 141.070 132.130 141.350 140.690 ;
        RECT 142.580 132.400 143.580 134.445 ;
        RECT 142.550 131.400 143.610 132.400 ;
        RECT 145.210 132.170 145.490 140.690 ;
        RECT 146.930 132.400 147.930 134.445 ;
        RECT 146.900 131.400 147.960 132.400 ;
        RECT 60.570 104.080 61.630 105.080 ;
        RECT 101.570 104.080 102.630 105.080 ;
        RECT 142.570 104.080 143.630 105.080 ;
        RECT 30.200 84.600 32.400 85.600 ;
        RECT 30.200 25.000 31.200 84.600 ;
        RECT 60.600 55.000 61.600 104.080 ;
        RECT 101.600 55.000 102.600 104.080 ;
        RECT 142.600 55.000 143.600 104.080 ;
        RECT 146.955 52.570 147.845 52.590 ;
        RECT 143.500 51.630 147.870 52.570 ;
        RECT 146.955 51.610 147.845 51.630 ;
        RECT 130.285 50.340 131.120 50.360 ;
        RECT 126.630 49.455 131.145 50.340 ;
        RECT 130.285 49.435 131.120 49.455 ;
        RECT 126.595 48.130 127.410 48.150 ;
        RECT 122.840 47.265 127.435 48.130 ;
        RECT 126.595 47.245 127.410 47.265 ;
        RECT 30.200 24.000 34.800 25.000 ;
        RECT 24.300 23.000 25.300 23.030 ;
        RECT 20.455 22.000 25.300 23.000 ;
        RECT 24.300 21.970 25.300 22.000 ;
        RECT 31.570 18.065 31.930 18.365 ;
        RECT 22.800 16.615 23.800 16.645 ;
        RECT 20.455 15.615 23.800 16.615 ;
        RECT 31.600 16.015 31.900 18.065 ;
        RECT 31.570 15.715 31.930 16.015 ;
        RECT 22.800 15.585 23.800 15.615 ;
        RECT 31.600 13.765 31.900 15.715 ;
        RECT 31.570 13.465 31.930 13.765 ;
        RECT 33.800 13.670 34.800 24.000 ;
        RECT 30.950 12.365 31.250 12.395 ;
        RECT 29.870 12.065 31.250 12.365 ;
        RECT 30.950 12.035 31.250 12.065 ;
        RECT 35.600 7.675 36.600 9.030 ;
        RECT 35.580 6.725 36.620 7.675 ;
        RECT 35.600 6.700 36.600 6.725 ;
      LAYER via2 ;
        RECT 51.840 222.160 52.120 222.440 ;
        RECT 55.520 222.040 55.800 222.320 ;
        RECT 59.200 222.040 59.480 222.320 ;
        RECT 62.880 222.040 63.160 222.320 ;
        RECT 66.560 222.040 66.840 222.320 ;
        RECT 70.240 222.040 70.520 222.320 ;
        RECT 73.920 222.040 74.200 222.320 ;
        RECT 77.600 222.040 77.880 222.320 ;
        RECT 81.280 222.040 81.560 222.320 ;
        RECT 84.960 222.040 85.240 222.320 ;
        RECT 88.640 222.040 88.920 222.320 ;
        RECT 32.470 214.470 33.130 215.130 ;
        RECT 40.160 214.710 40.440 214.990 ;
        RECT 40.560 214.710 40.840 214.990 ;
        RECT 40.960 214.710 41.240 214.990 ;
        RECT 41.360 214.710 41.640 214.990 ;
        RECT 41.760 214.710 42.040 214.990 ;
        RECT 40.160 209.270 40.440 209.550 ;
        RECT 40.560 209.270 40.840 209.550 ;
        RECT 40.960 209.270 41.240 209.550 ;
        RECT 41.360 209.270 41.640 209.550 ;
        RECT 41.760 209.270 42.040 209.550 ;
        RECT 55.160 211.990 55.440 212.270 ;
        RECT 55.560 211.990 55.840 212.270 ;
        RECT 55.960 211.990 56.240 212.270 ;
        RECT 56.360 211.990 56.640 212.270 ;
        RECT 56.760 211.990 57.040 212.270 ;
        RECT 40.160 203.830 40.440 204.110 ;
        RECT 40.560 203.830 40.840 204.110 ;
        RECT 40.960 203.830 41.240 204.110 ;
        RECT 41.360 203.830 41.640 204.110 ;
        RECT 41.760 203.830 42.040 204.110 ;
        RECT 42.170 202.130 42.450 202.410 ;
        RECT 42.630 200.090 42.910 200.370 ;
        RECT 40.160 198.390 40.440 198.670 ;
        RECT 40.560 198.390 40.840 198.670 ;
        RECT 40.960 198.390 41.240 198.670 ;
        RECT 41.360 198.390 41.640 198.670 ;
        RECT 41.760 198.390 42.040 198.670 ;
        RECT 40.160 192.950 40.440 193.230 ;
        RECT 40.560 192.950 40.840 193.230 ;
        RECT 40.960 192.950 41.240 193.230 ;
        RECT 41.360 192.950 41.640 193.230 ;
        RECT 41.760 192.950 42.040 193.230 ;
        RECT 41.710 189.210 41.990 189.490 ;
        RECT 40.160 187.510 40.440 187.790 ;
        RECT 40.560 187.510 40.840 187.790 ;
        RECT 40.960 187.510 41.240 187.790 ;
        RECT 41.360 187.510 41.640 187.790 ;
        RECT 41.760 187.510 42.040 187.790 ;
        RECT 40.160 182.070 40.440 182.350 ;
        RECT 40.560 182.070 40.840 182.350 ;
        RECT 40.960 182.070 41.240 182.350 ;
        RECT 41.360 182.070 41.640 182.350 ;
        RECT 41.760 182.070 42.040 182.350 ;
        RECT 40.160 176.630 40.440 176.910 ;
        RECT 40.560 176.630 40.840 176.910 ;
        RECT 40.960 176.630 41.240 176.910 ;
        RECT 41.360 176.630 41.640 176.910 ;
        RECT 41.760 176.630 42.040 176.910 ;
        RECT 45.850 200.090 46.130 200.370 ;
        RECT 48.150 202.130 48.430 202.410 ;
        RECT 40.160 171.190 40.440 171.470 ;
        RECT 40.560 171.190 40.840 171.470 ;
        RECT 40.960 171.190 41.240 171.470 ;
        RECT 41.360 171.190 41.640 171.470 ;
        RECT 41.760 171.190 42.040 171.470 ;
        RECT 40.160 165.750 40.440 166.030 ;
        RECT 40.560 165.750 40.840 166.030 ;
        RECT 40.960 165.750 41.240 166.030 ;
        RECT 41.360 165.750 41.640 166.030 ;
        RECT 41.760 165.750 42.040 166.030 ;
        RECT 44.010 181.730 44.290 182.010 ;
        RECT 46.310 197.370 46.590 197.650 ;
        RECT 50.450 197.370 50.730 197.650 ;
        RECT 48.150 196.010 48.430 196.290 ;
        RECT 46.770 191.250 47.050 191.530 ;
        RECT 40.160 160.310 40.440 160.590 ;
        RECT 40.560 160.310 40.840 160.590 ;
        RECT 40.960 160.310 41.240 160.590 ;
        RECT 41.360 160.310 41.640 160.590 ;
        RECT 41.760 160.310 42.040 160.590 ;
        RECT 40.160 154.870 40.440 155.150 ;
        RECT 40.560 154.870 40.840 155.150 ;
        RECT 40.960 154.870 41.240 155.150 ;
        RECT 41.360 154.870 41.640 155.150 ;
        RECT 41.760 154.870 42.040 155.150 ;
        RECT 41.250 153.170 41.530 153.450 ;
        RECT 40.160 149.430 40.440 149.710 ;
        RECT 40.560 149.430 40.840 149.710 ;
        RECT 40.960 149.430 41.240 149.710 ;
        RECT 41.360 149.430 41.640 149.710 ;
        RECT 41.760 149.430 42.040 149.710 ;
        RECT 40.160 143.990 40.440 144.270 ;
        RECT 40.560 143.990 40.840 144.270 ;
        RECT 40.960 143.990 41.240 144.270 ;
        RECT 41.360 143.990 41.640 144.270 ;
        RECT 41.760 143.990 42.040 144.270 ;
        RECT 55.160 206.550 55.440 206.830 ;
        RECT 55.560 206.550 55.840 206.830 ;
        RECT 55.960 206.550 56.240 206.830 ;
        RECT 56.360 206.550 56.640 206.830 ;
        RECT 56.760 206.550 57.040 206.830 ;
        RECT 55.160 201.110 55.440 201.390 ;
        RECT 55.560 201.110 55.840 201.390 ;
        RECT 55.960 201.110 56.240 201.390 ;
        RECT 56.360 201.110 56.640 201.390 ;
        RECT 56.760 201.110 57.040 201.390 ;
        RECT 48.610 181.730 48.890 182.010 ;
        RECT 47.690 175.610 47.970 175.890 ;
        RECT 52.290 186.490 52.570 186.770 ;
        RECT 55.160 195.670 55.440 195.950 ;
        RECT 55.560 195.670 55.840 195.950 ;
        RECT 55.960 195.670 56.240 195.950 ;
        RECT 56.360 195.670 56.640 195.950 ;
        RECT 56.760 195.670 57.040 195.950 ;
        RECT 55.050 193.970 55.330 194.250 ;
        RECT 53.670 188.530 53.950 188.810 ;
        RECT 70.160 214.710 70.440 214.990 ;
        RECT 70.560 214.710 70.840 214.990 ;
        RECT 70.960 214.710 71.240 214.990 ;
        RECT 71.360 214.710 71.640 214.990 ;
        RECT 71.760 214.710 72.040 214.990 ;
        RECT 121.760 221.040 122.040 221.320 ;
        RECT 125.440 221.040 125.720 221.320 ;
        RECT 129.120 221.040 129.400 221.320 ;
        RECT 132.800 221.040 133.080 221.320 ;
        RECT 136.480 221.040 136.760 221.320 ;
        RECT 140.160 221.040 140.440 221.320 ;
        RECT 143.840 221.040 144.120 221.320 ;
        RECT 147.520 221.040 147.800 221.320 ;
        RECT 100.160 214.710 100.440 214.990 ;
        RECT 100.560 214.710 100.840 214.990 ;
        RECT 100.960 214.710 101.240 214.990 ;
        RECT 101.360 214.710 101.640 214.990 ;
        RECT 101.760 214.710 102.040 214.990 ;
        RECT 57.810 194.650 58.090 194.930 ;
        RECT 55.160 190.230 55.440 190.510 ;
        RECT 55.560 190.230 55.840 190.510 ;
        RECT 55.960 190.230 56.240 190.510 ;
        RECT 56.360 190.230 56.640 190.510 ;
        RECT 56.760 190.230 57.040 190.510 ;
        RECT 50.910 178.330 51.190 178.610 ;
        RECT 55.160 184.790 55.440 185.070 ;
        RECT 55.560 184.790 55.840 185.070 ;
        RECT 55.960 184.790 56.240 185.070 ;
        RECT 56.360 184.790 56.640 185.070 ;
        RECT 56.760 184.790 57.040 185.070 ;
        RECT 53.670 175.610 53.950 175.890 ;
        RECT 55.160 179.350 55.440 179.630 ;
        RECT 55.560 179.350 55.840 179.630 ;
        RECT 55.960 179.350 56.240 179.630 ;
        RECT 56.360 179.350 56.640 179.630 ;
        RECT 56.760 179.350 57.040 179.630 ;
        RECT 55.160 173.910 55.440 174.190 ;
        RECT 55.560 173.910 55.840 174.190 ;
        RECT 55.960 173.910 56.240 174.190 ;
        RECT 56.360 173.910 56.640 174.190 ;
        RECT 56.760 173.910 57.040 174.190 ;
        RECT 59.190 196.690 59.470 196.970 ;
        RECT 60.110 195.330 60.390 195.610 ;
        RECT 61.030 175.610 61.310 175.890 ;
        RECT 55.160 168.470 55.440 168.750 ;
        RECT 55.560 168.470 55.840 168.750 ;
        RECT 55.960 168.470 56.240 168.750 ;
        RECT 56.360 168.470 56.640 168.750 ;
        RECT 56.760 168.470 57.040 168.750 ;
        RECT 55.160 163.030 55.440 163.310 ;
        RECT 55.560 163.030 55.840 163.310 ;
        RECT 55.960 163.030 56.240 163.310 ;
        RECT 56.360 163.030 56.640 163.310 ;
        RECT 56.760 163.030 57.040 163.310 ;
        RECT 55.160 157.590 55.440 157.870 ;
        RECT 55.560 157.590 55.840 157.870 ;
        RECT 55.960 157.590 56.240 157.870 ;
        RECT 56.360 157.590 56.640 157.870 ;
        RECT 56.760 157.590 57.040 157.870 ;
        RECT 70.160 209.270 70.440 209.550 ;
        RECT 70.560 209.270 70.840 209.550 ;
        RECT 70.960 209.270 71.240 209.550 ;
        RECT 71.360 209.270 71.640 209.550 ;
        RECT 71.760 209.270 72.040 209.550 ;
        RECT 73.910 204.850 74.190 205.130 ;
        RECT 70.160 203.830 70.440 204.110 ;
        RECT 70.560 203.830 70.840 204.110 ;
        RECT 70.960 203.830 71.240 204.110 ;
        RECT 71.360 203.830 71.640 204.110 ;
        RECT 71.760 203.830 72.040 204.110 ;
        RECT 67.470 196.690 67.750 196.970 ;
        RECT 69.310 193.970 69.590 194.250 ;
        RECT 67.930 190.570 68.210 190.850 ;
        RECT 70.160 198.390 70.440 198.670 ;
        RECT 70.560 198.390 70.840 198.670 ;
        RECT 70.960 198.390 71.240 198.670 ;
        RECT 71.360 198.390 71.640 198.670 ;
        RECT 71.760 198.390 72.040 198.670 ;
        RECT 70.160 192.950 70.440 193.230 ;
        RECT 70.560 192.950 70.840 193.230 ;
        RECT 70.960 192.950 71.240 193.230 ;
        RECT 71.360 192.950 71.640 193.230 ;
        RECT 71.760 192.950 72.040 193.230 ;
        RECT 74.370 191.930 74.650 192.210 ;
        RECT 70.160 187.510 70.440 187.790 ;
        RECT 70.560 187.510 70.840 187.790 ;
        RECT 70.960 187.510 71.240 187.790 ;
        RECT 71.360 187.510 71.640 187.790 ;
        RECT 71.760 187.510 72.040 187.790 ;
        RECT 70.160 182.070 70.440 182.350 ;
        RECT 70.560 182.070 70.840 182.350 ;
        RECT 70.960 182.070 71.240 182.350 ;
        RECT 71.360 182.070 71.640 182.350 ;
        RECT 71.760 182.070 72.040 182.350 ;
        RECT 70.160 176.630 70.440 176.910 ;
        RECT 70.560 176.630 70.840 176.910 ;
        RECT 70.960 176.630 71.240 176.910 ;
        RECT 71.360 176.630 71.640 176.910 ;
        RECT 71.760 176.630 72.040 176.910 ;
        RECT 70.160 171.190 70.440 171.470 ;
        RECT 70.560 171.190 70.840 171.470 ;
        RECT 70.960 171.190 71.240 171.470 ;
        RECT 71.360 171.190 71.640 171.470 ;
        RECT 71.760 171.190 72.040 171.470 ;
        RECT 63.790 161.330 64.070 161.610 ;
        RECT 66.550 156.570 66.830 156.850 ;
        RECT 70.160 165.750 70.440 166.030 ;
        RECT 70.560 165.750 70.840 166.030 ;
        RECT 70.960 165.750 71.240 166.030 ;
        RECT 71.360 165.750 71.640 166.030 ;
        RECT 71.760 165.750 72.040 166.030 ;
        RECT 69.770 164.730 70.050 165.010 ;
        RECT 72.070 161.330 72.350 161.610 ;
        RECT 70.160 160.310 70.440 160.590 ;
        RECT 70.560 160.310 70.840 160.590 ;
        RECT 70.960 160.310 71.240 160.590 ;
        RECT 71.360 160.310 71.640 160.590 ;
        RECT 71.760 160.310 72.040 160.590 ;
        RECT 68.390 155.890 68.670 156.170 ;
        RECT 53.670 151.130 53.950 151.410 ;
        RECT 55.160 152.150 55.440 152.430 ;
        RECT 55.560 152.150 55.840 152.430 ;
        RECT 55.960 152.150 56.240 152.430 ;
        RECT 56.360 152.150 56.640 152.430 ;
        RECT 56.760 152.150 57.040 152.430 ;
        RECT 70.160 154.870 70.440 155.150 ;
        RECT 70.560 154.870 70.840 155.150 ;
        RECT 70.960 154.870 71.240 155.150 ;
        RECT 71.360 154.870 71.640 155.150 ;
        RECT 71.760 154.870 72.040 155.150 ;
        RECT 73.450 157.250 73.730 157.530 ;
        RECT 74.370 166.770 74.650 167.050 ;
        RECT 74.370 162.010 74.650 162.290 ;
        RECT 72.530 153.170 72.810 153.450 ;
        RECT 55.050 147.730 55.330 148.010 ;
        RECT 55.160 146.710 55.440 146.990 ;
        RECT 55.560 146.710 55.840 146.990 ;
        RECT 55.960 146.710 56.240 146.990 ;
        RECT 56.360 146.710 56.640 146.990 ;
        RECT 56.760 146.710 57.040 146.990 ;
        RECT 70.160 149.430 70.440 149.710 ;
        RECT 70.560 149.430 70.840 149.710 ;
        RECT 70.960 149.430 71.240 149.710 ;
        RECT 71.360 149.430 71.640 149.710 ;
        RECT 71.760 149.430 72.040 149.710 ;
        RECT 71.150 148.410 71.430 148.690 ;
        RECT 55.160 141.270 55.440 141.550 ;
        RECT 55.560 141.270 55.840 141.550 ;
        RECT 55.960 141.270 56.240 141.550 ;
        RECT 56.360 141.270 56.640 141.550 ;
        RECT 56.760 141.270 57.040 141.550 ;
        RECT 76.210 149.090 76.490 149.370 ;
        RECT 78.510 187.170 78.790 187.450 ;
        RECT 80.810 202.810 81.090 203.090 ;
        RECT 80.350 190.570 80.630 190.850 ;
        RECT 80.810 180.370 81.090 180.650 ;
        RECT 78.970 178.330 79.250 178.610 ;
        RECT 85.160 211.990 85.440 212.270 ;
        RECT 85.560 211.990 85.840 212.270 ;
        RECT 85.960 211.990 86.240 212.270 ;
        RECT 86.360 211.990 86.640 212.270 ;
        RECT 86.760 211.990 87.040 212.270 ;
        RECT 81.730 202.130 82.010 202.410 ;
        RECT 82.190 198.730 82.470 199.010 ;
        RECT 85.870 207.570 86.150 207.850 ;
        RECT 85.160 206.550 85.440 206.830 ;
        RECT 85.560 206.550 85.840 206.830 ;
        RECT 85.960 206.550 86.240 206.830 ;
        RECT 86.360 206.550 86.640 206.830 ;
        RECT 86.760 206.550 87.040 206.830 ;
        RECT 82.650 182.410 82.930 182.690 ;
        RECT 78.970 157.250 79.250 157.530 ;
        RECT 81.270 175.610 81.550 175.890 ;
        RECT 81.730 172.210 82.010 172.490 ;
        RECT 81.270 169.490 81.550 169.770 ;
        RECT 81.270 157.930 81.550 158.210 ;
        RECT 82.650 181.050 82.930 181.330 ;
        RECT 84.030 200.090 84.310 200.370 ;
        RECT 85.160 201.110 85.440 201.390 ;
        RECT 85.560 201.110 85.840 201.390 ;
        RECT 85.960 201.110 86.240 201.390 ;
        RECT 86.360 201.110 86.640 201.390 ;
        RECT 86.760 201.110 87.040 201.390 ;
        RECT 92.310 204.850 92.590 205.130 ;
        RECT 89.090 202.130 89.370 202.410 ;
        RECT 89.090 201.450 89.370 201.730 ;
        RECT 86.330 199.410 86.610 199.690 ;
        RECT 85.160 195.670 85.440 195.950 ;
        RECT 85.560 195.670 85.840 195.950 ;
        RECT 85.960 195.670 86.240 195.950 ;
        RECT 86.360 195.670 86.640 195.950 ;
        RECT 86.760 195.670 87.040 195.950 ;
        RECT 85.160 190.230 85.440 190.510 ;
        RECT 85.560 190.230 85.840 190.510 ;
        RECT 85.960 190.230 86.240 190.510 ;
        RECT 86.360 190.230 86.640 190.510 ;
        RECT 86.760 190.230 87.040 190.510 ;
        RECT 89.090 195.330 89.370 195.610 ;
        RECT 90.930 200.090 91.210 200.370 ;
        RECT 91.390 198.730 91.670 199.010 ;
        RECT 86.790 185.810 87.070 186.090 ;
        RECT 85.160 184.790 85.440 185.070 ;
        RECT 85.560 184.790 85.840 185.070 ;
        RECT 85.960 184.790 86.240 185.070 ;
        RECT 86.360 184.790 86.640 185.070 ;
        RECT 86.760 184.790 87.040 185.070 ;
        RECT 84.490 183.090 84.770 183.370 ;
        RECT 85.160 179.350 85.440 179.630 ;
        RECT 85.560 179.350 85.840 179.630 ;
        RECT 85.960 179.350 86.240 179.630 ;
        RECT 86.360 179.350 86.640 179.630 ;
        RECT 86.760 179.350 87.040 179.630 ;
        RECT 84.490 176.290 84.770 176.570 ;
        RECT 85.160 173.910 85.440 174.190 ;
        RECT 85.560 173.910 85.840 174.190 ;
        RECT 85.960 173.910 86.240 174.190 ;
        RECT 86.360 173.910 86.640 174.190 ;
        RECT 86.760 173.910 87.040 174.190 ;
        RECT 85.870 171.530 86.150 171.810 ;
        RECT 83.570 165.410 83.850 165.690 ;
        RECT 85.160 168.470 85.440 168.750 ;
        RECT 85.560 168.470 85.840 168.750 ;
        RECT 85.960 168.470 86.240 168.750 ;
        RECT 86.360 168.470 86.640 168.750 ;
        RECT 86.760 168.470 87.040 168.750 ;
        RECT 87.710 170.170 87.990 170.450 ;
        RECT 87.710 168.810 87.990 169.090 ;
        RECT 85.160 163.030 85.440 163.310 ;
        RECT 85.560 163.030 85.840 163.310 ;
        RECT 85.960 163.030 86.240 163.310 ;
        RECT 86.360 163.030 86.640 163.310 ;
        RECT 86.760 163.030 87.040 163.310 ;
        RECT 85.870 161.330 86.150 161.610 ;
        RECT 83.570 157.250 83.850 157.530 ;
        RECT 77.130 149.770 77.410 150.050 ;
        RECT 70.160 143.990 70.440 144.270 ;
        RECT 70.560 143.990 70.840 144.270 ;
        RECT 70.960 143.990 71.240 144.270 ;
        RECT 71.360 143.990 71.640 144.270 ;
        RECT 71.760 143.990 72.040 144.270 ;
        RECT 76.210 145.690 76.490 145.970 ;
        RECT 85.160 157.590 85.440 157.870 ;
        RECT 85.560 157.590 85.840 157.870 ;
        RECT 85.960 157.590 86.240 157.870 ;
        RECT 86.360 157.590 86.640 157.870 ;
        RECT 86.760 157.590 87.040 157.870 ;
        RECT 81.270 155.210 81.550 155.490 ;
        RECT 80.810 154.530 81.090 154.810 ;
        RECT 83.110 154.530 83.390 154.810 ;
        RECT 81.730 153.850 82.010 154.130 ;
        RECT 79.890 152.490 80.170 152.770 ;
        RECT 82.190 152.490 82.470 152.770 ;
        RECT 80.810 151.810 81.090 152.090 ;
        RECT 82.190 151.810 82.470 152.090 ;
        RECT 83.570 151.810 83.850 152.090 ;
        RECT 80.350 150.450 80.630 150.730 ;
        RECT 78.970 148.410 79.250 148.690 ;
        RECT 80.810 147.050 81.090 147.330 ;
        RECT 60.580 133.400 61.580 134.400 ;
        RECT 64.930 133.400 65.930 134.400 ;
        RECT 85.410 154.530 85.690 154.810 ;
        RECT 85.160 152.150 85.440 152.430 ;
        RECT 85.560 152.150 85.840 152.430 ;
        RECT 85.960 152.150 86.240 152.430 ;
        RECT 86.360 152.150 86.640 152.430 ;
        RECT 86.760 152.150 87.040 152.430 ;
        RECT 87.710 148.410 87.990 148.690 ;
        RECT 82.190 142.970 82.470 143.250 ;
        RECT 85.160 146.710 85.440 146.990 ;
        RECT 85.560 146.710 85.840 146.990 ;
        RECT 85.960 146.710 86.240 146.990 ;
        RECT 86.360 146.710 86.640 146.990 ;
        RECT 86.760 146.710 87.040 146.990 ;
        RECT 88.630 164.050 88.910 164.330 ;
        RECT 88.630 155.210 88.910 155.490 ;
        RECT 91.390 189.890 91.670 190.170 ;
        RECT 100.160 209.270 100.440 209.550 ;
        RECT 100.560 209.270 100.840 209.550 ;
        RECT 100.960 209.270 101.240 209.550 ;
        RECT 101.360 209.270 101.640 209.550 ;
        RECT 101.760 209.270 102.040 209.550 ;
        RECT 102.430 208.250 102.710 208.530 ;
        RECT 92.310 183.770 92.590 184.050 ;
        RECT 94.610 190.570 94.890 190.850 ;
        RECT 92.310 174.930 92.590 175.210 ;
        RECT 90.930 173.570 91.210 173.850 ;
        RECT 90.930 172.890 91.210 173.170 ;
        RECT 90.010 168.130 90.290 168.410 ;
        RECT 92.770 173.570 93.050 173.850 ;
        RECT 95.070 185.130 95.350 185.410 ;
        RECT 94.150 176.290 94.430 176.570 ;
        RECT 95.530 179.690 95.810 179.970 ;
        RECT 95.990 179.010 96.270 179.290 ;
        RECT 94.150 173.570 94.430 173.850 ;
        RECT 94.150 171.530 94.430 171.810 ;
        RECT 93.230 168.130 93.510 168.410 ;
        RECT 90.010 163.370 90.290 163.650 ;
        RECT 92.310 153.850 92.590 154.130 ;
        RECT 90.010 150.450 90.290 150.730 ;
        RECT 91.850 149.770 92.130 150.050 ;
        RECT 92.310 149.090 92.590 149.370 ;
        RECT 90.930 145.690 91.210 145.970 ;
        RECT 97.830 202.810 98.110 203.090 ;
        RECT 98.290 197.370 98.570 197.650 ;
        RECT 96.910 185.130 97.190 185.410 ;
        RECT 100.160 203.830 100.440 204.110 ;
        RECT 100.560 203.830 100.840 204.110 ;
        RECT 100.960 203.830 101.240 204.110 ;
        RECT 101.360 203.830 101.640 204.110 ;
        RECT 101.760 203.830 102.040 204.110 ;
        RECT 101.970 201.450 102.250 201.730 ;
        RECT 100.160 198.390 100.440 198.670 ;
        RECT 100.560 198.390 100.840 198.670 ;
        RECT 100.960 198.390 101.240 198.670 ;
        RECT 101.360 198.390 101.640 198.670 ;
        RECT 101.760 198.390 102.040 198.670 ;
        RECT 102.890 195.330 103.170 195.610 ;
        RECT 102.430 193.970 102.710 194.250 ;
        RECT 99.210 189.890 99.490 190.170 ;
        RECT 95.990 172.890 96.270 173.170 ;
        RECT 97.370 166.770 97.650 167.050 ;
        RECT 100.160 192.950 100.440 193.230 ;
        RECT 100.560 192.950 100.840 193.230 ;
        RECT 100.960 192.950 101.240 193.230 ;
        RECT 101.360 192.950 101.640 193.230 ;
        RECT 101.760 192.950 102.040 193.230 ;
        RECT 106.570 207.570 106.850 207.850 ;
        RECT 100.160 187.510 100.440 187.790 ;
        RECT 100.560 187.510 100.840 187.790 ;
        RECT 100.960 187.510 101.240 187.790 ;
        RECT 101.360 187.510 101.640 187.790 ;
        RECT 101.760 187.510 102.040 187.790 ;
        RECT 100.130 184.450 100.410 184.730 ;
        RECT 101.510 183.770 101.790 184.050 ;
        RECT 100.160 182.070 100.440 182.350 ;
        RECT 100.560 182.070 100.840 182.350 ;
        RECT 100.960 182.070 101.240 182.350 ;
        RECT 101.360 182.070 101.640 182.350 ;
        RECT 101.760 182.070 102.040 182.350 ;
        RECT 101.970 178.330 102.250 178.610 ;
        RECT 100.160 176.630 100.440 176.910 ;
        RECT 100.560 176.630 100.840 176.910 ;
        RECT 100.960 176.630 101.240 176.910 ;
        RECT 101.360 176.630 101.640 176.910 ;
        RECT 101.760 176.630 102.040 176.910 ;
        RECT 98.290 162.690 98.570 162.970 ;
        RECT 103.350 179.010 103.630 179.290 ;
        RECT 101.510 172.210 101.790 172.490 ;
        RECT 100.160 171.190 100.440 171.470 ;
        RECT 100.560 171.190 100.840 171.470 ;
        RECT 100.960 171.190 101.240 171.470 ;
        RECT 101.360 171.190 101.640 171.470 ;
        RECT 101.760 171.190 102.040 171.470 ;
        RECT 104.270 176.290 104.550 176.570 ;
        RECT 104.270 174.930 104.550 175.210 ;
        RECT 102.890 170.850 103.170 171.130 ;
        RECT 103.810 170.170 104.090 170.450 ;
        RECT 99.670 166.770 99.950 167.050 ;
        RECT 100.160 165.750 100.440 166.030 ;
        RECT 100.560 165.750 100.840 166.030 ;
        RECT 100.960 165.750 101.240 166.030 ;
        RECT 101.360 165.750 101.640 166.030 ;
        RECT 101.760 165.750 102.040 166.030 ;
        RECT 99.210 164.050 99.490 164.330 ;
        RECT 97.370 158.610 97.650 158.890 ;
        RECT 101.510 163.370 101.790 163.650 ;
        RECT 100.160 160.310 100.440 160.590 ;
        RECT 100.560 160.310 100.840 160.590 ;
        RECT 100.960 160.310 101.240 160.590 ;
        RECT 101.360 160.310 101.640 160.590 ;
        RECT 101.760 160.310 102.040 160.590 ;
        RECT 100.590 159.290 100.870 159.570 ;
        RECT 95.070 153.170 95.350 153.450 ;
        RECT 98.290 151.810 98.570 152.090 ;
        RECT 100.160 154.870 100.440 155.150 ;
        RECT 100.560 154.870 100.840 155.150 ;
        RECT 100.960 154.870 101.240 155.150 ;
        RECT 101.360 154.870 101.640 155.150 ;
        RECT 101.760 154.870 102.040 155.150 ;
        RECT 101.050 151.810 101.330 152.090 ;
        RECT 100.160 149.430 100.440 149.710 ;
        RECT 100.560 149.430 100.840 149.710 ;
        RECT 100.960 149.430 101.240 149.710 ;
        RECT 101.360 149.430 101.640 149.710 ;
        RECT 101.760 149.430 102.040 149.710 ;
        RECT 100.130 146.370 100.410 146.650 ;
        RECT 85.160 141.270 85.440 141.550 ;
        RECT 85.560 141.270 85.840 141.550 ;
        RECT 85.960 141.270 86.240 141.550 ;
        RECT 86.360 141.270 86.640 141.550 ;
        RECT 86.760 141.270 87.040 141.550 ;
        RECT 106.570 201.450 106.850 201.730 ;
        RECT 106.570 195.330 106.850 195.610 ;
        RECT 106.110 190.570 106.390 190.850 ;
        RECT 107.030 189.890 107.310 190.170 ;
        RECT 106.570 183.770 106.850 184.050 ;
        RECT 108.410 182.410 108.690 182.690 ;
        RECT 107.490 176.290 107.770 176.570 ;
        RECT 107.030 168.810 107.310 169.090 ;
        RECT 107.030 167.450 107.310 167.730 ;
        RECT 112.550 210.290 112.830 210.570 ;
        RECT 115.160 211.990 115.440 212.270 ;
        RECT 115.560 211.990 115.840 212.270 ;
        RECT 115.960 211.990 116.240 212.270 ;
        RECT 116.360 211.990 116.640 212.270 ;
        RECT 116.760 211.990 117.040 212.270 ;
        RECT 112.550 206.890 112.830 207.170 ;
        RECT 115.160 206.550 115.440 206.830 ;
        RECT 115.560 206.550 115.840 206.830 ;
        RECT 115.960 206.550 116.240 206.830 ;
        RECT 116.360 206.550 116.640 206.830 ;
        RECT 116.760 206.550 117.040 206.830 ;
        RECT 115.160 201.110 115.440 201.390 ;
        RECT 115.560 201.110 115.840 201.390 ;
        RECT 115.960 201.110 116.240 201.390 ;
        RECT 116.360 201.110 116.640 201.390 ;
        RECT 116.760 201.110 117.040 201.390 ;
        RECT 112.550 200.770 112.830 201.050 ;
        RECT 113.470 197.370 113.750 197.650 ;
        RECT 117.150 197.370 117.430 197.650 ;
        RECT 115.160 195.670 115.440 195.950 ;
        RECT 115.560 195.670 115.840 195.950 ;
        RECT 115.960 195.670 116.240 195.950 ;
        RECT 116.360 195.670 116.640 195.950 ;
        RECT 116.760 195.670 117.040 195.950 ;
        RECT 115.160 190.230 115.440 190.510 ;
        RECT 115.560 190.230 115.840 190.510 ;
        RECT 115.960 190.230 116.240 190.510 ;
        RECT 116.360 190.230 116.640 190.510 ;
        RECT 116.760 190.230 117.040 190.510 ;
        RECT 117.610 191.250 117.890 191.530 ;
        RECT 110.250 183.770 110.530 184.050 ;
        RECT 110.710 181.050 110.990 181.330 ;
        RECT 109.790 174.930 110.070 175.210 ;
        RECT 106.570 153.850 106.850 154.130 ;
        RECT 107.490 153.170 107.770 153.450 ;
        RECT 111.630 179.690 111.910 179.970 ;
        RECT 110.710 164.730 110.990 165.010 ;
        RECT 107.950 149.090 108.230 149.370 ;
        RECT 113.470 182.410 113.750 182.690 ;
        RECT 113.010 170.850 113.290 171.130 ;
        RECT 113.010 166.090 113.290 166.370 ;
        RECT 116.690 185.810 116.970 186.090 ;
        RECT 115.160 184.790 115.440 185.070 ;
        RECT 115.560 184.790 115.840 185.070 ;
        RECT 115.960 184.790 116.240 185.070 ;
        RECT 116.360 184.790 116.640 185.070 ;
        RECT 116.760 184.790 117.040 185.070 ;
        RECT 116.230 180.370 116.510 180.650 ;
        RECT 115.160 179.350 115.440 179.630 ;
        RECT 115.560 179.350 115.840 179.630 ;
        RECT 115.960 179.350 116.240 179.630 ;
        RECT 116.360 179.350 116.640 179.630 ;
        RECT 116.760 179.350 117.040 179.630 ;
        RECT 115.160 173.910 115.440 174.190 ;
        RECT 115.560 173.910 115.840 174.190 ;
        RECT 115.960 173.910 116.240 174.190 ;
        RECT 116.360 173.910 116.640 174.190 ;
        RECT 116.760 173.910 117.040 174.190 ;
        RECT 114.390 173.570 114.670 173.850 ;
        RECT 110.710 161.330 110.990 161.610 ;
        RECT 111.170 155.210 111.450 155.490 ;
        RECT 112.090 153.850 112.370 154.130 ;
        RECT 100.160 143.990 100.440 144.270 ;
        RECT 100.560 143.990 100.840 144.270 ;
        RECT 100.960 143.990 101.240 144.270 ;
        RECT 101.360 143.990 101.640 144.270 ;
        RECT 101.760 143.990 102.040 144.270 ;
        RECT 101.580 133.400 102.580 134.400 ;
        RECT 111.630 149.090 111.910 149.370 ;
        RECT 111.630 146.370 111.910 146.650 ;
        RECT 113.470 161.330 113.750 161.610 ;
        RECT 113.010 149.770 113.290 150.050 ;
        RECT 115.160 168.470 115.440 168.750 ;
        RECT 115.560 168.470 115.840 168.750 ;
        RECT 115.960 168.470 116.240 168.750 ;
        RECT 116.360 168.470 116.640 168.750 ;
        RECT 116.760 168.470 117.040 168.750 ;
        RECT 118.990 210.290 119.270 210.570 ;
        RECT 118.990 191.930 119.270 192.210 ;
        RECT 123.130 210.970 123.410 211.250 ;
        RECT 120.370 199.410 120.650 199.690 ;
        RECT 119.450 181.730 119.730 182.010 ;
        RECT 119.910 181.050 120.190 181.330 ;
        RECT 118.070 166.090 118.350 166.370 ;
        RECT 118.070 164.050 118.350 164.330 ;
        RECT 115.160 163.030 115.440 163.310 ;
        RECT 115.560 163.030 115.840 163.310 ;
        RECT 115.960 163.030 116.240 163.310 ;
        RECT 116.360 163.030 116.640 163.310 ;
        RECT 116.760 163.030 117.040 163.310 ;
        RECT 115.160 157.590 115.440 157.870 ;
        RECT 115.560 157.590 115.840 157.870 ;
        RECT 115.960 157.590 116.240 157.870 ;
        RECT 116.360 157.590 116.640 157.870 ;
        RECT 116.760 157.590 117.040 157.870 ;
        RECT 116.230 155.890 116.510 156.170 ;
        RECT 115.310 155.210 115.590 155.490 ;
        RECT 114.390 153.850 114.670 154.130 ;
        RECT 115.160 152.150 115.440 152.430 ;
        RECT 115.560 152.150 115.840 152.430 ;
        RECT 115.960 152.150 116.240 152.430 ;
        RECT 116.360 152.150 116.640 152.430 ;
        RECT 116.760 152.150 117.040 152.430 ;
        RECT 113.930 149.090 114.210 149.370 ;
        RECT 115.160 146.710 115.440 146.990 ;
        RECT 115.560 146.710 115.840 146.990 ;
        RECT 115.960 146.710 116.240 146.990 ;
        RECT 116.360 146.710 116.640 146.990 ;
        RECT 116.760 146.710 117.040 146.990 ;
        RECT 115.310 145.690 115.590 145.970 ;
        RECT 118.530 162.010 118.810 162.290 ;
        RECT 130.160 214.710 130.440 214.990 ;
        RECT 130.560 214.710 130.840 214.990 ;
        RECT 130.960 214.710 131.240 214.990 ;
        RECT 131.360 214.710 131.640 214.990 ;
        RECT 131.760 214.710 132.040 214.990 ;
        RECT 127.730 210.970 128.010 211.250 ;
        RECT 126.350 208.250 126.630 208.530 ;
        RECT 126.350 207.570 126.630 207.850 ;
        RECT 130.160 209.270 130.440 209.550 ;
        RECT 130.560 209.270 130.840 209.550 ;
        RECT 130.960 209.270 131.240 209.550 ;
        RECT 131.360 209.270 131.640 209.550 ;
        RECT 131.760 209.270 132.040 209.550 ;
        RECT 133.710 208.250 133.990 208.530 ;
        RECT 127.730 205.530 128.010 205.810 ;
        RECT 130.160 203.830 130.440 204.110 ;
        RECT 130.560 203.830 130.840 204.110 ;
        RECT 130.960 203.830 131.240 204.110 ;
        RECT 131.360 203.830 131.640 204.110 ;
        RECT 131.760 203.830 132.040 204.110 ;
        RECT 123.130 193.970 123.410 194.250 ;
        RECT 122.210 185.810 122.490 186.090 ;
        RECT 122.210 181.730 122.490 182.010 ;
        RECT 122.210 181.050 122.490 181.330 ;
        RECT 120.830 178.330 121.110 178.610 ;
        RECT 120.370 175.610 120.650 175.890 ;
        RECT 119.910 172.890 120.190 173.170 ;
        RECT 118.990 148.410 119.270 148.690 ;
        RECT 121.750 174.930 122.030 175.210 ;
        RECT 120.830 149.770 121.110 150.050 ;
        RECT 123.130 155.890 123.410 156.170 ;
        RECT 124.970 200.090 125.250 200.370 ;
        RECT 124.970 177.650 125.250 177.930 ;
        RECT 127.270 180.370 127.550 180.650 ;
        RECT 124.510 151.810 124.790 152.090 ;
        RECT 125.890 159.290 126.170 159.570 ;
        RECT 125.890 158.610 126.170 158.890 ;
        RECT 126.350 155.890 126.630 156.170 ;
        RECT 127.730 156.570 128.010 156.850 ;
        RECT 130.160 198.390 130.440 198.670 ;
        RECT 130.560 198.390 130.840 198.670 ;
        RECT 130.960 198.390 131.240 198.670 ;
        RECT 131.360 198.390 131.640 198.670 ;
        RECT 131.760 198.390 132.040 198.670 ;
        RECT 131.870 193.970 132.150 194.250 ;
        RECT 130.160 192.950 130.440 193.230 ;
        RECT 130.560 192.950 130.840 193.230 ;
        RECT 130.960 192.950 131.240 193.230 ;
        RECT 131.360 192.950 131.640 193.230 ;
        RECT 131.760 192.950 132.040 193.230 ;
        RECT 145.160 211.990 145.440 212.270 ;
        RECT 145.560 211.990 145.840 212.270 ;
        RECT 145.960 211.990 146.240 212.270 ;
        RECT 146.360 211.990 146.640 212.270 ;
        RECT 146.760 211.990 147.040 212.270 ;
        RECT 145.160 206.550 145.440 206.830 ;
        RECT 145.560 206.550 145.840 206.830 ;
        RECT 145.960 206.550 146.240 206.830 ;
        RECT 146.360 206.550 146.640 206.830 ;
        RECT 146.760 206.550 147.040 206.830 ;
        RECT 128.650 189.210 128.930 189.490 ;
        RECT 130.030 188.530 130.310 188.810 ;
        RECT 130.160 187.510 130.440 187.790 ;
        RECT 130.560 187.510 130.840 187.790 ;
        RECT 130.960 187.510 131.240 187.790 ;
        RECT 131.360 187.510 131.640 187.790 ;
        RECT 131.760 187.510 132.040 187.790 ;
        RECT 132.790 187.850 133.070 188.130 ;
        RECT 130.030 186.490 130.310 186.770 ;
        RECT 130.490 184.450 130.770 184.730 ;
        RECT 131.870 183.770 132.150 184.050 ;
        RECT 133.250 186.490 133.530 186.770 ;
        RECT 130.160 182.070 130.440 182.350 ;
        RECT 130.560 182.070 130.840 182.350 ;
        RECT 130.960 182.070 131.240 182.350 ;
        RECT 131.360 182.070 131.640 182.350 ;
        RECT 131.760 182.070 132.040 182.350 ;
        RECT 130.160 176.630 130.440 176.910 ;
        RECT 130.560 176.630 130.840 176.910 ;
        RECT 130.960 176.630 131.240 176.910 ;
        RECT 131.360 176.630 131.640 176.910 ;
        RECT 131.760 176.630 132.040 176.910 ;
        RECT 130.160 171.190 130.440 171.470 ;
        RECT 130.560 171.190 130.840 171.470 ;
        RECT 130.960 171.190 131.240 171.470 ;
        RECT 131.360 171.190 131.640 171.470 ;
        RECT 131.760 171.190 132.040 171.470 ;
        RECT 130.160 165.750 130.440 166.030 ;
        RECT 130.560 165.750 130.840 166.030 ;
        RECT 130.960 165.750 131.240 166.030 ;
        RECT 131.360 165.750 131.640 166.030 ;
        RECT 131.760 165.750 132.040 166.030 ;
        RECT 131.410 161.330 131.690 161.610 ;
        RECT 130.160 160.310 130.440 160.590 ;
        RECT 130.560 160.310 130.840 160.590 ;
        RECT 130.960 160.310 131.240 160.590 ;
        RECT 131.360 160.310 131.640 160.590 ;
        RECT 131.760 160.310 132.040 160.590 ;
        RECT 134.630 186.490 134.910 186.770 ;
        RECT 133.250 179.690 133.530 179.970 ;
        RECT 134.630 179.690 134.910 179.970 ;
        RECT 136.930 196.690 137.210 196.970 ;
        RECT 136.470 193.970 136.750 194.250 ;
        RECT 149.810 202.810 150.090 203.090 ;
        RECT 138.310 187.850 138.590 188.130 ;
        RECT 133.250 169.490 133.530 169.770 ;
        RECT 133.250 156.570 133.530 156.850 ;
        RECT 130.160 154.870 130.440 155.150 ;
        RECT 130.560 154.870 130.840 155.150 ;
        RECT 130.960 154.870 131.240 155.150 ;
        RECT 131.360 154.870 131.640 155.150 ;
        RECT 131.760 154.870 132.040 155.150 ;
        RECT 131.870 153.170 132.150 153.450 ;
        RECT 139.690 186.490 139.970 186.770 ;
        RECT 138.770 185.810 139.050 186.090 ;
        RECT 137.390 183.090 137.670 183.370 ;
        RECT 136.930 180.370 137.210 180.650 ;
        RECT 140.150 183.770 140.430 184.050 ;
        RECT 139.690 179.690 139.970 179.970 ;
        RECT 140.150 166.770 140.430 167.050 ;
        RECT 141.530 186.490 141.810 186.770 ;
        RECT 141.530 181.050 141.810 181.330 ;
        RECT 145.160 201.110 145.440 201.390 ;
        RECT 145.560 201.110 145.840 201.390 ;
        RECT 145.960 201.110 146.240 201.390 ;
        RECT 146.360 201.110 146.640 201.390 ;
        RECT 146.760 201.110 147.040 201.390 ;
        RECT 145.160 195.670 145.440 195.950 ;
        RECT 145.560 195.670 145.840 195.950 ;
        RECT 145.960 195.670 146.240 195.950 ;
        RECT 146.360 195.670 146.640 195.950 ;
        RECT 146.760 195.670 147.040 195.950 ;
        RECT 145.160 190.230 145.440 190.510 ;
        RECT 145.560 190.230 145.840 190.510 ;
        RECT 145.960 190.230 146.240 190.510 ;
        RECT 146.360 190.230 146.640 190.510 ;
        RECT 146.760 190.230 147.040 190.510 ;
        RECT 143.830 185.810 144.110 186.090 ;
        RECT 145.160 184.790 145.440 185.070 ;
        RECT 145.560 184.790 145.840 185.070 ;
        RECT 145.960 184.790 146.240 185.070 ;
        RECT 146.360 184.790 146.640 185.070 ;
        RECT 146.760 184.790 147.040 185.070 ;
        RECT 145.160 179.350 145.440 179.630 ;
        RECT 145.560 179.350 145.840 179.630 ;
        RECT 145.960 179.350 146.240 179.630 ;
        RECT 146.360 179.350 146.640 179.630 ;
        RECT 146.760 179.350 147.040 179.630 ;
        RECT 145.160 173.910 145.440 174.190 ;
        RECT 145.560 173.910 145.840 174.190 ;
        RECT 145.960 173.910 146.240 174.190 ;
        RECT 146.360 173.910 146.640 174.190 ;
        RECT 146.760 173.910 147.040 174.190 ;
        RECT 145.160 168.470 145.440 168.750 ;
        RECT 145.560 168.470 145.840 168.750 ;
        RECT 145.960 168.470 146.240 168.750 ;
        RECT 146.360 168.470 146.640 168.750 ;
        RECT 146.760 168.470 147.040 168.750 ;
        RECT 127.730 150.450 128.010 150.730 ;
        RECT 115.160 141.270 115.440 141.550 ;
        RECT 115.560 141.270 115.840 141.550 ;
        RECT 115.960 141.270 116.240 141.550 ;
        RECT 116.360 141.270 116.640 141.550 ;
        RECT 116.760 141.270 117.040 141.550 ;
        RECT 105.930 133.400 106.930 134.400 ;
        RECT 125.430 147.730 125.710 148.010 ;
        RECT 130.160 149.430 130.440 149.710 ;
        RECT 130.560 149.430 130.840 149.710 ;
        RECT 130.960 149.430 131.240 149.710 ;
        RECT 131.360 149.430 131.640 149.710 ;
        RECT 131.760 149.430 132.040 149.710 ;
        RECT 140.610 161.330 140.890 161.610 ;
        RECT 145.160 163.030 145.440 163.310 ;
        RECT 145.560 163.030 145.840 163.310 ;
        RECT 145.960 163.030 146.240 163.310 ;
        RECT 146.360 163.030 146.640 163.310 ;
        RECT 146.760 163.030 147.040 163.310 ;
        RECT 141.070 156.570 141.350 156.850 ;
        RECT 140.610 151.130 140.890 151.410 ;
        RECT 145.160 157.590 145.440 157.870 ;
        RECT 145.560 157.590 145.840 157.870 ;
        RECT 145.960 157.590 146.240 157.870 ;
        RECT 146.360 157.590 146.640 157.870 ;
        RECT 146.760 157.590 147.040 157.870 ;
        RECT 145.160 152.150 145.440 152.430 ;
        RECT 145.560 152.150 145.840 152.430 ;
        RECT 145.960 152.150 146.240 152.430 ;
        RECT 146.360 152.150 146.640 152.430 ;
        RECT 146.760 152.150 147.040 152.430 ;
        RECT 130.160 143.990 130.440 144.270 ;
        RECT 130.560 143.990 130.840 144.270 ;
        RECT 130.960 143.990 131.240 144.270 ;
        RECT 131.360 143.990 131.640 144.270 ;
        RECT 131.760 143.990 132.040 144.270 ;
        RECT 145.160 146.710 145.440 146.990 ;
        RECT 145.560 146.710 145.840 146.990 ;
        RECT 145.960 146.710 146.240 146.990 ;
        RECT 146.360 146.710 146.640 146.990 ;
        RECT 146.760 146.710 147.040 146.990 ;
        RECT 145.160 141.270 145.440 141.550 ;
        RECT 145.560 141.270 145.840 141.550 ;
        RECT 145.960 141.270 146.240 141.550 ;
        RECT 146.360 141.270 146.640 141.550 ;
        RECT 146.760 141.270 147.040 141.550 ;
        RECT 142.580 133.400 143.580 134.400 ;
        RECT 146.930 133.400 147.930 134.400 ;
        RECT 146.955 51.655 147.845 52.545 ;
        RECT 130.285 49.480 131.120 50.315 ;
        RECT 126.595 47.290 127.410 48.105 ;
        RECT 20.500 22.000 21.500 23.000 ;
        RECT 20.500 15.615 21.500 16.615 ;
        RECT 35.625 6.725 36.575 7.675 ;
      LAYER met3 ;
        RECT 32.470 223.905 33.130 224.030 ;
        RECT 92.160 223.905 92.640 223.975 ;
        RECT 32.470 223.500 92.640 223.905 ;
        RECT 31.350 222.295 31.850 222.300 ;
        RECT 31.325 221.805 31.875 222.295 ;
        RECT 31.350 221.050 31.850 221.805 ;
        RECT 20.620 220.550 31.850 221.050 ;
        RECT 9.305 218.400 9.695 218.425 ;
        RECT 9.300 218.000 13.030 218.400 ;
        RECT 9.305 217.975 9.695 218.000 ;
        RECT 32.470 215.155 33.130 223.500 ;
        RECT 92.160 223.435 92.640 223.500 ;
        RECT 51.790 222.840 52.170 223.160 ;
        RECT 51.830 222.465 52.130 222.840 ;
        RECT 55.470 222.770 55.850 223.090 ;
        RECT 59.150 222.770 59.530 223.090 ;
        RECT 62.830 222.770 63.210 223.090 ;
        RECT 66.510 222.770 66.890 223.090 ;
        RECT 70.190 222.770 70.570 223.090 ;
        RECT 73.870 222.770 74.250 223.090 ;
        RECT 77.550 222.770 77.930 223.090 ;
        RECT 81.230 222.770 81.610 223.090 ;
        RECT 84.910 222.770 85.290 223.090 ;
        RECT 88.590 222.770 88.970 223.090 ;
        RECT 121.710 222.770 122.090 223.090 ;
        RECT 125.390 222.770 125.770 223.090 ;
        RECT 129.070 222.770 129.450 223.090 ;
        RECT 132.750 222.770 133.130 223.090 ;
        RECT 136.430 222.770 136.810 223.090 ;
        RECT 140.110 222.770 140.490 223.090 ;
        RECT 143.790 222.770 144.170 223.090 ;
        RECT 147.470 222.770 147.850 223.090 ;
        RECT 51.815 222.135 52.145 222.465 ;
        RECT 55.510 222.345 55.810 222.770 ;
        RECT 59.190 222.345 59.490 222.770 ;
        RECT 62.870 222.345 63.170 222.770 ;
        RECT 66.550 222.345 66.850 222.770 ;
        RECT 70.230 222.345 70.530 222.770 ;
        RECT 73.910 222.345 74.210 222.770 ;
        RECT 77.590 222.345 77.890 222.770 ;
        RECT 81.270 222.345 81.570 222.770 ;
        RECT 84.950 222.345 85.250 222.770 ;
        RECT 88.630 222.345 88.930 222.770 ;
        RECT 55.495 222.015 55.825 222.345 ;
        RECT 59.175 222.015 59.505 222.345 ;
        RECT 62.855 222.015 63.185 222.345 ;
        RECT 66.535 222.015 66.865 222.345 ;
        RECT 70.215 222.015 70.545 222.345 ;
        RECT 73.895 222.015 74.225 222.345 ;
        RECT 77.575 222.015 77.905 222.345 ;
        RECT 81.255 222.015 81.585 222.345 ;
        RECT 84.935 222.015 85.265 222.345 ;
        RECT 88.615 222.015 88.945 222.345 ;
        RECT 55.510 221.600 55.810 222.015 ;
        RECT 59.190 221.600 59.490 222.015 ;
        RECT 62.870 221.600 63.170 222.015 ;
        RECT 66.550 221.600 66.850 222.015 ;
        RECT 70.230 221.600 70.530 222.015 ;
        RECT 73.910 221.600 74.210 222.015 ;
        RECT 77.590 221.600 77.890 222.015 ;
        RECT 81.270 221.600 81.570 222.015 ;
        RECT 84.950 221.600 85.250 222.015 ;
        RECT 88.630 221.600 88.930 222.015 ;
        RECT 121.750 221.345 122.050 222.770 ;
        RECT 125.430 221.345 125.730 222.770 ;
        RECT 129.110 221.345 129.410 222.770 ;
        RECT 132.790 221.345 133.090 222.770 ;
        RECT 136.470 221.345 136.770 222.770 ;
        RECT 140.150 221.345 140.450 222.770 ;
        RECT 143.830 221.345 144.130 222.770 ;
        RECT 147.510 221.345 147.810 222.770 ;
        RECT 121.735 221.015 122.065 221.345 ;
        RECT 125.415 221.015 125.745 221.345 ;
        RECT 129.095 221.015 129.425 221.345 ;
        RECT 132.775 221.015 133.105 221.345 ;
        RECT 136.455 221.015 136.785 221.345 ;
        RECT 140.135 221.015 140.465 221.345 ;
        RECT 143.815 221.015 144.145 221.345 ;
        RECT 147.495 221.015 147.825 221.345 ;
        RECT 95.940 220.705 96.340 220.730 ;
        RECT 95.195 220.295 96.345 220.705 ;
        RECT 95.940 220.270 96.340 220.295 ;
        RECT 99.625 219.905 100.020 219.930 ;
        RECT 95.200 219.500 100.025 219.905 ;
        RECT 99.625 219.475 100.020 219.500 ;
        RECT 103.310 219.100 103.695 219.125 ;
        RECT 95.205 218.705 103.700 219.100 ;
        RECT 103.310 218.680 103.695 218.705 ;
        RECT 106.985 218.300 107.375 218.325 ;
        RECT 95.200 217.900 107.380 218.300 ;
        RECT 106.985 217.875 107.375 217.900 ;
        RECT 32.445 214.445 33.155 215.155 ;
        RECT 40.110 214.685 42.090 215.015 ;
        RECT 70.110 214.685 72.090 215.015 ;
        RECT 100.110 214.685 102.090 215.015 ;
        RECT 130.110 214.685 132.090 215.015 ;
        RECT 55.110 211.965 57.090 212.295 ;
        RECT 85.110 211.965 87.090 212.295 ;
        RECT 115.110 211.965 117.090 212.295 ;
        RECT 145.110 211.965 147.090 212.295 ;
        RECT 154.820 211.695 155.220 211.700 ;
        RECT 154.795 211.305 155.245 211.695 ;
        RECT 123.105 211.260 123.435 211.275 ;
        RECT 127.705 211.260 128.035 211.275 ;
        RECT 123.105 210.960 128.035 211.260 ;
        RECT 123.105 210.945 123.435 210.960 ;
        RECT 127.705 210.945 128.035 210.960 ;
        RECT 112.525 210.580 112.855 210.595 ;
        RECT 118.965 210.580 119.295 210.595 ;
        RECT 112.525 210.280 119.295 210.580 ;
        RECT 112.525 210.265 112.855 210.280 ;
        RECT 118.965 210.265 119.295 210.280 ;
        RECT 40.110 209.245 42.090 209.575 ;
        RECT 70.110 209.245 72.090 209.575 ;
        RECT 100.110 209.245 102.090 209.575 ;
        RECT 130.110 209.245 132.090 209.575 ;
        RECT 151.340 208.610 153.340 208.690 ;
        RECT 154.820 208.610 155.220 211.305 ;
        RECT 102.405 208.540 102.735 208.555 ;
        RECT 126.325 208.540 126.655 208.555 ;
        RECT 102.405 208.240 126.655 208.540 ;
        RECT 102.405 208.225 102.735 208.240 ;
        RECT 126.325 208.225 126.655 208.240 ;
        RECT 133.685 208.540 134.015 208.555 ;
        RECT 151.340 208.540 155.220 208.610 ;
        RECT 133.685 208.240 155.220 208.540 ;
        RECT 133.685 208.225 134.015 208.240 ;
        RECT 151.340 208.210 155.220 208.240 ;
        RECT 151.340 208.090 153.340 208.210 ;
        RECT 85.845 207.860 86.175 207.875 ;
        RECT 106.545 207.860 106.875 207.875 ;
        RECT 126.325 207.860 126.655 207.875 ;
        RECT 85.845 207.560 105.710 207.860 ;
        RECT 85.845 207.545 86.175 207.560 ;
        RECT 105.410 207.180 105.710 207.560 ;
        RECT 106.545 207.560 126.655 207.860 ;
        RECT 106.545 207.545 106.875 207.560 ;
        RECT 126.325 207.545 126.655 207.560 ;
        RECT 112.525 207.180 112.855 207.195 ;
        RECT 105.410 206.880 112.855 207.180 ;
        RECT 112.525 206.865 112.855 206.880 ;
        RECT 55.110 206.525 57.090 206.855 ;
        RECT 85.110 206.525 87.090 206.855 ;
        RECT 115.110 206.525 117.090 206.855 ;
        RECT 145.110 206.525 147.090 206.855 ;
        RECT 154.020 206.005 154.380 206.010 ;
        RECT 98.930 205.820 99.310 205.830 ;
        RECT 127.705 205.820 128.035 205.835 ;
        RECT 98.930 205.520 128.035 205.820 ;
        RECT 153.995 205.655 154.405 206.005 ;
        RECT 98.930 205.510 99.310 205.520 ;
        RECT 127.705 205.505 128.035 205.520 ;
        RECT 73.885 205.140 74.215 205.155 ;
        RECT 92.285 205.140 92.615 205.155 ;
        RECT 73.885 204.840 92.615 205.140 ;
        RECT 73.885 204.825 74.215 204.840 ;
        RECT 92.285 204.825 92.615 204.840 ;
        RECT 40.110 203.805 42.090 204.135 ;
        RECT 70.110 203.805 72.090 204.135 ;
        RECT 100.110 203.805 102.090 204.135 ;
        RECT 130.110 203.805 132.090 204.135 ;
        RECT 80.785 203.100 81.115 203.115 ;
        RECT 97.805 203.100 98.135 203.115 ;
        RECT 111.810 203.100 112.190 203.110 ;
        RECT 80.785 202.800 112.190 203.100 ;
        RECT 80.785 202.785 81.115 202.800 ;
        RECT 97.805 202.785 98.135 202.800 ;
        RECT 111.810 202.790 112.190 202.800 ;
        RECT 149.785 203.100 150.115 203.115 ;
        RECT 151.340 203.100 153.340 203.250 ;
        RECT 154.020 203.100 154.380 205.655 ;
        RECT 149.785 202.800 154.380 203.100 ;
        RECT 149.785 202.785 150.115 202.800 ;
        RECT 151.340 202.740 154.380 202.800 ;
        RECT 151.340 202.650 153.340 202.740 ;
        RECT 42.145 202.420 42.475 202.435 ;
        RECT 48.125 202.420 48.455 202.435 ;
        RECT 42.145 202.120 48.455 202.420 ;
        RECT 42.145 202.105 42.475 202.120 ;
        RECT 48.125 202.105 48.455 202.120 ;
        RECT 81.705 202.420 82.035 202.435 ;
        RECT 89.065 202.420 89.395 202.435 ;
        RECT 81.705 202.120 89.395 202.420 ;
        RECT 81.705 202.105 82.035 202.120 ;
        RECT 89.065 202.105 89.395 202.120 ;
        RECT 89.065 201.740 89.395 201.755 ;
        RECT 101.945 201.740 102.275 201.755 ;
        RECT 89.065 201.440 102.275 201.740 ;
        RECT 89.065 201.425 89.395 201.440 ;
        RECT 101.945 201.425 102.275 201.440 ;
        RECT 106.545 201.740 106.875 201.755 ;
        RECT 108.130 201.740 108.510 201.750 ;
        RECT 106.545 201.440 108.510 201.740 ;
        RECT 106.545 201.425 106.875 201.440 ;
        RECT 108.130 201.430 108.510 201.440 ;
        RECT 55.110 201.085 57.090 201.415 ;
        RECT 85.110 201.085 87.090 201.415 ;
        RECT 115.110 201.085 117.090 201.415 ;
        RECT 145.110 201.085 147.090 201.415 ;
        RECT 112.525 201.060 112.855 201.075 ;
        RECT 89.770 200.760 112.855 201.060 ;
        RECT 42.605 200.380 42.935 200.395 ;
        RECT 45.825 200.380 46.155 200.395 ;
        RECT 42.605 200.080 46.155 200.380 ;
        RECT 42.605 200.065 42.935 200.080 ;
        RECT 45.825 200.065 46.155 200.080 ;
        RECT 84.005 200.380 84.335 200.395 ;
        RECT 89.770 200.380 90.070 200.760 ;
        RECT 112.525 200.745 112.855 200.760 ;
        RECT 84.005 200.080 90.070 200.380 ;
        RECT 90.905 200.380 91.235 200.395 ;
        RECT 124.945 200.380 125.275 200.395 ;
        RECT 90.905 200.080 125.275 200.380 ;
        RECT 84.005 200.065 84.335 200.080 ;
        RECT 90.905 200.065 91.235 200.080 ;
        RECT 124.945 200.065 125.275 200.080 ;
        RECT 86.305 199.700 86.635 199.715 ;
        RECT 120.345 199.700 120.675 199.715 ;
        RECT 86.305 199.400 120.675 199.700 ;
        RECT 86.305 199.385 86.635 199.400 ;
        RECT 120.345 199.385 120.675 199.400 ;
        RECT 82.165 199.020 82.495 199.035 ;
        RECT 91.365 199.020 91.695 199.035 ;
        RECT 82.165 198.720 91.695 199.020 ;
        RECT 82.165 198.705 82.495 198.720 ;
        RECT 91.365 198.705 91.695 198.720 ;
        RECT 40.110 198.365 42.090 198.695 ;
        RECT 70.110 198.365 72.090 198.695 ;
        RECT 100.110 198.365 102.090 198.695 ;
        RECT 130.110 198.365 132.090 198.695 ;
        RECT 46.285 197.660 46.615 197.675 ;
        RECT 50.425 197.660 50.755 197.675 ;
        RECT 46.285 197.360 50.755 197.660 ;
        RECT 46.285 197.345 46.615 197.360 ;
        RECT 50.425 197.345 50.755 197.360 ;
        RECT 98.265 197.660 98.595 197.675 ;
        RECT 113.445 197.660 113.775 197.675 ;
        RECT 117.125 197.660 117.455 197.675 ;
        RECT 98.265 197.360 117.455 197.660 ;
        RECT 98.265 197.345 98.595 197.360 ;
        RECT 113.445 197.345 113.775 197.360 ;
        RECT 117.125 197.345 117.455 197.360 ;
        RECT 59.165 196.980 59.495 196.995 ;
        RECT 67.445 196.980 67.775 196.995 ;
        RECT 136.905 196.980 137.235 196.995 ;
        RECT 59.165 196.680 137.235 196.980 ;
        RECT 59.165 196.665 59.495 196.680 ;
        RECT 67.445 196.665 67.775 196.680 ;
        RECT 136.905 196.665 137.235 196.680 ;
        RECT 48.125 196.300 48.455 196.315 ;
        RECT 53.850 196.300 54.230 196.310 ;
        RECT 48.125 196.000 54.230 196.300 ;
        RECT 48.125 195.985 48.455 196.000 ;
        RECT 53.850 195.990 54.230 196.000 ;
        RECT 55.110 195.645 57.090 195.975 ;
        RECT 85.110 195.645 87.090 195.975 ;
        RECT 115.110 195.645 117.090 195.975 ;
        RECT 145.110 195.645 147.090 195.975 ;
        RECT 60.085 195.620 60.415 195.635 ;
        RECT 57.800 195.320 60.415 195.620 ;
        RECT 57.800 194.955 58.100 195.320 ;
        RECT 60.085 195.305 60.415 195.320 ;
        RECT 89.065 195.620 89.395 195.635 ;
        RECT 102.865 195.620 103.195 195.635 ;
        RECT 106.545 195.620 106.875 195.635 ;
        RECT 89.065 195.320 106.875 195.620 ;
        RECT 89.065 195.305 89.395 195.320 ;
        RECT 102.865 195.305 103.195 195.320 ;
        RECT 106.545 195.305 106.875 195.320 ;
        RECT 57.785 194.625 58.115 194.955 ;
        RECT 55.025 194.260 55.355 194.275 ;
        RECT 69.285 194.260 69.615 194.275 ;
        RECT 55.025 193.960 69.615 194.260 ;
        RECT 55.025 193.945 55.355 193.960 ;
        RECT 69.285 193.945 69.615 193.960 ;
        RECT 102.405 194.260 102.735 194.275 ;
        RECT 123.105 194.260 123.435 194.275 ;
        RECT 102.405 193.960 123.435 194.260 ;
        RECT 102.405 193.945 102.735 193.960 ;
        RECT 123.105 193.945 123.435 193.960 ;
        RECT 131.845 194.260 132.175 194.275 ;
        RECT 136.445 194.260 136.775 194.275 ;
        RECT 131.845 193.960 136.775 194.260 ;
        RECT 131.845 193.945 132.175 193.960 ;
        RECT 136.445 193.945 136.775 193.960 ;
        RECT 40.110 192.925 42.090 193.255 ;
        RECT 70.110 192.925 72.090 193.255 ;
        RECT 100.110 192.925 102.090 193.255 ;
        RECT 130.110 192.925 132.090 193.255 ;
        RECT 74.345 192.220 74.675 192.235 ;
        RECT 118.965 192.220 119.295 192.235 ;
        RECT 74.345 191.920 119.295 192.220 ;
        RECT 74.345 191.905 74.675 191.920 ;
        RECT 118.965 191.905 119.295 191.920 ;
        RECT 46.745 191.540 47.075 191.555 ;
        RECT 117.585 191.540 117.915 191.555 ;
        RECT 46.745 191.240 117.915 191.540 ;
        RECT 46.745 191.225 47.075 191.240 ;
        RECT 117.585 191.225 117.915 191.240 ;
        RECT 67.905 190.860 68.235 190.875 ;
        RECT 80.325 190.860 80.655 190.875 ;
        RECT 67.905 190.560 80.655 190.860 ;
        RECT 67.905 190.545 68.235 190.560 ;
        RECT 80.325 190.545 80.655 190.560 ;
        RECT 94.585 190.860 94.915 190.875 ;
        RECT 106.085 190.860 106.415 190.875 ;
        RECT 94.585 190.560 106.415 190.860 ;
        RECT 94.585 190.545 94.915 190.560 ;
        RECT 106.085 190.545 106.415 190.560 ;
        RECT 55.110 190.205 57.090 190.535 ;
        RECT 85.110 190.205 87.090 190.535 ;
        RECT 115.110 190.205 117.090 190.535 ;
        RECT 145.110 190.205 147.090 190.535 ;
        RECT 91.365 190.180 91.695 190.195 ;
        RECT 99.185 190.180 99.515 190.195 ;
        RECT 91.365 189.880 99.515 190.180 ;
        RECT 91.365 189.865 91.695 189.880 ;
        RECT 99.185 189.865 99.515 189.880 ;
        RECT 107.005 190.180 107.335 190.195 ;
        RECT 109.050 190.180 109.430 190.190 ;
        RECT 107.005 189.880 109.430 190.180 ;
        RECT 107.005 189.865 107.335 189.880 ;
        RECT 109.050 189.870 109.430 189.880 ;
        RECT 41.685 189.500 42.015 189.515 ;
        RECT 128.625 189.500 128.955 189.515 ;
        RECT 41.685 189.200 128.955 189.500 ;
        RECT 41.685 189.185 42.015 189.200 ;
        RECT 128.625 189.185 128.955 189.200 ;
        RECT 53.645 188.820 53.975 188.835 ;
        RECT 130.005 188.820 130.335 188.835 ;
        RECT 53.645 188.520 130.335 188.820 ;
        RECT 53.645 188.505 53.975 188.520 ;
        RECT 130.005 188.505 130.335 188.520 ;
        RECT 132.765 188.140 133.095 188.155 ;
        RECT 138.285 188.140 138.615 188.155 ;
        RECT 132.765 187.840 138.615 188.140 ;
        RECT 132.765 187.825 133.095 187.840 ;
        RECT 138.285 187.825 138.615 187.840 ;
        RECT 40.110 187.485 42.090 187.815 ;
        RECT 70.110 187.485 72.090 187.815 ;
        RECT 100.110 187.485 102.090 187.815 ;
        RECT 130.110 187.485 132.090 187.815 ;
        RECT 78.485 187.460 78.815 187.475 ;
        RECT 82.370 187.460 82.750 187.470 ;
        RECT 78.485 187.160 82.750 187.460 ;
        RECT 78.485 187.145 78.815 187.160 ;
        RECT 82.370 187.150 82.750 187.160 ;
        RECT 52.265 186.780 52.595 186.795 ;
        RECT 130.005 186.780 130.335 186.795 ;
        RECT 133.225 186.780 133.555 186.795 ;
        RECT 52.265 186.480 133.555 186.780 ;
        RECT 52.265 186.465 52.595 186.480 ;
        RECT 130.005 186.465 130.335 186.480 ;
        RECT 133.225 186.465 133.555 186.480 ;
        RECT 134.605 186.780 134.935 186.795 ;
        RECT 139.665 186.780 139.995 186.795 ;
        RECT 141.505 186.780 141.835 186.795 ;
        RECT 134.605 186.480 141.835 186.780 ;
        RECT 134.605 186.465 134.935 186.480 ;
        RECT 139.665 186.465 139.995 186.480 ;
        RECT 141.505 186.465 141.835 186.480 ;
        RECT 86.765 186.100 87.095 186.115 ;
        RECT 88.810 186.100 89.190 186.110 ;
        RECT 86.765 185.800 89.190 186.100 ;
        RECT 86.765 185.785 87.095 185.800 ;
        RECT 88.810 185.790 89.190 185.800 ;
        RECT 116.665 186.100 116.995 186.115 ;
        RECT 122.185 186.100 122.515 186.115 ;
        RECT 116.665 185.800 122.515 186.100 ;
        RECT 116.665 185.785 116.995 185.800 ;
        RECT 122.185 185.785 122.515 185.800 ;
        RECT 138.745 186.100 139.075 186.115 ;
        RECT 143.805 186.100 144.135 186.115 ;
        RECT 138.745 185.800 144.135 186.100 ;
        RECT 138.745 185.785 139.075 185.800 ;
        RECT 143.805 185.785 144.135 185.800 ;
        RECT 95.045 185.420 95.375 185.435 ;
        RECT 96.885 185.420 97.215 185.435 ;
        RECT 95.045 185.120 97.215 185.420 ;
        RECT 95.045 185.105 95.375 185.120 ;
        RECT 96.885 185.105 97.215 185.120 ;
        RECT 55.110 184.765 57.090 185.095 ;
        RECT 85.110 184.765 87.090 185.095 ;
        RECT 115.110 184.765 117.090 185.095 ;
        RECT 145.110 184.765 147.090 185.095 ;
        RECT 100.105 184.740 100.435 184.755 ;
        RECT 107.210 184.740 107.590 184.750 ;
        RECT 100.105 184.440 107.590 184.740 ;
        RECT 100.105 184.425 100.435 184.440 ;
        RECT 107.210 184.430 107.590 184.440 ;
        RECT 130.465 184.740 130.795 184.755 ;
        RECT 132.970 184.740 133.350 184.750 ;
        RECT 130.465 184.440 133.350 184.740 ;
        RECT 130.465 184.425 130.795 184.440 ;
        RECT 132.970 184.430 133.350 184.440 ;
        RECT 92.285 184.060 92.615 184.075 ;
        RECT 101.485 184.060 101.815 184.075 ;
        RECT 92.285 183.760 101.815 184.060 ;
        RECT 92.285 183.745 92.615 183.760 ;
        RECT 101.485 183.745 101.815 183.760 ;
        RECT 106.545 184.060 106.875 184.075 ;
        RECT 110.225 184.060 110.555 184.075 ;
        RECT 106.545 183.760 110.555 184.060 ;
        RECT 106.545 183.745 106.875 183.760 ;
        RECT 110.225 183.745 110.555 183.760 ;
        RECT 131.845 184.060 132.175 184.075 ;
        RECT 140.125 184.060 140.455 184.075 ;
        RECT 131.845 183.760 140.455 184.060 ;
        RECT 131.845 183.745 132.175 183.760 ;
        RECT 140.125 183.745 140.455 183.760 ;
        RECT 84.465 183.380 84.795 183.395 ;
        RECT 137.365 183.380 137.695 183.395 ;
        RECT 84.465 183.080 137.695 183.380 ;
        RECT 84.465 183.065 84.795 183.080 ;
        RECT 137.365 183.065 137.695 183.080 ;
        RECT 82.625 182.700 82.955 182.715 ;
        RECT 82.410 182.385 82.955 182.700 ;
        RECT 108.385 182.700 108.715 182.715 ;
        RECT 113.445 182.700 113.775 182.715 ;
        RECT 108.385 182.400 113.775 182.700 ;
        RECT 108.385 182.385 108.715 182.400 ;
        RECT 113.445 182.385 113.775 182.400 ;
        RECT 40.110 182.045 42.090 182.375 ;
        RECT 70.110 182.045 72.090 182.375 ;
        RECT 43.985 182.020 44.315 182.035 ;
        RECT 48.585 182.020 48.915 182.035 ;
        RECT 43.985 181.720 48.915 182.020 ;
        RECT 43.985 181.705 44.315 181.720 ;
        RECT 48.585 181.705 48.915 181.720 ;
        RECT 82.410 181.355 82.710 182.385 ;
        RECT 100.110 182.045 102.090 182.375 ;
        RECT 130.110 182.045 132.090 182.375 ;
        RECT 119.425 182.020 119.755 182.035 ;
        RECT 122.185 182.020 122.515 182.035 ;
        RECT 119.425 181.720 122.515 182.020 ;
        RECT 119.425 181.705 119.755 181.720 ;
        RECT 122.185 181.705 122.515 181.720 ;
        RECT 82.410 181.040 82.955 181.355 ;
        RECT 82.625 181.025 82.955 181.040 ;
        RECT 110.685 181.340 111.015 181.355 ;
        RECT 119.885 181.340 120.215 181.355 ;
        RECT 110.685 181.040 120.215 181.340 ;
        RECT 110.685 181.025 111.015 181.040 ;
        RECT 119.885 181.025 120.215 181.040 ;
        RECT 122.185 181.340 122.515 181.355 ;
        RECT 141.505 181.340 141.835 181.355 ;
        RECT 122.185 181.040 141.835 181.340 ;
        RECT 122.185 181.025 122.515 181.040 ;
        RECT 141.505 181.025 141.835 181.040 ;
        RECT 80.785 180.660 81.115 180.675 ;
        RECT 116.205 180.660 116.535 180.675 ;
        RECT 80.785 180.360 116.535 180.660 ;
        RECT 80.785 180.345 81.115 180.360 ;
        RECT 116.205 180.345 116.535 180.360 ;
        RECT 127.245 180.660 127.575 180.675 ;
        RECT 136.905 180.660 137.235 180.675 ;
        RECT 127.245 180.360 137.235 180.660 ;
        RECT 127.245 180.345 127.575 180.360 ;
        RECT 136.905 180.345 137.235 180.360 ;
        RECT 95.505 179.980 95.835 179.995 ;
        RECT 111.605 179.980 111.935 179.995 ;
        RECT 133.225 179.990 133.555 179.995 ;
        RECT 132.970 179.980 133.555 179.990 ;
        RECT 95.505 179.680 111.935 179.980 ;
        RECT 132.770 179.680 133.555 179.980 ;
        RECT 95.505 179.665 95.835 179.680 ;
        RECT 111.605 179.665 111.935 179.680 ;
        RECT 132.970 179.670 133.555 179.680 ;
        RECT 133.225 179.665 133.555 179.670 ;
        RECT 134.605 179.980 134.935 179.995 ;
        RECT 139.665 179.980 139.995 179.995 ;
        RECT 134.605 179.680 139.995 179.980 ;
        RECT 134.605 179.665 134.935 179.680 ;
        RECT 139.665 179.665 139.995 179.680 ;
        RECT 55.110 179.325 57.090 179.655 ;
        RECT 85.110 179.325 87.090 179.655 ;
        RECT 115.110 179.325 117.090 179.655 ;
        RECT 145.110 179.325 147.090 179.655 ;
        RECT 95.965 179.300 96.295 179.315 ;
        RECT 103.325 179.300 103.655 179.315 ;
        RECT 95.965 179.000 103.655 179.300 ;
        RECT 95.965 178.985 96.295 179.000 ;
        RECT 103.325 178.985 103.655 179.000 ;
        RECT 50.885 178.620 51.215 178.635 ;
        RECT 78.945 178.620 79.275 178.635 ;
        RECT 50.885 178.320 79.275 178.620 ;
        RECT 50.885 178.305 51.215 178.320 ;
        RECT 78.945 178.305 79.275 178.320 ;
        RECT 101.945 178.620 102.275 178.635 ;
        RECT 120.805 178.620 121.135 178.635 ;
        RECT 101.945 178.320 121.135 178.620 ;
        RECT 101.945 178.305 102.275 178.320 ;
        RECT 120.805 178.305 121.135 178.320 ;
        RECT 53.850 177.940 54.230 177.950 ;
        RECT 124.945 177.940 125.275 177.955 ;
        RECT 53.850 177.640 125.275 177.940 ;
        RECT 53.850 177.630 54.230 177.640 ;
        RECT 124.945 177.625 125.275 177.640 ;
        RECT 40.110 176.605 42.090 176.935 ;
        RECT 70.110 176.605 72.090 176.935 ;
        RECT 100.110 176.605 102.090 176.935 ;
        RECT 130.110 176.605 132.090 176.935 ;
        RECT 84.465 176.580 84.795 176.595 ;
        RECT 94.125 176.580 94.455 176.595 ;
        RECT 84.465 176.280 94.455 176.580 ;
        RECT 84.465 176.265 84.795 176.280 ;
        RECT 94.125 176.265 94.455 176.280 ;
        RECT 104.245 176.580 104.575 176.595 ;
        RECT 107.465 176.580 107.795 176.595 ;
        RECT 104.245 176.280 107.795 176.580 ;
        RECT 104.245 176.265 104.575 176.280 ;
        RECT 107.465 176.265 107.795 176.280 ;
        RECT 47.665 175.900 47.995 175.915 ;
        RECT 53.645 175.900 53.975 175.915 ;
        RECT 61.005 175.900 61.335 175.915 ;
        RECT 47.665 175.600 61.335 175.900 ;
        RECT 47.665 175.585 47.995 175.600 ;
        RECT 53.645 175.585 53.975 175.600 ;
        RECT 61.005 175.585 61.335 175.600 ;
        RECT 81.245 175.900 81.575 175.915 ;
        RECT 120.345 175.900 120.675 175.915 ;
        RECT 81.245 175.600 120.675 175.900 ;
        RECT 81.245 175.585 81.575 175.600 ;
        RECT 120.345 175.585 120.675 175.600 ;
        RECT 82.370 175.220 82.750 175.230 ;
        RECT 92.285 175.220 92.615 175.235 ;
        RECT 104.245 175.220 104.575 175.235 ;
        RECT 109.765 175.220 110.095 175.235 ;
        RECT 121.725 175.220 122.055 175.235 ;
        RECT 82.370 174.920 91.910 175.220 ;
        RECT 82.370 174.910 82.750 174.920 ;
        RECT 91.610 174.540 91.910 174.920 ;
        RECT 92.285 174.920 110.095 175.220 ;
        RECT 92.285 174.905 92.615 174.920 ;
        RECT 104.245 174.905 104.575 174.920 ;
        RECT 109.765 174.905 110.095 174.920 ;
        RECT 114.380 174.920 122.055 175.220 ;
        RECT 114.380 174.540 114.680 174.920 ;
        RECT 121.725 174.905 122.055 174.920 ;
        RECT 91.610 174.240 114.680 174.540 ;
        RECT 55.110 173.885 57.090 174.215 ;
        RECT 85.110 173.885 87.090 174.215 ;
        RECT 115.110 173.885 117.090 174.215 ;
        RECT 145.110 173.885 147.090 174.215 ;
        RECT 90.905 173.860 91.235 173.875 ;
        RECT 92.745 173.860 93.075 173.875 ;
        RECT 90.905 173.560 93.075 173.860 ;
        RECT 90.905 173.545 91.235 173.560 ;
        RECT 92.745 173.545 93.075 173.560 ;
        RECT 94.125 173.860 94.455 173.875 ;
        RECT 114.365 173.860 114.695 173.875 ;
        RECT 94.125 173.560 114.695 173.860 ;
        RECT 94.125 173.545 94.455 173.560 ;
        RECT 114.365 173.545 114.695 173.560 ;
        RECT 90.905 173.180 91.235 173.195 ;
        RECT 95.965 173.180 96.295 173.195 ;
        RECT 90.905 172.880 96.295 173.180 ;
        RECT 90.905 172.865 91.235 172.880 ;
        RECT 95.965 172.865 96.295 172.880 ;
        RECT 111.810 173.180 112.190 173.190 ;
        RECT 119.885 173.180 120.215 173.195 ;
        RECT 111.810 172.880 120.215 173.180 ;
        RECT 111.810 172.870 112.190 172.880 ;
        RECT 119.885 172.865 120.215 172.880 ;
        RECT 81.705 172.500 82.035 172.515 ;
        RECT 101.485 172.500 101.815 172.515 ;
        RECT 81.705 172.200 101.815 172.500 ;
        RECT 81.705 172.185 82.035 172.200 ;
        RECT 101.485 172.185 101.815 172.200 ;
        RECT 85.845 171.820 86.175 171.835 ;
        RECT 94.125 171.820 94.455 171.835 ;
        RECT 85.845 171.520 94.455 171.820 ;
        RECT 85.845 171.505 86.175 171.520 ;
        RECT 94.125 171.505 94.455 171.520 ;
        RECT 40.110 171.165 42.090 171.495 ;
        RECT 70.110 171.165 72.090 171.495 ;
        RECT 100.110 171.165 102.090 171.495 ;
        RECT 130.110 171.165 132.090 171.495 ;
        RECT 102.865 171.140 103.195 171.155 ;
        RECT 112.985 171.140 113.315 171.155 ;
        RECT 102.865 170.840 113.315 171.140 ;
        RECT 102.865 170.825 103.195 170.840 ;
        RECT 112.985 170.825 113.315 170.840 ;
        RECT 87.685 170.460 88.015 170.475 ;
        RECT 103.785 170.460 104.115 170.475 ;
        RECT 87.685 170.160 104.115 170.460 ;
        RECT 87.685 170.145 88.015 170.160 ;
        RECT 103.785 170.145 104.115 170.160 ;
        RECT 81.245 169.780 81.575 169.795 ;
        RECT 133.225 169.780 133.555 169.795 ;
        RECT 81.245 169.480 133.555 169.780 ;
        RECT 81.245 169.465 81.575 169.480 ;
        RECT 133.225 169.465 133.555 169.480 ;
        RECT 87.685 169.100 88.015 169.115 ;
        RECT 107.005 169.100 107.335 169.115 ;
        RECT 87.685 168.800 107.335 169.100 ;
        RECT 87.685 168.785 88.015 168.800 ;
        RECT 107.005 168.785 107.335 168.800 ;
        RECT 55.110 168.445 57.090 168.775 ;
        RECT 85.110 168.445 87.090 168.775 ;
        RECT 115.110 168.445 117.090 168.775 ;
        RECT 145.110 168.445 147.090 168.775 ;
        RECT 89.985 168.420 90.315 168.435 ;
        RECT 93.205 168.420 93.535 168.435 ;
        RECT 89.985 168.120 93.535 168.420 ;
        RECT 89.985 168.105 90.315 168.120 ;
        RECT 93.205 168.105 93.535 168.120 ;
        RECT 107.005 167.750 107.335 167.755 ;
        RECT 107.005 167.740 107.590 167.750 ;
        RECT 106.780 167.440 107.590 167.740 ;
        RECT 107.005 167.430 107.590 167.440 ;
        RECT 107.005 167.425 107.335 167.430 ;
        RECT 74.345 167.060 74.675 167.075 ;
        RECT 97.345 167.060 97.675 167.075 ;
        RECT 99.645 167.060 99.975 167.075 ;
        RECT 74.345 166.760 99.975 167.060 ;
        RECT 74.345 166.745 74.675 166.760 ;
        RECT 97.345 166.745 97.675 166.760 ;
        RECT 99.645 166.745 99.975 166.760 ;
        RECT 136.650 167.060 137.030 167.070 ;
        RECT 140.125 167.060 140.455 167.075 ;
        RECT 136.650 166.760 140.455 167.060 ;
        RECT 136.650 166.750 137.030 166.760 ;
        RECT 140.125 166.745 140.455 166.760 ;
        RECT 109.050 166.380 109.430 166.390 ;
        RECT 112.985 166.380 113.315 166.395 ;
        RECT 109.050 166.080 113.315 166.380 ;
        RECT 109.050 166.070 109.430 166.080 ;
        RECT 112.985 166.065 113.315 166.080 ;
        RECT 113.650 166.380 114.030 166.390 ;
        RECT 118.045 166.380 118.375 166.395 ;
        RECT 113.650 166.080 118.375 166.380 ;
        RECT 113.650 166.070 114.030 166.080 ;
        RECT 118.045 166.065 118.375 166.080 ;
        RECT 40.110 165.725 42.090 166.055 ;
        RECT 70.110 165.725 72.090 166.055 ;
        RECT 100.110 165.725 102.090 166.055 ;
        RECT 130.110 165.725 132.090 166.055 ;
        RECT 83.545 165.710 83.875 165.715 ;
        RECT 83.290 165.700 83.875 165.710 ;
        RECT 83.290 165.400 84.100 165.700 ;
        RECT 83.290 165.390 83.875 165.400 ;
        RECT 83.545 165.385 83.875 165.390 ;
        RECT 69.745 165.020 70.075 165.035 ;
        RECT 110.685 165.020 111.015 165.035 ;
        RECT 69.745 164.720 111.015 165.020 ;
        RECT 69.745 164.705 70.075 164.720 ;
        RECT 110.685 164.705 111.015 164.720 ;
        RECT 82.370 164.340 82.750 164.350 ;
        RECT 88.605 164.340 88.935 164.355 ;
        RECT 82.370 164.040 88.935 164.340 ;
        RECT 82.370 164.030 82.750 164.040 ;
        RECT 88.605 164.025 88.935 164.040 ;
        RECT 99.185 164.340 99.515 164.355 ;
        RECT 118.045 164.340 118.375 164.355 ;
        RECT 99.185 164.040 118.375 164.340 ;
        RECT 99.185 164.025 99.515 164.040 ;
        RECT 118.045 164.025 118.375 164.040 ;
        RECT 89.985 163.660 90.315 163.675 ;
        RECT 101.485 163.660 101.815 163.675 ;
        RECT 89.985 163.360 101.815 163.660 ;
        RECT 89.985 163.345 90.315 163.360 ;
        RECT 101.485 163.345 101.815 163.360 ;
        RECT 55.110 163.005 57.090 163.335 ;
        RECT 85.110 163.005 87.090 163.335 ;
        RECT 115.110 163.005 117.090 163.335 ;
        RECT 145.110 163.005 147.090 163.335 ;
        RECT 98.265 162.980 98.595 162.995 ;
        RECT 95.290 162.680 98.595 162.980 ;
        RECT 74.345 162.300 74.675 162.315 ;
        RECT 95.290 162.300 95.590 162.680 ;
        RECT 98.265 162.665 98.595 162.680 ;
        RECT 118.505 162.300 118.835 162.315 ;
        RECT 74.345 162.000 95.590 162.300 ;
        RECT 110.010 162.000 118.835 162.300 ;
        RECT 74.345 161.985 74.675 162.000 ;
        RECT 63.765 161.620 64.095 161.635 ;
        RECT 72.045 161.620 72.375 161.635 ;
        RECT 63.765 161.320 72.375 161.620 ;
        RECT 63.765 161.305 64.095 161.320 ;
        RECT 72.045 161.305 72.375 161.320 ;
        RECT 85.845 161.620 86.175 161.635 ;
        RECT 110.010 161.620 110.310 162.000 ;
        RECT 118.505 161.985 118.835 162.000 ;
        RECT 85.845 161.320 110.310 161.620 ;
        RECT 110.685 161.620 111.015 161.635 ;
        RECT 113.445 161.620 113.775 161.635 ;
        RECT 110.685 161.320 113.775 161.620 ;
        RECT 85.845 161.305 86.175 161.320 ;
        RECT 110.685 161.305 111.015 161.320 ;
        RECT 113.445 161.305 113.775 161.320 ;
        RECT 131.385 161.620 131.715 161.635 ;
        RECT 140.585 161.620 140.915 161.635 ;
        RECT 131.385 161.320 140.915 161.620 ;
        RECT 131.385 161.305 131.715 161.320 ;
        RECT 140.585 161.305 140.915 161.320 ;
        RECT 40.110 160.285 42.090 160.615 ;
        RECT 70.110 160.285 72.090 160.615 ;
        RECT 100.110 160.285 102.090 160.615 ;
        RECT 130.110 160.285 132.090 160.615 ;
        RECT 100.565 159.580 100.895 159.595 ;
        RECT 125.865 159.580 126.195 159.595 ;
        RECT 100.565 159.280 126.195 159.580 ;
        RECT 100.565 159.265 100.895 159.280 ;
        RECT 125.865 159.265 126.195 159.280 ;
        RECT 97.345 158.900 97.675 158.915 ;
        RECT 125.865 158.900 126.195 158.915 ;
        RECT 97.345 158.600 126.195 158.900 ;
        RECT 97.345 158.585 97.675 158.600 ;
        RECT 125.865 158.585 126.195 158.600 ;
        RECT 80.530 158.220 80.910 158.230 ;
        RECT 81.245 158.220 81.575 158.235 ;
        RECT 80.530 157.920 81.575 158.220 ;
        RECT 80.530 157.910 80.910 157.920 ;
        RECT 81.245 157.905 81.575 157.920 ;
        RECT 55.110 157.565 57.090 157.895 ;
        RECT 85.110 157.565 87.090 157.895 ;
        RECT 115.110 157.565 117.090 157.895 ;
        RECT 145.110 157.565 147.090 157.895 ;
        RECT 73.425 157.540 73.755 157.555 ;
        RECT 78.945 157.540 79.275 157.555 ;
        RECT 73.425 157.240 79.275 157.540 ;
        RECT 73.425 157.225 73.755 157.240 ;
        RECT 78.945 157.225 79.275 157.240 ;
        RECT 82.370 157.540 82.750 157.550 ;
        RECT 83.545 157.540 83.875 157.555 ;
        RECT 82.370 157.240 83.875 157.540 ;
        RECT 82.370 157.230 82.750 157.240 ;
        RECT 83.545 157.225 83.875 157.240 ;
        RECT 66.525 156.860 66.855 156.875 ;
        RECT 127.705 156.860 128.035 156.875 ;
        RECT 66.525 156.560 128.035 156.860 ;
        RECT 66.525 156.545 66.855 156.560 ;
        RECT 127.705 156.545 128.035 156.560 ;
        RECT 133.225 156.860 133.555 156.875 ;
        RECT 141.045 156.860 141.375 156.875 ;
        RECT 133.225 156.560 141.375 156.860 ;
        RECT 133.225 156.545 133.555 156.560 ;
        RECT 141.045 156.545 141.375 156.560 ;
        RECT 68.365 156.180 68.695 156.195 ;
        RECT 116.205 156.180 116.535 156.195 ;
        RECT 68.365 155.880 116.535 156.180 ;
        RECT 68.365 155.865 68.695 155.880 ;
        RECT 116.205 155.865 116.535 155.880 ;
        RECT 123.105 156.180 123.435 156.195 ;
        RECT 126.325 156.180 126.655 156.195 ;
        RECT 123.105 155.880 126.655 156.180 ;
        RECT 123.105 155.865 123.435 155.880 ;
        RECT 126.325 155.865 126.655 155.880 ;
        RECT 78.690 155.500 79.070 155.510 ;
        RECT 81.245 155.500 81.575 155.515 ;
        RECT 88.605 155.510 88.935 155.515 ;
        RECT 88.605 155.500 89.190 155.510 ;
        RECT 78.690 155.200 81.575 155.500 ;
        RECT 88.380 155.200 89.190 155.500 ;
        RECT 78.690 155.190 79.070 155.200 ;
        RECT 81.245 155.185 81.575 155.200 ;
        RECT 88.605 155.190 89.190 155.200 ;
        RECT 111.145 155.500 111.475 155.515 ;
        RECT 115.285 155.500 115.615 155.515 ;
        RECT 111.145 155.200 115.615 155.500 ;
        RECT 88.605 155.185 88.935 155.190 ;
        RECT 111.145 155.185 111.475 155.200 ;
        RECT 115.285 155.185 115.615 155.200 ;
        RECT 40.110 154.845 42.090 155.175 ;
        RECT 70.110 154.845 72.090 155.175 ;
        RECT 100.110 154.845 102.090 155.175 ;
        RECT 130.110 154.845 132.090 155.175 ;
        RECT 80.785 154.505 81.115 154.835 ;
        RECT 83.085 154.820 83.415 154.835 ;
        RECT 85.385 154.820 85.715 154.835 ;
        RECT 83.085 154.520 85.715 154.820 ;
        RECT 83.085 154.505 83.415 154.520 ;
        RECT 85.385 154.505 85.715 154.520 ;
        RECT 79.610 154.140 79.990 154.150 ;
        RECT 80.800 154.140 81.100 154.505 ;
        RECT 79.610 153.840 81.100 154.140 ;
        RECT 81.705 154.140 82.035 154.155 ;
        RECT 92.285 154.140 92.615 154.155 ;
        RECT 81.705 153.840 92.615 154.140 ;
        RECT 79.610 153.830 79.990 153.840 ;
        RECT 81.705 153.825 82.035 153.840 ;
        RECT 92.285 153.825 92.615 153.840 ;
        RECT 106.545 154.140 106.875 154.155 ;
        RECT 112.065 154.140 112.395 154.155 ;
        RECT 114.365 154.140 114.695 154.155 ;
        RECT 106.545 153.840 114.695 154.140 ;
        RECT 106.545 153.825 106.875 153.840 ;
        RECT 112.065 153.825 112.395 153.840 ;
        RECT 114.365 153.825 114.695 153.840 ;
        RECT 41.225 153.460 41.555 153.475 ;
        RECT 72.505 153.460 72.835 153.475 ;
        RECT 95.045 153.460 95.375 153.475 ;
        RECT 107.465 153.460 107.795 153.475 ;
        RECT 131.845 153.460 132.175 153.475 ;
        RECT 41.225 153.160 71.670 153.460 ;
        RECT 41.225 153.145 41.555 153.160 ;
        RECT 71.370 152.780 71.670 153.160 ;
        RECT 72.505 153.290 81.100 153.460 ;
        RECT 81.490 153.290 88.230 153.460 ;
        RECT 72.505 153.160 88.230 153.290 ;
        RECT 72.505 153.145 72.835 153.160 ;
        RECT 80.800 152.990 81.790 153.160 ;
        RECT 79.865 152.780 80.195 152.795 ;
        RECT 71.370 152.480 80.195 152.780 ;
        RECT 79.865 152.465 80.195 152.480 ;
        RECT 82.165 152.790 82.495 152.795 ;
        RECT 82.165 152.780 82.750 152.790 ;
        RECT 87.930 152.780 88.230 153.160 ;
        RECT 95.045 153.160 107.795 153.460 ;
        RECT 95.045 153.145 95.375 153.160 ;
        RECT 107.465 153.145 107.795 153.160 ;
        RECT 113.690 153.160 132.175 153.460 ;
        RECT 113.690 152.780 113.990 153.160 ;
        RECT 131.845 153.145 132.175 153.160 ;
        RECT 82.165 152.480 82.950 152.780 ;
        RECT 87.930 152.480 113.990 152.780 ;
        RECT 82.165 152.470 82.750 152.480 ;
        RECT 82.165 152.465 82.495 152.470 ;
        RECT 55.110 152.125 57.090 152.455 ;
        RECT 85.110 152.125 87.090 152.455 ;
        RECT 115.110 152.125 117.090 152.455 ;
        RECT 145.110 152.125 147.090 152.455 ;
        RECT 78.690 152.100 79.070 152.110 ;
        RECT 80.785 152.100 81.115 152.115 ;
        RECT 78.690 151.800 81.115 152.100 ;
        RECT 78.690 151.790 79.070 151.800 ;
        RECT 80.785 151.785 81.115 151.800 ;
        RECT 82.165 152.100 82.495 152.115 ;
        RECT 83.545 152.100 83.875 152.115 ;
        RECT 82.165 151.800 83.875 152.100 ;
        RECT 82.165 151.785 82.495 151.800 ;
        RECT 83.545 151.785 83.875 151.800 ;
        RECT 98.265 152.100 98.595 152.115 ;
        RECT 98.930 152.100 99.310 152.110 ;
        RECT 101.025 152.100 101.355 152.115 ;
        RECT 98.265 151.800 101.355 152.100 ;
        RECT 98.265 151.785 98.595 151.800 ;
        RECT 98.930 151.790 99.310 151.800 ;
        RECT 101.025 151.785 101.355 151.800 ;
        RECT 124.485 152.100 124.815 152.115 ;
        RECT 136.650 152.100 137.030 152.110 ;
        RECT 124.485 151.800 137.030 152.100 ;
        RECT 124.485 151.785 124.815 151.800 ;
        RECT 136.650 151.790 137.030 151.800 ;
        RECT 53.645 151.420 53.975 151.435 ;
        RECT 140.585 151.420 140.915 151.435 ;
        RECT 53.645 151.120 140.915 151.420 ;
        RECT 53.645 151.105 53.975 151.120 ;
        RECT 140.585 151.105 140.915 151.120 ;
        RECT 79.610 150.740 79.990 150.750 ;
        RECT 80.325 150.740 80.655 150.755 ;
        RECT 79.610 150.440 80.655 150.740 ;
        RECT 79.610 150.430 79.990 150.440 ;
        RECT 80.325 150.425 80.655 150.440 ;
        RECT 89.985 150.740 90.315 150.755 ;
        RECT 127.705 150.740 128.035 150.755 ;
        RECT 89.985 150.440 128.035 150.740 ;
        RECT 89.985 150.425 90.315 150.440 ;
        RECT 127.705 150.425 128.035 150.440 ;
        RECT 77.105 150.060 77.435 150.075 ;
        RECT 91.825 150.060 92.155 150.075 ;
        RECT 77.105 149.760 92.155 150.060 ;
        RECT 77.105 149.745 77.435 149.760 ;
        RECT 91.825 149.745 92.155 149.760 ;
        RECT 112.985 150.060 113.315 150.075 ;
        RECT 120.805 150.060 121.135 150.075 ;
        RECT 112.985 149.760 121.135 150.060 ;
        RECT 112.985 149.745 113.315 149.760 ;
        RECT 120.805 149.745 121.135 149.760 ;
        RECT 40.110 149.405 42.090 149.735 ;
        RECT 70.110 149.405 72.090 149.735 ;
        RECT 100.110 149.405 102.090 149.735 ;
        RECT 130.110 149.405 132.090 149.735 ;
        RECT 76.185 149.380 76.515 149.395 ;
        RECT 92.285 149.380 92.615 149.395 ;
        RECT 76.185 149.080 92.615 149.380 ;
        RECT 76.185 149.065 76.515 149.080 ;
        RECT 92.285 149.065 92.615 149.080 ;
        RECT 107.925 149.390 108.255 149.395 ;
        RECT 107.925 149.380 108.510 149.390 ;
        RECT 111.605 149.380 111.935 149.395 ;
        RECT 113.905 149.380 114.235 149.395 ;
        RECT 107.925 149.080 108.710 149.380 ;
        RECT 111.605 149.080 114.235 149.380 ;
        RECT 107.925 149.070 108.510 149.080 ;
        RECT 107.925 149.065 108.255 149.070 ;
        RECT 111.605 149.065 111.935 149.080 ;
        RECT 113.905 149.065 114.235 149.080 ;
        RECT 71.125 148.700 71.455 148.715 ;
        RECT 78.945 148.700 79.275 148.715 ;
        RECT 71.125 148.400 79.275 148.700 ;
        RECT 71.125 148.385 71.455 148.400 ;
        RECT 78.945 148.385 79.275 148.400 ;
        RECT 87.685 148.700 88.015 148.715 ;
        RECT 118.965 148.700 119.295 148.715 ;
        RECT 87.685 148.400 119.295 148.700 ;
        RECT 87.685 148.385 88.015 148.400 ;
        RECT 118.965 148.385 119.295 148.400 ;
        RECT 55.025 148.020 55.355 148.035 ;
        RECT 125.405 148.020 125.735 148.035 ;
        RECT 55.025 147.720 125.735 148.020 ;
        RECT 55.025 147.705 55.355 147.720 ;
        RECT 125.405 147.705 125.735 147.720 ;
        RECT 80.785 147.350 81.115 147.355 ;
        RECT 80.530 147.340 81.115 147.350 ;
        RECT 80.530 147.040 81.340 147.340 ;
        RECT 80.530 147.030 81.115 147.040 ;
        RECT 80.785 147.025 81.115 147.030 ;
        RECT 55.110 146.685 57.090 147.015 ;
        RECT 85.110 146.685 87.090 147.015 ;
        RECT 115.110 146.685 117.090 147.015 ;
        RECT 145.110 146.685 147.090 147.015 ;
        RECT 100.105 146.660 100.435 146.675 ;
        RECT 111.605 146.660 111.935 146.675 ;
        RECT 100.105 146.360 111.935 146.660 ;
        RECT 100.105 146.345 100.435 146.360 ;
        RECT 111.605 146.345 111.935 146.360 ;
        RECT 76.185 145.980 76.515 145.995 ;
        RECT 90.905 145.980 91.235 145.995 ;
        RECT 113.650 145.980 114.030 145.990 ;
        RECT 115.285 145.980 115.615 145.995 ;
        RECT 76.185 145.680 115.615 145.980 ;
        RECT 76.185 145.665 76.515 145.680 ;
        RECT 90.905 145.665 91.235 145.680 ;
        RECT 113.650 145.670 114.030 145.680 ;
        RECT 115.285 145.665 115.615 145.680 ;
        RECT 40.110 143.965 42.090 144.295 ;
        RECT 70.110 143.965 72.090 144.295 ;
        RECT 100.110 143.965 102.090 144.295 ;
        RECT 130.110 143.965 132.090 144.295 ;
        RECT 82.165 143.260 82.495 143.275 ;
        RECT 83.290 143.260 83.670 143.270 ;
        RECT 82.165 142.960 83.670 143.260 ;
        RECT 82.165 142.945 82.495 142.960 ;
        RECT 83.290 142.950 83.670 142.960 ;
        RECT 55.110 141.245 57.090 141.575 ;
        RECT 85.110 141.245 87.090 141.575 ;
        RECT 115.110 141.245 117.090 141.575 ;
        RECT 145.110 141.245 147.090 141.575 ;
        RECT 3.455 137.450 4.945 137.475 ;
        RECT 42.975 137.450 45.025 137.695 ;
        RECT 70.075 137.450 72.125 137.695 ;
        RECT 96.775 137.450 98.825 137.695 ;
        RECT 130.075 137.450 132.125 137.695 ;
        RECT 3.450 135.950 135.850 137.450 ;
        RECT 3.455 135.925 4.945 135.950 ;
        RECT 42.975 135.705 45.025 135.950 ;
        RECT 70.075 135.705 72.125 135.950 ;
        RECT 96.775 135.705 98.825 135.950 ;
        RECT 130.075 135.705 132.125 135.950 ;
        RECT 12.655 134.650 14.145 134.675 ;
        RECT 55.075 134.650 57.125 134.795 ;
        RECT 84.275 134.650 86.325 134.795 ;
        RECT 112.175 134.650 114.225 134.795 ;
        RECT 147.775 134.650 149.825 134.795 ;
        RECT 12.650 133.150 149.850 134.650 ;
        RECT 12.655 133.125 14.145 133.150 ;
        RECT 55.075 132.805 57.125 133.150 ;
        RECT 84.275 132.805 86.325 133.150 ;
        RECT 112.175 132.805 114.225 133.150 ;
        RECT 147.775 132.805 149.825 133.150 ;
        RECT 156.395 52.570 157.325 52.595 ;
        RECT 146.930 51.630 157.330 52.570 ;
        RECT 156.395 51.605 157.325 51.630 ;
        RECT 134.345 50.340 135.220 50.365 ;
        RECT 130.260 49.455 135.225 50.340 ;
        RECT 134.345 49.430 135.220 49.455 ;
        RECT 130.670 48.130 131.525 48.155 ;
        RECT 126.570 47.265 131.530 48.130 ;
        RECT 130.670 47.240 131.525 47.265 ;
        RECT 20.475 23.000 21.525 23.025 ;
        RECT 17.070 22.000 21.525 23.000 ;
        RECT 20.475 21.975 21.525 22.000 ;
        RECT 20.475 16.615 21.525 16.640 ;
        RECT 5.870 15.615 21.525 16.615 ;
        RECT 20.475 15.590 21.525 15.615 ;
        RECT 35.600 5.670 36.600 7.700 ;
      LAYER via3 ;
        RECT 31.355 221.805 31.845 222.295 ;
        RECT 20.650 220.550 21.150 221.050 ;
        RECT 9.305 218.005 9.695 218.395 ;
        RECT 12.600 218.000 13.000 218.400 ;
        RECT 92.160 223.465 92.640 223.945 ;
        RECT 51.820 222.840 52.140 223.160 ;
        RECT 55.500 222.770 55.820 223.090 ;
        RECT 59.180 222.770 59.500 223.090 ;
        RECT 62.860 222.770 63.180 223.090 ;
        RECT 66.540 222.770 66.860 223.090 ;
        RECT 70.220 222.770 70.540 223.090 ;
        RECT 73.900 222.770 74.220 223.090 ;
        RECT 77.580 222.770 77.900 223.090 ;
        RECT 81.260 222.770 81.580 223.090 ;
        RECT 84.940 222.770 85.260 223.090 ;
        RECT 88.620 222.770 88.940 223.090 ;
        RECT 121.740 222.770 122.060 223.090 ;
        RECT 125.420 222.770 125.740 223.090 ;
        RECT 129.100 222.770 129.420 223.090 ;
        RECT 132.780 222.770 133.100 223.090 ;
        RECT 136.460 222.770 136.780 223.090 ;
        RECT 140.140 222.770 140.460 223.090 ;
        RECT 143.820 222.770 144.140 223.090 ;
        RECT 147.500 222.770 147.820 223.090 ;
        RECT 95.940 220.300 96.340 220.700 ;
        RECT 99.625 219.505 100.020 219.900 ;
        RECT 103.310 218.710 103.695 219.095 ;
        RECT 106.985 217.905 107.375 218.295 ;
        RECT 40.140 214.690 40.460 215.010 ;
        RECT 40.540 214.690 40.860 215.010 ;
        RECT 40.940 214.690 41.260 215.010 ;
        RECT 41.340 214.690 41.660 215.010 ;
        RECT 41.740 214.690 42.060 215.010 ;
        RECT 70.140 214.690 70.460 215.010 ;
        RECT 70.540 214.690 70.860 215.010 ;
        RECT 70.940 214.690 71.260 215.010 ;
        RECT 71.340 214.690 71.660 215.010 ;
        RECT 71.740 214.690 72.060 215.010 ;
        RECT 100.140 214.690 100.460 215.010 ;
        RECT 100.540 214.690 100.860 215.010 ;
        RECT 100.940 214.690 101.260 215.010 ;
        RECT 101.340 214.690 101.660 215.010 ;
        RECT 101.740 214.690 102.060 215.010 ;
        RECT 130.140 214.690 130.460 215.010 ;
        RECT 130.540 214.690 130.860 215.010 ;
        RECT 130.940 214.690 131.260 215.010 ;
        RECT 131.340 214.690 131.660 215.010 ;
        RECT 131.740 214.690 132.060 215.010 ;
        RECT 55.140 211.970 55.460 212.290 ;
        RECT 55.540 211.970 55.860 212.290 ;
        RECT 55.940 211.970 56.260 212.290 ;
        RECT 56.340 211.970 56.660 212.290 ;
        RECT 56.740 211.970 57.060 212.290 ;
        RECT 85.140 211.970 85.460 212.290 ;
        RECT 85.540 211.970 85.860 212.290 ;
        RECT 85.940 211.970 86.260 212.290 ;
        RECT 86.340 211.970 86.660 212.290 ;
        RECT 86.740 211.970 87.060 212.290 ;
        RECT 115.140 211.970 115.460 212.290 ;
        RECT 115.540 211.970 115.860 212.290 ;
        RECT 115.940 211.970 116.260 212.290 ;
        RECT 116.340 211.970 116.660 212.290 ;
        RECT 116.740 211.970 117.060 212.290 ;
        RECT 145.140 211.970 145.460 212.290 ;
        RECT 145.540 211.970 145.860 212.290 ;
        RECT 145.940 211.970 146.260 212.290 ;
        RECT 146.340 211.970 146.660 212.290 ;
        RECT 146.740 211.970 147.060 212.290 ;
        RECT 154.825 211.305 155.215 211.695 ;
        RECT 40.140 209.250 40.460 209.570 ;
        RECT 40.540 209.250 40.860 209.570 ;
        RECT 40.940 209.250 41.260 209.570 ;
        RECT 41.340 209.250 41.660 209.570 ;
        RECT 41.740 209.250 42.060 209.570 ;
        RECT 70.140 209.250 70.460 209.570 ;
        RECT 70.540 209.250 70.860 209.570 ;
        RECT 70.940 209.250 71.260 209.570 ;
        RECT 71.340 209.250 71.660 209.570 ;
        RECT 71.740 209.250 72.060 209.570 ;
        RECT 100.140 209.250 100.460 209.570 ;
        RECT 100.540 209.250 100.860 209.570 ;
        RECT 100.940 209.250 101.260 209.570 ;
        RECT 101.340 209.250 101.660 209.570 ;
        RECT 101.740 209.250 102.060 209.570 ;
        RECT 130.140 209.250 130.460 209.570 ;
        RECT 130.540 209.250 130.860 209.570 ;
        RECT 130.940 209.250 131.260 209.570 ;
        RECT 131.340 209.250 131.660 209.570 ;
        RECT 131.740 209.250 132.060 209.570 ;
        RECT 55.140 206.530 55.460 206.850 ;
        RECT 55.540 206.530 55.860 206.850 ;
        RECT 55.940 206.530 56.260 206.850 ;
        RECT 56.340 206.530 56.660 206.850 ;
        RECT 56.740 206.530 57.060 206.850 ;
        RECT 85.140 206.530 85.460 206.850 ;
        RECT 85.540 206.530 85.860 206.850 ;
        RECT 85.940 206.530 86.260 206.850 ;
        RECT 86.340 206.530 86.660 206.850 ;
        RECT 86.740 206.530 87.060 206.850 ;
        RECT 115.140 206.530 115.460 206.850 ;
        RECT 115.540 206.530 115.860 206.850 ;
        RECT 115.940 206.530 116.260 206.850 ;
        RECT 116.340 206.530 116.660 206.850 ;
        RECT 116.740 206.530 117.060 206.850 ;
        RECT 145.140 206.530 145.460 206.850 ;
        RECT 145.540 206.530 145.860 206.850 ;
        RECT 145.940 206.530 146.260 206.850 ;
        RECT 146.340 206.530 146.660 206.850 ;
        RECT 146.740 206.530 147.060 206.850 ;
        RECT 98.960 205.510 99.280 205.830 ;
        RECT 154.025 205.655 154.375 206.005 ;
        RECT 40.140 203.810 40.460 204.130 ;
        RECT 40.540 203.810 40.860 204.130 ;
        RECT 40.940 203.810 41.260 204.130 ;
        RECT 41.340 203.810 41.660 204.130 ;
        RECT 41.740 203.810 42.060 204.130 ;
        RECT 70.140 203.810 70.460 204.130 ;
        RECT 70.540 203.810 70.860 204.130 ;
        RECT 70.940 203.810 71.260 204.130 ;
        RECT 71.340 203.810 71.660 204.130 ;
        RECT 71.740 203.810 72.060 204.130 ;
        RECT 100.140 203.810 100.460 204.130 ;
        RECT 100.540 203.810 100.860 204.130 ;
        RECT 100.940 203.810 101.260 204.130 ;
        RECT 101.340 203.810 101.660 204.130 ;
        RECT 101.740 203.810 102.060 204.130 ;
        RECT 130.140 203.810 130.460 204.130 ;
        RECT 130.540 203.810 130.860 204.130 ;
        RECT 130.940 203.810 131.260 204.130 ;
        RECT 131.340 203.810 131.660 204.130 ;
        RECT 131.740 203.810 132.060 204.130 ;
        RECT 111.840 202.790 112.160 203.110 ;
        RECT 108.160 201.430 108.480 201.750 ;
        RECT 55.140 201.090 55.460 201.410 ;
        RECT 55.540 201.090 55.860 201.410 ;
        RECT 55.940 201.090 56.260 201.410 ;
        RECT 56.340 201.090 56.660 201.410 ;
        RECT 56.740 201.090 57.060 201.410 ;
        RECT 85.140 201.090 85.460 201.410 ;
        RECT 85.540 201.090 85.860 201.410 ;
        RECT 85.940 201.090 86.260 201.410 ;
        RECT 86.340 201.090 86.660 201.410 ;
        RECT 86.740 201.090 87.060 201.410 ;
        RECT 115.140 201.090 115.460 201.410 ;
        RECT 115.540 201.090 115.860 201.410 ;
        RECT 115.940 201.090 116.260 201.410 ;
        RECT 116.340 201.090 116.660 201.410 ;
        RECT 116.740 201.090 117.060 201.410 ;
        RECT 145.140 201.090 145.460 201.410 ;
        RECT 145.540 201.090 145.860 201.410 ;
        RECT 145.940 201.090 146.260 201.410 ;
        RECT 146.340 201.090 146.660 201.410 ;
        RECT 146.740 201.090 147.060 201.410 ;
        RECT 40.140 198.370 40.460 198.690 ;
        RECT 40.540 198.370 40.860 198.690 ;
        RECT 40.940 198.370 41.260 198.690 ;
        RECT 41.340 198.370 41.660 198.690 ;
        RECT 41.740 198.370 42.060 198.690 ;
        RECT 70.140 198.370 70.460 198.690 ;
        RECT 70.540 198.370 70.860 198.690 ;
        RECT 70.940 198.370 71.260 198.690 ;
        RECT 71.340 198.370 71.660 198.690 ;
        RECT 71.740 198.370 72.060 198.690 ;
        RECT 100.140 198.370 100.460 198.690 ;
        RECT 100.540 198.370 100.860 198.690 ;
        RECT 100.940 198.370 101.260 198.690 ;
        RECT 101.340 198.370 101.660 198.690 ;
        RECT 101.740 198.370 102.060 198.690 ;
        RECT 130.140 198.370 130.460 198.690 ;
        RECT 130.540 198.370 130.860 198.690 ;
        RECT 130.940 198.370 131.260 198.690 ;
        RECT 131.340 198.370 131.660 198.690 ;
        RECT 131.740 198.370 132.060 198.690 ;
        RECT 53.880 195.990 54.200 196.310 ;
        RECT 55.140 195.650 55.460 195.970 ;
        RECT 55.540 195.650 55.860 195.970 ;
        RECT 55.940 195.650 56.260 195.970 ;
        RECT 56.340 195.650 56.660 195.970 ;
        RECT 56.740 195.650 57.060 195.970 ;
        RECT 85.140 195.650 85.460 195.970 ;
        RECT 85.540 195.650 85.860 195.970 ;
        RECT 85.940 195.650 86.260 195.970 ;
        RECT 86.340 195.650 86.660 195.970 ;
        RECT 86.740 195.650 87.060 195.970 ;
        RECT 115.140 195.650 115.460 195.970 ;
        RECT 115.540 195.650 115.860 195.970 ;
        RECT 115.940 195.650 116.260 195.970 ;
        RECT 116.340 195.650 116.660 195.970 ;
        RECT 116.740 195.650 117.060 195.970 ;
        RECT 145.140 195.650 145.460 195.970 ;
        RECT 145.540 195.650 145.860 195.970 ;
        RECT 145.940 195.650 146.260 195.970 ;
        RECT 146.340 195.650 146.660 195.970 ;
        RECT 146.740 195.650 147.060 195.970 ;
        RECT 40.140 192.930 40.460 193.250 ;
        RECT 40.540 192.930 40.860 193.250 ;
        RECT 40.940 192.930 41.260 193.250 ;
        RECT 41.340 192.930 41.660 193.250 ;
        RECT 41.740 192.930 42.060 193.250 ;
        RECT 70.140 192.930 70.460 193.250 ;
        RECT 70.540 192.930 70.860 193.250 ;
        RECT 70.940 192.930 71.260 193.250 ;
        RECT 71.340 192.930 71.660 193.250 ;
        RECT 71.740 192.930 72.060 193.250 ;
        RECT 100.140 192.930 100.460 193.250 ;
        RECT 100.540 192.930 100.860 193.250 ;
        RECT 100.940 192.930 101.260 193.250 ;
        RECT 101.340 192.930 101.660 193.250 ;
        RECT 101.740 192.930 102.060 193.250 ;
        RECT 130.140 192.930 130.460 193.250 ;
        RECT 130.540 192.930 130.860 193.250 ;
        RECT 130.940 192.930 131.260 193.250 ;
        RECT 131.340 192.930 131.660 193.250 ;
        RECT 131.740 192.930 132.060 193.250 ;
        RECT 55.140 190.210 55.460 190.530 ;
        RECT 55.540 190.210 55.860 190.530 ;
        RECT 55.940 190.210 56.260 190.530 ;
        RECT 56.340 190.210 56.660 190.530 ;
        RECT 56.740 190.210 57.060 190.530 ;
        RECT 85.140 190.210 85.460 190.530 ;
        RECT 85.540 190.210 85.860 190.530 ;
        RECT 85.940 190.210 86.260 190.530 ;
        RECT 86.340 190.210 86.660 190.530 ;
        RECT 86.740 190.210 87.060 190.530 ;
        RECT 115.140 190.210 115.460 190.530 ;
        RECT 115.540 190.210 115.860 190.530 ;
        RECT 115.940 190.210 116.260 190.530 ;
        RECT 116.340 190.210 116.660 190.530 ;
        RECT 116.740 190.210 117.060 190.530 ;
        RECT 145.140 190.210 145.460 190.530 ;
        RECT 145.540 190.210 145.860 190.530 ;
        RECT 145.940 190.210 146.260 190.530 ;
        RECT 146.340 190.210 146.660 190.530 ;
        RECT 146.740 190.210 147.060 190.530 ;
        RECT 109.080 189.870 109.400 190.190 ;
        RECT 40.140 187.490 40.460 187.810 ;
        RECT 40.540 187.490 40.860 187.810 ;
        RECT 40.940 187.490 41.260 187.810 ;
        RECT 41.340 187.490 41.660 187.810 ;
        RECT 41.740 187.490 42.060 187.810 ;
        RECT 70.140 187.490 70.460 187.810 ;
        RECT 70.540 187.490 70.860 187.810 ;
        RECT 70.940 187.490 71.260 187.810 ;
        RECT 71.340 187.490 71.660 187.810 ;
        RECT 71.740 187.490 72.060 187.810 ;
        RECT 100.140 187.490 100.460 187.810 ;
        RECT 100.540 187.490 100.860 187.810 ;
        RECT 100.940 187.490 101.260 187.810 ;
        RECT 101.340 187.490 101.660 187.810 ;
        RECT 101.740 187.490 102.060 187.810 ;
        RECT 130.140 187.490 130.460 187.810 ;
        RECT 130.540 187.490 130.860 187.810 ;
        RECT 130.940 187.490 131.260 187.810 ;
        RECT 131.340 187.490 131.660 187.810 ;
        RECT 131.740 187.490 132.060 187.810 ;
        RECT 82.400 187.150 82.720 187.470 ;
        RECT 88.840 185.790 89.160 186.110 ;
        RECT 55.140 184.770 55.460 185.090 ;
        RECT 55.540 184.770 55.860 185.090 ;
        RECT 55.940 184.770 56.260 185.090 ;
        RECT 56.340 184.770 56.660 185.090 ;
        RECT 56.740 184.770 57.060 185.090 ;
        RECT 85.140 184.770 85.460 185.090 ;
        RECT 85.540 184.770 85.860 185.090 ;
        RECT 85.940 184.770 86.260 185.090 ;
        RECT 86.340 184.770 86.660 185.090 ;
        RECT 86.740 184.770 87.060 185.090 ;
        RECT 115.140 184.770 115.460 185.090 ;
        RECT 115.540 184.770 115.860 185.090 ;
        RECT 115.940 184.770 116.260 185.090 ;
        RECT 116.340 184.770 116.660 185.090 ;
        RECT 116.740 184.770 117.060 185.090 ;
        RECT 145.140 184.770 145.460 185.090 ;
        RECT 145.540 184.770 145.860 185.090 ;
        RECT 145.940 184.770 146.260 185.090 ;
        RECT 146.340 184.770 146.660 185.090 ;
        RECT 146.740 184.770 147.060 185.090 ;
        RECT 107.240 184.430 107.560 184.750 ;
        RECT 133.000 184.430 133.320 184.750 ;
        RECT 40.140 182.050 40.460 182.370 ;
        RECT 40.540 182.050 40.860 182.370 ;
        RECT 40.940 182.050 41.260 182.370 ;
        RECT 41.340 182.050 41.660 182.370 ;
        RECT 41.740 182.050 42.060 182.370 ;
        RECT 70.140 182.050 70.460 182.370 ;
        RECT 70.540 182.050 70.860 182.370 ;
        RECT 70.940 182.050 71.260 182.370 ;
        RECT 71.340 182.050 71.660 182.370 ;
        RECT 71.740 182.050 72.060 182.370 ;
        RECT 100.140 182.050 100.460 182.370 ;
        RECT 100.540 182.050 100.860 182.370 ;
        RECT 100.940 182.050 101.260 182.370 ;
        RECT 101.340 182.050 101.660 182.370 ;
        RECT 101.740 182.050 102.060 182.370 ;
        RECT 130.140 182.050 130.460 182.370 ;
        RECT 130.540 182.050 130.860 182.370 ;
        RECT 130.940 182.050 131.260 182.370 ;
        RECT 131.340 182.050 131.660 182.370 ;
        RECT 131.740 182.050 132.060 182.370 ;
        RECT 133.000 179.670 133.320 179.990 ;
        RECT 55.140 179.330 55.460 179.650 ;
        RECT 55.540 179.330 55.860 179.650 ;
        RECT 55.940 179.330 56.260 179.650 ;
        RECT 56.340 179.330 56.660 179.650 ;
        RECT 56.740 179.330 57.060 179.650 ;
        RECT 85.140 179.330 85.460 179.650 ;
        RECT 85.540 179.330 85.860 179.650 ;
        RECT 85.940 179.330 86.260 179.650 ;
        RECT 86.340 179.330 86.660 179.650 ;
        RECT 86.740 179.330 87.060 179.650 ;
        RECT 115.140 179.330 115.460 179.650 ;
        RECT 115.540 179.330 115.860 179.650 ;
        RECT 115.940 179.330 116.260 179.650 ;
        RECT 116.340 179.330 116.660 179.650 ;
        RECT 116.740 179.330 117.060 179.650 ;
        RECT 145.140 179.330 145.460 179.650 ;
        RECT 145.540 179.330 145.860 179.650 ;
        RECT 145.940 179.330 146.260 179.650 ;
        RECT 146.340 179.330 146.660 179.650 ;
        RECT 146.740 179.330 147.060 179.650 ;
        RECT 53.880 177.630 54.200 177.950 ;
        RECT 40.140 176.610 40.460 176.930 ;
        RECT 40.540 176.610 40.860 176.930 ;
        RECT 40.940 176.610 41.260 176.930 ;
        RECT 41.340 176.610 41.660 176.930 ;
        RECT 41.740 176.610 42.060 176.930 ;
        RECT 70.140 176.610 70.460 176.930 ;
        RECT 70.540 176.610 70.860 176.930 ;
        RECT 70.940 176.610 71.260 176.930 ;
        RECT 71.340 176.610 71.660 176.930 ;
        RECT 71.740 176.610 72.060 176.930 ;
        RECT 100.140 176.610 100.460 176.930 ;
        RECT 100.540 176.610 100.860 176.930 ;
        RECT 100.940 176.610 101.260 176.930 ;
        RECT 101.340 176.610 101.660 176.930 ;
        RECT 101.740 176.610 102.060 176.930 ;
        RECT 130.140 176.610 130.460 176.930 ;
        RECT 130.540 176.610 130.860 176.930 ;
        RECT 130.940 176.610 131.260 176.930 ;
        RECT 131.340 176.610 131.660 176.930 ;
        RECT 131.740 176.610 132.060 176.930 ;
        RECT 82.400 174.910 82.720 175.230 ;
        RECT 55.140 173.890 55.460 174.210 ;
        RECT 55.540 173.890 55.860 174.210 ;
        RECT 55.940 173.890 56.260 174.210 ;
        RECT 56.340 173.890 56.660 174.210 ;
        RECT 56.740 173.890 57.060 174.210 ;
        RECT 85.140 173.890 85.460 174.210 ;
        RECT 85.540 173.890 85.860 174.210 ;
        RECT 85.940 173.890 86.260 174.210 ;
        RECT 86.340 173.890 86.660 174.210 ;
        RECT 86.740 173.890 87.060 174.210 ;
        RECT 115.140 173.890 115.460 174.210 ;
        RECT 115.540 173.890 115.860 174.210 ;
        RECT 115.940 173.890 116.260 174.210 ;
        RECT 116.340 173.890 116.660 174.210 ;
        RECT 116.740 173.890 117.060 174.210 ;
        RECT 145.140 173.890 145.460 174.210 ;
        RECT 145.540 173.890 145.860 174.210 ;
        RECT 145.940 173.890 146.260 174.210 ;
        RECT 146.340 173.890 146.660 174.210 ;
        RECT 146.740 173.890 147.060 174.210 ;
        RECT 111.840 172.870 112.160 173.190 ;
        RECT 40.140 171.170 40.460 171.490 ;
        RECT 40.540 171.170 40.860 171.490 ;
        RECT 40.940 171.170 41.260 171.490 ;
        RECT 41.340 171.170 41.660 171.490 ;
        RECT 41.740 171.170 42.060 171.490 ;
        RECT 70.140 171.170 70.460 171.490 ;
        RECT 70.540 171.170 70.860 171.490 ;
        RECT 70.940 171.170 71.260 171.490 ;
        RECT 71.340 171.170 71.660 171.490 ;
        RECT 71.740 171.170 72.060 171.490 ;
        RECT 100.140 171.170 100.460 171.490 ;
        RECT 100.540 171.170 100.860 171.490 ;
        RECT 100.940 171.170 101.260 171.490 ;
        RECT 101.340 171.170 101.660 171.490 ;
        RECT 101.740 171.170 102.060 171.490 ;
        RECT 130.140 171.170 130.460 171.490 ;
        RECT 130.540 171.170 130.860 171.490 ;
        RECT 130.940 171.170 131.260 171.490 ;
        RECT 131.340 171.170 131.660 171.490 ;
        RECT 131.740 171.170 132.060 171.490 ;
        RECT 55.140 168.450 55.460 168.770 ;
        RECT 55.540 168.450 55.860 168.770 ;
        RECT 55.940 168.450 56.260 168.770 ;
        RECT 56.340 168.450 56.660 168.770 ;
        RECT 56.740 168.450 57.060 168.770 ;
        RECT 85.140 168.450 85.460 168.770 ;
        RECT 85.540 168.450 85.860 168.770 ;
        RECT 85.940 168.450 86.260 168.770 ;
        RECT 86.340 168.450 86.660 168.770 ;
        RECT 86.740 168.450 87.060 168.770 ;
        RECT 115.140 168.450 115.460 168.770 ;
        RECT 115.540 168.450 115.860 168.770 ;
        RECT 115.940 168.450 116.260 168.770 ;
        RECT 116.340 168.450 116.660 168.770 ;
        RECT 116.740 168.450 117.060 168.770 ;
        RECT 145.140 168.450 145.460 168.770 ;
        RECT 145.540 168.450 145.860 168.770 ;
        RECT 145.940 168.450 146.260 168.770 ;
        RECT 146.340 168.450 146.660 168.770 ;
        RECT 146.740 168.450 147.060 168.770 ;
        RECT 107.240 167.430 107.560 167.750 ;
        RECT 136.680 166.750 137.000 167.070 ;
        RECT 109.080 166.070 109.400 166.390 ;
        RECT 113.680 166.070 114.000 166.390 ;
        RECT 40.140 165.730 40.460 166.050 ;
        RECT 40.540 165.730 40.860 166.050 ;
        RECT 40.940 165.730 41.260 166.050 ;
        RECT 41.340 165.730 41.660 166.050 ;
        RECT 41.740 165.730 42.060 166.050 ;
        RECT 70.140 165.730 70.460 166.050 ;
        RECT 70.540 165.730 70.860 166.050 ;
        RECT 70.940 165.730 71.260 166.050 ;
        RECT 71.340 165.730 71.660 166.050 ;
        RECT 71.740 165.730 72.060 166.050 ;
        RECT 100.140 165.730 100.460 166.050 ;
        RECT 100.540 165.730 100.860 166.050 ;
        RECT 100.940 165.730 101.260 166.050 ;
        RECT 101.340 165.730 101.660 166.050 ;
        RECT 101.740 165.730 102.060 166.050 ;
        RECT 130.140 165.730 130.460 166.050 ;
        RECT 130.540 165.730 130.860 166.050 ;
        RECT 130.940 165.730 131.260 166.050 ;
        RECT 131.340 165.730 131.660 166.050 ;
        RECT 131.740 165.730 132.060 166.050 ;
        RECT 83.320 165.390 83.640 165.710 ;
        RECT 82.400 164.030 82.720 164.350 ;
        RECT 55.140 163.010 55.460 163.330 ;
        RECT 55.540 163.010 55.860 163.330 ;
        RECT 55.940 163.010 56.260 163.330 ;
        RECT 56.340 163.010 56.660 163.330 ;
        RECT 56.740 163.010 57.060 163.330 ;
        RECT 85.140 163.010 85.460 163.330 ;
        RECT 85.540 163.010 85.860 163.330 ;
        RECT 85.940 163.010 86.260 163.330 ;
        RECT 86.340 163.010 86.660 163.330 ;
        RECT 86.740 163.010 87.060 163.330 ;
        RECT 115.140 163.010 115.460 163.330 ;
        RECT 115.540 163.010 115.860 163.330 ;
        RECT 115.940 163.010 116.260 163.330 ;
        RECT 116.340 163.010 116.660 163.330 ;
        RECT 116.740 163.010 117.060 163.330 ;
        RECT 145.140 163.010 145.460 163.330 ;
        RECT 145.540 163.010 145.860 163.330 ;
        RECT 145.940 163.010 146.260 163.330 ;
        RECT 146.340 163.010 146.660 163.330 ;
        RECT 146.740 163.010 147.060 163.330 ;
        RECT 40.140 160.290 40.460 160.610 ;
        RECT 40.540 160.290 40.860 160.610 ;
        RECT 40.940 160.290 41.260 160.610 ;
        RECT 41.340 160.290 41.660 160.610 ;
        RECT 41.740 160.290 42.060 160.610 ;
        RECT 70.140 160.290 70.460 160.610 ;
        RECT 70.540 160.290 70.860 160.610 ;
        RECT 70.940 160.290 71.260 160.610 ;
        RECT 71.340 160.290 71.660 160.610 ;
        RECT 71.740 160.290 72.060 160.610 ;
        RECT 100.140 160.290 100.460 160.610 ;
        RECT 100.540 160.290 100.860 160.610 ;
        RECT 100.940 160.290 101.260 160.610 ;
        RECT 101.340 160.290 101.660 160.610 ;
        RECT 101.740 160.290 102.060 160.610 ;
        RECT 130.140 160.290 130.460 160.610 ;
        RECT 130.540 160.290 130.860 160.610 ;
        RECT 130.940 160.290 131.260 160.610 ;
        RECT 131.340 160.290 131.660 160.610 ;
        RECT 131.740 160.290 132.060 160.610 ;
        RECT 80.560 157.910 80.880 158.230 ;
        RECT 55.140 157.570 55.460 157.890 ;
        RECT 55.540 157.570 55.860 157.890 ;
        RECT 55.940 157.570 56.260 157.890 ;
        RECT 56.340 157.570 56.660 157.890 ;
        RECT 56.740 157.570 57.060 157.890 ;
        RECT 85.140 157.570 85.460 157.890 ;
        RECT 85.540 157.570 85.860 157.890 ;
        RECT 85.940 157.570 86.260 157.890 ;
        RECT 86.340 157.570 86.660 157.890 ;
        RECT 86.740 157.570 87.060 157.890 ;
        RECT 115.140 157.570 115.460 157.890 ;
        RECT 115.540 157.570 115.860 157.890 ;
        RECT 115.940 157.570 116.260 157.890 ;
        RECT 116.340 157.570 116.660 157.890 ;
        RECT 116.740 157.570 117.060 157.890 ;
        RECT 145.140 157.570 145.460 157.890 ;
        RECT 145.540 157.570 145.860 157.890 ;
        RECT 145.940 157.570 146.260 157.890 ;
        RECT 146.340 157.570 146.660 157.890 ;
        RECT 146.740 157.570 147.060 157.890 ;
        RECT 82.400 157.230 82.720 157.550 ;
        RECT 78.720 155.190 79.040 155.510 ;
        RECT 88.840 155.190 89.160 155.510 ;
        RECT 40.140 154.850 40.460 155.170 ;
        RECT 40.540 154.850 40.860 155.170 ;
        RECT 40.940 154.850 41.260 155.170 ;
        RECT 41.340 154.850 41.660 155.170 ;
        RECT 41.740 154.850 42.060 155.170 ;
        RECT 70.140 154.850 70.460 155.170 ;
        RECT 70.540 154.850 70.860 155.170 ;
        RECT 70.940 154.850 71.260 155.170 ;
        RECT 71.340 154.850 71.660 155.170 ;
        RECT 71.740 154.850 72.060 155.170 ;
        RECT 100.140 154.850 100.460 155.170 ;
        RECT 100.540 154.850 100.860 155.170 ;
        RECT 100.940 154.850 101.260 155.170 ;
        RECT 101.340 154.850 101.660 155.170 ;
        RECT 101.740 154.850 102.060 155.170 ;
        RECT 130.140 154.850 130.460 155.170 ;
        RECT 130.540 154.850 130.860 155.170 ;
        RECT 130.940 154.850 131.260 155.170 ;
        RECT 131.340 154.850 131.660 155.170 ;
        RECT 131.740 154.850 132.060 155.170 ;
        RECT 79.640 153.830 79.960 154.150 ;
        RECT 82.400 152.470 82.720 152.790 ;
        RECT 55.140 152.130 55.460 152.450 ;
        RECT 55.540 152.130 55.860 152.450 ;
        RECT 55.940 152.130 56.260 152.450 ;
        RECT 56.340 152.130 56.660 152.450 ;
        RECT 56.740 152.130 57.060 152.450 ;
        RECT 85.140 152.130 85.460 152.450 ;
        RECT 85.540 152.130 85.860 152.450 ;
        RECT 85.940 152.130 86.260 152.450 ;
        RECT 86.340 152.130 86.660 152.450 ;
        RECT 86.740 152.130 87.060 152.450 ;
        RECT 115.140 152.130 115.460 152.450 ;
        RECT 115.540 152.130 115.860 152.450 ;
        RECT 115.940 152.130 116.260 152.450 ;
        RECT 116.340 152.130 116.660 152.450 ;
        RECT 116.740 152.130 117.060 152.450 ;
        RECT 145.140 152.130 145.460 152.450 ;
        RECT 145.540 152.130 145.860 152.450 ;
        RECT 145.940 152.130 146.260 152.450 ;
        RECT 146.340 152.130 146.660 152.450 ;
        RECT 146.740 152.130 147.060 152.450 ;
        RECT 78.720 151.790 79.040 152.110 ;
        RECT 98.960 151.790 99.280 152.110 ;
        RECT 136.680 151.790 137.000 152.110 ;
        RECT 79.640 150.430 79.960 150.750 ;
        RECT 40.140 149.410 40.460 149.730 ;
        RECT 40.540 149.410 40.860 149.730 ;
        RECT 40.940 149.410 41.260 149.730 ;
        RECT 41.340 149.410 41.660 149.730 ;
        RECT 41.740 149.410 42.060 149.730 ;
        RECT 70.140 149.410 70.460 149.730 ;
        RECT 70.540 149.410 70.860 149.730 ;
        RECT 70.940 149.410 71.260 149.730 ;
        RECT 71.340 149.410 71.660 149.730 ;
        RECT 71.740 149.410 72.060 149.730 ;
        RECT 100.140 149.410 100.460 149.730 ;
        RECT 100.540 149.410 100.860 149.730 ;
        RECT 100.940 149.410 101.260 149.730 ;
        RECT 101.340 149.410 101.660 149.730 ;
        RECT 101.740 149.410 102.060 149.730 ;
        RECT 130.140 149.410 130.460 149.730 ;
        RECT 130.540 149.410 130.860 149.730 ;
        RECT 130.940 149.410 131.260 149.730 ;
        RECT 131.340 149.410 131.660 149.730 ;
        RECT 131.740 149.410 132.060 149.730 ;
        RECT 108.160 149.070 108.480 149.390 ;
        RECT 80.560 147.030 80.880 147.350 ;
        RECT 55.140 146.690 55.460 147.010 ;
        RECT 55.540 146.690 55.860 147.010 ;
        RECT 55.940 146.690 56.260 147.010 ;
        RECT 56.340 146.690 56.660 147.010 ;
        RECT 56.740 146.690 57.060 147.010 ;
        RECT 85.140 146.690 85.460 147.010 ;
        RECT 85.540 146.690 85.860 147.010 ;
        RECT 85.940 146.690 86.260 147.010 ;
        RECT 86.340 146.690 86.660 147.010 ;
        RECT 86.740 146.690 87.060 147.010 ;
        RECT 115.140 146.690 115.460 147.010 ;
        RECT 115.540 146.690 115.860 147.010 ;
        RECT 115.940 146.690 116.260 147.010 ;
        RECT 116.340 146.690 116.660 147.010 ;
        RECT 116.740 146.690 117.060 147.010 ;
        RECT 145.140 146.690 145.460 147.010 ;
        RECT 145.540 146.690 145.860 147.010 ;
        RECT 145.940 146.690 146.260 147.010 ;
        RECT 146.340 146.690 146.660 147.010 ;
        RECT 146.740 146.690 147.060 147.010 ;
        RECT 113.680 145.670 114.000 145.990 ;
        RECT 40.140 143.970 40.460 144.290 ;
        RECT 40.540 143.970 40.860 144.290 ;
        RECT 40.940 143.970 41.260 144.290 ;
        RECT 41.340 143.970 41.660 144.290 ;
        RECT 41.740 143.970 42.060 144.290 ;
        RECT 70.140 143.970 70.460 144.290 ;
        RECT 70.540 143.970 70.860 144.290 ;
        RECT 70.940 143.970 71.260 144.290 ;
        RECT 71.340 143.970 71.660 144.290 ;
        RECT 71.740 143.970 72.060 144.290 ;
        RECT 100.140 143.970 100.460 144.290 ;
        RECT 100.540 143.970 100.860 144.290 ;
        RECT 100.940 143.970 101.260 144.290 ;
        RECT 101.340 143.970 101.660 144.290 ;
        RECT 101.740 143.970 102.060 144.290 ;
        RECT 130.140 143.970 130.460 144.290 ;
        RECT 130.540 143.970 130.860 144.290 ;
        RECT 130.940 143.970 131.260 144.290 ;
        RECT 131.340 143.970 131.660 144.290 ;
        RECT 131.740 143.970 132.060 144.290 ;
        RECT 83.320 142.950 83.640 143.270 ;
        RECT 55.140 141.250 55.460 141.570 ;
        RECT 55.540 141.250 55.860 141.570 ;
        RECT 55.940 141.250 56.260 141.570 ;
        RECT 56.340 141.250 56.660 141.570 ;
        RECT 56.740 141.250 57.060 141.570 ;
        RECT 85.140 141.250 85.460 141.570 ;
        RECT 85.540 141.250 85.860 141.570 ;
        RECT 85.940 141.250 86.260 141.570 ;
        RECT 86.340 141.250 86.660 141.570 ;
        RECT 86.740 141.250 87.060 141.570 ;
        RECT 115.140 141.250 115.460 141.570 ;
        RECT 115.540 141.250 115.860 141.570 ;
        RECT 115.940 141.250 116.260 141.570 ;
        RECT 116.340 141.250 116.660 141.570 ;
        RECT 116.740 141.250 117.060 141.570 ;
        RECT 145.140 141.250 145.460 141.570 ;
        RECT 145.540 141.250 145.860 141.570 ;
        RECT 145.940 141.250 146.260 141.570 ;
        RECT 146.340 141.250 146.660 141.570 ;
        RECT 146.740 141.250 147.060 141.570 ;
        RECT 3.455 135.955 4.945 137.445 ;
        RECT 43.005 135.705 44.995 137.695 ;
        RECT 70.105 135.705 72.095 137.695 ;
        RECT 96.805 135.705 98.795 137.695 ;
        RECT 130.105 135.705 132.095 137.695 ;
        RECT 12.655 133.155 14.145 134.645 ;
        RECT 55.105 132.805 57.095 134.795 ;
        RECT 84.305 132.805 86.295 134.795 ;
        RECT 112.205 132.805 114.195 134.795 ;
        RECT 147.805 132.805 149.795 134.795 ;
        RECT 156.395 51.635 157.325 52.565 ;
        RECT 134.345 49.460 135.220 50.335 ;
        RECT 130.670 47.270 131.525 48.125 ;
        RECT 17.100 22.000 18.100 23.000 ;
        RECT 5.900 15.615 6.900 16.615 ;
        RECT 35.600 5.700 36.600 6.700 ;
      LAYER met4 ;
        RECT 3.990 220.800 4.290 224.760 ;
        RECT 7.670 222.300 7.970 224.760 ;
        RECT 11.350 222.300 11.650 224.760 ;
        RECT 15.030 222.300 15.330 224.760 ;
        RECT 18.710 222.300 19.010 224.760 ;
        RECT 22.390 222.300 22.690 224.760 ;
        RECT 26.070 222.300 26.370 224.760 ;
        RECT 29.750 222.300 30.050 224.760 ;
        RECT 33.430 222.300 33.730 224.760 ;
        RECT 37.110 222.300 37.410 224.760 ;
        RECT 40.790 222.300 41.090 224.760 ;
        RECT 44.470 222.300 44.770 224.760 ;
        RECT 48.150 222.300 48.450 224.760 ;
        RECT 51.830 223.165 52.130 224.760 ;
        RECT 51.815 222.835 52.145 223.165 ;
        RECT 55.510 223.095 55.810 224.760 ;
        RECT 59.190 223.095 59.490 224.760 ;
        RECT 62.870 223.095 63.170 224.760 ;
        RECT 66.550 223.095 66.850 224.760 ;
        RECT 70.230 223.095 70.530 224.760 ;
        RECT 73.910 223.095 74.210 224.760 ;
        RECT 77.590 223.095 77.890 224.760 ;
        RECT 81.270 223.095 81.570 224.760 ;
        RECT 84.950 223.095 85.250 224.760 ;
        RECT 88.630 223.095 88.930 224.760 ;
        RECT 92.310 224.540 92.610 224.760 ;
        RECT 92.160 223.950 92.640 224.540 ;
        RECT 92.155 223.460 92.645 223.950 ;
        RECT 55.495 222.765 55.825 223.095 ;
        RECT 59.175 222.765 59.505 223.095 ;
        RECT 62.855 222.765 63.185 223.095 ;
        RECT 66.535 222.765 66.865 223.095 ;
        RECT 70.215 222.765 70.545 223.095 ;
        RECT 73.895 222.765 74.225 223.095 ;
        RECT 77.575 222.765 77.905 223.095 ;
        RECT 81.255 222.765 81.585 223.095 ;
        RECT 84.935 222.765 85.265 223.095 ;
        RECT 88.615 222.765 88.945 223.095 ;
        RECT 55.510 222.700 55.810 222.765 ;
        RECT 59.190 222.700 59.490 222.765 ;
        RECT 62.870 222.700 63.170 222.765 ;
        RECT 66.550 222.700 66.850 222.765 ;
        RECT 70.230 222.700 70.530 222.765 ;
        RECT 73.910 222.700 74.210 222.765 ;
        RECT 77.590 222.700 77.890 222.765 ;
        RECT 81.270 222.700 81.570 222.765 ;
        RECT 84.950 222.700 85.250 222.765 ;
        RECT 7.400 222.190 19.010 222.300 ;
        RECT 7.400 221.050 19.000 222.190 ;
        RECT 22.200 221.800 30.100 222.300 ;
        RECT 31.350 221.800 48.700 222.300 ;
        RECT 20.645 221.050 21.155 221.055 ;
        RECT 7.400 220.800 21.155 221.050 ;
        RECT 3.990 220.760 21.155 220.800 ;
        RECT 3.990 220.500 10.500 220.760 ;
        RECT 7.400 219.600 10.500 220.500 ;
        RECT 12.000 220.550 21.155 220.760 ;
        RECT 12.000 219.600 19.000 220.550 ;
        RECT 20.645 220.545 21.155 220.550 ;
        RECT 22.200 219.600 23.000 221.800 ;
        RECT 95.990 220.705 96.290 224.760 ;
        RECT 95.935 220.295 96.345 220.705 ;
        RECT 95.990 220.200 96.290 220.295 ;
        RECT 99.670 219.905 99.970 224.760 ;
        RECT 12.595 218.400 13.005 218.405 ;
        RECT 22.400 218.400 22.800 219.600 ;
        RECT 99.620 219.500 100.025 219.905 ;
        RECT 99.670 219.400 99.970 219.500 ;
        RECT 103.350 219.100 103.650 224.760 ;
        RECT 103.305 218.705 103.700 219.100 ;
        RECT 103.350 218.600 103.650 218.705 ;
        RECT 2.500 218.000 9.700 218.400 ;
        RECT 12.595 218.000 22.800 218.400 ;
        RECT 107.030 218.300 107.330 224.760 ;
        RECT 110.710 224.270 111.010 224.760 ;
        RECT 114.390 224.270 114.690 224.760 ;
        RECT 118.070 224.270 118.370 224.760 ;
        RECT 121.750 223.095 122.050 224.760 ;
        RECT 125.430 223.095 125.730 224.760 ;
        RECT 129.110 223.095 129.410 224.760 ;
        RECT 132.790 223.095 133.090 224.760 ;
        RECT 136.470 223.095 136.770 224.760 ;
        RECT 140.150 223.095 140.450 224.760 ;
        RECT 143.830 223.095 144.130 224.760 ;
        RECT 147.510 223.095 147.810 224.760 ;
        RECT 121.735 222.765 122.065 223.095 ;
        RECT 125.415 222.765 125.745 223.095 ;
        RECT 129.095 222.765 129.425 223.095 ;
        RECT 132.775 222.765 133.105 223.095 ;
        RECT 136.455 222.765 136.785 223.095 ;
        RECT 140.135 222.765 140.465 223.095 ;
        RECT 143.815 222.765 144.145 223.095 ;
        RECT 147.495 222.765 147.825 223.095 ;
        RECT 151.190 221.280 151.490 224.760 ;
        RECT 151.190 220.980 153.000 221.280 ;
        RECT 12.595 217.995 13.005 218.000 ;
        RECT 106.980 217.900 107.380 218.300 ;
        RECT 107.030 217.800 107.330 217.900 ;
        RECT 40.100 143.200 42.100 215.090 ;
        RECT 53.875 195.985 54.205 196.315 ;
        RECT 53.890 177.955 54.190 195.985 ;
        RECT 53.875 177.625 54.205 177.955 ;
        RECT 40.100 141.200 45.000 143.200 ;
        RECT 40.100 141.170 42.100 141.200 ;
        RECT 2.500 135.950 4.950 137.450 ;
        RECT 43.000 135.700 45.000 141.200 ;
        RECT 12.000 133.150 14.150 134.650 ;
        RECT 55.100 132.800 57.100 215.090 ;
        RECT 70.100 135.700 72.100 215.090 ;
        RECT 82.395 187.145 82.725 187.475 ;
        RECT 82.410 175.235 82.710 187.145 ;
        RECT 82.395 174.905 82.725 175.235 ;
        RECT 82.410 164.355 82.710 174.905 ;
        RECT 83.315 165.385 83.645 165.715 ;
        RECT 82.395 164.025 82.725 164.355 ;
        RECT 80.555 157.905 80.885 158.235 ;
        RECT 78.715 155.185 79.045 155.515 ;
        RECT 78.730 152.115 79.030 155.185 ;
        RECT 79.635 153.825 79.965 154.155 ;
        RECT 78.715 151.785 79.045 152.115 ;
        RECT 79.650 150.755 79.950 153.825 ;
        RECT 79.635 150.425 79.965 150.755 ;
        RECT 80.570 147.355 80.870 157.905 ;
        RECT 82.395 157.225 82.725 157.555 ;
        RECT 82.410 152.795 82.710 157.225 ;
        RECT 82.395 152.465 82.725 152.795 ;
        RECT 80.555 147.025 80.885 147.355 ;
        RECT 83.330 143.275 83.630 165.385 ;
        RECT 85.100 144.000 87.100 215.090 ;
        RECT 98.955 205.505 99.285 205.835 ;
        RECT 88.835 185.785 89.165 186.115 ;
        RECT 88.850 155.515 89.150 185.785 ;
        RECT 88.835 155.185 89.165 155.515 ;
        RECT 98.970 152.115 99.270 205.505 ;
        RECT 98.955 151.785 99.285 152.115 ;
        RECT 83.315 142.945 83.645 143.275 ;
        RECT 84.300 142.000 87.600 144.000 ;
        RECT 100.100 143.170 102.100 215.090 ;
        RECT 111.835 202.785 112.165 203.115 ;
        RECT 108.155 201.425 108.485 201.755 ;
        RECT 107.235 184.425 107.565 184.755 ;
        RECT 107.250 167.755 107.550 184.425 ;
        RECT 107.235 167.425 107.565 167.755 ;
        RECT 108.170 149.395 108.470 201.425 ;
        RECT 109.075 189.865 109.405 190.195 ;
        RECT 109.090 166.395 109.390 189.865 ;
        RECT 111.850 173.195 112.150 202.785 ;
        RECT 111.835 172.865 112.165 173.195 ;
        RECT 109.075 166.065 109.405 166.395 ;
        RECT 113.675 166.065 114.005 166.395 ;
        RECT 108.155 149.065 108.485 149.395 ;
        RECT 113.690 145.995 113.990 166.065 ;
        RECT 113.675 145.665 114.005 145.995 ;
        RECT 115.100 143.570 117.100 215.090 ;
        RECT 84.300 141.170 87.100 142.000 ;
        RECT 96.800 141.170 102.100 143.170 ;
        RECT 112.200 141.570 117.100 143.570 ;
        RECT 84.300 132.800 86.300 141.170 ;
        RECT 96.800 135.700 98.800 141.170 ;
        RECT 112.200 132.800 114.200 141.570 ;
        RECT 115.100 141.170 117.100 141.570 ;
        RECT 130.100 135.700 132.100 215.090 ;
        RECT 132.995 184.425 133.325 184.755 ;
        RECT 133.010 179.995 133.310 184.425 ;
        RECT 132.995 179.665 133.325 179.995 ;
        RECT 136.675 166.745 137.005 167.075 ;
        RECT 136.690 152.115 136.990 166.745 ;
        RECT 136.675 151.785 137.005 152.115 ;
        RECT 145.100 143.570 147.100 215.090 ;
        RECT 152.700 210.120 153.000 220.980 ;
        RECT 154.870 211.700 155.170 224.760 ;
        RECT 154.820 211.300 155.220 211.700 ;
        RECT 152.700 209.820 154.350 210.120 ;
        RECT 154.050 206.010 154.350 209.820 ;
        RECT 154.020 205.650 154.380 206.010 ;
        RECT 145.100 141.570 149.800 143.570 ;
        RECT 145.100 141.170 147.100 141.570 ;
        RECT 147.800 132.800 149.800 141.570 ;
        RECT 17.095 23.000 18.105 23.005 ;
        RECT 12.000 22.000 18.105 23.000 ;
        RECT 17.095 21.995 18.105 22.000 ;
        RECT 5.895 16.615 6.905 16.620 ;
        RECT 2.500 15.615 6.905 16.615 ;
        RECT 5.895 15.610 6.905 15.615 ;
        RECT 35.595 5.695 36.605 6.705 ;
        RECT 35.600 3.800 36.600 5.695 ;
        RECT 130.665 4.135 131.530 48.130 ;
        RECT 35.600 3.600 89.900 3.800 ;
        RECT 35.600 3.000 90.920 3.600 ;
        RECT 112.270 3.270 131.530 4.135 ;
        RECT 134.340 3.860 135.225 50.340 ;
        RECT 156.390 4.230 157.330 52.570 ;
        RECT 35.600 2.800 89.900 3.000 ;
        RECT 46.160 1.000 46.760 1.400 ;
        RECT 90.320 1.000 90.920 3.000 ;
        RECT 112.400 1.000 113.000 3.270 ;
        RECT 134.480 1.000 135.080 3.860 ;
        RECT 156.560 1.000 157.160 4.230 ;
  END
END tt_um_algofoogle_tt06_grab_bag
END LIBRARY

