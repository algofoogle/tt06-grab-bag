magic
tech sky130A
magscale 1 2
timestamp 1713537803
<< pwell >>
rect -225 2441 225 2527
rect -225 -2441 -139 2441
rect 139 -2441 225 2441
rect -225 -2527 225 -2441
<< psubdiff >>
rect -199 2467 -85 2501
rect -51 2467 -17 2501
rect 17 2467 51 2501
rect 85 2467 199 2501
rect -199 2397 -165 2467
rect 165 2397 199 2467
rect -199 2329 -165 2363
rect -199 2261 -165 2295
rect -199 2193 -165 2227
rect -199 2125 -165 2159
rect -199 2057 -165 2091
rect -199 1989 -165 2023
rect -199 1921 -165 1955
rect -199 1853 -165 1887
rect -199 1785 -165 1819
rect -199 1717 -165 1751
rect -199 1649 -165 1683
rect -199 1581 -165 1615
rect -199 1513 -165 1547
rect -199 1445 -165 1479
rect -199 1377 -165 1411
rect -199 1309 -165 1343
rect -199 1241 -165 1275
rect -199 1173 -165 1207
rect -199 1105 -165 1139
rect -199 1037 -165 1071
rect -199 969 -165 1003
rect -199 901 -165 935
rect -199 833 -165 867
rect -199 765 -165 799
rect -199 697 -165 731
rect -199 629 -165 663
rect -199 561 -165 595
rect -199 493 -165 527
rect -199 425 -165 459
rect -199 357 -165 391
rect -199 289 -165 323
rect -199 221 -165 255
rect -199 153 -165 187
rect -199 85 -165 119
rect -199 17 -165 51
rect -199 -51 -165 -17
rect -199 -119 -165 -85
rect -199 -187 -165 -153
rect -199 -255 -165 -221
rect -199 -323 -165 -289
rect -199 -391 -165 -357
rect -199 -459 -165 -425
rect -199 -527 -165 -493
rect -199 -595 -165 -561
rect -199 -663 -165 -629
rect -199 -731 -165 -697
rect -199 -799 -165 -765
rect -199 -867 -165 -833
rect -199 -935 -165 -901
rect -199 -1003 -165 -969
rect -199 -1071 -165 -1037
rect -199 -1139 -165 -1105
rect -199 -1207 -165 -1173
rect -199 -1275 -165 -1241
rect -199 -1343 -165 -1309
rect -199 -1411 -165 -1377
rect -199 -1479 -165 -1445
rect -199 -1547 -165 -1513
rect -199 -1615 -165 -1581
rect -199 -1683 -165 -1649
rect -199 -1751 -165 -1717
rect -199 -1819 -165 -1785
rect -199 -1887 -165 -1853
rect -199 -1955 -165 -1921
rect -199 -2023 -165 -1989
rect -199 -2091 -165 -2057
rect -199 -2159 -165 -2125
rect -199 -2227 -165 -2193
rect -199 -2295 -165 -2261
rect -199 -2363 -165 -2329
rect 165 2329 199 2363
rect 165 2261 199 2295
rect 165 2193 199 2227
rect 165 2125 199 2159
rect 165 2057 199 2091
rect 165 1989 199 2023
rect 165 1921 199 1955
rect 165 1853 199 1887
rect 165 1785 199 1819
rect 165 1717 199 1751
rect 165 1649 199 1683
rect 165 1581 199 1615
rect 165 1513 199 1547
rect 165 1445 199 1479
rect 165 1377 199 1411
rect 165 1309 199 1343
rect 165 1241 199 1275
rect 165 1173 199 1207
rect 165 1105 199 1139
rect 165 1037 199 1071
rect 165 969 199 1003
rect 165 901 199 935
rect 165 833 199 867
rect 165 765 199 799
rect 165 697 199 731
rect 165 629 199 663
rect 165 561 199 595
rect 165 493 199 527
rect 165 425 199 459
rect 165 357 199 391
rect 165 289 199 323
rect 165 221 199 255
rect 165 153 199 187
rect 165 85 199 119
rect 165 17 199 51
rect 165 -51 199 -17
rect 165 -119 199 -85
rect 165 -187 199 -153
rect 165 -255 199 -221
rect 165 -323 199 -289
rect 165 -391 199 -357
rect 165 -459 199 -425
rect 165 -527 199 -493
rect 165 -595 199 -561
rect 165 -663 199 -629
rect 165 -731 199 -697
rect 165 -799 199 -765
rect 165 -867 199 -833
rect 165 -935 199 -901
rect 165 -1003 199 -969
rect 165 -1071 199 -1037
rect 165 -1139 199 -1105
rect 165 -1207 199 -1173
rect 165 -1275 199 -1241
rect 165 -1343 199 -1309
rect 165 -1411 199 -1377
rect 165 -1479 199 -1445
rect 165 -1547 199 -1513
rect 165 -1615 199 -1581
rect 165 -1683 199 -1649
rect 165 -1751 199 -1717
rect 165 -1819 199 -1785
rect 165 -1887 199 -1853
rect 165 -1955 199 -1921
rect 165 -2023 199 -1989
rect 165 -2091 199 -2057
rect 165 -2159 199 -2125
rect 165 -2227 199 -2193
rect 165 -2295 199 -2261
rect 165 -2363 199 -2329
rect -199 -2467 -165 -2397
rect 165 -2467 199 -2397
rect -199 -2501 -85 -2467
rect -51 -2501 -17 -2467
rect 17 -2501 51 -2467
rect 85 -2501 199 -2467
<< psubdiffcont >>
rect -85 2467 -51 2501
rect -17 2467 17 2501
rect 51 2467 85 2501
rect -199 2363 -165 2397
rect -199 2295 -165 2329
rect -199 2227 -165 2261
rect -199 2159 -165 2193
rect -199 2091 -165 2125
rect -199 2023 -165 2057
rect -199 1955 -165 1989
rect -199 1887 -165 1921
rect -199 1819 -165 1853
rect -199 1751 -165 1785
rect -199 1683 -165 1717
rect -199 1615 -165 1649
rect -199 1547 -165 1581
rect -199 1479 -165 1513
rect -199 1411 -165 1445
rect -199 1343 -165 1377
rect -199 1275 -165 1309
rect -199 1207 -165 1241
rect -199 1139 -165 1173
rect -199 1071 -165 1105
rect -199 1003 -165 1037
rect -199 935 -165 969
rect -199 867 -165 901
rect -199 799 -165 833
rect -199 731 -165 765
rect -199 663 -165 697
rect -199 595 -165 629
rect -199 527 -165 561
rect -199 459 -165 493
rect -199 391 -165 425
rect -199 323 -165 357
rect -199 255 -165 289
rect -199 187 -165 221
rect -199 119 -165 153
rect -199 51 -165 85
rect -199 -17 -165 17
rect -199 -85 -165 -51
rect -199 -153 -165 -119
rect -199 -221 -165 -187
rect -199 -289 -165 -255
rect -199 -357 -165 -323
rect -199 -425 -165 -391
rect -199 -493 -165 -459
rect -199 -561 -165 -527
rect -199 -629 -165 -595
rect -199 -697 -165 -663
rect -199 -765 -165 -731
rect -199 -833 -165 -799
rect -199 -901 -165 -867
rect -199 -969 -165 -935
rect -199 -1037 -165 -1003
rect -199 -1105 -165 -1071
rect -199 -1173 -165 -1139
rect -199 -1241 -165 -1207
rect -199 -1309 -165 -1275
rect -199 -1377 -165 -1343
rect -199 -1445 -165 -1411
rect -199 -1513 -165 -1479
rect -199 -1581 -165 -1547
rect -199 -1649 -165 -1615
rect -199 -1717 -165 -1683
rect -199 -1785 -165 -1751
rect -199 -1853 -165 -1819
rect -199 -1921 -165 -1887
rect -199 -1989 -165 -1955
rect -199 -2057 -165 -2023
rect -199 -2125 -165 -2091
rect -199 -2193 -165 -2159
rect -199 -2261 -165 -2227
rect -199 -2329 -165 -2295
rect -199 -2397 -165 -2363
rect 165 2363 199 2397
rect 165 2295 199 2329
rect 165 2227 199 2261
rect 165 2159 199 2193
rect 165 2091 199 2125
rect 165 2023 199 2057
rect 165 1955 199 1989
rect 165 1887 199 1921
rect 165 1819 199 1853
rect 165 1751 199 1785
rect 165 1683 199 1717
rect 165 1615 199 1649
rect 165 1547 199 1581
rect 165 1479 199 1513
rect 165 1411 199 1445
rect 165 1343 199 1377
rect 165 1275 199 1309
rect 165 1207 199 1241
rect 165 1139 199 1173
rect 165 1071 199 1105
rect 165 1003 199 1037
rect 165 935 199 969
rect 165 867 199 901
rect 165 799 199 833
rect 165 731 199 765
rect 165 663 199 697
rect 165 595 199 629
rect 165 527 199 561
rect 165 459 199 493
rect 165 391 199 425
rect 165 323 199 357
rect 165 255 199 289
rect 165 187 199 221
rect 165 119 199 153
rect 165 51 199 85
rect 165 -17 199 17
rect 165 -85 199 -51
rect 165 -153 199 -119
rect 165 -221 199 -187
rect 165 -289 199 -255
rect 165 -357 199 -323
rect 165 -425 199 -391
rect 165 -493 199 -459
rect 165 -561 199 -527
rect 165 -629 199 -595
rect 165 -697 199 -663
rect 165 -765 199 -731
rect 165 -833 199 -799
rect 165 -901 199 -867
rect 165 -969 199 -935
rect 165 -1037 199 -1003
rect 165 -1105 199 -1071
rect 165 -1173 199 -1139
rect 165 -1241 199 -1207
rect 165 -1309 199 -1275
rect 165 -1377 199 -1343
rect 165 -1445 199 -1411
rect 165 -1513 199 -1479
rect 165 -1581 199 -1547
rect 165 -1649 199 -1615
rect 165 -1717 199 -1683
rect 165 -1785 199 -1751
rect 165 -1853 199 -1819
rect 165 -1921 199 -1887
rect 165 -1989 199 -1955
rect 165 -2057 199 -2023
rect 165 -2125 199 -2091
rect 165 -2193 199 -2159
rect 165 -2261 199 -2227
rect 165 -2329 199 -2295
rect 165 -2397 199 -2363
rect -85 -2501 -51 -2467
rect -17 -2501 17 -2467
rect 51 -2501 85 -2467
<< xpolycontact >>
rect -69 1939 69 2371
rect -69 -2371 69 -1939
<< ppolyres >>
rect -69 -1939 69 1939
<< locali >>
rect -199 2467 -85 2501
rect -51 2467 -17 2501
rect 17 2467 51 2501
rect 85 2467 199 2501
rect -199 2397 -165 2467
rect 165 2397 199 2467
rect -199 2329 -165 2363
rect -199 2261 -165 2295
rect -199 2193 -165 2227
rect -199 2125 -165 2159
rect -199 2057 -165 2091
rect -199 1989 -165 2023
rect -199 1921 -165 1955
rect 165 2329 199 2363
rect 165 2261 199 2295
rect 165 2193 199 2227
rect 165 2125 199 2159
rect 165 2057 199 2091
rect 165 1989 199 2023
rect -199 1853 -165 1887
rect -199 1785 -165 1819
rect -199 1717 -165 1751
rect -199 1649 -165 1683
rect -199 1581 -165 1615
rect -199 1513 -165 1547
rect -199 1445 -165 1479
rect -199 1377 -165 1411
rect -199 1309 -165 1343
rect -199 1241 -165 1275
rect -199 1173 -165 1207
rect -199 1105 -165 1139
rect -199 1037 -165 1071
rect -199 969 -165 1003
rect -199 901 -165 935
rect -199 833 -165 867
rect -199 765 -165 799
rect -199 697 -165 731
rect -199 629 -165 663
rect -199 561 -165 595
rect -199 493 -165 527
rect -199 425 -165 459
rect -199 357 -165 391
rect -199 289 -165 323
rect -199 221 -165 255
rect -199 153 -165 187
rect -199 85 -165 119
rect -199 17 -165 51
rect -199 -51 -165 -17
rect -199 -119 -165 -85
rect -199 -187 -165 -153
rect -199 -255 -165 -221
rect -199 -323 -165 -289
rect -199 -391 -165 -357
rect -199 -459 -165 -425
rect -199 -527 -165 -493
rect -199 -595 -165 -561
rect -199 -663 -165 -629
rect -199 -731 -165 -697
rect -199 -799 -165 -765
rect -199 -867 -165 -833
rect -199 -935 -165 -901
rect -199 -1003 -165 -969
rect -199 -1071 -165 -1037
rect -199 -1139 -165 -1105
rect -199 -1207 -165 -1173
rect -199 -1275 -165 -1241
rect -199 -1343 -165 -1309
rect -199 -1411 -165 -1377
rect -199 -1479 -165 -1445
rect -199 -1547 -165 -1513
rect -199 -1615 -165 -1581
rect -199 -1683 -165 -1649
rect -199 -1751 -165 -1717
rect -199 -1819 -165 -1785
rect -199 -1887 -165 -1853
rect -199 -1955 -165 -1921
rect 165 1921 199 1955
rect 165 1853 199 1887
rect 165 1785 199 1819
rect 165 1717 199 1751
rect 165 1649 199 1683
rect 165 1581 199 1615
rect 165 1513 199 1547
rect 165 1445 199 1479
rect 165 1377 199 1411
rect 165 1309 199 1343
rect 165 1241 199 1275
rect 165 1173 199 1207
rect 165 1105 199 1139
rect 165 1037 199 1071
rect 165 969 199 1003
rect 165 901 199 935
rect 165 833 199 867
rect 165 765 199 799
rect 165 697 199 731
rect 165 629 199 663
rect 165 561 199 595
rect 165 493 199 527
rect 165 425 199 459
rect 165 357 199 391
rect 165 289 199 323
rect 165 221 199 255
rect 165 153 199 187
rect 165 85 199 119
rect 165 17 199 51
rect 165 -51 199 -17
rect 165 -119 199 -85
rect 165 -187 199 -153
rect 165 -255 199 -221
rect 165 -323 199 -289
rect 165 -391 199 -357
rect 165 -459 199 -425
rect 165 -527 199 -493
rect 165 -595 199 -561
rect 165 -663 199 -629
rect 165 -731 199 -697
rect 165 -799 199 -765
rect 165 -867 199 -833
rect 165 -935 199 -901
rect 165 -1003 199 -969
rect 165 -1071 199 -1037
rect 165 -1139 199 -1105
rect 165 -1207 199 -1173
rect 165 -1275 199 -1241
rect 165 -1343 199 -1309
rect 165 -1411 199 -1377
rect 165 -1479 199 -1445
rect 165 -1547 199 -1513
rect 165 -1615 199 -1581
rect 165 -1683 199 -1649
rect 165 -1751 199 -1717
rect 165 -1819 199 -1785
rect 165 -1887 199 -1853
rect -199 -2023 -165 -1989
rect -199 -2091 -165 -2057
rect -199 -2159 -165 -2125
rect -199 -2227 -165 -2193
rect -199 -2295 -165 -2261
rect -199 -2363 -165 -2329
rect 165 -1955 199 -1921
rect 165 -2023 199 -1989
rect 165 -2091 199 -2057
rect 165 -2159 199 -2125
rect 165 -2227 199 -2193
rect 165 -2295 199 -2261
rect 165 -2363 199 -2329
rect -199 -2467 -165 -2397
rect 165 -2467 199 -2397
rect -199 -2501 -85 -2467
rect -51 -2501 -17 -2467
rect 17 -2501 51 -2467
rect 85 -2501 199 -2467
<< viali >>
rect -53 1957 53 2351
rect -53 -2352 53 -1958
<< metal1 >>
rect -59 2351 59 2365
rect -59 1957 -53 2351
rect 53 1957 59 2351
rect -59 1944 59 1957
rect -59 -1958 59 -1944
rect -59 -2352 -53 -1958
rect 53 -2352 59 -1958
rect -59 -2365 59 -2352
<< properties >>
string FIXED_BBOX -182 -2484 182 2484
string GDS_END 12450
string GDS_FILE /home/anton/projects/tt06-grab-bag/gds/tt_um_algofoogle_tt06_grab_bag.gds
string GDS_START 158
<< end >>
