magic
tech sky130A
magscale 1 2
timestamp 1713537803
<< pwell >>
rect -225 4476 225 4562
rect -225 -4476 -139 4476
rect 139 -4476 225 4476
rect -225 -4562 225 -4476
<< psubdiff >>
rect -199 4502 -85 4536
rect -51 4502 -17 4536
rect 17 4502 51 4536
rect 85 4502 199 4536
rect -199 4437 -165 4502
rect 165 4437 199 4502
rect -199 4369 -165 4403
rect -199 4301 -165 4335
rect -199 4233 -165 4267
rect -199 4165 -165 4199
rect -199 4097 -165 4131
rect -199 4029 -165 4063
rect -199 3961 -165 3995
rect -199 3893 -165 3927
rect -199 3825 -165 3859
rect -199 3757 -165 3791
rect -199 3689 -165 3723
rect -199 3621 -165 3655
rect -199 3553 -165 3587
rect -199 3485 -165 3519
rect -199 3417 -165 3451
rect -199 3349 -165 3383
rect -199 3281 -165 3315
rect -199 3213 -165 3247
rect -199 3145 -165 3179
rect -199 3077 -165 3111
rect -199 3009 -165 3043
rect -199 2941 -165 2975
rect -199 2873 -165 2907
rect -199 2805 -165 2839
rect -199 2737 -165 2771
rect -199 2669 -165 2703
rect -199 2601 -165 2635
rect -199 2533 -165 2567
rect -199 2465 -165 2499
rect -199 2397 -165 2431
rect -199 2329 -165 2363
rect -199 2261 -165 2295
rect -199 2193 -165 2227
rect -199 2125 -165 2159
rect -199 2057 -165 2091
rect -199 1989 -165 2023
rect -199 1921 -165 1955
rect -199 1853 -165 1887
rect -199 1785 -165 1819
rect -199 1717 -165 1751
rect -199 1649 -165 1683
rect -199 1581 -165 1615
rect -199 1513 -165 1547
rect -199 1445 -165 1479
rect -199 1377 -165 1411
rect -199 1309 -165 1343
rect -199 1241 -165 1275
rect -199 1173 -165 1207
rect -199 1105 -165 1139
rect -199 1037 -165 1071
rect -199 969 -165 1003
rect -199 901 -165 935
rect -199 833 -165 867
rect -199 765 -165 799
rect -199 697 -165 731
rect -199 629 -165 663
rect -199 561 -165 595
rect -199 493 -165 527
rect -199 425 -165 459
rect -199 357 -165 391
rect -199 289 -165 323
rect -199 221 -165 255
rect -199 153 -165 187
rect -199 85 -165 119
rect -199 17 -165 51
rect -199 -51 -165 -17
rect -199 -119 -165 -85
rect -199 -187 -165 -153
rect -199 -255 -165 -221
rect -199 -323 -165 -289
rect -199 -391 -165 -357
rect -199 -459 -165 -425
rect -199 -527 -165 -493
rect -199 -595 -165 -561
rect -199 -663 -165 -629
rect -199 -731 -165 -697
rect -199 -799 -165 -765
rect -199 -867 -165 -833
rect -199 -935 -165 -901
rect -199 -1003 -165 -969
rect -199 -1071 -165 -1037
rect -199 -1139 -165 -1105
rect -199 -1207 -165 -1173
rect -199 -1275 -165 -1241
rect -199 -1343 -165 -1309
rect -199 -1411 -165 -1377
rect -199 -1479 -165 -1445
rect -199 -1547 -165 -1513
rect -199 -1615 -165 -1581
rect -199 -1683 -165 -1649
rect -199 -1751 -165 -1717
rect -199 -1819 -165 -1785
rect -199 -1887 -165 -1853
rect -199 -1955 -165 -1921
rect -199 -2023 -165 -1989
rect -199 -2091 -165 -2057
rect -199 -2159 -165 -2125
rect -199 -2227 -165 -2193
rect -199 -2295 -165 -2261
rect -199 -2363 -165 -2329
rect -199 -2431 -165 -2397
rect -199 -2499 -165 -2465
rect -199 -2567 -165 -2533
rect -199 -2635 -165 -2601
rect -199 -2703 -165 -2669
rect -199 -2771 -165 -2737
rect -199 -2839 -165 -2805
rect -199 -2907 -165 -2873
rect -199 -2975 -165 -2941
rect -199 -3043 -165 -3009
rect -199 -3111 -165 -3077
rect -199 -3179 -165 -3145
rect -199 -3247 -165 -3213
rect -199 -3315 -165 -3281
rect -199 -3383 -165 -3349
rect -199 -3451 -165 -3417
rect -199 -3519 -165 -3485
rect -199 -3587 -165 -3553
rect -199 -3655 -165 -3621
rect -199 -3723 -165 -3689
rect -199 -3791 -165 -3757
rect -199 -3859 -165 -3825
rect -199 -3927 -165 -3893
rect -199 -3995 -165 -3961
rect -199 -4063 -165 -4029
rect -199 -4131 -165 -4097
rect -199 -4199 -165 -4165
rect -199 -4267 -165 -4233
rect -199 -4335 -165 -4301
rect -199 -4403 -165 -4369
rect 165 4369 199 4403
rect 165 4301 199 4335
rect 165 4233 199 4267
rect 165 4165 199 4199
rect 165 4097 199 4131
rect 165 4029 199 4063
rect 165 3961 199 3995
rect 165 3893 199 3927
rect 165 3825 199 3859
rect 165 3757 199 3791
rect 165 3689 199 3723
rect 165 3621 199 3655
rect 165 3553 199 3587
rect 165 3485 199 3519
rect 165 3417 199 3451
rect 165 3349 199 3383
rect 165 3281 199 3315
rect 165 3213 199 3247
rect 165 3145 199 3179
rect 165 3077 199 3111
rect 165 3009 199 3043
rect 165 2941 199 2975
rect 165 2873 199 2907
rect 165 2805 199 2839
rect 165 2737 199 2771
rect 165 2669 199 2703
rect 165 2601 199 2635
rect 165 2533 199 2567
rect 165 2465 199 2499
rect 165 2397 199 2431
rect 165 2329 199 2363
rect 165 2261 199 2295
rect 165 2193 199 2227
rect 165 2125 199 2159
rect 165 2057 199 2091
rect 165 1989 199 2023
rect 165 1921 199 1955
rect 165 1853 199 1887
rect 165 1785 199 1819
rect 165 1717 199 1751
rect 165 1649 199 1683
rect 165 1581 199 1615
rect 165 1513 199 1547
rect 165 1445 199 1479
rect 165 1377 199 1411
rect 165 1309 199 1343
rect 165 1241 199 1275
rect 165 1173 199 1207
rect 165 1105 199 1139
rect 165 1037 199 1071
rect 165 969 199 1003
rect 165 901 199 935
rect 165 833 199 867
rect 165 765 199 799
rect 165 697 199 731
rect 165 629 199 663
rect 165 561 199 595
rect 165 493 199 527
rect 165 425 199 459
rect 165 357 199 391
rect 165 289 199 323
rect 165 221 199 255
rect 165 153 199 187
rect 165 85 199 119
rect 165 17 199 51
rect 165 -51 199 -17
rect 165 -119 199 -85
rect 165 -187 199 -153
rect 165 -255 199 -221
rect 165 -323 199 -289
rect 165 -391 199 -357
rect 165 -459 199 -425
rect 165 -527 199 -493
rect 165 -595 199 -561
rect 165 -663 199 -629
rect 165 -731 199 -697
rect 165 -799 199 -765
rect 165 -867 199 -833
rect 165 -935 199 -901
rect 165 -1003 199 -969
rect 165 -1071 199 -1037
rect 165 -1139 199 -1105
rect 165 -1207 199 -1173
rect 165 -1275 199 -1241
rect 165 -1343 199 -1309
rect 165 -1411 199 -1377
rect 165 -1479 199 -1445
rect 165 -1547 199 -1513
rect 165 -1615 199 -1581
rect 165 -1683 199 -1649
rect 165 -1751 199 -1717
rect 165 -1819 199 -1785
rect 165 -1887 199 -1853
rect 165 -1955 199 -1921
rect 165 -2023 199 -1989
rect 165 -2091 199 -2057
rect 165 -2159 199 -2125
rect 165 -2227 199 -2193
rect 165 -2295 199 -2261
rect 165 -2363 199 -2329
rect 165 -2431 199 -2397
rect 165 -2499 199 -2465
rect 165 -2567 199 -2533
rect 165 -2635 199 -2601
rect 165 -2703 199 -2669
rect 165 -2771 199 -2737
rect 165 -2839 199 -2805
rect 165 -2907 199 -2873
rect 165 -2975 199 -2941
rect 165 -3043 199 -3009
rect 165 -3111 199 -3077
rect 165 -3179 199 -3145
rect 165 -3247 199 -3213
rect 165 -3315 199 -3281
rect 165 -3383 199 -3349
rect 165 -3451 199 -3417
rect 165 -3519 199 -3485
rect 165 -3587 199 -3553
rect 165 -3655 199 -3621
rect 165 -3723 199 -3689
rect 165 -3791 199 -3757
rect 165 -3859 199 -3825
rect 165 -3927 199 -3893
rect 165 -3995 199 -3961
rect 165 -4063 199 -4029
rect 165 -4131 199 -4097
rect 165 -4199 199 -4165
rect 165 -4267 199 -4233
rect 165 -4335 199 -4301
rect 165 -4403 199 -4369
rect -199 -4502 -165 -4437
rect 165 -4502 199 -4437
rect -199 -4536 -85 -4502
rect -51 -4536 -17 -4502
rect 17 -4536 51 -4502
rect 85 -4536 199 -4502
<< psubdiffcont >>
rect -85 4502 -51 4536
rect -17 4502 17 4536
rect 51 4502 85 4536
rect -199 4403 -165 4437
rect -199 4335 -165 4369
rect -199 4267 -165 4301
rect -199 4199 -165 4233
rect -199 4131 -165 4165
rect -199 4063 -165 4097
rect -199 3995 -165 4029
rect -199 3927 -165 3961
rect -199 3859 -165 3893
rect -199 3791 -165 3825
rect -199 3723 -165 3757
rect -199 3655 -165 3689
rect -199 3587 -165 3621
rect -199 3519 -165 3553
rect -199 3451 -165 3485
rect -199 3383 -165 3417
rect -199 3315 -165 3349
rect -199 3247 -165 3281
rect -199 3179 -165 3213
rect -199 3111 -165 3145
rect -199 3043 -165 3077
rect -199 2975 -165 3009
rect -199 2907 -165 2941
rect -199 2839 -165 2873
rect -199 2771 -165 2805
rect -199 2703 -165 2737
rect -199 2635 -165 2669
rect -199 2567 -165 2601
rect -199 2499 -165 2533
rect -199 2431 -165 2465
rect -199 2363 -165 2397
rect -199 2295 -165 2329
rect -199 2227 -165 2261
rect -199 2159 -165 2193
rect -199 2091 -165 2125
rect -199 2023 -165 2057
rect -199 1955 -165 1989
rect -199 1887 -165 1921
rect -199 1819 -165 1853
rect -199 1751 -165 1785
rect -199 1683 -165 1717
rect -199 1615 -165 1649
rect -199 1547 -165 1581
rect -199 1479 -165 1513
rect -199 1411 -165 1445
rect -199 1343 -165 1377
rect -199 1275 -165 1309
rect -199 1207 -165 1241
rect -199 1139 -165 1173
rect -199 1071 -165 1105
rect -199 1003 -165 1037
rect -199 935 -165 969
rect -199 867 -165 901
rect -199 799 -165 833
rect -199 731 -165 765
rect -199 663 -165 697
rect -199 595 -165 629
rect -199 527 -165 561
rect -199 459 -165 493
rect -199 391 -165 425
rect -199 323 -165 357
rect -199 255 -165 289
rect -199 187 -165 221
rect -199 119 -165 153
rect -199 51 -165 85
rect -199 -17 -165 17
rect -199 -85 -165 -51
rect -199 -153 -165 -119
rect -199 -221 -165 -187
rect -199 -289 -165 -255
rect -199 -357 -165 -323
rect -199 -425 -165 -391
rect -199 -493 -165 -459
rect -199 -561 -165 -527
rect -199 -629 -165 -595
rect -199 -697 -165 -663
rect -199 -765 -165 -731
rect -199 -833 -165 -799
rect -199 -901 -165 -867
rect -199 -969 -165 -935
rect -199 -1037 -165 -1003
rect -199 -1105 -165 -1071
rect -199 -1173 -165 -1139
rect -199 -1241 -165 -1207
rect -199 -1309 -165 -1275
rect -199 -1377 -165 -1343
rect -199 -1445 -165 -1411
rect -199 -1513 -165 -1479
rect -199 -1581 -165 -1547
rect -199 -1649 -165 -1615
rect -199 -1717 -165 -1683
rect -199 -1785 -165 -1751
rect -199 -1853 -165 -1819
rect -199 -1921 -165 -1887
rect -199 -1989 -165 -1955
rect -199 -2057 -165 -2023
rect -199 -2125 -165 -2091
rect -199 -2193 -165 -2159
rect -199 -2261 -165 -2227
rect -199 -2329 -165 -2295
rect -199 -2397 -165 -2363
rect -199 -2465 -165 -2431
rect -199 -2533 -165 -2499
rect -199 -2601 -165 -2567
rect -199 -2669 -165 -2635
rect -199 -2737 -165 -2703
rect -199 -2805 -165 -2771
rect -199 -2873 -165 -2839
rect -199 -2941 -165 -2907
rect -199 -3009 -165 -2975
rect -199 -3077 -165 -3043
rect -199 -3145 -165 -3111
rect -199 -3213 -165 -3179
rect -199 -3281 -165 -3247
rect -199 -3349 -165 -3315
rect -199 -3417 -165 -3383
rect -199 -3485 -165 -3451
rect -199 -3553 -165 -3519
rect -199 -3621 -165 -3587
rect -199 -3689 -165 -3655
rect -199 -3757 -165 -3723
rect -199 -3825 -165 -3791
rect -199 -3893 -165 -3859
rect -199 -3961 -165 -3927
rect -199 -4029 -165 -3995
rect -199 -4097 -165 -4063
rect -199 -4165 -165 -4131
rect -199 -4233 -165 -4199
rect -199 -4301 -165 -4267
rect -199 -4369 -165 -4335
rect -199 -4437 -165 -4403
rect 165 4403 199 4437
rect 165 4335 199 4369
rect 165 4267 199 4301
rect 165 4199 199 4233
rect 165 4131 199 4165
rect 165 4063 199 4097
rect 165 3995 199 4029
rect 165 3927 199 3961
rect 165 3859 199 3893
rect 165 3791 199 3825
rect 165 3723 199 3757
rect 165 3655 199 3689
rect 165 3587 199 3621
rect 165 3519 199 3553
rect 165 3451 199 3485
rect 165 3383 199 3417
rect 165 3315 199 3349
rect 165 3247 199 3281
rect 165 3179 199 3213
rect 165 3111 199 3145
rect 165 3043 199 3077
rect 165 2975 199 3009
rect 165 2907 199 2941
rect 165 2839 199 2873
rect 165 2771 199 2805
rect 165 2703 199 2737
rect 165 2635 199 2669
rect 165 2567 199 2601
rect 165 2499 199 2533
rect 165 2431 199 2465
rect 165 2363 199 2397
rect 165 2295 199 2329
rect 165 2227 199 2261
rect 165 2159 199 2193
rect 165 2091 199 2125
rect 165 2023 199 2057
rect 165 1955 199 1989
rect 165 1887 199 1921
rect 165 1819 199 1853
rect 165 1751 199 1785
rect 165 1683 199 1717
rect 165 1615 199 1649
rect 165 1547 199 1581
rect 165 1479 199 1513
rect 165 1411 199 1445
rect 165 1343 199 1377
rect 165 1275 199 1309
rect 165 1207 199 1241
rect 165 1139 199 1173
rect 165 1071 199 1105
rect 165 1003 199 1037
rect 165 935 199 969
rect 165 867 199 901
rect 165 799 199 833
rect 165 731 199 765
rect 165 663 199 697
rect 165 595 199 629
rect 165 527 199 561
rect 165 459 199 493
rect 165 391 199 425
rect 165 323 199 357
rect 165 255 199 289
rect 165 187 199 221
rect 165 119 199 153
rect 165 51 199 85
rect 165 -17 199 17
rect 165 -85 199 -51
rect 165 -153 199 -119
rect 165 -221 199 -187
rect 165 -289 199 -255
rect 165 -357 199 -323
rect 165 -425 199 -391
rect 165 -493 199 -459
rect 165 -561 199 -527
rect 165 -629 199 -595
rect 165 -697 199 -663
rect 165 -765 199 -731
rect 165 -833 199 -799
rect 165 -901 199 -867
rect 165 -969 199 -935
rect 165 -1037 199 -1003
rect 165 -1105 199 -1071
rect 165 -1173 199 -1139
rect 165 -1241 199 -1207
rect 165 -1309 199 -1275
rect 165 -1377 199 -1343
rect 165 -1445 199 -1411
rect 165 -1513 199 -1479
rect 165 -1581 199 -1547
rect 165 -1649 199 -1615
rect 165 -1717 199 -1683
rect 165 -1785 199 -1751
rect 165 -1853 199 -1819
rect 165 -1921 199 -1887
rect 165 -1989 199 -1955
rect 165 -2057 199 -2023
rect 165 -2125 199 -2091
rect 165 -2193 199 -2159
rect 165 -2261 199 -2227
rect 165 -2329 199 -2295
rect 165 -2397 199 -2363
rect 165 -2465 199 -2431
rect 165 -2533 199 -2499
rect 165 -2601 199 -2567
rect 165 -2669 199 -2635
rect 165 -2737 199 -2703
rect 165 -2805 199 -2771
rect 165 -2873 199 -2839
rect 165 -2941 199 -2907
rect 165 -3009 199 -2975
rect 165 -3077 199 -3043
rect 165 -3145 199 -3111
rect 165 -3213 199 -3179
rect 165 -3281 199 -3247
rect 165 -3349 199 -3315
rect 165 -3417 199 -3383
rect 165 -3485 199 -3451
rect 165 -3553 199 -3519
rect 165 -3621 199 -3587
rect 165 -3689 199 -3655
rect 165 -3757 199 -3723
rect 165 -3825 199 -3791
rect 165 -3893 199 -3859
rect 165 -3961 199 -3927
rect 165 -4029 199 -3995
rect 165 -4097 199 -4063
rect 165 -4165 199 -4131
rect 165 -4233 199 -4199
rect 165 -4301 199 -4267
rect 165 -4369 199 -4335
rect 165 -4437 199 -4403
rect -85 -4536 -51 -4502
rect -17 -4536 17 -4502
rect 51 -4536 85 -4502
<< xpolycontact >>
rect -69 3974 69 4406
rect -69 -4406 69 -3974
<< ppolyres >>
rect -69 -3974 69 3974
<< locali >>
rect -199 4502 -85 4536
rect -51 4502 -17 4536
rect 17 4502 51 4536
rect 85 4502 199 4536
rect -199 4437 -165 4502
rect 165 4437 199 4502
rect -199 4369 -165 4403
rect -199 4301 -165 4335
rect -199 4233 -165 4267
rect -199 4165 -165 4199
rect -199 4097 -165 4131
rect -199 4029 -165 4063
rect -199 3961 -165 3995
rect 165 4369 199 4403
rect 165 4301 199 4335
rect 165 4233 199 4267
rect 165 4165 199 4199
rect 165 4097 199 4131
rect 165 4029 199 4063
rect -199 3893 -165 3927
rect -199 3825 -165 3859
rect -199 3757 -165 3791
rect -199 3689 -165 3723
rect -199 3621 -165 3655
rect -199 3553 -165 3587
rect -199 3485 -165 3519
rect -199 3417 -165 3451
rect -199 3349 -165 3383
rect -199 3281 -165 3315
rect -199 3213 -165 3247
rect -199 3145 -165 3179
rect -199 3077 -165 3111
rect -199 3009 -165 3043
rect -199 2941 -165 2975
rect -199 2873 -165 2907
rect -199 2805 -165 2839
rect -199 2737 -165 2771
rect -199 2669 -165 2703
rect -199 2601 -165 2635
rect -199 2533 -165 2567
rect -199 2465 -165 2499
rect -199 2397 -165 2431
rect -199 2329 -165 2363
rect -199 2261 -165 2295
rect -199 2193 -165 2227
rect -199 2125 -165 2159
rect -199 2057 -165 2091
rect -199 1989 -165 2023
rect -199 1921 -165 1955
rect -199 1853 -165 1887
rect -199 1785 -165 1819
rect -199 1717 -165 1751
rect -199 1649 -165 1683
rect -199 1581 -165 1615
rect -199 1513 -165 1547
rect -199 1445 -165 1479
rect -199 1377 -165 1411
rect -199 1309 -165 1343
rect -199 1241 -165 1275
rect -199 1173 -165 1207
rect -199 1105 -165 1139
rect -199 1037 -165 1071
rect -199 969 -165 1003
rect -199 901 -165 935
rect -199 833 -165 867
rect -199 765 -165 799
rect -199 697 -165 731
rect -199 629 -165 663
rect -199 561 -165 595
rect -199 493 -165 527
rect -199 425 -165 459
rect -199 357 -165 391
rect -199 289 -165 323
rect -199 221 -165 255
rect -199 153 -165 187
rect -199 85 -165 119
rect -199 17 -165 51
rect -199 -51 -165 -17
rect -199 -119 -165 -85
rect -199 -187 -165 -153
rect -199 -255 -165 -221
rect -199 -323 -165 -289
rect -199 -391 -165 -357
rect -199 -459 -165 -425
rect -199 -527 -165 -493
rect -199 -595 -165 -561
rect -199 -663 -165 -629
rect -199 -731 -165 -697
rect -199 -799 -165 -765
rect -199 -867 -165 -833
rect -199 -935 -165 -901
rect -199 -1003 -165 -969
rect -199 -1071 -165 -1037
rect -199 -1139 -165 -1105
rect -199 -1207 -165 -1173
rect -199 -1275 -165 -1241
rect -199 -1343 -165 -1309
rect -199 -1411 -165 -1377
rect -199 -1479 -165 -1445
rect -199 -1547 -165 -1513
rect -199 -1615 -165 -1581
rect -199 -1683 -165 -1649
rect -199 -1751 -165 -1717
rect -199 -1819 -165 -1785
rect -199 -1887 -165 -1853
rect -199 -1955 -165 -1921
rect -199 -2023 -165 -1989
rect -199 -2091 -165 -2057
rect -199 -2159 -165 -2125
rect -199 -2227 -165 -2193
rect -199 -2295 -165 -2261
rect -199 -2363 -165 -2329
rect -199 -2431 -165 -2397
rect -199 -2499 -165 -2465
rect -199 -2567 -165 -2533
rect -199 -2635 -165 -2601
rect -199 -2703 -165 -2669
rect -199 -2771 -165 -2737
rect -199 -2839 -165 -2805
rect -199 -2907 -165 -2873
rect -199 -2975 -165 -2941
rect -199 -3043 -165 -3009
rect -199 -3111 -165 -3077
rect -199 -3179 -165 -3145
rect -199 -3247 -165 -3213
rect -199 -3315 -165 -3281
rect -199 -3383 -165 -3349
rect -199 -3451 -165 -3417
rect -199 -3519 -165 -3485
rect -199 -3587 -165 -3553
rect -199 -3655 -165 -3621
rect -199 -3723 -165 -3689
rect -199 -3791 -165 -3757
rect -199 -3859 -165 -3825
rect -199 -3927 -165 -3893
rect -199 -3995 -165 -3961
rect 165 3961 199 3995
rect 165 3893 199 3927
rect 165 3825 199 3859
rect 165 3757 199 3791
rect 165 3689 199 3723
rect 165 3621 199 3655
rect 165 3553 199 3587
rect 165 3485 199 3519
rect 165 3417 199 3451
rect 165 3349 199 3383
rect 165 3281 199 3315
rect 165 3213 199 3247
rect 165 3145 199 3179
rect 165 3077 199 3111
rect 165 3009 199 3043
rect 165 2941 199 2975
rect 165 2873 199 2907
rect 165 2805 199 2839
rect 165 2737 199 2771
rect 165 2669 199 2703
rect 165 2601 199 2635
rect 165 2533 199 2567
rect 165 2465 199 2499
rect 165 2397 199 2431
rect 165 2329 199 2363
rect 165 2261 199 2295
rect 165 2193 199 2227
rect 165 2125 199 2159
rect 165 2057 199 2091
rect 165 1989 199 2023
rect 165 1921 199 1955
rect 165 1853 199 1887
rect 165 1785 199 1819
rect 165 1717 199 1751
rect 165 1649 199 1683
rect 165 1581 199 1615
rect 165 1513 199 1547
rect 165 1445 199 1479
rect 165 1377 199 1411
rect 165 1309 199 1343
rect 165 1241 199 1275
rect 165 1173 199 1207
rect 165 1105 199 1139
rect 165 1037 199 1071
rect 165 969 199 1003
rect 165 901 199 935
rect 165 833 199 867
rect 165 765 199 799
rect 165 697 199 731
rect 165 629 199 663
rect 165 561 199 595
rect 165 493 199 527
rect 165 425 199 459
rect 165 357 199 391
rect 165 289 199 323
rect 165 221 199 255
rect 165 153 199 187
rect 165 85 199 119
rect 165 17 199 51
rect 165 -51 199 -17
rect 165 -119 199 -85
rect 165 -187 199 -153
rect 165 -255 199 -221
rect 165 -323 199 -289
rect 165 -391 199 -357
rect 165 -459 199 -425
rect 165 -527 199 -493
rect 165 -595 199 -561
rect 165 -663 199 -629
rect 165 -731 199 -697
rect 165 -799 199 -765
rect 165 -867 199 -833
rect 165 -935 199 -901
rect 165 -1003 199 -969
rect 165 -1071 199 -1037
rect 165 -1139 199 -1105
rect 165 -1207 199 -1173
rect 165 -1275 199 -1241
rect 165 -1343 199 -1309
rect 165 -1411 199 -1377
rect 165 -1479 199 -1445
rect 165 -1547 199 -1513
rect 165 -1615 199 -1581
rect 165 -1683 199 -1649
rect 165 -1751 199 -1717
rect 165 -1819 199 -1785
rect 165 -1887 199 -1853
rect 165 -1955 199 -1921
rect 165 -2023 199 -1989
rect 165 -2091 199 -2057
rect 165 -2159 199 -2125
rect 165 -2227 199 -2193
rect 165 -2295 199 -2261
rect 165 -2363 199 -2329
rect 165 -2431 199 -2397
rect 165 -2499 199 -2465
rect 165 -2567 199 -2533
rect 165 -2635 199 -2601
rect 165 -2703 199 -2669
rect 165 -2771 199 -2737
rect 165 -2839 199 -2805
rect 165 -2907 199 -2873
rect 165 -2975 199 -2941
rect 165 -3043 199 -3009
rect 165 -3111 199 -3077
rect 165 -3179 199 -3145
rect 165 -3247 199 -3213
rect 165 -3315 199 -3281
rect 165 -3383 199 -3349
rect 165 -3451 199 -3417
rect 165 -3519 199 -3485
rect 165 -3587 199 -3553
rect 165 -3655 199 -3621
rect 165 -3723 199 -3689
rect 165 -3791 199 -3757
rect 165 -3859 199 -3825
rect 165 -3927 199 -3893
rect -199 -4063 -165 -4029
rect -199 -4131 -165 -4097
rect -199 -4199 -165 -4165
rect -199 -4267 -165 -4233
rect -199 -4335 -165 -4301
rect -199 -4403 -165 -4369
rect 165 -3995 199 -3961
rect 165 -4063 199 -4029
rect 165 -4131 199 -4097
rect 165 -4199 199 -4165
rect 165 -4267 199 -4233
rect 165 -4335 199 -4301
rect 165 -4403 199 -4369
rect -199 -4502 -165 -4437
rect 165 -4502 199 -4437
rect -199 -4536 -85 -4502
rect -51 -4536 -17 -4502
rect 17 -4536 51 -4502
rect 85 -4536 199 -4502
<< viali >>
rect -53 3992 53 4386
rect -53 -4387 53 -3993
<< metal1 >>
rect -59 4386 59 4400
rect -59 3992 -53 4386
rect 53 3992 59 4386
rect -59 3979 59 3992
rect -59 -3993 59 -3979
rect -59 -4387 -53 -3993
rect 53 -4387 59 -3993
rect -59 -4400 59 -4387
<< properties >>
string FIXED_BBOX -182 -4519 182 4519
string GDS_END 32492
string GDS_FILE /home/anton/projects/tt06-grab-bag/gds/tt_um_algofoogle_tt06_grab_bag.gds
string GDS_START 12520
<< end >>
