Cosimulation of my VGA digital test block with 3 R2R DACs, using Verilator and d_cosim in ngspice-42

*.lib /home/matt/work/asic-workshop/shuttle-2404/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.lib /home/anton/.volare/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* https://sourceforge.net/p/ngspice/ngspice/ci/master/tree/examples/xspice/verilator/

* The digital portion of the circuit is specified in compiled Verilog.
* list the inputs and outputs.
* NOTE: We name bus signals individually, in the order they're defined in the Verilog:
adut 
+ [ clk rst_n in7 in6 in5 in4 in3 in2 in1 in0 ]
+ [
+ hsync vsync hblank vblank
+ r7 r6 r5 r4 r3 r2 r1 r0
+ g7 g6 g5 g4 g3 g2 g1 g0
+ b7 b6 b5 b4 b3 b2 b1 b0
+ dr7 dg7 db7
+ dr6 dg6 db6
+] null dut
.model dut d_cosim simulation="./spicewrap.so"
* Debug outputs:
*+ m7 m6 m5 m4 m3 m2 m1 m0
*+ o_reset o_visible
*+ c7 c6 c5 c4 c3 c2 c1 c0
*+ o_clk
*+ x7 x6 x5 x4 x3 x2 x1 x0
*+ o_clk2 o_zero o_one


* connect the driver to the R2R dac
* had to edit spice exported by xschem to add the subckt and ends

.include "../xschem/simulation/r2r.spice" 
.include "../xschem/simulation/dacboost.spice" 
*.include "../mag/r2r.spice" 

xr2r_R rdac r7 r6 r5 r4 r3 r2 r1 r0 GND GND r2r
xr2r_G gdac g7 g6 g5 g4 g3 g2 g1 g0 GND GND r2r
xr2r_B bdac b7 b6 b5 b4 b3 b2 b1 b0 GND GND r2r

xr2r_Rhz rdachz r7 r6 r5 r4 r3 r2 r1 r0 GND GND r2r
xr2r_Ghz gdachz g7 g6 g5 g4 g3 g2 g1 g0 GND GND r2r
xr2r_Bhz bdachz b7 b6 b5 b4 b3 b2 b1 b0 GND GND r2r

xr2r_Rhhz rdachhz r7 r6 r5 r4 r3 r2 r1 r0 GND GND r2r
xr2r_Ghhz gdachhz g7 g6 g5 g4 g3 g2 g1 g0 GND GND r2r
xr2r_Bhhz bdachhz b7 b6 b5 b4 b3 b2 b1 b0 GND GND r2r

xr2r_Rxhz rdacxhz r7 r6 r5 r4 r3 r2 r1 r0 GND GND r2r
xr2r_Gxhz gdacxhz g7 g6 g5 g4 g3 g2 g1 g0 GND GND r2r
xr2r_Bxhz bdacxhz b7 b6 b5 b4 b3 b2 b1 b0 GND GND r2r

xdacboost_r rout rdac vcc GND dacboost
xdacboost_g gout gdac vcc GND dacboost
xdacboost_b bout bdac vcc GND dacboost

* Simulate tt output path load...
*NOTE: According to @tnt it is better to model 2.5pF (to GND)
* either side of the resistor, but because the digital model
* has zero impedance (I think), I will be more conservative
* and do it with 5pF just at the final output node...
*Cr1 red             GND 2.5p
Rr1 rout            routpin 500
Cr2 routpin         GND 5p

*Cg1 green           GND 2.5p
Rg1 gout            goutpin 500
Cg2 goutpin         GND 5p

*Cb1 blue            GND 2.5p
Rb1 bout            boutpin 500
Cb2 boutpin         GND 5p

Rrhz1 rdachz        rdachzpin 500
Crhz2 rdachzpin     GND 5p
Rghz1 gdachz        gdachzpin 500
Cghz2 gdachzpin     GND 5p
Rbhz1 bdachz        bdachzpin 500
Cbhz2 bdachzpin     GND 5p

Rrhhz1 rdachhz        rdachhzpin 5500
Crhhz2 rdachhzpin     GND 5p
Rghhz1 gdachhz        gdachhzpin 5500
Cghhz2 gdachhzpin     GND 5p
Rbhhz1 bdachhz        bdachhzpin 5500
Cbhhz2 bdachhzpin     GND 5p

Rrxhz1 rdacxhz        rdacxhzpin 65500
Crxhz2 rdacxhzpin     GND 7p
Rgxhz1 gdacxhz        gdacxhzpin 65500
Cgxhz2 gdacxhzpin     GND 7p
Rbxhz1 bdacxhz        bdacxhzpin 65500
Cbxhz2 bdacxhzpin     GND 7p


**** End of the ADC and its subcircuits.  Begin test circuit ****

.param vcc=1.8
vcc vcc 0 {vcc}

* Digital clock signal

aclock 0 clk clock
.model clock d_osc cntl_array=[-1 1] freq_array=[25Meg 25Meg]

* reset signal

Vreset rst_n GND PULSE 1.8 0 40n 1n 1n 120n 34m ;256u

* DAC input value
.param rise=    1n
.param fall=    1n
.param h0=  40n-1n
.param h1=  80n-1n
.param h2= 160n-1n
.param h3= 320n-1n
.param h4= 640n-1n
.param h5=1280n-1n
.param h6=2560n-1n
.param h7=5120n-1n

* --- Mode 3: XOR ---
* Vin0 in0 GND dc 0.0 ; PULSE    0.0  1.8    2u {rise} {fall} {h0}    80n
* Vin1 in1 GND dc 0.0 ; PULSE    0.0  1.8    2u {rise} {fall} {h1}   160n
* Vin2 in2 GND dc 0.0 ; PULSE    0.0  1.8    2u {rise} {fall} {h2}   320n
* Vin3 in3 GND dc 0.0 ; PULSE    0.0  1.8    2u {rise} {fall} {h3}   640n
* Vin4 in4 GND dc 1.8 ; PULSE    1.8  0.0    2u {rise} {fall} {h4}  1280n
* Vin5 in5 GND dc 1.8 ; PULSE    1.8  0.0    2u {rise} {fall} {h5}  2560n
* Vin6 in6 GND dc 0.0 ; PULSE    0.0  1.8    2u {rise} {fall} {h6}  5120n
* Vin7 in7 GND dc 0.0 ; PULSE    0.0  1.8    2u {rise} {fall} {h7} 10240n

* --- Mode 1: RAMP ---
Vin0 in0 GND dc 0.0 ; Primary...
Vin1 in1 GND dc 0.0 ; ...= 0 (Red primary, Green secondary, Blue fade)
Vin2 in2 GND dc 0.0 ; Divider...
Vin3 in3 GND dc 0.0 ; ...= 0 (none)
Vin4 in4 GND dc 1.8 ; Mode...
Vin5 in5 GND dc 0.0 ; ...
Vin6 in6 GND dc 0.0 ; ...= 001 (ramp tests)
Vin7 in7 GND dc 0.0 ; Timing = 0 (standard VGA)


.control
  tran 8n 16.8m 0 8n UIC
  * let r_digi = (r7/2)+(r6/4)+(r5/8)+(r4/16)+(r3/32)+(r2/64)+(r1/128)+(r0/256)
  * let g_digi = (g7/2)+(g6/4)+(g5/8)+(g4/16)+(g3/32)+(g2/64)+(g1/128)+(g0/256)
  * let b_digi = (b7/2)+(b6/4)+(b5/8)+(b4/16)+(b3/32)+(b2/64)+(b1/128)+(b0/256)
  * let in_digi = (in7/2)+(in6/4)+(in5/8)+(in4/16)+(in3/32)+(in2/64)+(in1/128)+(in0/256)
  * let s_in0 = in0 + 2
  * let s_in1 = in1 + 4
  * let s_in2 = in2 + 6
  * let s_in3 = in3 + 8
  * let s_in4 = in4 + 10
  * let s_in5 = in5 + 12
  * let s_in6 = in6 + 14
  * let s_in7 = in7 + 16
  * set color2=rgb:F/0/0
  * set color3=rgb:0/F/0
  * set color4=rgb:0/0/F
  * plot in_digi s_in0 s_in1 s_in2 s_in3 s_in4 s_in5 s_in6 s_in7 title 'Digital inputs'
  * plot r_digi g_digi b_digi title 'Digital block outputs'
  * plot red_pin_out green_pin_out blue_pin_out title 'Analog DAC outputs'

  * dac = normal DAC hiZ output into dacboost.
  * out = dacboost output, before TT pin.
  * outpin = dacboost output, after TT pin.
  * dachzpin = unbuffered DAC output, after TT pin.
  * dachhzpin = weak digital drive unbuffered DAC output, after TT pin.
  write mixed.raw
  + v(rdac)
  + v(gdac)
  + v(bdac)
  + v(rdachzpin)
  + v(gdachzpin)
  + v(bdachzpin)
  + v(rdachhzpin)
  + v(gdachhzpin)
  + v(bdachhzpin)
  + v(rdacxhzpin)
  + v(gdacxhzpin)
  + v(bdacxhzpin)
  + v(rout)
  + v(gout)
  + v(bout)
  + v(routpin)
  + v(goutpin)
  + v(boutpin)
  + v(hsync)
  + v(vsync)
  + v(hblank)
  + v(vblank)
  quit
.endc
.end
